magic
tech sky130B
magscale 1 2
timestamp 1680008677
<< viali >>
rect 2421 57477 2455 57511
rect 4077 57477 4111 57511
rect 4997 57477 5031 57511
rect 7573 57477 7607 57511
rect 9229 57477 9263 57511
rect 10149 57477 10183 57511
rect 12725 57477 12759 57511
rect 16957 57477 16991 57511
rect 17877 57477 17911 57511
rect 20453 57477 20487 57511
rect 22109 57477 22143 57511
rect 23029 57477 23063 57511
rect 25605 57477 25639 57511
rect 27261 57477 27295 57511
rect 28181 57477 28215 57511
rect 29837 57477 29871 57511
rect 30757 57477 30791 57511
rect 32413 57477 32447 57511
rect 33333 57477 33367 57511
rect 34989 57477 35023 57511
rect 35909 57477 35943 57511
rect 37565 57477 37599 57511
rect 38485 57477 38519 57511
rect 41061 57477 41095 57511
rect 42717 57477 42751 57511
rect 43637 57477 43671 57511
rect 45293 57477 45327 57511
rect 47869 57477 47903 57511
rect 50445 57477 50479 57511
rect 53941 57477 53975 57511
rect 55597 57477 55631 57511
rect 56425 57477 56459 57511
rect 57161 57477 57195 57511
rect 6561 57409 6595 57443
rect 11713 57409 11747 57443
rect 14289 57409 14323 57443
rect 15209 57409 15243 57443
rect 19441 57409 19475 57443
rect 24593 57409 24627 57443
rect 40049 57409 40083 57443
rect 46121 57409 46155 57443
rect 48697 57409 48731 57443
rect 51273 57409 51307 57443
rect 52929 57409 52963 57443
rect 58173 57409 58207 57443
rect 14565 57341 14599 57375
rect 2605 57273 2639 57307
rect 17141 57273 17175 57307
rect 56609 57273 56643 57307
rect 4169 57205 4203 57239
rect 5089 57205 5123 57239
rect 6745 57205 6779 57239
rect 7665 57205 7699 57239
rect 9321 57205 9355 57239
rect 10241 57205 10275 57239
rect 11897 57205 11931 57239
rect 12817 57205 12851 57239
rect 15393 57205 15427 57239
rect 17969 57205 18003 57239
rect 19625 57205 19659 57239
rect 20545 57205 20579 57239
rect 22201 57205 22235 57239
rect 23121 57205 23155 57239
rect 24777 57205 24811 57239
rect 25697 57205 25731 57239
rect 27353 57205 27387 57239
rect 28273 57205 28307 57239
rect 29929 57205 29963 57239
rect 30849 57205 30883 57239
rect 32505 57205 32539 57239
rect 33425 57205 33459 57239
rect 35081 57205 35115 57239
rect 36001 57205 36035 57239
rect 37657 57205 37691 57239
rect 38577 57205 38611 57239
rect 40233 57205 40267 57239
rect 41153 57205 41187 57239
rect 42809 57205 42843 57239
rect 43729 57205 43763 57239
rect 45385 57205 45419 57239
rect 46305 57205 46339 57239
rect 47961 57205 47995 57239
rect 48881 57205 48915 57239
rect 50537 57205 50571 57239
rect 51457 57205 51491 57239
rect 53113 57205 53147 57239
rect 54033 57205 54067 57239
rect 55689 57205 55723 57239
rect 57253 57205 57287 57239
rect 58265 57205 58299 57239
rect 56057 56797 56091 56831
rect 56793 56797 56827 56831
rect 57805 56797 57839 56831
rect 57069 56729 57103 56763
rect 58173 56729 58207 56763
rect 56241 56661 56275 56695
rect 55873 56389 55907 56423
rect 56609 56389 56643 56423
rect 57345 56389 57379 56423
rect 1593 56321 1627 56355
rect 58173 56321 58207 56355
rect 1869 56253 1903 56287
rect 58357 56253 58391 56287
rect 57529 56185 57563 56219
rect 55965 56117 55999 56151
rect 56701 56117 56735 56151
rect 58265 55845 58299 55879
rect 1593 55709 1627 55743
rect 57437 55709 57471 55743
rect 58081 55709 58115 55743
rect 1869 55641 1903 55675
rect 57529 55573 57563 55607
rect 58265 55369 58299 55403
rect 1685 55233 1719 55267
rect 58081 55233 58115 55267
rect 1961 55029 1995 55063
rect 57437 54621 57471 54655
rect 1685 54553 1719 54587
rect 2053 54553 2087 54587
rect 58173 54553 58207 54587
rect 57529 54485 57563 54519
rect 58265 54485 58299 54519
rect 1685 54145 1719 54179
rect 58081 54145 58115 54179
rect 1961 53941 1995 53975
rect 58265 53941 58299 53975
rect 1685 53465 1719 53499
rect 58173 53465 58207 53499
rect 58357 53465 58391 53499
rect 1961 53397 1995 53431
rect 1685 53057 1719 53091
rect 48237 53057 48271 53091
rect 48421 53057 48455 53091
rect 48789 53057 48823 53091
rect 58081 53057 58115 53091
rect 48697 52989 48731 53023
rect 1961 52853 1995 52887
rect 48053 52853 48087 52887
rect 58265 52853 58299 52887
rect 47685 52649 47719 52683
rect 41797 52445 41831 52479
rect 42165 52445 42199 52479
rect 42349 52445 42383 52479
rect 42441 52445 42475 52479
rect 42533 52445 42567 52479
rect 47869 52445 47903 52479
rect 48053 52445 48087 52479
rect 48421 52445 48455 52479
rect 48513 52445 48547 52479
rect 57897 52445 57931 52479
rect 1685 52377 1719 52411
rect 2053 52377 2087 52411
rect 58173 52377 58207 52411
rect 42717 52309 42751 52343
rect 57345 52037 57379 52071
rect 1593 51969 1627 52003
rect 48237 51969 48271 52003
rect 48421 51969 48455 52003
rect 48789 51969 48823 52003
rect 58081 51969 58115 52003
rect 47777 51901 47811 51935
rect 48697 51901 48731 51935
rect 57529 51833 57563 51867
rect 1777 51765 1811 51799
rect 58265 51765 58299 51799
rect 47409 51493 47443 51527
rect 36921 51357 36955 51391
rect 37069 51357 37103 51391
rect 37289 51357 37323 51391
rect 37427 51357 37461 51391
rect 46857 51357 46891 51391
rect 47277 51357 47311 51391
rect 48421 51357 48455 51391
rect 48697 51357 48731 51391
rect 48789 51357 48823 51391
rect 49065 51357 49099 51391
rect 49249 51357 49283 51391
rect 57345 51357 57379 51391
rect 1685 51289 1719 51323
rect 2053 51289 2087 51323
rect 37197 51289 37231 51323
rect 47041 51289 47075 51323
rect 47133 51289 47167 51323
rect 47961 51289 47995 51323
rect 58173 51289 58207 51323
rect 37565 51221 37599 51255
rect 57529 51221 57563 51255
rect 58265 51221 58299 51255
rect 49709 50949 49743 50983
rect 49801 50949 49835 50983
rect 1685 50881 1719 50915
rect 48053 50881 48087 50915
rect 48237 50881 48271 50915
rect 48605 50881 48639 50915
rect 49433 50881 49467 50915
rect 49526 50881 49560 50915
rect 49898 50881 49932 50915
rect 58173 50881 58207 50915
rect 47593 50813 47627 50847
rect 48513 50813 48547 50847
rect 1961 50677 1995 50711
rect 49065 50677 49099 50711
rect 50077 50677 50111 50711
rect 58265 50677 58299 50711
rect 49065 50337 49099 50371
rect 49433 50337 49467 50371
rect 48973 50269 49007 50303
rect 49341 50269 49375 50303
rect 1685 50201 1719 50235
rect 48329 50201 48363 50235
rect 58173 50201 58207 50235
rect 1961 50133 1995 50167
rect 58265 50133 58299 50167
rect 1685 49793 1719 49827
rect 43085 49793 43119 49827
rect 43269 49793 43303 49827
rect 43637 49793 43671 49827
rect 58173 49793 58207 49827
rect 1961 49725 1995 49759
rect 42625 49725 42659 49759
rect 43545 49725 43579 49759
rect 58357 49725 58391 49759
rect 30205 49181 30239 49215
rect 30481 49181 30515 49215
rect 30573 49181 30607 49215
rect 1685 49113 1719 49147
rect 30389 49113 30423 49147
rect 57989 49113 58023 49147
rect 1961 49045 1995 49079
rect 30757 49045 30791 49079
rect 58081 49045 58115 49079
rect 10241 48773 10275 48807
rect 1685 48705 1719 48739
rect 9965 48705 9999 48739
rect 10149 48705 10183 48739
rect 10338 48705 10372 48739
rect 30757 48705 30791 48739
rect 31033 48705 31067 48739
rect 31125 48705 31159 48739
rect 31401 48705 31435 48739
rect 31585 48705 31619 48739
rect 58081 48705 58115 48739
rect 1777 48501 1811 48535
rect 10517 48501 10551 48535
rect 30389 48501 30423 48535
rect 58265 48501 58299 48535
rect 31033 48093 31067 48127
rect 31181 48093 31215 48127
rect 31401 48093 31435 48127
rect 31498 48093 31532 48127
rect 34897 48093 34931 48127
rect 35173 48093 35207 48127
rect 35265 48093 35299 48127
rect 57161 48093 57195 48127
rect 57897 48093 57931 48127
rect 1685 48025 1719 48059
rect 31309 48025 31343 48059
rect 35081 48025 35115 48059
rect 58173 48025 58207 48059
rect 1777 47957 1811 47991
rect 31677 47957 31711 47991
rect 35449 47957 35483 47991
rect 57345 47957 57379 47991
rect 31125 47685 31159 47719
rect 40969 47685 41003 47719
rect 41613 47685 41647 47719
rect 41705 47685 41739 47719
rect 1593 47617 1627 47651
rect 30757 47617 30791 47651
rect 30850 47617 30884 47651
rect 31033 47617 31067 47651
rect 31263 47617 31297 47651
rect 41337 47617 41371 47651
rect 41485 47617 41519 47651
rect 41802 47617 41836 47651
rect 57253 47617 57287 47651
rect 58081 47617 58115 47651
rect 1777 47413 1811 47447
rect 31401 47413 31435 47447
rect 41981 47413 42015 47447
rect 57437 47413 57471 47447
rect 58265 47413 58299 47447
rect 58265 47141 58299 47175
rect 58081 47005 58115 47039
rect 1685 46937 1719 46971
rect 1869 46937 1903 46971
rect 33149 46597 33183 46631
rect 1593 46529 1627 46563
rect 32321 46529 32355 46563
rect 32505 46529 32539 46563
rect 32597 46529 32631 46563
rect 32689 46529 32723 46563
rect 58173 46529 58207 46563
rect 1777 46325 1811 46359
rect 32873 46325 32907 46359
rect 58265 46325 58299 46359
rect 37013 46121 37047 46155
rect 1593 45917 1627 45951
rect 36461 45917 36495 45951
rect 36829 45917 36863 45951
rect 57897 45917 57931 45951
rect 36645 45849 36679 45883
rect 36737 45849 36771 45883
rect 58173 45849 58207 45883
rect 1777 45781 1811 45815
rect 35633 45509 35667 45543
rect 1593 45441 1627 45475
rect 32321 45441 32355 45475
rect 32414 45441 32448 45475
rect 32597 45441 32631 45475
rect 32689 45441 32723 45475
rect 32786 45441 32820 45475
rect 35357 45441 35391 45475
rect 35541 45441 35575 45475
rect 35725 45441 35759 45475
rect 58173 45441 58207 45475
rect 34989 45373 35023 45407
rect 1777 45237 1811 45271
rect 32965 45237 32999 45271
rect 35909 45237 35943 45271
rect 58265 45237 58299 45271
rect 49157 44897 49191 44931
rect 49341 44897 49375 44931
rect 49065 44829 49099 44863
rect 49433 44829 49467 44863
rect 57253 44829 57287 44863
rect 57897 44829 57931 44863
rect 1685 44761 1719 44795
rect 1869 44761 1903 44795
rect 58173 44761 58207 44795
rect 48697 44693 48731 44727
rect 57345 44693 57379 44727
rect 41981 44421 42015 44455
rect 1593 44353 1627 44387
rect 41429 44353 41463 44387
rect 58081 44353 58115 44387
rect 1777 44149 1811 44183
rect 58265 44149 58299 44183
rect 41337 43741 41371 43775
rect 41613 43741 41647 43775
rect 41705 43741 41739 43775
rect 42625 43741 42659 43775
rect 58081 43741 58115 43775
rect 1685 43673 1719 43707
rect 1869 43673 1903 43707
rect 41521 43673 41555 43707
rect 42441 43673 42475 43707
rect 42901 43673 42935 43707
rect 41889 43605 41923 43639
rect 42809 43605 42843 43639
rect 58265 43605 58299 43639
rect 1593 43265 1627 43299
rect 58081 43265 58115 43299
rect 1777 43061 1811 43095
rect 58265 43061 58299 43095
rect 57989 42653 58023 42687
rect 1685 42585 1719 42619
rect 1777 42517 1811 42551
rect 58265 42517 58299 42551
rect 28089 42245 28123 42279
rect 28181 42245 28215 42279
rect 1685 42177 1719 42211
rect 27905 42177 27939 42211
rect 28273 42177 28307 42211
rect 58357 42177 58391 42211
rect 1777 41973 1811 42007
rect 28457 41973 28491 42007
rect 26985 41701 27019 41735
rect 1593 41565 1627 41599
rect 26433 41565 26467 41599
rect 26709 41565 26743 41599
rect 26853 41565 26887 41599
rect 58357 41565 58391 41599
rect 26617 41497 26651 41531
rect 1777 41429 1811 41463
rect 1593 41089 1627 41123
rect 1777 40885 1811 40919
rect 9689 40613 9723 40647
rect 1869 40545 1903 40579
rect 9137 40477 9171 40511
rect 9413 40477 9447 40511
rect 9557 40477 9591 40511
rect 31401 40477 31435 40511
rect 40233 40477 40267 40511
rect 40325 40477 40359 40511
rect 40509 40477 40543 40511
rect 40601 40477 40635 40511
rect 1685 40409 1719 40443
rect 9321 40409 9355 40443
rect 31217 40409 31251 40443
rect 40049 40409 40083 40443
rect 31493 40341 31527 40375
rect 1685 40069 1719 40103
rect 58357 39865 58391 39899
rect 1777 39797 1811 39831
rect 7941 39525 7975 39559
rect 7389 39389 7423 39423
rect 7665 39389 7699 39423
rect 7809 39389 7843 39423
rect 1685 39321 1719 39355
rect 7573 39321 7607 39355
rect 1777 39253 1811 39287
rect 32965 38981 32999 39015
rect 1685 38913 1719 38947
rect 32689 38913 32723 38947
rect 32873 38913 32907 38947
rect 33057 38913 33091 38947
rect 1869 38777 1903 38811
rect 33241 38709 33275 38743
rect 58357 38709 58391 38743
rect 5273 38437 5307 38471
rect 33425 38369 33459 38403
rect 4721 38301 4755 38335
rect 4905 38301 4939 38335
rect 4997 38301 5031 38335
rect 5094 38301 5128 38335
rect 33149 38301 33183 38335
rect 1685 38233 1719 38267
rect 1777 38165 1811 38199
rect 32965 37893 32999 37927
rect 1685 37825 1719 37859
rect 32689 37825 32723 37859
rect 32873 37825 32907 37859
rect 33062 37825 33096 37859
rect 1869 37689 1903 37723
rect 33241 37621 33275 37655
rect 1869 37281 1903 37315
rect 57897 37213 57931 37247
rect 58173 37213 58207 37247
rect 1685 37145 1719 37179
rect 1685 36737 1719 36771
rect 3617 36737 3651 36771
rect 3709 36737 3743 36771
rect 3985 36737 4019 36771
rect 4261 36737 4295 36771
rect 4445 36737 4479 36771
rect 19717 36737 19751 36771
rect 58081 36737 58115 36771
rect 21465 36669 21499 36703
rect 1869 36601 1903 36635
rect 3249 36533 3283 36567
rect 58265 36533 58299 36567
rect 58173 36193 58207 36227
rect 1593 36125 1627 36159
rect 19901 36125 19935 36159
rect 20177 36125 20211 36159
rect 20269 36125 20303 36159
rect 30389 36125 30423 36159
rect 30665 36125 30699 36159
rect 31033 36125 31067 36159
rect 31401 36125 31435 36159
rect 57897 36125 57931 36159
rect 20085 36057 20119 36091
rect 1777 35989 1811 36023
rect 20453 35989 20487 36023
rect 30481 35989 30515 36023
rect 3249 35785 3283 35819
rect 58173 35717 58207 35751
rect 1685 35649 1719 35683
rect 2421 35649 2455 35683
rect 2697 35649 2731 35683
rect 2881 35649 2915 35683
rect 2973 35649 3007 35683
rect 3065 35649 3099 35683
rect 28181 35649 28215 35683
rect 28273 35649 28307 35683
rect 28457 35649 28491 35683
rect 28549 35649 28583 35683
rect 29101 35649 29135 35683
rect 33241 35649 33275 35683
rect 33333 35649 33367 35683
rect 33517 35649 33551 35683
rect 33609 35649 33643 35683
rect 29377 35581 29411 35615
rect 1869 35513 1903 35547
rect 58357 35513 58391 35547
rect 27997 35445 28031 35479
rect 33057 35445 33091 35479
rect 31033 35241 31067 35275
rect 32413 35173 32447 35207
rect 32965 35173 32999 35207
rect 30481 35037 30515 35071
rect 30849 35037 30883 35071
rect 31861 35037 31895 35071
rect 32229 35037 32263 35071
rect 32873 35037 32907 35071
rect 33149 35037 33183 35071
rect 42257 35037 42291 35071
rect 42717 35037 42751 35071
rect 57897 35037 57931 35071
rect 1685 34969 1719 35003
rect 30665 34969 30699 35003
rect 30757 34969 30791 35003
rect 32045 34969 32079 35003
rect 32137 34969 32171 35003
rect 58173 34969 58207 35003
rect 1777 34901 1811 34935
rect 33333 34901 33367 34935
rect 1777 34697 1811 34731
rect 33425 34697 33459 34731
rect 41153 34697 41187 34731
rect 58265 34697 58299 34731
rect 33793 34629 33827 34663
rect 41705 34629 41739 34663
rect 41797 34629 41831 34663
rect 1685 34561 1719 34595
rect 24317 34561 24351 34595
rect 24685 34561 24719 34595
rect 32505 34561 32539 34595
rect 32653 34561 32687 34595
rect 32781 34561 32815 34595
rect 32873 34561 32907 34595
rect 32970 34561 33004 34595
rect 41521 34561 41555 34595
rect 41889 34561 41923 34595
rect 43269 34561 43303 34595
rect 43637 34561 43671 34595
rect 43729 34561 43763 34595
rect 58081 34561 58115 34595
rect 34161 34493 34195 34527
rect 34345 34493 34379 34527
rect 43177 34493 43211 34527
rect 33149 34425 33183 34459
rect 33931 34425 33965 34459
rect 34069 34425 34103 34459
rect 42073 34425 42107 34459
rect 42717 34357 42751 34391
rect 35265 34153 35299 34187
rect 4537 34085 4571 34119
rect 42809 34085 42843 34119
rect 1869 34017 1903 34051
rect 34897 34017 34931 34051
rect 47961 34017 47995 34051
rect 3985 33949 4019 33983
rect 4261 33949 4295 33983
rect 4358 33949 4392 33983
rect 33885 33949 33919 33983
rect 34069 33949 34103 33983
rect 34161 33949 34195 33983
rect 35081 33949 35115 33983
rect 42993 33949 43027 33983
rect 43085 33949 43119 33983
rect 43269 33949 43303 33983
rect 43361 33949 43395 33983
rect 47869 33949 47903 33983
rect 48237 33949 48271 33983
rect 48329 33949 48363 33983
rect 57897 33949 57931 33983
rect 1685 33881 1719 33915
rect 4169 33881 4203 33915
rect 47225 33881 47259 33915
rect 58173 33881 58207 33915
rect 33983 33813 34017 33847
rect 33241 33609 33275 33643
rect 1869 33541 1903 33575
rect 1685 33473 1719 33507
rect 33241 33473 33275 33507
rect 33609 33473 33643 33507
rect 34161 33473 34195 33507
rect 34713 33473 34747 33507
rect 58081 33473 58115 33507
rect 58265 33269 58299 33303
rect 27905 32861 27939 32895
rect 57897 32861 57931 32895
rect 1685 32793 1719 32827
rect 28365 32793 28399 32827
rect 58173 32793 58207 32827
rect 1777 32725 1811 32759
rect 2237 32453 2271 32487
rect 2329 32453 2363 32487
rect 3065 32453 3099 32487
rect 3617 32453 3651 32487
rect 28273 32453 28307 32487
rect 37565 32453 37599 32487
rect 2053 32385 2087 32419
rect 2421 32385 2455 32419
rect 3341 32385 3375 32419
rect 3434 32385 3468 32419
rect 3709 32385 3743 32419
rect 3806 32385 3840 32419
rect 27905 32385 27939 32419
rect 27998 32385 28032 32419
rect 28181 32385 28215 32419
rect 28411 32385 28445 32419
rect 29009 32385 29043 32419
rect 29285 32385 29319 32419
rect 58081 32385 58115 32419
rect 29561 32317 29595 32351
rect 3985 32249 4019 32283
rect 28549 32249 28583 32283
rect 29101 32249 29135 32283
rect 2605 32181 2639 32215
rect 37841 32181 37875 32215
rect 58265 32181 58299 32215
rect 2513 31977 2547 32011
rect 28181 31977 28215 32011
rect 37105 31977 37139 32011
rect 1869 31909 1903 31943
rect 27353 31909 27387 31943
rect 57253 31841 57287 31875
rect 1685 31773 1719 31807
rect 2421 31773 2455 31807
rect 27629 31773 27663 31807
rect 27813 31773 27847 31807
rect 27905 31773 27939 31807
rect 27997 31773 28031 31807
rect 36461 31773 36495 31807
rect 36609 31773 36643 31807
rect 36737 31773 36771 31807
rect 36829 31773 36863 31807
rect 36967 31773 37001 31807
rect 56977 31773 57011 31807
rect 57897 31773 57931 31807
rect 58173 31705 58207 31739
rect 2605 31433 2639 31467
rect 48237 31365 48271 31399
rect 2053 31297 2087 31331
rect 2237 31297 2271 31331
rect 2329 31297 2363 31331
rect 2421 31297 2455 31331
rect 48053 31297 48087 31331
rect 48329 31297 48363 31331
rect 58081 31297 58115 31331
rect 47869 31093 47903 31127
rect 58265 31093 58299 31127
rect 48145 30889 48179 30923
rect 1685 30685 1719 30719
rect 28273 30685 28307 30719
rect 28366 30685 28400 30719
rect 28738 30685 28772 30719
rect 29745 30685 29779 30719
rect 29838 30685 29872 30719
rect 30251 30685 30285 30719
rect 31585 30685 31619 30719
rect 47593 30685 47627 30719
rect 47777 30685 47811 30719
rect 47961 30685 47995 30719
rect 28549 30617 28583 30651
rect 28641 30617 28675 30651
rect 30021 30617 30055 30651
rect 30113 30617 30147 30651
rect 32137 30617 32171 30651
rect 47869 30617 47903 30651
rect 58173 30617 58207 30651
rect 1777 30549 1811 30583
rect 28917 30549 28951 30583
rect 30389 30549 30423 30583
rect 58265 30549 58299 30583
rect 1685 30277 1719 30311
rect 1869 30277 1903 30311
rect 2789 30277 2823 30311
rect 17141 30277 17175 30311
rect 22845 30277 22879 30311
rect 2605 30209 2639 30243
rect 2881 30209 2915 30243
rect 16865 30209 16899 30243
rect 17049 30209 17083 30243
rect 17233 30209 17267 30243
rect 22753 30209 22787 30243
rect 22937 30209 22971 30243
rect 23075 30209 23109 30243
rect 23213 30209 23247 30243
rect 30297 30209 30331 30243
rect 30389 30209 30423 30243
rect 30757 30209 30791 30243
rect 31217 30209 31251 30243
rect 31493 30209 31527 30243
rect 58081 30209 58115 30243
rect 17417 30073 17451 30107
rect 22569 30073 22603 30107
rect 2421 30005 2455 30039
rect 58265 30005 58299 30039
rect 32689 29801 32723 29835
rect 1869 29733 1903 29767
rect 28549 29733 28583 29767
rect 29837 29733 29871 29767
rect 32597 29733 32631 29767
rect 32321 29665 32355 29699
rect 58173 29665 58207 29699
rect 1685 29597 1719 29631
rect 23213 29597 23247 29631
rect 23857 29597 23891 29631
rect 28457 29597 28491 29631
rect 28733 29597 28767 29631
rect 29745 29597 29779 29631
rect 30021 29597 30055 29631
rect 32781 29597 32815 29631
rect 33057 29597 33091 29631
rect 57897 29597 57931 29631
rect 2421 29529 2455 29563
rect 28181 29529 28215 29563
rect 29193 29529 29227 29563
rect 2513 29461 2547 29495
rect 30205 29461 30239 29495
rect 32965 29461 32999 29495
rect 2622 29257 2656 29291
rect 22477 29257 22511 29291
rect 22753 29257 22787 29291
rect 24317 29257 24351 29291
rect 2237 29189 2271 29223
rect 2329 29189 2363 29223
rect 2053 29121 2087 29155
rect 2426 29121 2460 29155
rect 22109 29121 22143 29155
rect 23213 29121 23247 29155
rect 23489 29121 23523 29155
rect 23765 29121 23799 29155
rect 24501 29121 24535 29155
rect 28457 29121 28491 29155
rect 28641 29121 28675 29155
rect 28733 29121 28767 29155
rect 28825 29121 28859 29155
rect 29653 29121 29687 29155
rect 31309 29121 31343 29155
rect 31585 29121 31619 29155
rect 58081 29121 58115 29155
rect 22201 29053 22235 29087
rect 29929 29053 29963 29087
rect 31493 29053 31527 29087
rect 28181 28985 28215 29019
rect 58265 28985 58299 29019
rect 22293 28917 22327 28951
rect 29009 28917 29043 28951
rect 31309 28917 31343 28951
rect 31769 28917 31803 28951
rect 28917 28713 28951 28747
rect 49065 28645 49099 28679
rect 23121 28577 23155 28611
rect 24041 28577 24075 28611
rect 25722 28577 25756 28611
rect 58173 28577 58207 28611
rect 1685 28509 1719 28543
rect 23489 28509 23523 28543
rect 23581 28509 23615 28543
rect 25237 28509 25271 28543
rect 28641 28509 28675 28543
rect 28825 28509 28859 28543
rect 28917 28509 28951 28543
rect 29837 28509 29871 28543
rect 31585 28509 31619 28543
rect 31769 28509 31803 28543
rect 42257 28509 42291 28543
rect 42441 28509 42475 28543
rect 48421 28509 48455 28543
rect 48569 28509 48603 28543
rect 48927 28509 48961 28543
rect 57897 28509 57931 28543
rect 23029 28441 23063 28475
rect 25605 28441 25639 28475
rect 30205 28441 30239 28475
rect 48697 28441 48731 28475
rect 48789 28441 48823 28475
rect 1777 28373 1811 28407
rect 25513 28373 25547 28407
rect 25881 28373 25915 28407
rect 29101 28373 29135 28407
rect 31861 28373 31895 28407
rect 42533 28373 42567 28407
rect 24317 28169 24351 28203
rect 25605 28169 25639 28203
rect 29101 28169 29135 28203
rect 31401 28169 31435 28203
rect 1685 28101 1719 28135
rect 31125 28101 31159 28135
rect 23213 28033 23247 28067
rect 23397 28033 23431 28067
rect 23765 28033 23799 28067
rect 24501 28033 24535 28067
rect 25053 28033 25087 28067
rect 25513 28033 25547 28067
rect 25605 28033 25639 28067
rect 27169 28033 27203 28067
rect 28549 28033 28583 28067
rect 28733 28033 28767 28067
rect 28825 28033 28859 28067
rect 28917 28033 28951 28067
rect 29653 28033 29687 28067
rect 30757 28033 30791 28067
rect 30850 28033 30884 28067
rect 31033 28033 31067 28067
rect 31222 28033 31256 28067
rect 58081 28033 58115 28067
rect 27353 27965 27387 27999
rect 29929 27965 29963 27999
rect 26065 27897 26099 27931
rect 1777 27829 1811 27863
rect 58265 27829 58299 27863
rect 30297 27557 30331 27591
rect 32505 27557 32539 27591
rect 49617 27557 49651 27591
rect 58173 27489 58207 27523
rect 1685 27421 1719 27455
rect 23121 27421 23155 27455
rect 23489 27421 23523 27455
rect 23581 27421 23615 27455
rect 24041 27421 24075 27455
rect 25421 27421 25455 27455
rect 26617 27421 26651 27455
rect 26801 27421 26835 27455
rect 26985 27421 27019 27455
rect 27077 27421 27111 27455
rect 27445 27421 27479 27455
rect 27721 27421 27755 27455
rect 27997 27421 28031 27455
rect 28135 27421 28169 27455
rect 30481 27421 30515 27455
rect 30665 27421 30699 27455
rect 30849 27421 30883 27455
rect 32229 27421 32263 27455
rect 32321 27421 32355 27455
rect 32965 27421 32999 27455
rect 33517 27421 33551 27455
rect 33977 27421 34011 27455
rect 49065 27421 49099 27455
rect 49438 27421 49472 27455
rect 57897 27421 57931 27455
rect 23029 27353 23063 27387
rect 25789 27353 25823 27387
rect 26709 27353 26743 27387
rect 27905 27353 27939 27387
rect 49249 27353 49283 27387
rect 49341 27353 49375 27387
rect 1777 27285 1811 27319
rect 26433 27285 26467 27319
rect 28273 27285 28307 27319
rect 33726 27285 33760 27319
rect 26065 27081 26099 27115
rect 26249 27081 26283 27115
rect 26341 27081 26375 27115
rect 31033 27081 31067 27115
rect 1685 27013 1719 27047
rect 26157 27013 26191 27047
rect 26525 27013 26559 27047
rect 58173 27013 58207 27047
rect 2421 26945 2455 26979
rect 23029 26945 23063 26979
rect 23397 26945 23431 26979
rect 23489 26945 23523 26979
rect 24869 26945 24903 26979
rect 25053 26945 25087 26979
rect 25145 26945 25179 26979
rect 25238 26945 25272 26979
rect 27997 26945 28031 26979
rect 28549 26945 28583 26979
rect 30481 26945 30515 26979
rect 30665 26945 30699 26979
rect 30757 26945 30791 26979
rect 30849 26945 30883 26979
rect 32781 26945 32815 26979
rect 32965 26945 32999 26979
rect 33149 26945 33183 26979
rect 22937 26877 22971 26911
rect 23949 26877 23983 26911
rect 1869 26809 1903 26843
rect 25513 26809 25547 26843
rect 32597 26809 32631 26843
rect 2513 26741 2547 26775
rect 58265 26741 58299 26775
rect 23489 26537 23523 26571
rect 30665 26537 30699 26571
rect 25053 26469 25087 26503
rect 49617 26469 49651 26503
rect 28365 26401 28399 26435
rect 31493 26401 31527 26435
rect 58173 26401 58207 26435
rect 1593 26333 1627 26367
rect 25237 26333 25271 26367
rect 25461 26333 25495 26367
rect 25605 26333 25639 26367
rect 26525 26333 26559 26367
rect 27905 26333 27939 26367
rect 29745 26333 29779 26367
rect 29929 26333 29963 26367
rect 30021 26333 30055 26367
rect 30113 26333 30147 26367
rect 31585 26333 31619 26367
rect 32045 26333 32079 26367
rect 47869 26333 47903 26367
rect 47962 26333 47996 26367
rect 48237 26333 48271 26367
rect 48334 26333 48368 26367
rect 48973 26333 49007 26367
rect 49121 26333 49155 26367
rect 49438 26333 49472 26367
rect 57897 26333 57931 26367
rect 1869 26265 1903 26299
rect 23397 26265 23431 26299
rect 25339 26265 25373 26299
rect 26341 26265 26375 26299
rect 26893 26265 26927 26299
rect 48145 26265 48179 26299
rect 49249 26265 49283 26299
rect 49341 26265 49375 26299
rect 30297 26197 30331 26231
rect 48513 26197 48547 26231
rect 24593 25993 24627 26027
rect 21189 25925 21223 25959
rect 22937 25925 22971 25959
rect 23489 25925 23523 25959
rect 28549 25925 28583 25959
rect 43545 25925 43579 25959
rect 43637 25925 43671 25959
rect 58173 25925 58207 25959
rect 1593 25857 1627 25891
rect 21005 25857 21039 25891
rect 21465 25857 21499 25891
rect 23029 25857 23063 25891
rect 23397 25857 23431 25891
rect 24501 25857 24535 25891
rect 27169 25857 27203 25891
rect 28181 25857 28215 25891
rect 30113 25857 30147 25891
rect 30205 25857 30239 25891
rect 30389 25857 30423 25891
rect 37657 25857 37691 25891
rect 38577 25857 38611 25891
rect 43269 25857 43303 25891
rect 43417 25857 43451 25891
rect 43775 25857 43809 25891
rect 1777 25789 1811 25823
rect 23949 25789 23983 25823
rect 27445 25789 27479 25823
rect 30573 25789 30607 25823
rect 37841 25789 37875 25823
rect 38853 25789 38887 25823
rect 43913 25653 43947 25687
rect 58265 25653 58299 25687
rect 2697 25449 2731 25483
rect 23489 25449 23523 25483
rect 37933 25449 37967 25483
rect 22753 25381 22787 25415
rect 23305 25313 23339 25347
rect 24961 25313 24995 25347
rect 28641 25313 28675 25347
rect 1593 25245 1627 25279
rect 2513 25245 2547 25279
rect 2667 25245 2701 25279
rect 23213 25245 23247 25279
rect 24685 25245 24719 25279
rect 27169 25245 27203 25279
rect 27353 25245 27387 25279
rect 27537 25245 27571 25279
rect 28181 25245 28215 25279
rect 28273 25245 28307 25279
rect 28457 25245 28491 25279
rect 29745 25245 29779 25279
rect 37289 25245 37323 25279
rect 37437 25245 37471 25279
rect 37657 25245 37691 25279
rect 37795 25245 37829 25279
rect 46029 25245 46063 25279
rect 46177 25245 46211 25279
rect 46397 25245 46431 25279
rect 46494 25245 46528 25279
rect 47133 25245 47167 25279
rect 47226 25245 47260 25279
rect 47409 25245 47443 25279
rect 47501 25245 47535 25279
rect 47598 25245 47632 25279
rect 48421 25245 48455 25279
rect 57897 25245 57931 25279
rect 1869 25177 1903 25211
rect 22753 25177 22787 25211
rect 27445 25177 27479 25211
rect 37565 25177 37599 25211
rect 46305 25177 46339 25211
rect 48237 25177 48271 25211
rect 58173 25177 58207 25211
rect 27721 25109 27755 25143
rect 31033 25109 31067 25143
rect 46673 25109 46707 25143
rect 47777 25109 47811 25143
rect 48513 25109 48547 25143
rect 24225 24905 24259 24939
rect 38025 24905 38059 24939
rect 22293 24837 22327 24871
rect 25605 24837 25639 24871
rect 30481 24837 30515 24871
rect 47777 24837 47811 24871
rect 1593 24769 1627 24803
rect 2513 24769 2547 24803
rect 2606 24769 2640 24803
rect 22109 24769 22143 24803
rect 23305 24769 23339 24803
rect 23581 24769 23615 24803
rect 24041 24769 24075 24803
rect 24593 24769 24627 24803
rect 25237 24769 25271 24803
rect 27537 24769 27571 24803
rect 27721 24769 27755 24803
rect 27813 24769 27847 24803
rect 27997 24769 28031 24803
rect 28089 24769 28123 24803
rect 28733 24769 28767 24803
rect 37473 24769 37507 24803
rect 37657 24769 37691 24803
rect 37749 24769 37783 24803
rect 37841 24769 37875 24803
rect 47961 24769 47995 24803
rect 58081 24769 58115 24803
rect 1777 24701 1811 24735
rect 22385 24701 22419 24735
rect 2881 24633 2915 24667
rect 58265 24633 58299 24667
rect 48053 24565 48087 24599
rect 2697 24361 2731 24395
rect 28825 24361 28859 24395
rect 30389 24361 30423 24395
rect 47685 24361 47719 24395
rect 1593 24157 1627 24191
rect 2513 24157 2547 24191
rect 2667 24157 2701 24191
rect 23121 24157 23155 24191
rect 23489 24157 23523 24191
rect 24041 24157 24075 24191
rect 28181 24157 28215 24191
rect 28274 24157 28308 24191
rect 28457 24157 28491 24191
rect 28549 24157 28583 24191
rect 28646 24157 28680 24191
rect 29745 24157 29779 24191
rect 29838 24157 29872 24191
rect 30251 24157 30285 24191
rect 37289 24157 37323 24191
rect 37473 24157 37507 24191
rect 37657 24157 37691 24191
rect 40785 24157 40819 24191
rect 47041 24157 47075 24191
rect 47189 24157 47223 24191
rect 47547 24157 47581 24191
rect 57897 24157 57931 24191
rect 1869 24089 1903 24123
rect 23029 24089 23063 24123
rect 23581 24089 23615 24123
rect 30021 24089 30055 24123
rect 30113 24089 30147 24123
rect 37565 24089 37599 24123
rect 47317 24089 47351 24123
rect 47409 24089 47443 24123
rect 58173 24089 58207 24123
rect 37841 24021 37875 24055
rect 40969 24021 41003 24055
rect 16129 23817 16163 23851
rect 24409 23817 24443 23851
rect 36829 23817 36863 23851
rect 1593 23681 1627 23715
rect 15761 23681 15795 23715
rect 15915 23681 15949 23715
rect 23489 23681 23523 23715
rect 23765 23681 23799 23715
rect 24041 23681 24075 23715
rect 24409 23681 24443 23715
rect 34161 23681 34195 23715
rect 34345 23681 34379 23715
rect 36645 23681 36679 23715
rect 38393 23681 38427 23715
rect 39129 23681 39163 23715
rect 40233 23681 40267 23715
rect 40969 23681 41003 23715
rect 41705 23681 41739 23715
rect 41889 23681 41923 23715
rect 58081 23681 58115 23715
rect 1777 23613 1811 23647
rect 39313 23545 39347 23579
rect 41153 23545 41187 23579
rect 58265 23545 58299 23579
rect 34161 23477 34195 23511
rect 38577 23477 38611 23511
rect 40417 23477 40451 23511
rect 41797 23477 41831 23511
rect 36645 23273 36679 23307
rect 40233 23273 40267 23307
rect 42901 23273 42935 23307
rect 2881 23205 2915 23239
rect 38025 23205 38059 23239
rect 56517 23205 56551 23239
rect 37105 23137 37139 23171
rect 37197 23137 37231 23171
rect 51549 23137 51583 23171
rect 1593 23069 1627 23103
rect 2513 23069 2547 23103
rect 2667 23069 2701 23103
rect 29745 23069 29779 23103
rect 30481 23069 30515 23103
rect 30665 23069 30699 23103
rect 33241 23069 33275 23103
rect 33977 23069 34011 23103
rect 34897 23069 34931 23103
rect 35909 23069 35943 23103
rect 37841 23069 37875 23103
rect 39129 23069 39163 23103
rect 39221 23069 39255 23103
rect 39313 23069 39347 23103
rect 39497 23069 39531 23103
rect 40049 23069 40083 23103
rect 40785 23069 40819 23103
rect 41889 23069 41923 23103
rect 41981 23069 42015 23103
rect 42073 23069 42107 23103
rect 42257 23069 42291 23103
rect 42717 23069 42751 23103
rect 48237 23069 48271 23103
rect 48605 23069 48639 23103
rect 51733 23069 51767 23103
rect 56149 23069 56183 23103
rect 56333 23069 56367 23103
rect 56977 23069 57011 23103
rect 57897 23069 57931 23103
rect 1869 23001 1903 23035
rect 30573 23001 30607 23035
rect 37013 23001 37047 23035
rect 48421 23001 48455 23035
rect 48513 23001 48547 23035
rect 57253 23001 57287 23035
rect 58173 23001 58207 23035
rect 29929 22933 29963 22967
rect 33425 22933 33459 22967
rect 34161 22933 34195 22967
rect 35081 22933 35115 22967
rect 36093 22933 36127 22967
rect 38853 22933 38887 22967
rect 40969 22933 41003 22967
rect 41613 22933 41647 22967
rect 48789 22933 48823 22967
rect 51917 22933 51951 22967
rect 2513 22729 2547 22763
rect 33149 22729 33183 22763
rect 33793 22729 33827 22763
rect 37657 22729 37691 22763
rect 40509 22729 40543 22763
rect 42809 22729 42843 22763
rect 45477 22729 45511 22763
rect 46581 22729 46615 22763
rect 46673 22729 46707 22763
rect 49893 22729 49927 22763
rect 51641 22729 51675 22763
rect 58265 22729 58299 22763
rect 22385 22661 22419 22695
rect 24133 22661 24167 22695
rect 34713 22661 34747 22695
rect 38752 22661 38786 22695
rect 2237 22593 2271 22627
rect 29561 22593 29595 22627
rect 30297 22593 30331 22627
rect 32781 22593 32815 22627
rect 33609 22593 33643 22627
rect 34897 22593 34931 22627
rect 35541 22593 35575 22627
rect 35797 22593 35831 22627
rect 37473 22593 37507 22627
rect 38485 22593 38519 22627
rect 40325 22593 40359 22627
rect 41613 22593 41647 22627
rect 41705 22593 41739 22627
rect 41797 22593 41831 22627
rect 41981 22593 42015 22627
rect 42625 22593 42659 22627
rect 43361 22593 43395 22627
rect 44353 22593 44387 22627
rect 48780 22593 48814 22627
rect 51089 22593 51123 22627
rect 51273 22593 51307 22627
rect 51365 22593 51399 22627
rect 51457 22593 51491 22627
rect 53113 22593 53147 22627
rect 56241 22593 56275 22627
rect 58081 22593 58115 22627
rect 31033 22525 31067 22559
rect 32689 22525 32723 22559
rect 44097 22525 44131 22559
rect 46765 22525 46799 22559
rect 48513 22525 48547 22559
rect 52929 22525 52963 22559
rect 56517 22525 56551 22559
rect 31401 22457 31435 22491
rect 36921 22457 36955 22491
rect 29745 22389 29779 22423
rect 30481 22389 30515 22423
rect 31493 22389 31527 22423
rect 35081 22389 35115 22423
rect 39865 22389 39899 22423
rect 41337 22389 41371 22423
rect 43545 22389 43579 22423
rect 46213 22389 46247 22423
rect 53297 22389 53331 22423
rect 2697 22185 2731 22219
rect 29101 22185 29135 22219
rect 31585 22185 31619 22219
rect 32229 22185 32263 22219
rect 35449 22185 35483 22219
rect 48881 22185 48915 22219
rect 53113 22185 53147 22219
rect 54125 22185 54159 22219
rect 58265 22185 58299 22219
rect 22201 22117 22235 22151
rect 38761 22117 38795 22151
rect 47133 22117 47167 22151
rect 1777 22049 1811 22083
rect 42073 22049 42107 22083
rect 43453 22049 43487 22083
rect 47685 22049 47719 22083
rect 1593 21981 1627 22015
rect 2513 21981 2547 22015
rect 2606 21981 2640 22015
rect 22017 21981 22051 22015
rect 22477 21981 22511 22015
rect 26249 21981 26283 22015
rect 27997 21981 28031 22015
rect 28917 21981 28951 22015
rect 30297 21981 30331 22015
rect 31217 21981 31251 22015
rect 31401 21981 31435 22015
rect 32045 21981 32079 22015
rect 32781 21981 32815 22015
rect 33517 21981 33551 22015
rect 35705 21981 35739 22015
rect 35817 21981 35851 22015
rect 35930 21978 35964 22012
rect 36093 21981 36127 22015
rect 36553 21981 36587 22015
rect 37289 21981 37323 22015
rect 37933 21981 37967 22015
rect 39037 21981 39071 22015
rect 39126 21975 39160 22009
rect 39242 21981 39276 22015
rect 39405 21981 39439 22015
rect 40049 21981 40083 22015
rect 41337 21981 41371 22015
rect 42349 21981 42383 22015
rect 45201 21981 45235 22015
rect 48605 21981 48639 22015
rect 48697 21981 48731 22015
rect 51733 21981 51767 22015
rect 53573 21981 53607 22015
rect 53941 21981 53975 22015
rect 55873 21981 55907 22015
rect 57713 21981 57747 22015
rect 57989 21981 58023 22015
rect 58081 21981 58115 22015
rect 31033 21913 31067 21947
rect 38117 21913 38151 21947
rect 38301 21913 38335 21947
rect 40969 21913 41003 21947
rect 41153 21913 41187 21947
rect 44189 21913 44223 21947
rect 44373 21913 44407 21947
rect 45446 21913 45480 21947
rect 47501 21913 47535 21947
rect 47593 21913 47627 21947
rect 52000 21913 52034 21947
rect 53757 21913 53791 21947
rect 53849 21913 53883 21947
rect 56118 21913 56152 21947
rect 57897 21913 57931 21947
rect 26433 21845 26467 21879
rect 28181 21845 28215 21879
rect 30481 21845 30515 21879
rect 31309 21845 31343 21879
rect 32965 21845 32999 21879
rect 33701 21845 33735 21879
rect 36737 21845 36771 21879
rect 37381 21845 37415 21879
rect 40233 21845 40267 21879
rect 44557 21845 44591 21879
rect 46581 21845 46615 21879
rect 57253 21845 57287 21879
rect 24777 21641 24811 21675
rect 28273 21641 28307 21675
rect 30297 21641 30331 21675
rect 30941 21641 30975 21675
rect 35265 21641 35299 21675
rect 36737 21641 36771 21675
rect 41705 21641 41739 21675
rect 45569 21641 45603 21675
rect 54309 21641 54343 21675
rect 55689 21641 55723 21675
rect 23305 21573 23339 21607
rect 23397 21573 23431 21607
rect 23949 21573 23983 21607
rect 41521 21573 41555 21607
rect 44741 21573 44775 21607
rect 53196 21573 53230 21607
rect 1593 21505 1627 21539
rect 22109 21505 22143 21539
rect 23765 21505 23799 21539
rect 23857 21505 23891 21539
rect 24685 21505 24719 21539
rect 26341 21505 26375 21539
rect 27813 21505 27847 21539
rect 28917 21505 28951 21539
rect 29929 21505 29963 21539
rect 31125 21505 31159 21539
rect 31309 21505 31343 21539
rect 32321 21505 32355 21539
rect 33324 21505 33358 21539
rect 35081 21505 35115 21539
rect 35817 21505 35851 21539
rect 36553 21505 36587 21539
rect 37473 21505 37507 21539
rect 38209 21505 38243 21539
rect 39129 21505 39163 21539
rect 39385 21505 39419 21539
rect 41337 21505 41371 21539
rect 42625 21505 42659 21539
rect 42881 21505 42915 21539
rect 44557 21505 44591 21539
rect 45937 21505 45971 21539
rect 48789 21505 48823 21539
rect 48973 21505 49007 21539
rect 55413 21505 55447 21539
rect 55505 21505 55539 21539
rect 56405 21505 56439 21539
rect 58081 21505 58115 21539
rect 1777 21437 1811 21471
rect 22661 21437 22695 21471
rect 29009 21437 29043 21471
rect 29285 21437 29319 21471
rect 29837 21437 29871 21471
rect 31217 21437 31251 21471
rect 31401 21437 31435 21471
rect 33057 21437 33091 21471
rect 46029 21437 46063 21471
rect 46213 21437 46247 21471
rect 52929 21437 52963 21471
rect 56149 21437 56183 21471
rect 28181 21369 28215 21403
rect 37657 21369 37691 21403
rect 44925 21369 44959 21403
rect 26525 21301 26559 21335
rect 32505 21301 32539 21335
rect 34437 21301 34471 21335
rect 36001 21301 36035 21335
rect 38393 21301 38427 21335
rect 40509 21301 40543 21335
rect 44005 21301 44039 21335
rect 48789 21301 48823 21335
rect 57529 21301 57563 21335
rect 58265 21301 58299 21335
rect 23213 21097 23247 21131
rect 23949 21097 23983 21131
rect 25421 21097 25455 21131
rect 27353 21097 27387 21131
rect 31125 21097 31159 21131
rect 33057 21097 33091 21131
rect 33701 21097 33735 21131
rect 36277 21097 36311 21131
rect 36921 21097 36955 21131
rect 37657 21097 37691 21131
rect 43637 21097 43671 21131
rect 45201 21097 45235 21131
rect 49801 21097 49835 21131
rect 55781 21097 55815 21131
rect 58265 21097 58299 21131
rect 28549 21029 28583 21063
rect 29101 21029 29135 21063
rect 1777 20961 1811 20995
rect 34897 20961 34931 20995
rect 39017 20961 39051 20995
rect 56885 20961 56919 20995
rect 1593 20893 1627 20927
rect 22017 20893 22051 20927
rect 22477 20893 22511 20927
rect 23029 20893 23063 20927
rect 23765 20893 23799 20927
rect 25237 20893 25271 20927
rect 25973 20893 26007 20927
rect 27905 20893 27939 20927
rect 28089 20893 28123 20927
rect 28825 20893 28859 20927
rect 28917 20893 28951 20927
rect 29745 20893 29779 20927
rect 31677 20893 31711 20927
rect 33517 20893 33551 20927
rect 35164 20893 35198 20927
rect 36737 20893 36771 20927
rect 37473 20893 37507 20927
rect 38209 20893 38243 20927
rect 39221 20893 39255 20927
rect 40049 20893 40083 20927
rect 40785 20893 40819 20927
rect 41521 20893 41555 20927
rect 42625 20893 42659 20927
rect 43913 20893 43947 20927
rect 44005 20893 44039 20927
rect 44097 20893 44131 20927
rect 44281 20893 44315 20927
rect 45477 20893 45511 20927
rect 45569 20893 45603 20927
rect 45661 20893 45695 20927
rect 45845 20893 45879 20927
rect 48421 20893 48455 20927
rect 48688 20893 48722 20927
rect 55965 20893 55999 20927
rect 56425 20893 56459 20927
rect 57141 20893 57175 20927
rect 22201 20825 22235 20859
rect 26240 20825 26274 20859
rect 28733 20825 28767 20859
rect 30012 20825 30046 20859
rect 31944 20825 31978 20859
rect 38945 20825 38979 20859
rect 39129 20825 39163 20859
rect 41797 20825 41831 20859
rect 42809 20825 42843 20859
rect 56057 20825 56091 20859
rect 56149 20825 56183 20859
rect 56287 20825 56321 20859
rect 27997 20757 28031 20791
rect 38393 20757 38427 20791
rect 40233 20757 40267 20791
rect 40969 20757 41003 20791
rect 42993 20757 43027 20791
rect 26617 20553 26651 20587
rect 29285 20553 29319 20587
rect 37657 20553 37691 20587
rect 46121 20553 46155 20587
rect 47961 20553 47995 20587
rect 48973 20553 49007 20587
rect 49157 20553 49191 20587
rect 51457 20553 51491 20587
rect 53113 20553 53147 20587
rect 23673 20485 23707 20519
rect 28172 20485 28206 20519
rect 38669 20485 38703 20519
rect 40018 20485 40052 20519
rect 56149 20485 56183 20519
rect 1593 20417 1627 20451
rect 24317 20417 24351 20451
rect 24409 20417 24443 20451
rect 24685 20417 24719 20451
rect 24777 20417 24811 20451
rect 26249 20417 26283 20451
rect 27169 20417 27203 20451
rect 30021 20417 30055 20451
rect 32597 20417 32631 20451
rect 33333 20417 33367 20451
rect 33600 20417 33634 20451
rect 35265 20417 35299 20451
rect 36737 20417 36771 20451
rect 37473 20417 37507 20451
rect 38945 20417 38979 20451
rect 39037 20417 39071 20451
rect 39129 20417 39163 20451
rect 39313 20417 39347 20451
rect 39773 20417 39807 20451
rect 41705 20417 41739 20451
rect 42625 20417 42659 20451
rect 42809 20417 42843 20451
rect 43269 20417 43303 20451
rect 43536 20417 43570 20451
rect 45201 20417 45235 20451
rect 45937 20417 45971 20451
rect 47958 20417 47992 20451
rect 48329 20417 48363 20451
rect 49154 20417 49188 20451
rect 50077 20417 50111 20451
rect 50333 20417 50367 20451
rect 52193 20417 52227 20451
rect 52377 20417 52411 20451
rect 53110 20417 53144 20451
rect 56057 20417 56091 20451
rect 56241 20417 56275 20451
rect 56359 20417 56393 20451
rect 56517 20417 56551 20451
rect 58173 20417 58207 20451
rect 1777 20349 1811 20383
rect 26341 20349 26375 20383
rect 27905 20349 27939 20383
rect 30297 20349 30331 20383
rect 31677 20349 31711 20383
rect 36553 20349 36587 20383
rect 48421 20349 48455 20383
rect 49617 20349 49651 20383
rect 53573 20349 53607 20383
rect 32781 20281 32815 20315
rect 42717 20281 42751 20315
rect 47777 20281 47811 20315
rect 49525 20281 49559 20315
rect 52193 20281 52227 20315
rect 27353 20213 27387 20247
rect 34713 20213 34747 20247
rect 35449 20213 35483 20247
rect 36921 20213 36955 20247
rect 41153 20213 41187 20247
rect 41889 20213 41923 20247
rect 44649 20213 44683 20247
rect 45385 20213 45419 20247
rect 52929 20213 52963 20247
rect 53481 20213 53515 20247
rect 55873 20213 55907 20247
rect 58265 20213 58299 20247
rect 28457 20009 28491 20043
rect 31217 20009 31251 20043
rect 36921 20009 36955 20043
rect 40417 20009 40451 20043
rect 42901 20009 42935 20043
rect 53849 20009 53883 20043
rect 56241 20009 56275 20043
rect 22017 19941 22051 19975
rect 30481 19941 30515 19975
rect 31953 19941 31987 19975
rect 34345 19941 34379 19975
rect 53389 19941 53423 19975
rect 1777 19873 1811 19907
rect 28633 19873 28667 19907
rect 28825 19873 28859 19907
rect 28917 19873 28951 19907
rect 35265 19873 35299 19907
rect 37565 19873 37599 19907
rect 45385 19873 45419 19907
rect 48053 19873 48087 19907
rect 50905 19873 50939 19907
rect 54493 19873 54527 19907
rect 55873 19873 55907 19907
rect 58173 19873 58207 19907
rect 1593 19805 1627 19839
rect 21833 19805 21867 19839
rect 22293 19805 22327 19839
rect 24685 19805 24719 19839
rect 24869 19805 24903 19839
rect 25421 19805 25455 19839
rect 26341 19805 26375 19839
rect 28722 19805 28756 19839
rect 30297 19805 30331 19839
rect 31033 19805 31067 19839
rect 31769 19805 31803 19839
rect 32965 19805 32999 19839
rect 33232 19805 33266 19839
rect 36550 19805 36584 19839
rect 37007 19805 37041 19839
rect 37657 19805 37691 19839
rect 38485 19805 38519 19839
rect 39221 19805 39255 19839
rect 40233 19805 40267 19839
rect 40877 19805 40911 19839
rect 41613 19805 41647 19839
rect 43177 19805 43211 19839
rect 43269 19805 43303 19839
rect 43361 19805 43395 19839
rect 43545 19805 43579 19839
rect 44281 19805 44315 19839
rect 44373 19805 44407 19839
rect 44465 19805 44499 19839
rect 44649 19805 44683 19839
rect 45201 19805 45235 19839
rect 47777 19805 47811 19839
rect 47869 19805 47903 19839
rect 48145 19805 48179 19839
rect 48513 19805 48547 19839
rect 49065 19805 49099 19839
rect 49157 19805 49191 19839
rect 50534 19805 50568 19839
rect 50997 19805 51031 19839
rect 52009 19805 52043 19839
rect 54030 19805 54064 19839
rect 54401 19805 54435 19839
rect 56057 19805 56091 19839
rect 57897 19805 57931 19839
rect 2605 19737 2639 19771
rect 26608 19737 26642 19771
rect 35817 19737 35851 19771
rect 40049 19737 40083 19771
rect 52254 19737 52288 19771
rect 2697 19669 2731 19703
rect 24685 19669 24719 19703
rect 27721 19669 27755 19703
rect 35449 19669 35483 19703
rect 35541 19669 35575 19703
rect 35633 19669 35667 19703
rect 36369 19669 36403 19703
rect 36553 19669 36587 19703
rect 38025 19669 38059 19703
rect 38669 19669 38703 19703
rect 39405 19669 39439 19703
rect 41061 19669 41095 19703
rect 41797 19669 41831 19703
rect 44005 19669 44039 19703
rect 49341 19669 49375 19703
rect 50353 19669 50387 19703
rect 50537 19669 50571 19703
rect 54033 19669 54067 19703
rect 20637 19465 20671 19499
rect 21373 19465 21407 19499
rect 26525 19465 26559 19499
rect 28457 19465 28491 19499
rect 34621 19465 34655 19499
rect 35265 19465 35299 19499
rect 36093 19465 36127 19499
rect 36185 19465 36219 19499
rect 37571 19465 37605 19499
rect 37657 19465 37691 19499
rect 39589 19465 39623 19499
rect 40233 19465 40267 19499
rect 40969 19465 41003 19499
rect 41153 19465 41187 19499
rect 44189 19465 44223 19499
rect 46581 19465 46615 19499
rect 49709 19465 49743 19499
rect 50261 19465 50295 19499
rect 52101 19465 52135 19499
rect 54309 19465 54343 19499
rect 57161 19465 57195 19499
rect 1869 19397 1903 19431
rect 24409 19397 24443 19431
rect 36369 19397 36403 19431
rect 38476 19397 38510 19431
rect 43821 19397 43855 19431
rect 44005 19397 44039 19431
rect 44916 19397 44950 19431
rect 46857 19397 46891 19431
rect 46949 19397 46983 19431
rect 48596 19397 48630 19431
rect 1593 19329 1627 19363
rect 20453 19329 20487 19363
rect 21189 19329 21223 19363
rect 22017 19329 22051 19363
rect 22845 19329 22879 19363
rect 23121 19329 23155 19363
rect 24041 19329 24075 19363
rect 24134 19329 24168 19363
rect 26341 19329 26375 19363
rect 27353 19329 27387 19363
rect 28273 19329 28307 19363
rect 33241 19329 33275 19363
rect 33508 19329 33542 19363
rect 35081 19329 35115 19363
rect 36001 19329 36035 19363
rect 37473 19329 37507 19363
rect 37749 19329 37783 19363
rect 38209 19329 38243 19363
rect 40049 19329 40083 19363
rect 41094 19329 41128 19363
rect 42625 19329 42659 19363
rect 44649 19329 44683 19363
rect 46765 19329 46799 19363
rect 47087 19329 47121 19363
rect 48329 19329 48363 19363
rect 50169 19329 50203 19363
rect 50353 19329 50387 19363
rect 52009 19329 52043 19363
rect 52193 19329 52227 19363
rect 52929 19329 52963 19363
rect 53185 19329 53219 19363
rect 55781 19329 55815 19363
rect 56037 19329 56071 19363
rect 58173 19329 58207 19363
rect 23305 19261 23339 19295
rect 27445 19261 27479 19295
rect 41613 19261 41647 19295
rect 47225 19261 47259 19295
rect 22937 19193 22971 19227
rect 35817 19193 35851 19227
rect 58357 19193 58391 19227
rect 22201 19125 22235 19159
rect 27721 19125 27755 19159
rect 41521 19125 41555 19159
rect 42809 19125 42843 19159
rect 46029 19125 46063 19159
rect 21097 18921 21131 18955
rect 23213 18921 23247 18955
rect 27077 18921 27111 18955
rect 29745 18921 29779 18955
rect 35173 18921 35207 18955
rect 36553 18921 36587 18955
rect 38393 18921 38427 18955
rect 40233 18921 40267 18955
rect 44557 18921 44591 18955
rect 47317 18921 47351 18955
rect 33517 18853 33551 18887
rect 37381 18853 37415 18887
rect 20913 18785 20947 18819
rect 21925 18785 21959 18819
rect 25881 18785 25915 18819
rect 41705 18785 41739 18819
rect 43821 18785 43855 18819
rect 48513 18785 48547 18819
rect 49065 18785 49099 18819
rect 55689 18785 55723 18819
rect 58173 18785 58207 18819
rect 1593 18717 1627 18751
rect 20821 18717 20855 18751
rect 21649 18717 21683 18751
rect 24777 18717 24811 18751
rect 25053 18717 25087 18751
rect 25237 18717 25271 18751
rect 25697 18717 25731 18751
rect 26893 18717 26927 18751
rect 27629 18717 27663 18751
rect 29929 18717 29963 18751
rect 30205 18717 30239 18751
rect 32321 18717 32355 18751
rect 32505 18717 32539 18751
rect 33333 18717 33367 18751
rect 34069 18717 34103 18751
rect 34989 18717 35023 18751
rect 35725 18717 35759 18751
rect 35909 18717 35943 18751
rect 37197 18717 37231 18751
rect 38669 18717 38703 18751
rect 38761 18717 38795 18751
rect 38853 18717 38887 18751
rect 39037 18717 39071 18751
rect 40049 18717 40083 18751
rect 41429 18717 41463 18751
rect 41981 18717 42015 18751
rect 42073 18717 42107 18751
rect 42717 18717 42751 18751
rect 43637 18717 43671 18751
rect 44373 18717 44407 18751
rect 48605 18717 48639 18751
rect 48973 18717 49007 18751
rect 55873 18717 55907 18751
rect 56062 18717 56096 18751
rect 56977 18717 57011 18751
rect 57897 18717 57931 18751
rect 1869 18649 1903 18683
rect 35817 18649 35851 18683
rect 36369 18649 36403 18683
rect 46949 18649 46983 18683
rect 47133 18649 47167 18683
rect 47961 18649 47995 18683
rect 55689 18649 55723 18683
rect 55965 18649 55999 18683
rect 57253 18649 57287 18683
rect 24593 18581 24627 18615
rect 27813 18581 27847 18615
rect 30113 18581 30147 18615
rect 32413 18581 32447 18615
rect 34253 18581 34287 18615
rect 36569 18581 36603 18615
rect 36737 18581 36771 18615
rect 43177 18581 43211 18615
rect 43545 18581 43579 18615
rect 29653 18377 29687 18411
rect 34897 18377 34931 18411
rect 36829 18377 36863 18411
rect 39129 18377 39163 18411
rect 40325 18377 40359 18411
rect 45017 18377 45051 18411
rect 45385 18377 45419 18411
rect 50905 18377 50939 18411
rect 55873 18377 55907 18411
rect 36093 18309 36127 18343
rect 56701 18309 56735 18343
rect 56977 18309 57011 18343
rect 1593 18241 1627 18275
rect 24225 18241 24259 18275
rect 25513 18241 25547 18275
rect 26341 18241 26375 18275
rect 28733 18241 28767 18275
rect 29469 18241 29503 18275
rect 30205 18241 30239 18275
rect 30389 18241 30423 18275
rect 32413 18241 32447 18275
rect 33149 18241 33183 18275
rect 33885 18241 33919 18275
rect 34713 18241 34747 18275
rect 35909 18241 35943 18275
rect 36645 18241 36679 18275
rect 37473 18241 37507 18275
rect 38209 18241 38243 18275
rect 38945 18241 38979 18275
rect 40147 18241 40181 18275
rect 40877 18241 40911 18275
rect 41705 18241 41739 18275
rect 41889 18241 41923 18275
rect 44005 18241 44039 18275
rect 44373 18241 44407 18275
rect 48421 18241 48455 18275
rect 48789 18241 48823 18275
rect 48973 18241 49007 18275
rect 49433 18241 49467 18275
rect 55781 18241 55815 18275
rect 55965 18241 55999 18275
rect 56885 18241 56919 18275
rect 57074 18263 57108 18297
rect 58081 18241 58115 18275
rect 1777 18173 1811 18207
rect 24409 18173 24443 18207
rect 25329 18173 25363 18207
rect 25697 18173 25731 18207
rect 35725 18173 35759 18207
rect 43913 18173 43947 18207
rect 44465 18173 44499 18207
rect 45477 18173 45511 18207
rect 45661 18173 45695 18207
rect 48513 18173 48547 18207
rect 2421 18105 2455 18139
rect 34069 18105 34103 18139
rect 38393 18105 38427 18139
rect 41061 18105 41095 18139
rect 58265 18105 58299 18139
rect 24961 18037 24995 18071
rect 26341 18037 26375 18071
rect 28917 18037 28951 18071
rect 30205 18037 30239 18071
rect 32597 18037 32631 18071
rect 33333 18037 33367 18071
rect 37657 18037 37691 18071
rect 42073 18037 42107 18071
rect 43453 18037 43487 18071
rect 47869 18037 47903 18071
rect 56701 18037 56735 18071
rect 2421 17833 2455 17867
rect 38669 17833 38703 17867
rect 39405 17833 39439 17867
rect 43637 17833 43671 17867
rect 46305 17833 46339 17867
rect 49065 17833 49099 17867
rect 58265 17833 58299 17867
rect 24685 17765 24719 17799
rect 29929 17765 29963 17799
rect 34253 17765 34287 17799
rect 36921 17765 36955 17799
rect 28457 17697 28491 17731
rect 28917 17697 28951 17731
rect 36001 17697 36035 17731
rect 36277 17697 36311 17731
rect 40417 17697 40451 17731
rect 47409 17697 47443 17731
rect 47961 17697 47995 17731
rect 56885 17697 56919 17731
rect 1593 17629 1627 17663
rect 17877 17629 17911 17663
rect 18061 17629 18095 17663
rect 20545 17629 20579 17663
rect 21281 17629 21315 17663
rect 21465 17629 21499 17663
rect 24593 17629 24627 17663
rect 24869 17629 24903 17663
rect 25789 17629 25823 17663
rect 25973 17629 26007 17663
rect 26157 17629 26191 17663
rect 26801 17629 26835 17663
rect 28549 17629 28583 17663
rect 29745 17629 29779 17663
rect 30481 17629 30515 17663
rect 31493 17629 31527 17663
rect 31677 17629 31711 17663
rect 32137 17629 32171 17663
rect 32873 17629 32907 17663
rect 34897 17629 34931 17663
rect 35909 17629 35943 17663
rect 36737 17629 36771 17663
rect 37473 17629 37507 17663
rect 38485 17629 38519 17663
rect 39221 17629 39255 17663
rect 40141 17629 40175 17663
rect 40233 17629 40267 17663
rect 41061 17629 41095 17663
rect 42257 17629 42291 17663
rect 44281 17629 44315 17663
rect 44649 17629 44683 17663
rect 45661 17629 45695 17663
rect 46121 17629 46155 17663
rect 48053 17629 48087 17663
rect 48421 17629 48455 17663
rect 48605 17629 48639 17663
rect 49065 17629 49099 17663
rect 49249 17629 49283 17663
rect 51917 17629 51951 17663
rect 52101 17629 52135 17663
rect 56241 17629 56275 17663
rect 56425 17629 56459 17663
rect 1869 17561 1903 17595
rect 26065 17561 26099 17595
rect 26893 17561 26927 17595
rect 33140 17561 33174 17595
rect 42524 17561 42558 17595
rect 45293 17561 45327 17595
rect 56333 17561 56367 17595
rect 57130 17561 57164 17595
rect 18061 17493 18095 17527
rect 20729 17493 20763 17527
rect 21373 17493 21407 17527
rect 25053 17493 25087 17527
rect 26341 17493 26375 17527
rect 30665 17493 30699 17527
rect 31585 17493 31619 17527
rect 32321 17493 32355 17527
rect 35081 17493 35115 17527
rect 37657 17493 37691 17527
rect 41245 17493 41279 17527
rect 52009 17493 52043 17527
rect 20361 17289 20395 17323
rect 21005 17289 21039 17323
rect 22201 17289 22235 17323
rect 24133 17289 24167 17323
rect 31677 17289 31711 17323
rect 32505 17289 32539 17323
rect 39589 17289 39623 17323
rect 41613 17289 41647 17323
rect 42625 17289 42659 17323
rect 51733 17289 51767 17323
rect 51917 17289 51951 17323
rect 58265 17289 58299 17323
rect 23765 17221 23799 17255
rect 29000 17221 29034 17255
rect 33784 17221 33818 17255
rect 46397 17221 46431 17255
rect 56241 17221 56275 17255
rect 58173 17221 58207 17255
rect 1593 17153 1627 17187
rect 17601 17153 17635 17187
rect 18337 17153 18371 17187
rect 19993 17153 20027 17187
rect 20821 17153 20855 17187
rect 22017 17153 22051 17187
rect 22937 17153 22971 17187
rect 24225 17153 24259 17187
rect 25145 17153 25179 17187
rect 25513 17153 25547 17187
rect 26341 17153 26375 17187
rect 26617 17153 26651 17187
rect 27353 17153 27387 17187
rect 27445 17153 27479 17187
rect 27629 17153 27663 17187
rect 27721 17153 27755 17187
rect 30665 17153 30699 17187
rect 31493 17153 31527 17187
rect 32321 17153 32355 17187
rect 33517 17153 33551 17187
rect 35449 17153 35483 17187
rect 36001 17153 36035 17187
rect 36277 17153 36311 17187
rect 36645 17153 36679 17187
rect 37473 17153 37507 17187
rect 38577 17153 38611 17187
rect 38761 17153 38795 17187
rect 39405 17153 39439 17187
rect 40141 17153 40175 17187
rect 41429 17153 41463 17187
rect 42901 17153 42935 17187
rect 42993 17153 43027 17187
rect 43085 17153 43119 17187
rect 43269 17153 43303 17187
rect 43821 17153 43855 17187
rect 44097 17153 44131 17187
rect 44741 17153 44775 17187
rect 46121 17153 46155 17187
rect 48789 17153 48823 17187
rect 48881 17153 48915 17187
rect 49157 17153 49191 17187
rect 51914 17153 51948 17187
rect 55965 17153 55999 17187
rect 56149 17153 56183 17187
rect 56333 17153 56367 17187
rect 57069 17153 57103 17187
rect 23949 17119 23983 17153
rect 1777 17085 1811 17119
rect 20085 17085 20119 17119
rect 25605 17085 25639 17119
rect 26525 17085 26559 17119
rect 28733 17085 28767 17119
rect 35909 17085 35943 17119
rect 45477 17085 45511 17119
rect 49249 17085 49283 17119
rect 52377 17085 52411 17119
rect 57345 17085 57379 17119
rect 24961 17017 24995 17051
rect 34897 17017 34931 17051
rect 40325 17017 40359 17051
rect 52285 17017 52319 17051
rect 17785 16949 17819 16983
rect 18521 16949 18555 16983
rect 23121 16949 23155 16983
rect 26157 16949 26191 16983
rect 27169 16949 27203 16983
rect 30113 16949 30147 16983
rect 30849 16949 30883 16983
rect 37657 16949 37691 16983
rect 38945 16949 38979 16983
rect 48237 16949 48271 16983
rect 56517 16949 56551 16983
rect 16681 16745 16715 16779
rect 36921 16745 36955 16779
rect 37473 16745 37507 16779
rect 39497 16745 39531 16779
rect 48513 16745 48547 16779
rect 51089 16745 51123 16779
rect 58265 16745 58299 16779
rect 26617 16677 26651 16711
rect 27629 16677 27663 16711
rect 36185 16677 36219 16711
rect 43545 16677 43579 16711
rect 53205 16677 53239 16711
rect 17233 16609 17267 16643
rect 20085 16609 20119 16643
rect 22201 16609 22235 16643
rect 25513 16609 25547 16643
rect 26488 16609 26522 16643
rect 26709 16609 26743 16643
rect 29745 16609 29779 16643
rect 38117 16609 38151 16643
rect 40693 16609 40727 16643
rect 45201 16609 45235 16643
rect 48789 16609 48823 16643
rect 56057 16609 56091 16643
rect 56425 16609 56459 16643
rect 56885 16609 56919 16643
rect 1593 16541 1627 16575
rect 16497 16541 16531 16575
rect 17509 16541 17543 16575
rect 20361 16541 20395 16575
rect 22468 16541 22502 16575
rect 25053 16541 25087 16575
rect 25329 16541 25363 16575
rect 25697 16541 25731 16575
rect 26341 16541 26375 16575
rect 27537 16541 27571 16575
rect 27813 16541 27847 16575
rect 28917 16541 28951 16575
rect 31861 16541 31895 16575
rect 33701 16541 33735 16575
rect 34897 16541 34931 16575
rect 35270 16541 35304 16575
rect 36001 16541 36035 16575
rect 36737 16541 36771 16575
rect 37473 16541 37507 16575
rect 37657 16541 37691 16575
rect 40417 16541 40451 16575
rect 44281 16541 44315 16575
rect 44373 16541 44407 16575
rect 44465 16541 44499 16575
rect 44649 16541 44683 16575
rect 48881 16541 48915 16575
rect 51825 16541 51859 16575
rect 52092 16541 52126 16575
rect 54677 16541 54711 16575
rect 54861 16541 54895 16575
rect 56241 16541 56275 16575
rect 57141 16541 57175 16575
rect 1869 16473 1903 16507
rect 21741 16473 21775 16507
rect 27077 16473 27111 16507
rect 30012 16473 30046 16507
rect 32128 16473 32162 16507
rect 35081 16473 35115 16507
rect 35173 16473 35207 16507
rect 38362 16473 38396 16507
rect 43177 16473 43211 16507
rect 43361 16473 43395 16507
rect 44005 16473 44039 16507
rect 45446 16473 45480 16507
rect 47133 16473 47167 16507
rect 47317 16473 47351 16507
rect 48421 16473 48455 16507
rect 50813 16473 50847 16507
rect 18797 16405 18831 16439
rect 23581 16405 23615 16439
rect 27997 16405 28031 16439
rect 29101 16405 29135 16439
rect 31125 16405 31159 16439
rect 33241 16405 33275 16439
rect 33885 16405 33919 16439
rect 35466 16405 35500 16439
rect 40049 16405 40083 16439
rect 40509 16405 40543 16439
rect 46581 16405 46615 16439
rect 47501 16405 47535 16439
rect 49065 16405 49099 16439
rect 54769 16405 54803 16439
rect 16221 16201 16255 16235
rect 23581 16201 23615 16235
rect 28095 16201 28129 16235
rect 31769 16201 31803 16235
rect 34621 16201 34655 16235
rect 37565 16201 37599 16235
rect 41613 16201 41647 16235
rect 43637 16201 43671 16235
rect 45477 16201 45511 16235
rect 49157 16201 49191 16235
rect 53665 16201 53699 16235
rect 55597 16201 55631 16235
rect 25973 16133 26007 16167
rect 29000 16133 29034 16167
rect 31401 16133 31435 16167
rect 31617 16133 31651 16167
rect 32934 16133 32968 16167
rect 38936 16133 38970 16167
rect 53481 16133 53515 16167
rect 54462 16133 54496 16167
rect 58173 16133 58207 16167
rect 1593 16065 1627 16099
rect 16037 16065 16071 16099
rect 19625 16065 19659 16099
rect 22477 16065 22511 16099
rect 22569 16065 22603 16099
rect 24041 16065 24075 16099
rect 24225 16065 24259 16099
rect 24593 16065 24627 16099
rect 27997 16065 28031 16099
rect 28181 16065 28215 16099
rect 28273 16065 28307 16099
rect 30573 16065 30607 16099
rect 30777 16055 30811 16089
rect 32689 16065 32723 16099
rect 34529 16065 34563 16099
rect 34713 16065 34747 16099
rect 35449 16065 35483 16099
rect 36737 16065 36771 16099
rect 36921 16065 36955 16099
rect 37841 16065 37875 16099
rect 37933 16065 37967 16099
rect 38025 16065 38059 16099
rect 38209 16065 38243 16099
rect 43453 16065 43487 16099
rect 44189 16065 44223 16099
rect 46765 16065 46799 16099
rect 47777 16065 47811 16099
rect 48044 16065 48078 16099
rect 50077 16065 50111 16099
rect 50344 16065 50378 16099
rect 53757 16065 53791 16099
rect 1777 15997 1811 16031
rect 17049 15997 17083 16031
rect 17325 15997 17359 16031
rect 19901 15997 19935 16031
rect 22293 15997 22327 16031
rect 22385 15997 22419 16031
rect 23121 15997 23155 16031
rect 25495 15997 25529 16031
rect 25973 15997 26007 16031
rect 26065 15997 26099 16031
rect 28733 15997 28767 16031
rect 38669 15997 38703 16031
rect 41705 15997 41739 16031
rect 41889 15997 41923 16031
rect 46857 15997 46891 16031
rect 46949 15997 46983 16031
rect 54217 15997 54251 16031
rect 23397 15929 23431 15963
rect 34069 15929 34103 15963
rect 36737 15929 36771 15963
rect 58357 15929 58391 15963
rect 18429 15861 18463 15895
rect 21189 15861 21223 15895
rect 22109 15861 22143 15895
rect 30113 15861 30147 15895
rect 30941 15861 30975 15895
rect 31585 15861 31619 15895
rect 35633 15861 35667 15895
rect 40049 15861 40083 15895
rect 41245 15861 41279 15895
rect 46397 15861 46431 15895
rect 51457 15861 51491 15895
rect 53481 15861 53515 15895
rect 14565 15657 14599 15691
rect 23673 15657 23707 15691
rect 25053 15657 25087 15691
rect 31125 15657 31159 15691
rect 32229 15657 32263 15691
rect 32965 15657 32999 15691
rect 51825 15657 51859 15691
rect 17785 15589 17819 15623
rect 20269 15589 20303 15623
rect 42073 15589 42107 15623
rect 46949 15589 46983 15623
rect 11437 15521 11471 15555
rect 11805 15521 11839 15555
rect 14841 15521 14875 15555
rect 14933 15521 14967 15555
rect 15853 15521 15887 15555
rect 15945 15521 15979 15555
rect 17509 15521 17543 15555
rect 21649 15521 21683 15555
rect 22293 15521 22327 15555
rect 30021 15521 30055 15555
rect 31677 15521 31711 15555
rect 38853 15521 38887 15555
rect 40693 15521 40727 15555
rect 42993 15521 43027 15555
rect 45569 15521 45603 15555
rect 1593 15453 1627 15487
rect 11345 15453 11379 15487
rect 11713 15453 11747 15487
rect 14749 15453 14783 15487
rect 15025 15453 15059 15487
rect 15761 15453 15795 15487
rect 16037 15453 16071 15487
rect 17417 15453 17451 15487
rect 21373 15453 21407 15487
rect 21465 15453 21499 15487
rect 21557 15453 21591 15487
rect 23489 15453 23523 15487
rect 28181 15453 28215 15487
rect 28917 15453 28951 15487
rect 29929 15453 29963 15487
rect 30757 15453 30791 15487
rect 30941 15453 30975 15487
rect 31953 15453 31987 15487
rect 32781 15453 32815 15487
rect 33609 15453 33643 15487
rect 33793 15453 33827 15487
rect 33977 15453 34011 15487
rect 40960 15453 40994 15487
rect 45836 15453 45870 15487
rect 47501 15453 47535 15487
rect 47685 15453 47719 15487
rect 47869 15453 47903 15487
rect 48145 15453 48179 15487
rect 50626 15453 50660 15487
rect 50997 15453 51031 15487
rect 51089 15453 51123 15487
rect 51733 15453 51767 15487
rect 57897 15453 57931 15487
rect 1869 15385 1903 15419
rect 10701 15385 10735 15419
rect 18245 15385 18279 15419
rect 18429 15385 18463 15419
rect 19993 15385 20027 15419
rect 22661 15385 22695 15419
rect 23029 15385 23063 15419
rect 25329 15385 25363 15419
rect 25513 15385 25547 15419
rect 25605 15385 25639 15419
rect 38577 15385 38611 15419
rect 43260 15385 43294 15419
rect 47777 15385 47811 15419
rect 47987 15385 48021 15419
rect 51549 15385 51583 15419
rect 58173 15385 58207 15419
rect 15577 15317 15611 15351
rect 18613 15317 18647 15351
rect 20453 15317 20487 15351
rect 21189 15317 21223 15351
rect 22477 15317 22511 15351
rect 22569 15317 22603 15351
rect 28365 15317 28399 15351
rect 29101 15317 29135 15351
rect 30297 15317 30331 15351
rect 31861 15317 31895 15351
rect 32045 15317 32079 15351
rect 38209 15317 38243 15351
rect 38669 15317 38703 15351
rect 44373 15317 44407 15351
rect 50445 15317 50479 15351
rect 50629 15317 50663 15351
rect 15117 15113 15151 15147
rect 20453 15113 20487 15147
rect 23397 15113 23431 15147
rect 28641 15113 28675 15147
rect 30113 15113 30147 15147
rect 32505 15113 32539 15147
rect 43545 15113 43579 15147
rect 43913 15113 43947 15147
rect 48145 15113 48179 15147
rect 50261 15113 50295 15147
rect 22293 15045 22327 15079
rect 22753 15045 22787 15079
rect 33885 15045 33919 15079
rect 33977 15045 34011 15079
rect 45201 15045 45235 15079
rect 51089 15045 51123 15079
rect 54953 15045 54987 15079
rect 1593 14977 1627 15011
rect 15301 14977 15335 15011
rect 17693 14977 17727 15011
rect 17785 14977 17819 15011
rect 18429 14977 18463 15011
rect 20269 14977 20303 15011
rect 21005 14977 21039 15011
rect 23213 14977 23247 15011
rect 24869 14977 24903 15011
rect 25881 14977 25915 15011
rect 26157 14977 26191 15011
rect 28457 14977 28491 15011
rect 29377 14977 29411 15011
rect 29929 14977 29963 15011
rect 31125 14977 31159 15011
rect 32321 14977 32355 15011
rect 33609 14977 33643 15011
rect 34437 14977 34471 15011
rect 37657 14977 37691 15011
rect 37924 14977 37958 15011
rect 39957 14977 39991 15011
rect 40224 14977 40258 15011
rect 44925 14977 44959 15011
rect 47961 14977 47995 15011
rect 50169 14977 50203 15011
rect 50353 14977 50387 15011
rect 50813 14977 50847 15011
rect 54493 14977 54527 15011
rect 54769 14977 54803 15011
rect 58081 14977 58115 15011
rect 1777 14909 1811 14943
rect 15393 14909 15427 14943
rect 15485 14909 15519 14943
rect 15577 14909 15611 14943
rect 22017 14909 22051 14943
rect 22385 14909 22419 14943
rect 22477 14909 22511 14943
rect 25237 14909 25271 14943
rect 25329 14909 25363 14943
rect 26525 14909 26559 14943
rect 33793 14909 33827 14943
rect 44005 14909 44039 14943
rect 44097 14909 44131 14943
rect 47777 14909 47811 14943
rect 18613 14841 18647 14875
rect 25973 14841 26007 14875
rect 31309 14841 31343 14875
rect 17969 14773 18003 14807
rect 21189 14773 21223 14807
rect 29377 14773 29411 14807
rect 34621 14773 34655 14807
rect 39037 14773 39071 14807
rect 41337 14773 41371 14807
rect 58265 14773 58299 14807
rect 16313 14569 16347 14603
rect 25237 14569 25271 14603
rect 29101 14569 29135 14603
rect 31125 14569 31159 14603
rect 31769 14569 31803 14603
rect 32321 14569 32355 14603
rect 33517 14569 33551 14603
rect 35725 14569 35759 14603
rect 40509 14569 40543 14603
rect 16129 14501 16163 14535
rect 17693 14501 17727 14535
rect 20085 14501 20119 14535
rect 21281 14501 21315 14535
rect 33057 14501 33091 14535
rect 34253 14501 34287 14535
rect 26893 14433 26927 14467
rect 40969 14433 41003 14467
rect 41153 14433 41187 14467
rect 1593 14365 1627 14399
rect 15025 14365 15059 14399
rect 17509 14365 17543 14399
rect 20269 14365 20303 14399
rect 21097 14365 21131 14399
rect 23673 14365 23707 14399
rect 25053 14365 25087 14399
rect 26709 14365 26743 14399
rect 28273 14365 28307 14399
rect 28457 14365 28491 14399
rect 28917 14365 28951 14399
rect 29745 14365 29779 14399
rect 31585 14365 31619 14399
rect 32321 14365 32355 14399
rect 32505 14365 32539 14399
rect 33241 14365 33275 14399
rect 33333 14365 33367 14399
rect 33609 14365 33643 14399
rect 34069 14365 34103 14399
rect 34897 14365 34931 14399
rect 35633 14365 35667 14399
rect 49617 14365 49651 14399
rect 49801 14365 49835 14399
rect 50353 14365 50387 14399
rect 57897 14365 57931 14399
rect 1869 14297 1903 14331
rect 14841 14297 14875 14331
rect 15853 14297 15887 14331
rect 20493 14297 20527 14331
rect 20637 14297 20671 14331
rect 28365 14297 28399 14331
rect 29990 14297 30024 14331
rect 40233 14297 40267 14331
rect 40877 14297 40911 14331
rect 49709 14297 49743 14331
rect 50598 14297 50632 14331
rect 58173 14297 58207 14331
rect 15117 14229 15151 14263
rect 20361 14229 20395 14263
rect 23857 14229 23891 14263
rect 26249 14229 26283 14263
rect 26617 14229 26651 14263
rect 35081 14229 35115 14263
rect 51733 14229 51767 14263
rect 15577 14025 15611 14059
rect 21373 14025 21407 14059
rect 26617 14025 26651 14059
rect 27721 14025 27755 14059
rect 29101 14025 29135 14059
rect 30665 14025 30699 14059
rect 31499 14025 31533 14059
rect 31585 14025 31619 14059
rect 32321 14025 32355 14059
rect 35357 14025 35391 14059
rect 37841 14025 37875 14059
rect 50445 14025 50479 14059
rect 15117 13957 15151 13991
rect 24326 13957 24360 13991
rect 49893 13957 49927 13991
rect 1593 13889 1627 13923
rect 21189 13889 21223 13923
rect 23949 13889 23983 13923
rect 24593 13889 24627 13923
rect 25237 13889 25271 13923
rect 25504 13889 25538 13923
rect 27537 13889 27571 13923
rect 29377 13889 29411 13923
rect 29469 13889 29503 13923
rect 29561 13889 29595 13923
rect 29745 13889 29779 13923
rect 30481 13889 30515 13923
rect 31401 13889 31435 13923
rect 31677 13889 31711 13923
rect 32505 13889 32539 13923
rect 32597 13889 32631 13923
rect 32873 13889 32907 13923
rect 33333 13889 33367 13923
rect 33517 13889 33551 13923
rect 33977 13889 34011 13923
rect 34233 13889 34267 13923
rect 42625 13889 42659 13923
rect 42892 13889 42926 13923
rect 50442 13889 50476 13923
rect 56425 13889 56459 13923
rect 57069 13889 57103 13923
rect 58081 13889 58115 13923
rect 1777 13821 1811 13855
rect 37933 13821 37967 13855
rect 38117 13821 38151 13855
rect 50905 13821 50939 13855
rect 56241 13821 56275 13855
rect 57345 13821 57379 13855
rect 15393 13753 15427 13787
rect 32781 13753 32815 13787
rect 50261 13753 50295 13787
rect 50813 13753 50847 13787
rect 58265 13753 58299 13787
rect 24317 13685 24351 13719
rect 33425 13685 33459 13719
rect 37473 13685 37507 13719
rect 44005 13685 44039 13719
rect 56609 13685 56643 13719
rect 16221 13481 16255 13515
rect 21281 13481 21315 13515
rect 30297 13481 30331 13515
rect 32873 13481 32907 13515
rect 33701 13481 33735 13515
rect 37565 13481 37599 13515
rect 55689 13481 55723 13515
rect 58173 13481 58207 13515
rect 16037 13413 16071 13447
rect 27077 13413 27111 13447
rect 50353 13413 50387 13447
rect 15761 13345 15795 13379
rect 25237 13345 25271 13379
rect 27629 13345 27663 13379
rect 56793 13345 56827 13379
rect 1593 13277 1627 13311
rect 21097 13277 21131 13311
rect 23673 13277 23707 13311
rect 27537 13277 27571 13311
rect 30113 13277 30147 13311
rect 30849 13277 30883 13311
rect 32689 13277 32723 13311
rect 33957 13277 33991 13311
rect 34069 13277 34103 13311
rect 34161 13277 34195 13311
rect 34345 13277 34379 13311
rect 36185 13277 36219 13311
rect 36452 13277 36486 13311
rect 41797 13277 41831 13311
rect 50537 13277 50571 13311
rect 50629 13277 50663 13311
rect 55873 13277 55907 13311
rect 56333 13277 56367 13311
rect 57049 13277 57083 13311
rect 1869 13209 1903 13243
rect 25504 13209 25538 13243
rect 27445 13209 27479 13243
rect 32505 13209 32539 13243
rect 46857 13209 46891 13243
rect 50905 13209 50939 13243
rect 50997 13209 51031 13243
rect 55965 13209 55999 13243
rect 56057 13209 56091 13243
rect 56175 13209 56209 13243
rect 23857 13141 23891 13175
rect 26617 13141 26651 13175
rect 31033 13141 31067 13175
rect 43085 13141 43119 13175
rect 48145 13141 48179 13175
rect 51273 13141 51307 13175
rect 23305 12937 23339 12971
rect 25513 12937 25547 12971
rect 26157 12937 26191 12971
rect 29837 12937 29871 12971
rect 58265 12937 58299 12971
rect 30573 12869 30607 12903
rect 30665 12869 30699 12903
rect 33793 12869 33827 12903
rect 49433 12869 49467 12903
rect 51181 12869 51215 12903
rect 55781 12869 55815 12903
rect 55873 12869 55907 12903
rect 57161 12869 57195 12903
rect 1593 12801 1627 12835
rect 24133 12801 24167 12835
rect 24389 12801 24423 12835
rect 25973 12801 26007 12835
rect 29653 12801 29687 12835
rect 30389 12801 30423 12835
rect 30809 12801 30843 12835
rect 37841 12801 37875 12835
rect 42993 12801 43027 12835
rect 51641 12801 51675 12835
rect 55597 12801 55631 12835
rect 55965 12801 55999 12835
rect 56701 12801 56735 12835
rect 58081 12801 58115 12835
rect 1777 12733 1811 12767
rect 23397 12733 23431 12767
rect 23489 12733 23523 12767
rect 35541 12733 35575 12767
rect 37933 12733 37967 12767
rect 38117 12733 38151 12767
rect 43085 12733 43119 12767
rect 43269 12733 43303 12767
rect 51917 12733 51951 12767
rect 22937 12665 22971 12699
rect 30941 12665 30975 12699
rect 37473 12597 37507 12631
rect 42625 12597 42659 12631
rect 56149 12597 56183 12631
rect 13185 12393 13219 12427
rect 22753 12393 22787 12427
rect 29101 12393 29135 12427
rect 58173 12393 58207 12427
rect 13553 12257 13587 12291
rect 23857 12257 23891 12291
rect 24593 12257 24627 12291
rect 30849 12257 30883 12291
rect 42165 12257 42199 12291
rect 43361 12257 43395 12291
rect 50353 12257 50387 12291
rect 56057 12257 56091 12291
rect 56793 12257 56827 12291
rect 1593 12189 1627 12223
rect 13369 12189 13403 12223
rect 13461 12189 13495 12223
rect 13645 12189 13679 12223
rect 22569 12189 22603 12223
rect 23673 12189 23707 12223
rect 28917 12189 28951 12223
rect 30665 12189 30699 12223
rect 30941 12189 30975 12223
rect 31217 12189 31251 12223
rect 31861 12189 31895 12223
rect 36369 12189 36403 12223
rect 41889 12189 41923 12223
rect 43085 12189 43119 12223
rect 49433 12189 49467 12223
rect 49617 12189 49651 12223
rect 55873 12189 55907 12223
rect 1869 12121 1903 12155
rect 24838 12121 24872 12155
rect 36636 12121 36670 12155
rect 49801 12121 49835 12155
rect 50598 12121 50632 12155
rect 57038 12121 57072 12155
rect 23305 12053 23339 12087
rect 23765 12053 23799 12087
rect 25973 12053 26007 12087
rect 37749 12053 37783 12087
rect 41521 12053 41555 12087
rect 41981 12053 42015 12087
rect 42717 12053 42751 12087
rect 43177 12053 43211 12087
rect 51733 12053 51767 12087
rect 13093 11849 13127 11883
rect 24041 11849 24075 11883
rect 25329 11849 25363 11883
rect 27353 11849 27387 11883
rect 30941 11849 30975 11883
rect 32413 11849 32447 11883
rect 37473 11849 37507 11883
rect 37841 11849 37875 11883
rect 42993 11849 43027 11883
rect 56701 11849 56735 11883
rect 23949 11781 23983 11815
rect 31401 11781 31435 11815
rect 37933 11781 37967 11815
rect 40868 11781 40902 11815
rect 46213 11781 46247 11815
rect 1593 11713 1627 11747
rect 17877 11713 17911 11747
rect 17969 11713 18003 11747
rect 25145 11713 25179 11747
rect 27169 11713 27203 11747
rect 29828 11713 29862 11747
rect 31585 11713 31619 11747
rect 32597 11713 32631 11747
rect 32781 11713 32815 11747
rect 34897 11713 34931 11747
rect 35541 11713 35575 11747
rect 35808 11713 35842 11747
rect 42809 11713 42843 11747
rect 44364 11713 44398 11747
rect 45937 11713 45971 11747
rect 49157 11713 49191 11747
rect 49525 11713 49559 11747
rect 56517 11713 56551 11747
rect 58081 11713 58115 11747
rect 1777 11645 1811 11679
rect 13277 11645 13311 11679
rect 13369 11645 13403 11679
rect 13461 11645 13495 11679
rect 13553 11645 13587 11679
rect 17693 11645 17727 11679
rect 18061 11645 18095 11679
rect 18153 11645 18187 11679
rect 29561 11645 29595 11679
rect 31769 11645 31803 11679
rect 34713 11645 34747 11679
rect 38025 11645 38059 11679
rect 40601 11645 40635 11679
rect 44097 11645 44131 11679
rect 49065 11645 49099 11679
rect 49617 11645 49651 11679
rect 56333 11645 56367 11679
rect 48605 11577 48639 11611
rect 35081 11509 35115 11543
rect 36921 11509 36955 11543
rect 41981 11509 42015 11543
rect 45477 11509 45511 11543
rect 58265 11509 58299 11543
rect 13553 11305 13587 11339
rect 15485 11305 15519 11339
rect 17233 11305 17267 11339
rect 19901 11305 19935 11339
rect 23305 11305 23339 11339
rect 29745 11305 29779 11339
rect 45201 11305 45235 11339
rect 48789 11305 48823 11339
rect 13369 11237 13403 11271
rect 17049 11237 17083 11271
rect 19717 11237 19751 11271
rect 24777 11237 24811 11271
rect 31401 11237 31435 11271
rect 36553 11237 36587 11271
rect 38117 11237 38151 11271
rect 43085 11237 43119 11271
rect 57253 11237 57287 11271
rect 14289 11169 14323 11203
rect 14473 11169 14507 11203
rect 14565 11169 14599 11203
rect 14657 11169 14691 11203
rect 23857 11169 23891 11203
rect 32137 11169 32171 11203
rect 37473 11169 37507 11203
rect 41705 11169 41739 11203
rect 45845 11169 45879 11203
rect 46765 11169 46799 11203
rect 58173 11169 58207 11203
rect 1593 11101 1627 11135
rect 13093 11101 13127 11135
rect 14749 11101 14783 11135
rect 15393 11101 15427 11135
rect 23673 11101 23707 11135
rect 23765 11101 23799 11135
rect 24593 11101 24627 11135
rect 28825 11101 28859 11135
rect 30021 11101 30055 11135
rect 30113 11101 30147 11135
rect 30205 11098 30239 11132
rect 30389 11101 30423 11135
rect 31309 11101 31343 11135
rect 31953 11101 31987 11135
rect 32413 11101 32447 11135
rect 32781 11101 32815 11135
rect 33701 11101 33735 11135
rect 33793 11101 33827 11135
rect 33885 11101 33919 11135
rect 34069 11101 34103 11135
rect 35173 11101 35207 11135
rect 35440 11101 35474 11135
rect 37381 11101 37415 11135
rect 38301 11101 38335 11135
rect 38393 11101 38427 11135
rect 38577 11101 38611 11135
rect 38669 11101 38703 11135
rect 39129 11101 39163 11135
rect 39313 11101 39347 11135
rect 41972 11101 42006 11135
rect 45661 11101 45695 11135
rect 46489 11101 46523 11135
rect 48237 11101 48271 11135
rect 48605 11101 48639 11135
rect 57897 11101 57931 11135
rect 1869 11033 1903 11067
rect 16773 11033 16807 11067
rect 19441 11033 19475 11067
rect 29009 11033 29043 11067
rect 45569 11033 45603 11067
rect 48421 11033 48455 11067
rect 48513 11033 48547 11067
rect 57069 11033 57103 11067
rect 29193 10965 29227 10999
rect 33425 10965 33459 10999
rect 39497 10965 39531 10999
rect 12909 10761 12943 10795
rect 13829 10761 13863 10795
rect 23489 10761 23523 10795
rect 25697 10761 25731 10795
rect 30389 10761 30423 10795
rect 35449 10761 35483 10795
rect 35817 10761 35851 10795
rect 46397 10761 46431 10795
rect 46765 10761 46799 10795
rect 32956 10693 32990 10727
rect 38476 10693 38510 10727
rect 44824 10693 44858 10727
rect 1593 10625 1627 10659
rect 12449 10625 12483 10659
rect 13369 10625 13403 10659
rect 23213 10625 23247 10659
rect 23857 10625 23891 10659
rect 28181 10625 28215 10659
rect 28273 10625 28307 10659
rect 28365 10625 28399 10659
rect 28549 10625 28583 10659
rect 29265 10625 29299 10659
rect 35081 10625 35115 10659
rect 35909 10625 35943 10659
rect 38209 10625 38243 10659
rect 40141 10625 40175 10659
rect 56333 10625 56367 10659
rect 56517 10625 56551 10659
rect 56609 10625 56643 10659
rect 57069 10625 57103 10659
rect 58081 10635 58115 10669
rect 58265 10625 58299 10659
rect 1777 10557 1811 10591
rect 23949 10557 23983 10591
rect 24041 10557 24075 10591
rect 25789 10557 25823 10591
rect 25973 10557 26007 10591
rect 29009 10557 29043 10591
rect 32689 10557 32723 10591
rect 36093 10557 36127 10591
rect 44557 10557 44591 10591
rect 46857 10557 46891 10591
rect 46949 10557 46983 10591
rect 57345 10557 57379 10591
rect 12817 10489 12851 10523
rect 13645 10489 13679 10523
rect 27905 10489 27939 10523
rect 58173 10489 58207 10523
rect 25329 10421 25363 10455
rect 34069 10421 34103 10455
rect 39589 10421 39623 10455
rect 40233 10421 40267 10455
rect 45937 10421 45971 10455
rect 56333 10421 56367 10455
rect 12357 10217 12391 10251
rect 32689 10217 32723 10251
rect 38577 10217 38611 10251
rect 46581 10217 46615 10251
rect 58173 10217 58207 10251
rect 23581 10149 23615 10183
rect 27261 10149 27295 10183
rect 28273 10149 28307 10183
rect 56057 10149 56091 10183
rect 12541 10081 12575 10115
rect 12633 10081 12667 10115
rect 35633 10081 35667 10115
rect 39037 10081 39071 10115
rect 39129 10081 39163 10115
rect 56793 10081 56827 10115
rect 1593 10013 1627 10047
rect 12725 10013 12759 10047
rect 12817 10013 12851 10047
rect 24593 10013 24627 10047
rect 24860 10013 24894 10047
rect 27077 10013 27111 10047
rect 28089 10013 28123 10047
rect 36369 10013 36403 10047
rect 38945 10013 38979 10047
rect 45201 10013 45235 10047
rect 56333 10013 56367 10047
rect 57049 10013 57083 10047
rect 1869 9945 1903 9979
rect 23397 9945 23431 9979
rect 31217 9945 31251 9979
rect 34897 9945 34931 9979
rect 36737 9945 36771 9979
rect 45468 9945 45502 9979
rect 56057 9945 56091 9979
rect 25973 9877 26007 9911
rect 56241 9877 56275 9911
rect 25329 9673 25363 9707
rect 30481 9673 30515 9707
rect 45385 9673 45419 9707
rect 56517 9673 56551 9707
rect 23121 9605 23155 9639
rect 32597 9605 32631 9639
rect 32781 9605 32815 9639
rect 36277 9605 36311 9639
rect 45753 9605 45787 9639
rect 1593 9537 1627 9571
rect 12541 9537 12575 9571
rect 12633 9537 12667 9571
rect 23949 9537 23983 9571
rect 24205 9537 24239 9571
rect 26341 9537 26375 9571
rect 27169 9537 27203 9571
rect 27436 9537 27470 9571
rect 30297 9537 30331 9571
rect 30481 9537 30515 9571
rect 31037 9537 31071 9571
rect 31217 9537 31251 9571
rect 31309 9537 31343 9571
rect 31585 9537 31619 9571
rect 32413 9537 32447 9571
rect 33241 9537 33275 9571
rect 33425 9537 33459 9571
rect 34069 9537 34103 9571
rect 34336 9537 34370 9571
rect 36369 9537 36403 9571
rect 39037 9537 39071 9571
rect 39129 9537 39163 9571
rect 39313 9537 39347 9571
rect 39405 9537 39439 9571
rect 44189 9537 44223 9571
rect 56425 9537 56459 9571
rect 56609 9537 56643 9571
rect 57069 9537 57103 9571
rect 1777 9469 1811 9503
rect 12357 9469 12391 9503
rect 12725 9469 12759 9503
rect 12817 9469 12851 9503
rect 13369 9469 13403 9503
rect 13829 9469 13863 9503
rect 23213 9469 23247 9503
rect 23305 9469 23339 9503
rect 31401 9469 31435 9503
rect 31769 9469 31803 9503
rect 36461 9469 36495 9503
rect 44465 9469 44499 9503
rect 45845 9469 45879 9503
rect 46029 9469 46063 9503
rect 57345 9469 57379 9503
rect 13645 9401 13679 9435
rect 22753 9401 22787 9435
rect 26525 9401 26559 9435
rect 28549 9401 28583 9435
rect 33609 9401 33643 9435
rect 35909 9401 35943 9435
rect 35449 9333 35483 9367
rect 38853 9333 38887 9367
rect 12265 9129 12299 9163
rect 26617 9129 26651 9163
rect 31033 9129 31067 9163
rect 44097 9129 44131 9163
rect 58173 9129 58207 9163
rect 12541 8993 12575 9027
rect 25697 8993 25731 9027
rect 27169 8993 27203 9027
rect 36737 8993 36771 9027
rect 41245 8993 41279 9027
rect 56793 8993 56827 9027
rect 1593 8925 1627 8959
rect 12449 8925 12483 8959
rect 12633 8925 12667 8959
rect 12725 8925 12759 8959
rect 22937 8925 22971 8959
rect 23029 8925 23063 8959
rect 23213 8925 23247 8959
rect 25421 8925 25455 8959
rect 26433 8925 26467 8959
rect 29009 8925 29043 8959
rect 29193 8925 29227 8959
rect 30021 8925 30055 8959
rect 30113 8925 30147 8959
rect 30205 8925 30239 8959
rect 30389 8925 30423 8959
rect 30849 8925 30883 8959
rect 31585 8925 31619 8959
rect 31677 8925 31711 8959
rect 35541 8925 35575 8959
rect 35817 8925 35851 8959
rect 35909 8925 35943 8959
rect 41061 8925 41095 8959
rect 44005 8925 44039 8959
rect 57049 8925 57083 8959
rect 1869 8857 1903 8891
rect 27436 8857 27470 8891
rect 36277 8857 36311 8891
rect 25053 8789 25087 8823
rect 25513 8789 25547 8823
rect 28549 8789 28583 8823
rect 29101 8789 29135 8823
rect 29745 8789 29779 8823
rect 40693 8789 40727 8823
rect 41153 8789 41187 8823
rect 12173 8585 12207 8619
rect 27905 8585 27939 8619
rect 28273 8585 28307 8619
rect 29469 8585 29503 8619
rect 31585 8585 31619 8619
rect 41429 8585 41463 8619
rect 58265 8585 58299 8619
rect 13645 8517 13679 8551
rect 33609 8517 33643 8551
rect 33701 8517 33735 8551
rect 35909 8517 35943 8551
rect 36277 8517 36311 8551
rect 47961 8517 47995 8551
rect 48053 8517 48087 8551
rect 1593 8449 1627 8483
rect 10793 8449 10827 8483
rect 10885 8449 10919 8483
rect 12357 8449 12391 8483
rect 12449 8449 12483 8483
rect 13277 8449 13311 8483
rect 24225 8449 24259 8483
rect 24492 8449 24526 8483
rect 29285 8449 29319 8483
rect 30297 8449 30331 8483
rect 33333 8449 33367 8483
rect 33426 8449 33460 8483
rect 33839 8449 33873 8483
rect 34713 8449 34747 8483
rect 34805 8449 34839 8483
rect 34989 8449 35023 8483
rect 35081 8449 35115 8483
rect 35817 8449 35851 8483
rect 37473 8449 37507 8483
rect 40049 8449 40083 8483
rect 40316 8449 40350 8483
rect 42625 8449 42659 8483
rect 42892 8449 42926 8483
rect 47777 8449 47811 8483
rect 48145 8449 48179 8483
rect 48973 8449 49007 8483
rect 58081 8449 58115 8483
rect 1777 8381 1811 8415
rect 10609 8381 10643 8415
rect 10977 8381 11011 8415
rect 11069 8381 11103 8415
rect 12541 8381 12575 8415
rect 12633 8381 12667 8415
rect 28365 8381 28399 8415
rect 28549 8381 28583 8415
rect 30021 8381 30055 8415
rect 35541 8381 35575 8415
rect 37657 8381 37691 8415
rect 25605 8313 25639 8347
rect 34529 8313 34563 8347
rect 36461 8313 36495 8347
rect 48329 8313 48363 8347
rect 48789 8313 48823 8347
rect 33977 8245 34011 8279
rect 44005 8245 44039 8279
rect 10517 8041 10551 8075
rect 13461 8041 13495 8075
rect 22845 8041 22879 8075
rect 27905 8041 27939 8075
rect 31493 8041 31527 8075
rect 42993 8041 43027 8075
rect 48881 8041 48915 8075
rect 10333 7973 10367 8007
rect 12357 7973 12391 8007
rect 12541 7973 12575 8007
rect 13277 7973 13311 8007
rect 36737 7973 36771 8007
rect 38117 7973 38151 8007
rect 10977 7905 11011 7939
rect 11161 7905 11195 7939
rect 11253 7905 11287 7939
rect 12081 7905 12115 7939
rect 13001 7905 13035 7939
rect 23397 7905 23431 7939
rect 28549 7905 28583 7939
rect 43545 7905 43579 7939
rect 47501 7905 47535 7939
rect 58173 7905 58207 7939
rect 1593 7837 1627 7871
rect 11345 7837 11379 7871
rect 11437 7837 11471 7871
rect 27445 7837 27479 7871
rect 30205 7837 30239 7871
rect 30298 7837 30332 7871
rect 30670 7837 30704 7871
rect 31677 7837 31711 7871
rect 31769 7837 31803 7871
rect 31953 7837 31987 7871
rect 32045 7837 32079 7871
rect 33885 7837 33919 7871
rect 35541 7837 35575 7871
rect 35817 7837 35851 7871
rect 37197 7837 37231 7871
rect 37473 7837 37507 7871
rect 37565 7837 37599 7871
rect 43361 7837 43395 7871
rect 46029 7837 46063 7871
rect 46305 7837 46339 7871
rect 46397 7837 46431 7871
rect 56977 7837 57011 7871
rect 57161 7837 57195 7871
rect 57897 7837 57931 7871
rect 1869 7769 1903 7803
rect 10057 7769 10091 7803
rect 27077 7769 27111 7803
rect 27261 7769 27295 7803
rect 28273 7769 28307 7803
rect 30481 7769 30515 7803
rect 30573 7769 30607 7803
rect 34161 7769 34195 7803
rect 35909 7769 35943 7803
rect 36277 7769 36311 7803
rect 37933 7769 37967 7803
rect 46213 7769 46247 7803
rect 47768 7769 47802 7803
rect 23213 7701 23247 7735
rect 23305 7701 23339 7735
rect 28365 7701 28399 7735
rect 30849 7701 30883 7735
rect 43453 7701 43487 7735
rect 46581 7701 46615 7735
rect 57069 7701 57103 7735
rect 11161 7497 11195 7531
rect 12265 7497 12299 7531
rect 20545 7497 20579 7531
rect 29929 7497 29963 7531
rect 39313 7497 39347 7531
rect 44833 7497 44867 7531
rect 46857 7497 46891 7531
rect 48145 7497 48179 7531
rect 56517 7497 56551 7531
rect 10701 7429 10735 7463
rect 11805 7429 11839 7463
rect 28641 7429 28675 7463
rect 33793 7429 33827 7463
rect 37841 7429 37875 7463
rect 56333 7429 56367 7463
rect 1593 7361 1627 7395
rect 24133 7361 24167 7395
rect 24400 7361 24434 7395
rect 31217 7361 31251 7395
rect 31401 7361 31435 7395
rect 32413 7361 32447 7395
rect 32781 7361 32815 7395
rect 37473 7361 37507 7395
rect 37749 7361 37783 7395
rect 38209 7361 38243 7395
rect 45109 7361 45143 7395
rect 45201 7361 45235 7395
rect 45293 7361 45327 7395
rect 45477 7361 45511 7395
rect 46581 7361 46615 7395
rect 47961 7361 47995 7395
rect 55597 7361 55631 7395
rect 55781 7361 55815 7395
rect 55873 7361 55907 7395
rect 56609 7361 56643 7395
rect 57069 7361 57103 7395
rect 58081 7361 58115 7395
rect 1777 7293 1811 7327
rect 20085 7293 20119 7327
rect 31125 7293 31159 7327
rect 31309 7293 31343 7327
rect 35541 7293 35575 7327
rect 39129 7293 39163 7327
rect 39497 7293 39531 7327
rect 47777 7293 47811 7327
rect 57345 7293 57379 7327
rect 10977 7225 11011 7259
rect 12081 7225 12115 7259
rect 20361 7225 20395 7259
rect 30941 7225 30975 7259
rect 38393 7225 38427 7259
rect 58265 7225 58299 7259
rect 25513 7157 25547 7191
rect 39681 7157 39715 7191
rect 55597 7157 55631 7191
rect 56333 7157 56367 7191
rect 20913 6953 20947 6987
rect 24961 6953 24995 6987
rect 31401 6953 31435 6987
rect 39221 6953 39255 6987
rect 40969 6953 41003 6987
rect 47685 6953 47719 6987
rect 58081 6953 58115 6987
rect 19809 6885 19843 6919
rect 20729 6885 20763 6919
rect 45201 6885 45235 6919
rect 25605 6817 25639 6851
rect 27537 6817 27571 6851
rect 29009 6817 29043 6851
rect 30665 6817 30699 6851
rect 30849 6817 30883 6851
rect 32321 6817 32355 6851
rect 37933 6817 37967 6851
rect 38025 6817 38059 6851
rect 43821 6817 43855 6851
rect 1593 6749 1627 6783
rect 27813 6749 27847 6783
rect 30573 6749 30607 6783
rect 30757 6749 30791 6783
rect 31401 6749 31435 6783
rect 31585 6749 31619 6783
rect 32505 6749 32539 6783
rect 32781 6749 32815 6783
rect 33977 6749 34011 6783
rect 35633 6749 35667 6783
rect 38669 6749 38703 6783
rect 39037 6749 39071 6783
rect 40417 6749 40451 6783
rect 40785 6749 40819 6783
rect 43637 6749 43671 6783
rect 44465 6749 44499 6783
rect 44649 6749 44683 6783
rect 45377 6727 45411 6761
rect 45469 6749 45503 6783
rect 45646 6749 45680 6783
rect 45753 6749 45787 6783
rect 46121 6749 46155 6783
rect 47869 6749 47903 6783
rect 47961 6749 47995 6783
rect 56701 6749 56735 6783
rect 56968 6749 57002 6783
rect 1869 6681 1903 6715
rect 19533 6681 19567 6715
rect 20453 6681 20487 6715
rect 25421 6681 25455 6715
rect 33793 6681 33827 6715
rect 35878 6681 35912 6715
rect 37841 6681 37875 6715
rect 43729 6681 43763 6715
rect 46857 6681 46891 6715
rect 47685 6681 47719 6715
rect 55873 6681 55907 6715
rect 19993 6613 20027 6647
rect 25329 6613 25363 6647
rect 30389 6613 30423 6647
rect 31769 6613 31803 6647
rect 32689 6613 32723 6647
rect 34069 6613 34103 6647
rect 37013 6613 37047 6647
rect 37473 6613 37507 6647
rect 38853 6613 38887 6647
rect 40601 6613 40635 6647
rect 43269 6613 43303 6647
rect 44557 6613 44591 6647
rect 47317 6613 47351 6647
rect 48145 6613 48179 6647
rect 55965 6613 55999 6647
rect 10425 6409 10459 6443
rect 28365 6409 28399 6443
rect 34713 6409 34747 6443
rect 39221 6409 39255 6443
rect 39865 6409 39899 6443
rect 40509 6409 40543 6443
rect 44281 6409 44315 6443
rect 46213 6409 46247 6443
rect 55321 6409 55355 6443
rect 58265 6409 58299 6443
rect 25237 6341 25271 6375
rect 27537 6341 27571 6375
rect 29929 6341 29963 6375
rect 1593 6273 1627 6307
rect 27629 6273 27663 6307
rect 28641 6273 28675 6307
rect 28733 6273 28767 6307
rect 28825 6273 28859 6307
rect 29009 6273 29043 6307
rect 29653 6273 29687 6307
rect 29837 6273 29871 6307
rect 30665 6273 30699 6307
rect 30757 6273 30791 6307
rect 32597 6273 32631 6307
rect 32781 6273 32815 6307
rect 34529 6273 34563 6307
rect 35449 6273 35483 6307
rect 35541 6273 35575 6307
rect 35909 6273 35943 6307
rect 37473 6273 37507 6307
rect 38485 6273 38519 6307
rect 39129 6273 39163 6307
rect 39313 6273 39347 6307
rect 39773 6273 39807 6307
rect 39957 6273 39991 6307
rect 40417 6273 40451 6307
rect 40601 6273 40635 6307
rect 42901 6273 42935 6307
rect 43168 6273 43202 6307
rect 44833 6273 44867 6307
rect 45017 6273 45051 6307
rect 45109 6273 45143 6307
rect 46029 6273 46063 6307
rect 46397 6273 46431 6307
rect 46673 6273 46707 6307
rect 55137 6273 55171 6307
rect 55321 6273 55355 6307
rect 55781 6273 55815 6307
rect 56048 6273 56082 6307
rect 58081 6273 58115 6307
rect 58357 6273 58391 6307
rect 1777 6205 1811 6239
rect 10609 6205 10643 6239
rect 10701 6205 10735 6239
rect 10793 6205 10827 6239
rect 10885 6205 10919 6239
rect 20729 6205 20763 6239
rect 25329 6205 25363 6239
rect 25513 6205 25547 6239
rect 27813 6205 27847 6239
rect 30573 6205 30607 6239
rect 30849 6205 30883 6239
rect 34345 6205 34379 6239
rect 35173 6205 35207 6239
rect 37657 6205 37691 6239
rect 45569 6205 45603 6239
rect 21005 6137 21039 6171
rect 21189 6137 21223 6171
rect 30389 6137 30423 6171
rect 36277 6137 36311 6171
rect 38669 6137 38703 6171
rect 24869 6069 24903 6103
rect 27169 6069 27203 6103
rect 32965 6069 32999 6103
rect 46489 6069 46523 6103
rect 57161 6069 57195 6103
rect 58081 6069 58115 6103
rect 11069 5865 11103 5899
rect 17785 5865 17819 5899
rect 23121 5865 23155 5899
rect 26801 5865 26835 5899
rect 30941 5865 30975 5899
rect 40233 5865 40267 5899
rect 45385 5865 45419 5899
rect 45569 5865 45603 5899
rect 46121 5865 46155 5899
rect 46765 5865 46799 5899
rect 56241 5865 56275 5899
rect 10885 5797 10919 5831
rect 20269 5797 20303 5831
rect 20453 5797 20487 5831
rect 10149 5729 10183 5763
rect 10609 5729 10643 5763
rect 18061 5729 18095 5763
rect 30021 5729 30055 5763
rect 36737 5729 36771 5763
rect 56793 5729 56827 5763
rect 1593 5661 1627 5695
rect 9413 5661 9447 5695
rect 9505 5661 9539 5695
rect 9689 5661 9723 5695
rect 17969 5661 18003 5695
rect 18153 5661 18187 5695
rect 18245 5661 18279 5695
rect 19993 5661 20027 5695
rect 25421 5661 25455 5695
rect 27721 5661 27755 5695
rect 30205 5661 30239 5695
rect 30481 5661 30515 5695
rect 31125 5661 31159 5695
rect 31401 5661 31435 5695
rect 32781 5661 32815 5695
rect 32873 5661 32907 5695
rect 32965 5661 32999 5695
rect 33149 5661 33183 5695
rect 34161 5661 34195 5695
rect 35541 5661 35575 5695
rect 35817 5661 35851 5695
rect 35909 5661 35943 5695
rect 37197 5661 37231 5695
rect 39129 5661 39163 5695
rect 40049 5661 40083 5695
rect 43085 5661 43119 5695
rect 46029 5661 46063 5695
rect 46213 5661 46247 5695
rect 46673 5661 46707 5695
rect 56149 5661 56183 5695
rect 56333 5661 56367 5695
rect 57060 5661 57094 5695
rect 1869 5593 1903 5627
rect 22845 5593 22879 5627
rect 25688 5593 25722 5627
rect 27905 5593 27939 5627
rect 34345 5593 34379 5627
rect 36277 5593 36311 5627
rect 37473 5593 37507 5627
rect 38209 5593 38243 5627
rect 38393 5593 38427 5627
rect 38945 5593 38979 5627
rect 43821 5593 43855 5627
rect 45201 5593 45235 5627
rect 45401 5593 45435 5627
rect 28089 5525 28123 5559
rect 30389 5525 30423 5559
rect 31309 5525 31343 5559
rect 32505 5525 32539 5559
rect 58173 5525 58207 5559
rect 22661 5321 22695 5355
rect 25513 5321 25547 5355
rect 26341 5321 26375 5355
rect 26433 5321 26467 5355
rect 29193 5321 29227 5355
rect 40509 5321 40543 5355
rect 41245 5321 41279 5355
rect 58265 5321 58299 5355
rect 24400 5253 24434 5287
rect 26065 5253 26099 5287
rect 26249 5253 26283 5287
rect 31125 5253 31159 5287
rect 34621 5253 34655 5287
rect 43453 5253 43487 5287
rect 45201 5253 45235 5287
rect 57345 5253 57379 5287
rect 1593 5185 1627 5219
rect 19809 5185 19843 5219
rect 21005 5185 21039 5219
rect 24133 5185 24167 5219
rect 26617 5185 26651 5219
rect 27813 5185 27847 5219
rect 30297 5185 30331 5219
rect 31309 5185 31343 5219
rect 32597 5185 32631 5219
rect 35541 5185 35575 5219
rect 35817 5185 35851 5219
rect 35909 5185 35943 5219
rect 36277 5185 36311 5219
rect 36737 5185 36771 5219
rect 37565 5185 37599 5219
rect 39129 5185 39163 5219
rect 39396 5185 39430 5219
rect 41061 5185 41095 5219
rect 41797 5185 41831 5219
rect 43269 5185 43303 5219
rect 45109 5185 45143 5219
rect 45293 5185 45327 5219
rect 46305 5185 46339 5219
rect 55505 5185 55539 5219
rect 56149 5185 56183 5219
rect 57069 5185 57103 5219
rect 58081 5185 58115 5219
rect 1777 5117 1811 5151
rect 19993 5117 20027 5151
rect 21281 5117 21315 5151
rect 22753 5117 22787 5151
rect 22845 5117 22879 5151
rect 28089 5117 28123 5151
rect 31493 5117 31527 5151
rect 32321 5117 32355 5151
rect 37841 5117 37875 5151
rect 43085 5117 43119 5151
rect 56425 5117 56459 5151
rect 33701 5049 33735 5083
rect 41981 5049 42015 5083
rect 46489 5049 46523 5083
rect 55689 5049 55723 5083
rect 22293 4981 22327 5015
rect 30389 4981 30423 5015
rect 34713 4981 34747 5015
rect 17877 4777 17911 4811
rect 22201 4777 22235 4811
rect 27721 4777 27755 4811
rect 39497 4777 39531 4811
rect 42165 4777 42199 4811
rect 43545 4777 43579 4811
rect 45937 4777 45971 4811
rect 48697 4777 48731 4811
rect 11805 4709 11839 4743
rect 17693 4709 17727 4743
rect 40049 4709 40083 4743
rect 46765 4709 46799 4743
rect 10701 4641 10735 4675
rect 17417 4641 17451 4675
rect 22845 4641 22879 4675
rect 37197 4641 37231 4675
rect 38025 4641 38059 4675
rect 39129 4641 39163 4675
rect 40509 4641 40543 4675
rect 40693 4641 40727 4675
rect 56885 4641 56919 4675
rect 1593 4573 1627 4607
rect 18521 4573 18555 4607
rect 19441 4573 19475 4607
rect 20361 4573 20395 4607
rect 21097 4573 21131 4607
rect 22661 4573 22695 4607
rect 24593 4573 24627 4607
rect 24860 4573 24894 4607
rect 26617 4573 26651 4607
rect 27261 4573 27295 4607
rect 27997 4573 28031 4607
rect 28089 4573 28123 4607
rect 28181 4573 28215 4607
rect 28365 4573 28399 4607
rect 31033 4573 31067 4607
rect 31953 4573 31987 4607
rect 32045 4573 32079 4607
rect 32137 4573 32171 4607
rect 32321 4573 32355 4607
rect 32873 4573 32907 4607
rect 33609 4573 33643 4607
rect 35173 4573 35207 4607
rect 35909 4573 35943 4607
rect 36001 4573 36035 4607
rect 37013 4573 37047 4607
rect 37841 4573 37875 4607
rect 39313 4573 39347 4607
rect 41981 4573 42015 4607
rect 43453 4573 43487 4607
rect 47225 4573 47259 4607
rect 48053 4573 48087 4607
rect 48201 4573 48235 4607
rect 48329 4573 48363 4607
rect 48421 4573 48455 4607
rect 48557 4573 48591 4607
rect 55965 4573 55999 4607
rect 1869 4505 1903 4539
rect 10517 4505 10551 4539
rect 11621 4505 11655 4539
rect 19717 4505 19751 4539
rect 20637 4505 20671 4539
rect 21373 4505 21407 4539
rect 21925 4505 21959 4539
rect 23489 4505 23523 4539
rect 31217 4505 31251 4539
rect 33057 4505 33091 4539
rect 33793 4505 33827 4539
rect 35357 4505 35391 4539
rect 41337 4505 41371 4539
rect 42809 4505 42843 4539
rect 45845 4505 45879 4539
rect 46581 4505 46615 4539
rect 56241 4505 56275 4539
rect 57130 4505 57164 4539
rect 22569 4437 22603 4471
rect 23765 4437 23799 4471
rect 25973 4437 26007 4471
rect 28825 4437 28859 4471
rect 31677 4437 31711 4471
rect 36185 4437 36219 4471
rect 36645 4437 36679 4471
rect 37105 4437 37139 4471
rect 40417 4437 40451 4471
rect 41429 4437 41463 4471
rect 42901 4437 42935 4471
rect 47409 4437 47443 4471
rect 58265 4437 58299 4471
rect 12173 4233 12207 4267
rect 25237 4233 25271 4267
rect 25605 4233 25639 4267
rect 31769 4233 31803 4267
rect 45017 4233 45051 4267
rect 9137 4165 9171 4199
rect 10977 4165 11011 4199
rect 15761 4165 15795 4199
rect 27537 4165 27571 4199
rect 28549 4165 28583 4199
rect 36645 4165 36679 4199
rect 45661 4165 45695 4199
rect 46397 4165 46431 4199
rect 50537 4165 50571 4199
rect 51273 4165 51307 4199
rect 52009 4165 52043 4199
rect 54585 4165 54619 4199
rect 55321 4165 55355 4199
rect 8309 4097 8343 4131
rect 8493 4097 8527 4131
rect 10149 4097 10183 4131
rect 11161 4097 11195 4131
rect 12633 4097 12667 4131
rect 17325 4097 17359 4131
rect 19165 4097 19199 4131
rect 19441 4097 19475 4131
rect 20085 4097 20119 4131
rect 22477 4097 22511 4131
rect 23397 4097 23431 4131
rect 24317 4097 24351 4131
rect 24593 4097 24627 4131
rect 29193 4097 29227 4131
rect 29460 4097 29494 4131
rect 31401 4097 31435 4131
rect 31585 4097 31619 4131
rect 32321 4097 32355 4131
rect 34713 4097 34747 4131
rect 35633 4097 35667 4131
rect 37473 4097 37507 4131
rect 37749 4097 37783 4131
rect 38393 4097 38427 4131
rect 39313 4097 39347 4131
rect 40233 4097 40267 4131
rect 41061 4097 41095 4131
rect 41797 4097 41831 4131
rect 42717 4097 42751 4131
rect 42901 4097 42935 4131
rect 43361 4097 43395 4131
rect 44097 4097 44131 4131
rect 44925 4097 44959 4131
rect 45845 4097 45879 4131
rect 47777 4097 47811 4131
rect 48237 4095 48271 4129
rect 48513 4097 48547 4131
rect 48605 4097 48639 4131
rect 48881 4097 48915 4131
rect 49157 4097 49191 4131
rect 49801 4097 49835 4131
rect 51457 4097 51491 4131
rect 53021 4097 53055 4131
rect 55505 4097 55539 4131
rect 56057 4097 56091 4131
rect 57161 4097 57195 4131
rect 57345 4097 57379 4131
rect 58081 4097 58115 4131
rect 9965 4029 9999 4063
rect 10057 4029 10091 4063
rect 10241 4029 10275 4063
rect 11713 4029 11747 4063
rect 17509 4029 17543 4063
rect 22753 4029 22787 4063
rect 23581 4029 23615 4063
rect 25697 4029 25731 4063
rect 25789 4029 25823 4063
rect 27629 4029 27663 4063
rect 27721 4029 27755 4063
rect 32597 4029 32631 4063
rect 34897 4029 34931 4063
rect 35817 4029 35851 4063
rect 38669 4029 38703 4063
rect 39497 4029 39531 4063
rect 41981 4029 42015 4063
rect 49985 4029 50019 4063
rect 53205 4029 53239 4063
rect 56333 4029 56367 4063
rect 9781 3961 9815 3995
rect 11989 3961 12023 3995
rect 20361 3961 20395 3995
rect 26617 3961 26651 3995
rect 41245 3961 41279 3995
rect 43545 3961 43579 3995
rect 44281 3961 44315 3995
rect 46581 3961 46615 3995
rect 54769 3961 54803 3995
rect 58265 3961 58299 3995
rect 9229 3893 9263 3927
rect 12817 3893 12851 3927
rect 15853 3893 15887 3927
rect 18613 3893 18647 3927
rect 20545 3893 20579 3927
rect 27169 3893 27203 3927
rect 30573 3893 30607 3927
rect 33701 3893 33735 3927
rect 36737 3893 36771 3927
rect 40417 3893 40451 3927
rect 50629 3893 50663 3927
rect 52101 3893 52135 3927
rect 57253 3893 57287 3927
rect 8493 3689 8527 3723
rect 9689 3689 9723 3723
rect 12909 3689 12943 3723
rect 14473 3689 14507 3723
rect 15301 3689 15335 3723
rect 16037 3689 16071 3723
rect 27261 3689 27295 3723
rect 32045 3689 32079 3723
rect 37657 3689 37691 3723
rect 44189 3689 44223 3723
rect 47593 3689 47627 3723
rect 50537 3689 50571 3723
rect 53481 3689 53515 3723
rect 54217 3689 54251 3723
rect 57805 3689 57839 3723
rect 7849 3621 7883 3655
rect 10977 3621 11011 3655
rect 20637 3621 20671 3655
rect 20821 3621 20855 3655
rect 22845 3621 22879 3655
rect 52101 3621 52135 3655
rect 9873 3553 9907 3587
rect 10057 3553 10091 3587
rect 10149 3553 10183 3587
rect 11161 3553 11195 3587
rect 22201 3553 22235 3587
rect 25881 3553 25915 3587
rect 30481 3553 30515 3587
rect 33149 3553 33183 3587
rect 35081 3553 35115 3587
rect 36277 3553 36311 3587
rect 42625 3553 42659 3587
rect 52837 3553 52871 3587
rect 57437 3553 57471 3587
rect 7113 3485 7147 3519
rect 9954 3485 9988 3519
rect 16589 3485 16623 3519
rect 17509 3485 17543 3519
rect 18429 3485 18463 3519
rect 19441 3485 19475 3519
rect 19717 3485 19751 3519
rect 21925 3485 21959 3519
rect 23397 3485 23431 3519
rect 23857 3485 23891 3519
rect 24961 3485 24995 3519
rect 26148 3485 26182 3519
rect 30297 3485 30331 3519
rect 31033 3485 31067 3519
rect 31217 3485 31251 3519
rect 31309 3485 31343 3519
rect 31401 3485 31435 3519
rect 32229 3485 32263 3519
rect 32505 3485 32539 3519
rect 32965 3485 32999 3519
rect 33885 3485 33919 3519
rect 34897 3485 34931 3519
rect 36533 3485 36567 3519
rect 39405 3485 39439 3519
rect 42533 3485 42567 3519
rect 42901 3485 42935 3519
rect 42993 3485 43027 3519
rect 43545 3485 43579 3519
rect 43693 3485 43727 3519
rect 43913 3485 43947 3519
rect 44051 3485 44085 3519
rect 45293 3485 45327 3519
rect 46949 3485 46983 3519
rect 47097 3485 47131 3519
rect 47414 3485 47448 3519
rect 48145 3485 48179 3519
rect 48605 3485 48639 3519
rect 48789 3485 48823 3519
rect 49157 3485 49191 3519
rect 49249 3485 49283 3519
rect 50353 3485 50387 3519
rect 51365 3485 51399 3519
rect 52653 3485 52687 3519
rect 54125 3485 54159 3519
rect 54769 3485 54803 3519
rect 54953 3485 54987 3519
rect 55597 3485 55631 3519
rect 57621 3485 57655 3519
rect 6929 3417 6963 3451
rect 7665 3417 7699 3451
rect 8401 3417 8435 3451
rect 10701 3417 10735 3451
rect 11713 3417 11747 3451
rect 12817 3417 12851 3451
rect 13553 3417 13587 3451
rect 14381 3417 14415 3451
rect 15209 3417 15243 3451
rect 15945 3417 15979 3451
rect 16865 3417 16899 3451
rect 17785 3417 17819 3451
rect 18705 3417 18739 3451
rect 20361 3417 20395 3451
rect 23029 3417 23063 3451
rect 23131 3417 23165 3451
rect 25237 3417 25271 3451
rect 29009 3417 29043 3451
rect 30205 3417 30239 3451
rect 32413 3417 32447 3451
rect 34161 3417 34195 3451
rect 38577 3417 38611 3451
rect 40141 3417 40175 3451
rect 40877 3417 40911 3451
rect 41889 3417 41923 3451
rect 43821 3417 43855 3451
rect 46305 3417 46339 3451
rect 47225 3417 47259 3451
rect 47317 3417 47351 3451
rect 51181 3417 51215 3451
rect 51917 3417 51951 3451
rect 53389 3417 53423 3451
rect 54861 3417 54895 3451
rect 55842 3417 55876 3451
rect 11805 3349 11839 3383
rect 13645 3349 13679 3383
rect 23213 3349 23247 3383
rect 23949 3349 23983 3383
rect 28273 3349 28307 3383
rect 29101 3349 29135 3383
rect 29837 3349 29871 3383
rect 31585 3349 31619 3383
rect 40233 3349 40267 3383
rect 40969 3349 41003 3383
rect 45385 3349 45419 3383
rect 46397 3349 46431 3383
rect 56977 3349 57011 3383
rect 7665 3145 7699 3179
rect 12173 3145 12207 3179
rect 13829 3145 13863 3179
rect 15301 3145 15335 3179
rect 25789 3145 25823 3179
rect 26617 3145 26651 3179
rect 41797 3145 41831 3179
rect 43913 3145 43947 3179
rect 44649 3145 44683 3179
rect 46857 3145 46891 3179
rect 48513 3145 48547 3179
rect 53113 3145 53147 3179
rect 54585 3145 54619 3179
rect 55321 3145 55355 3179
rect 56977 3145 57011 3179
rect 6009 3077 6043 3111
rect 8309 3077 8343 3111
rect 9689 3077 9723 3111
rect 18705 3077 18739 3111
rect 24676 3077 24710 3111
rect 34437 3077 34471 3111
rect 38577 3077 38611 3111
rect 40693 3077 40727 3111
rect 42809 3077 42843 3111
rect 42901 3077 42935 3111
rect 46029 3077 46063 3111
rect 46213 3077 46247 3111
rect 50261 3077 50295 3111
rect 5825 3009 5859 3043
rect 6837 3009 6871 3043
rect 7573 3009 7607 3043
rect 9045 3009 9079 3043
rect 9229 3009 9263 3043
rect 10977 3009 11011 3043
rect 11161 3009 11195 3043
rect 13001 3009 13035 3043
rect 13737 3009 13771 3043
rect 14473 3009 14507 3043
rect 15209 3009 15243 3043
rect 15853 3009 15887 3043
rect 17509 3009 17543 3043
rect 18429 3009 18463 3043
rect 19349 3009 19383 3043
rect 19625 3009 19659 3043
rect 21281 3009 21315 3043
rect 22293 3009 22327 3043
rect 22569 3009 22603 3043
rect 23489 3009 23523 3043
rect 24409 3009 24443 3043
rect 26249 3009 26283 3043
rect 26433 3009 26467 3043
rect 27169 3009 27203 3043
rect 28641 3009 28675 3043
rect 29929 3009 29963 3043
rect 30849 3009 30883 3043
rect 32321 3009 32355 3043
rect 33241 3009 33275 3043
rect 34161 3009 34195 3043
rect 35081 3009 35115 3043
rect 36001 3009 36035 3043
rect 37473 3009 37507 3043
rect 38393 3009 38427 3043
rect 38669 3009 38703 3043
rect 38813 3009 38847 3043
rect 39497 3009 39531 3043
rect 40509 3009 40543 3043
rect 41705 3009 41739 3043
rect 42625 3009 42659 3043
rect 43045 3009 43079 3043
rect 43821 3009 43855 3043
rect 44465 3009 44499 3043
rect 45293 3009 45327 3043
rect 45477 3009 45511 3043
rect 46765 3009 46799 3043
rect 47869 3009 47903 3043
rect 48017 3009 48051 3043
rect 48145 3009 48179 3043
rect 48237 3009 48271 3043
rect 48375 3009 48409 3043
rect 49157 3009 49191 3043
rect 50077 3009 50111 3043
rect 50813 3009 50847 3043
rect 51549 3009 51583 3043
rect 52929 3009 52963 3043
rect 53757 3009 53791 3043
rect 54401 3009 54435 3043
rect 55229 3009 55263 3043
rect 55965 3009 55999 3043
rect 56609 3009 56643 3043
rect 56793 3009 56827 3043
rect 58173 3009 58207 3043
rect 8493 2941 8527 2975
rect 10149 2941 10183 2975
rect 11713 2941 11747 2975
rect 13185 2941 13219 2975
rect 14657 2941 14691 2975
rect 16129 2941 16163 2975
rect 17785 2941 17819 2975
rect 20269 2941 20303 2975
rect 22845 2941 22879 2975
rect 23765 2941 23799 2975
rect 27353 2941 27387 2975
rect 29285 2941 29319 2975
rect 30205 2941 30239 2975
rect 31033 2941 31067 2975
rect 32505 2941 32539 2975
rect 33425 2941 33459 2975
rect 35265 2941 35299 2975
rect 36185 2941 36219 2975
rect 37657 2941 37691 2975
rect 39681 2941 39715 2975
rect 51733 2941 51767 2975
rect 9965 2873 9999 2907
rect 11989 2873 12023 2907
rect 20545 2873 20579 2907
rect 20729 2873 20763 2907
rect 38945 2873 38979 2907
rect 43177 2873 43211 2907
rect 53941 2873 53975 2907
rect 58357 2873 58391 2907
rect 6929 2805 6963 2839
rect 17049 2805 17083 2839
rect 21373 2805 21407 2839
rect 49249 2805 49283 2839
rect 50905 2805 50939 2839
rect 56057 2805 56091 2839
rect 7757 2601 7791 2635
rect 10333 2601 10367 2635
rect 12173 2601 12207 2635
rect 13645 2601 13679 2635
rect 22109 2601 22143 2635
rect 24593 2601 24627 2635
rect 41429 2601 41463 2635
rect 42993 2601 43027 2635
rect 44465 2601 44499 2635
rect 45385 2601 45419 2635
rect 46121 2601 46155 2635
rect 48605 2601 48639 2635
rect 49341 2601 49375 2635
rect 50537 2601 50571 2635
rect 51641 2601 51675 2635
rect 53113 2601 53147 2635
rect 7113 2533 7147 2567
rect 8585 2533 8619 2567
rect 9689 2533 9723 2567
rect 13001 2533 13035 2567
rect 14473 2533 14507 2567
rect 46949 2533 46983 2567
rect 55781 2533 55815 2567
rect 56517 2533 56551 2567
rect 58357 2533 58391 2567
rect 6009 2465 6043 2499
rect 15209 2465 15243 2499
rect 21281 2465 21315 2499
rect 54309 2465 54343 2499
rect 57345 2465 57379 2499
rect 7665 2397 7699 2431
rect 9505 2397 9539 2431
rect 10977 2397 11011 2431
rect 14933 2397 14967 2431
rect 15853 2397 15887 2431
rect 17049 2397 17083 2431
rect 17509 2397 17543 2431
rect 17785 2397 17819 2431
rect 18429 2397 18463 2431
rect 19625 2397 19659 2431
rect 20085 2397 20119 2431
rect 21005 2397 21039 2431
rect 22017 2397 22051 2431
rect 22661 2397 22695 2431
rect 23581 2397 23615 2431
rect 24961 2397 24995 2431
rect 25237 2397 25271 2431
rect 26157 2397 26191 2431
rect 27169 2397 27203 2431
rect 28733 2397 28767 2431
rect 30205 2397 30239 2431
rect 31125 2397 31159 2431
rect 32321 2397 32355 2431
rect 33241 2397 33275 2431
rect 34897 2397 34931 2431
rect 35817 2397 35851 2431
rect 37473 2397 37507 2431
rect 38393 2397 38427 2431
rect 40049 2397 40083 2431
rect 43637 2397 43671 2431
rect 47961 2397 47995 2431
rect 48109 2397 48143 2431
rect 48329 2397 48363 2431
rect 48426 2397 48460 2431
rect 51457 2397 51491 2431
rect 54033 2397 54067 2431
rect 57069 2397 57103 2431
rect 5825 2329 5859 2363
rect 6929 2329 6963 2363
rect 8401 2329 8435 2363
rect 10241 2329 10275 2363
rect 12081 2329 12115 2363
rect 12817 2329 12851 2363
rect 13553 2329 13587 2363
rect 16129 2329 16163 2363
rect 18705 2329 18739 2363
rect 20361 2329 20395 2363
rect 22937 2329 22971 2363
rect 23857 2329 23891 2363
rect 25513 2329 25547 2363
rect 26433 2329 26467 2363
rect 27445 2329 27479 2363
rect 29009 2329 29043 2363
rect 30481 2329 30515 2363
rect 31401 2329 31435 2363
rect 32597 2329 32631 2363
rect 33517 2329 33551 2363
rect 35173 2329 35207 2363
rect 36093 2329 36127 2363
rect 37749 2329 37783 2363
rect 38669 2329 38703 2363
rect 40325 2329 40359 2363
rect 41153 2329 41187 2363
rect 42717 2329 42751 2363
rect 44373 2329 44407 2363
rect 45293 2329 45327 2363
rect 46029 2329 46063 2363
rect 46765 2329 46799 2363
rect 48237 2329 48271 2363
rect 49249 2329 49283 2363
rect 50445 2329 50479 2363
rect 53021 2329 53055 2363
rect 55597 2329 55631 2363
rect 56333 2329 56367 2363
rect 58173 2329 58207 2363
rect 11069 2261 11103 2295
rect 28089 2261 28123 2295
rect 43729 2261 43763 2295
<< metal1 >>
rect 16390 59100 16396 59152
rect 16448 59140 16454 59152
rect 16942 59140 16948 59152
rect 16448 59112 16948 59140
rect 16448 59100 16454 59112
rect 16942 59100 16948 59112
rect 17000 59100 17006 59152
rect 18966 59100 18972 59152
rect 19024 59140 19030 59152
rect 19426 59140 19432 59152
rect 19024 59112 19432 59140
rect 19024 59100 19030 59112
rect 19426 59100 19432 59112
rect 19484 59100 19490 59152
rect 21542 59100 21548 59152
rect 21600 59140 21606 59152
rect 22094 59140 22100 59152
rect 21600 59112 22100 59140
rect 21600 59100 21606 59112
rect 22094 59100 22100 59112
rect 22152 59100 22158 59152
rect 36998 59100 37004 59152
rect 37056 59140 37062 59152
rect 37550 59140 37556 59152
rect 37056 59112 37556 59140
rect 37056 59100 37062 59112
rect 37550 59100 37556 59112
rect 37608 59100 37614 59152
rect 39574 59100 39580 59152
rect 39632 59140 39638 59152
rect 40034 59140 40040 59152
rect 39632 59112 40040 59140
rect 39632 59100 39638 59112
rect 40034 59100 40040 59112
rect 40092 59100 40098 59152
rect 55030 59100 55036 59152
rect 55088 59140 55094 59152
rect 55582 59140 55588 59152
rect 55088 59112 55588 59140
rect 55088 59100 55094 59112
rect 55582 59100 55588 59112
rect 55640 59100 55646 59152
rect 56778 57944 56784 57996
rect 56836 57984 56842 57996
rect 58986 57984 58992 57996
rect 56836 57956 58992 57984
rect 56836 57944 56842 57956
rect 58986 57944 58992 57956
rect 59044 57944 59050 57996
rect 1104 57690 58880 57712
rect 1104 57638 19574 57690
rect 19626 57638 19638 57690
rect 19690 57638 19702 57690
rect 19754 57638 19766 57690
rect 19818 57638 19830 57690
rect 19882 57638 50294 57690
rect 50346 57638 50358 57690
rect 50410 57638 50422 57690
rect 50474 57638 50486 57690
rect 50538 57638 50550 57690
rect 50602 57638 58880 57690
rect 1104 57616 58880 57638
rect 2222 57468 2228 57520
rect 2280 57508 2286 57520
rect 2409 57511 2467 57517
rect 2409 57508 2421 57511
rect 2280 57480 2421 57508
rect 2280 57468 2286 57480
rect 2409 57477 2421 57480
rect 2455 57477 2467 57511
rect 2409 57471 2467 57477
rect 3510 57468 3516 57520
rect 3568 57508 3574 57520
rect 4065 57511 4123 57517
rect 4065 57508 4077 57511
rect 3568 57480 4077 57508
rect 3568 57468 3574 57480
rect 4065 57477 4077 57480
rect 4111 57477 4123 57511
rect 4065 57471 4123 57477
rect 4798 57468 4804 57520
rect 4856 57508 4862 57520
rect 4985 57511 5043 57517
rect 4985 57508 4997 57511
rect 4856 57480 4997 57508
rect 4856 57468 4862 57480
rect 4985 57477 4997 57480
rect 5031 57477 5043 57511
rect 4985 57471 5043 57477
rect 7374 57468 7380 57520
rect 7432 57508 7438 57520
rect 7561 57511 7619 57517
rect 7561 57508 7573 57511
rect 7432 57480 7573 57508
rect 7432 57468 7438 57480
rect 7561 57477 7573 57480
rect 7607 57477 7619 57511
rect 7561 57471 7619 57477
rect 8662 57468 8668 57520
rect 8720 57508 8726 57520
rect 9217 57511 9275 57517
rect 9217 57508 9229 57511
rect 8720 57480 9229 57508
rect 8720 57468 8726 57480
rect 9217 57477 9229 57480
rect 9263 57477 9275 57511
rect 9217 57471 9275 57477
rect 9950 57468 9956 57520
rect 10008 57508 10014 57520
rect 10137 57511 10195 57517
rect 10137 57508 10149 57511
rect 10008 57480 10149 57508
rect 10008 57468 10014 57480
rect 10137 57477 10149 57480
rect 10183 57477 10195 57511
rect 10137 57471 10195 57477
rect 12526 57468 12532 57520
rect 12584 57508 12590 57520
rect 12713 57511 12771 57517
rect 12713 57508 12725 57511
rect 12584 57480 12725 57508
rect 12584 57468 12590 57480
rect 12713 57477 12725 57480
rect 12759 57477 12771 57511
rect 12713 57471 12771 57477
rect 16942 57468 16948 57520
rect 17000 57468 17006 57520
rect 17678 57468 17684 57520
rect 17736 57508 17742 57520
rect 17865 57511 17923 57517
rect 17865 57508 17877 57511
rect 17736 57480 17877 57508
rect 17736 57468 17742 57480
rect 17865 57477 17877 57480
rect 17911 57477 17923 57511
rect 17865 57471 17923 57477
rect 20254 57468 20260 57520
rect 20312 57508 20318 57520
rect 20441 57511 20499 57517
rect 20441 57508 20453 57511
rect 20312 57480 20453 57508
rect 20312 57468 20318 57480
rect 20441 57477 20453 57480
rect 20487 57477 20499 57511
rect 20441 57471 20499 57477
rect 22094 57468 22100 57520
rect 22152 57468 22158 57520
rect 22830 57468 22836 57520
rect 22888 57508 22894 57520
rect 23017 57511 23075 57517
rect 23017 57508 23029 57511
rect 22888 57480 23029 57508
rect 22888 57468 22894 57480
rect 23017 57477 23029 57480
rect 23063 57477 23075 57511
rect 23017 57471 23075 57477
rect 25406 57468 25412 57520
rect 25464 57508 25470 57520
rect 25593 57511 25651 57517
rect 25593 57508 25605 57511
rect 25464 57480 25605 57508
rect 25464 57468 25470 57480
rect 25593 57477 25605 57480
rect 25639 57477 25651 57511
rect 25593 57471 25651 57477
rect 26694 57468 26700 57520
rect 26752 57508 26758 57520
rect 27249 57511 27307 57517
rect 27249 57508 27261 57511
rect 26752 57480 27261 57508
rect 26752 57468 26758 57480
rect 27249 57477 27261 57480
rect 27295 57477 27307 57511
rect 27249 57471 27307 57477
rect 27982 57468 27988 57520
rect 28040 57508 28046 57520
rect 28169 57511 28227 57517
rect 28169 57508 28181 57511
rect 28040 57480 28181 57508
rect 28040 57468 28046 57480
rect 28169 57477 28181 57480
rect 28215 57477 28227 57511
rect 28169 57471 28227 57477
rect 29270 57468 29276 57520
rect 29328 57508 29334 57520
rect 29825 57511 29883 57517
rect 29825 57508 29837 57511
rect 29328 57480 29837 57508
rect 29328 57468 29334 57480
rect 29825 57477 29837 57480
rect 29871 57477 29883 57511
rect 29825 57471 29883 57477
rect 30558 57468 30564 57520
rect 30616 57508 30622 57520
rect 30745 57511 30803 57517
rect 30745 57508 30757 57511
rect 30616 57480 30757 57508
rect 30616 57468 30622 57480
rect 30745 57477 30757 57480
rect 30791 57477 30803 57511
rect 30745 57471 30803 57477
rect 31846 57468 31852 57520
rect 31904 57508 31910 57520
rect 32401 57511 32459 57517
rect 32401 57508 32413 57511
rect 31904 57480 32413 57508
rect 31904 57468 31910 57480
rect 32401 57477 32413 57480
rect 32447 57477 32459 57511
rect 32401 57471 32459 57477
rect 33134 57468 33140 57520
rect 33192 57508 33198 57520
rect 33321 57511 33379 57517
rect 33321 57508 33333 57511
rect 33192 57480 33333 57508
rect 33192 57468 33198 57480
rect 33321 57477 33333 57480
rect 33367 57477 33379 57511
rect 33321 57471 33379 57477
rect 34514 57468 34520 57520
rect 34572 57508 34578 57520
rect 34977 57511 35035 57517
rect 34977 57508 34989 57511
rect 34572 57480 34989 57508
rect 34572 57468 34578 57480
rect 34977 57477 34989 57480
rect 35023 57477 35035 57511
rect 34977 57471 35035 57477
rect 35894 57468 35900 57520
rect 35952 57468 35958 57520
rect 37550 57468 37556 57520
rect 37608 57468 37614 57520
rect 38286 57468 38292 57520
rect 38344 57508 38350 57520
rect 38473 57511 38531 57517
rect 38473 57508 38485 57511
rect 38344 57480 38485 57508
rect 38344 57468 38350 57480
rect 38473 57477 38485 57480
rect 38519 57477 38531 57511
rect 38473 57471 38531 57477
rect 40862 57468 40868 57520
rect 40920 57508 40926 57520
rect 41049 57511 41107 57517
rect 41049 57508 41061 57511
rect 40920 57480 41061 57508
rect 40920 57468 40926 57480
rect 41049 57477 41061 57480
rect 41095 57477 41107 57511
rect 41049 57471 41107 57477
rect 42150 57468 42156 57520
rect 42208 57508 42214 57520
rect 42705 57511 42763 57517
rect 42705 57508 42717 57511
rect 42208 57480 42717 57508
rect 42208 57468 42214 57480
rect 42705 57477 42717 57480
rect 42751 57477 42763 57511
rect 42705 57471 42763 57477
rect 43438 57468 43444 57520
rect 43496 57508 43502 57520
rect 43625 57511 43683 57517
rect 43625 57508 43637 57511
rect 43496 57480 43637 57508
rect 43496 57468 43502 57480
rect 43625 57477 43637 57480
rect 43671 57477 43683 57511
rect 43625 57471 43683 57477
rect 44726 57468 44732 57520
rect 44784 57508 44790 57520
rect 45281 57511 45339 57517
rect 45281 57508 45293 57511
rect 44784 57480 45293 57508
rect 44784 57468 44790 57480
rect 45281 57477 45293 57480
rect 45327 57477 45339 57511
rect 45281 57471 45339 57477
rect 47302 57468 47308 57520
rect 47360 57508 47366 57520
rect 47857 57511 47915 57517
rect 47857 57508 47869 57511
rect 47360 57480 47869 57508
rect 47360 57468 47366 57480
rect 47857 57477 47869 57480
rect 47903 57477 47915 57511
rect 47857 57471 47915 57477
rect 49878 57468 49884 57520
rect 49936 57508 49942 57520
rect 50433 57511 50491 57517
rect 50433 57508 50445 57511
rect 49936 57480 50445 57508
rect 49936 57468 49942 57480
rect 50433 57477 50445 57480
rect 50479 57477 50491 57511
rect 50433 57471 50491 57477
rect 53834 57468 53840 57520
rect 53892 57508 53898 57520
rect 53929 57511 53987 57517
rect 53929 57508 53941 57511
rect 53892 57480 53941 57508
rect 53892 57468 53898 57480
rect 53929 57477 53941 57480
rect 53975 57477 53987 57511
rect 53929 57471 53987 57477
rect 55582 57468 55588 57520
rect 55640 57468 55646 57520
rect 56318 57468 56324 57520
rect 56376 57508 56382 57520
rect 56413 57511 56471 57517
rect 56413 57508 56425 57511
rect 56376 57480 56425 57508
rect 56376 57468 56382 57480
rect 56413 57477 56425 57480
rect 56459 57477 56471 57511
rect 56413 57471 56471 57477
rect 57149 57511 57207 57517
rect 57149 57477 57161 57511
rect 57195 57508 57207 57511
rect 58986 57508 58992 57520
rect 57195 57480 58992 57508
rect 57195 57477 57207 57480
rect 57149 57471 57207 57477
rect 58986 57468 58992 57480
rect 59044 57468 59050 57520
rect 6086 57400 6092 57452
rect 6144 57440 6150 57452
rect 6549 57443 6607 57449
rect 6549 57440 6561 57443
rect 6144 57412 6561 57440
rect 6144 57400 6150 57412
rect 6549 57409 6561 57412
rect 6595 57409 6607 57443
rect 6549 57403 6607 57409
rect 11238 57400 11244 57452
rect 11296 57440 11302 57452
rect 11701 57443 11759 57449
rect 11701 57440 11713 57443
rect 11296 57412 11713 57440
rect 11296 57400 11302 57412
rect 11701 57409 11713 57412
rect 11747 57409 11759 57443
rect 11701 57403 11759 57409
rect 13814 57400 13820 57452
rect 13872 57440 13878 57452
rect 14277 57443 14335 57449
rect 14277 57440 14289 57443
rect 13872 57412 14289 57440
rect 13872 57400 13878 57412
rect 14277 57409 14289 57412
rect 14323 57409 14335 57443
rect 14277 57403 14335 57409
rect 15194 57400 15200 57452
rect 15252 57400 15258 57452
rect 19426 57400 19432 57452
rect 19484 57400 19490 57452
rect 24118 57400 24124 57452
rect 24176 57440 24182 57452
rect 24581 57443 24639 57449
rect 24581 57440 24593 57443
rect 24176 57412 24593 57440
rect 24176 57400 24182 57412
rect 24581 57409 24593 57412
rect 24627 57409 24639 57443
rect 24581 57403 24639 57409
rect 40034 57400 40040 57452
rect 40092 57400 40098 57452
rect 46014 57400 46020 57452
rect 46072 57440 46078 57452
rect 46109 57443 46167 57449
rect 46109 57440 46121 57443
rect 46072 57412 46121 57440
rect 46072 57400 46078 57412
rect 46109 57409 46121 57412
rect 46155 57409 46167 57443
rect 46109 57403 46167 57409
rect 48590 57400 48596 57452
rect 48648 57440 48654 57452
rect 48685 57443 48743 57449
rect 48685 57440 48697 57443
rect 48648 57412 48697 57440
rect 48648 57400 48654 57412
rect 48685 57409 48697 57412
rect 48731 57409 48743 57443
rect 48685 57403 48743 57409
rect 51166 57400 51172 57452
rect 51224 57440 51230 57452
rect 51261 57443 51319 57449
rect 51261 57440 51273 57443
rect 51224 57412 51273 57440
rect 51224 57400 51230 57412
rect 51261 57409 51273 57412
rect 51307 57409 51319 57443
rect 51261 57403 51319 57409
rect 52454 57400 52460 57452
rect 52512 57440 52518 57452
rect 52917 57443 52975 57449
rect 52917 57440 52929 57443
rect 52512 57412 52929 57440
rect 52512 57400 52518 57412
rect 52917 57409 52929 57412
rect 52963 57409 52975 57443
rect 52917 57403 52975 57409
rect 58161 57443 58219 57449
rect 58161 57409 58173 57443
rect 58207 57440 58219 57443
rect 58894 57440 58900 57452
rect 58207 57412 58900 57440
rect 58207 57409 58219 57412
rect 58161 57403 58219 57409
rect 58894 57400 58900 57412
rect 58952 57400 58958 57452
rect 14553 57375 14611 57381
rect 14553 57341 14565 57375
rect 14599 57372 14611 57375
rect 26878 57372 26884 57384
rect 14599 57344 26884 57372
rect 14599 57341 14611 57344
rect 14553 57335 14611 57341
rect 26878 57332 26884 57344
rect 26936 57332 26942 57384
rect 2593 57307 2651 57313
rect 2593 57273 2605 57307
rect 2639 57304 2651 57307
rect 3418 57304 3424 57316
rect 2639 57276 3424 57304
rect 2639 57273 2651 57276
rect 2593 57267 2651 57273
rect 3418 57264 3424 57276
rect 3476 57264 3482 57316
rect 17126 57264 17132 57316
rect 17184 57264 17190 57316
rect 52638 57264 52644 57316
rect 52696 57304 52702 57316
rect 56597 57307 56655 57313
rect 56597 57304 56609 57307
rect 52696 57276 56609 57304
rect 52696 57264 52702 57276
rect 56597 57273 56609 57276
rect 56643 57273 56655 57307
rect 56597 57267 56655 57273
rect 56686 57264 56692 57316
rect 56744 57304 56750 57316
rect 58802 57304 58808 57316
rect 56744 57276 58808 57304
rect 56744 57264 56750 57276
rect 58802 57264 58808 57276
rect 58860 57264 58866 57316
rect 3970 57196 3976 57248
rect 4028 57236 4034 57248
rect 4157 57239 4215 57245
rect 4157 57236 4169 57239
rect 4028 57208 4169 57236
rect 4028 57196 4034 57208
rect 4157 57205 4169 57208
rect 4203 57205 4215 57239
rect 4157 57199 4215 57205
rect 4706 57196 4712 57248
rect 4764 57236 4770 57248
rect 5077 57239 5135 57245
rect 5077 57236 5089 57239
rect 4764 57208 5089 57236
rect 4764 57196 4770 57208
rect 5077 57205 5089 57208
rect 5123 57205 5135 57239
rect 5077 57199 5135 57205
rect 6730 57196 6736 57248
rect 6788 57196 6794 57248
rect 7374 57196 7380 57248
rect 7432 57236 7438 57248
rect 7653 57239 7711 57245
rect 7653 57236 7665 57239
rect 7432 57208 7665 57236
rect 7432 57196 7438 57208
rect 7653 57205 7665 57208
rect 7699 57205 7711 57239
rect 7653 57199 7711 57205
rect 9122 57196 9128 57248
rect 9180 57236 9186 57248
rect 9309 57239 9367 57245
rect 9309 57236 9321 57239
rect 9180 57208 9321 57236
rect 9180 57196 9186 57208
rect 9309 57205 9321 57208
rect 9355 57205 9367 57239
rect 9309 57199 9367 57205
rect 9950 57196 9956 57248
rect 10008 57236 10014 57248
rect 10229 57239 10287 57245
rect 10229 57236 10241 57239
rect 10008 57208 10241 57236
rect 10008 57196 10014 57208
rect 10229 57205 10241 57208
rect 10275 57205 10287 57239
rect 10229 57199 10287 57205
rect 11882 57196 11888 57248
rect 11940 57196 11946 57248
rect 12802 57196 12808 57248
rect 12860 57196 12866 57248
rect 15378 57196 15384 57248
rect 15436 57196 15442 57248
rect 17954 57196 17960 57248
rect 18012 57196 18018 57248
rect 19613 57239 19671 57245
rect 19613 57205 19625 57239
rect 19659 57236 19671 57239
rect 19978 57236 19984 57248
rect 19659 57208 19984 57236
rect 19659 57205 19671 57208
rect 19613 57199 19671 57205
rect 19978 57196 19984 57208
rect 20036 57196 20042 57248
rect 20162 57196 20168 57248
rect 20220 57236 20226 57248
rect 20533 57239 20591 57245
rect 20533 57236 20545 57239
rect 20220 57208 20545 57236
rect 20220 57196 20226 57208
rect 20533 57205 20545 57208
rect 20579 57205 20591 57239
rect 20533 57199 20591 57205
rect 22186 57196 22192 57248
rect 22244 57196 22250 57248
rect 22646 57196 22652 57248
rect 22704 57236 22710 57248
rect 23109 57239 23167 57245
rect 23109 57236 23121 57239
rect 22704 57208 23121 57236
rect 22704 57196 22710 57208
rect 23109 57205 23121 57208
rect 23155 57205 23167 57239
rect 23109 57199 23167 57205
rect 24762 57196 24768 57248
rect 24820 57196 24826 57248
rect 25682 57196 25688 57248
rect 25740 57196 25746 57248
rect 26694 57196 26700 57248
rect 26752 57236 26758 57248
rect 27341 57239 27399 57245
rect 27341 57236 27353 57239
rect 26752 57208 27353 57236
rect 26752 57196 26758 57208
rect 27341 57205 27353 57208
rect 27387 57205 27399 57239
rect 27341 57199 27399 57205
rect 27982 57196 27988 57248
rect 28040 57236 28046 57248
rect 28261 57239 28319 57245
rect 28261 57236 28273 57239
rect 28040 57208 28273 57236
rect 28040 57196 28046 57208
rect 28261 57205 28273 57208
rect 28307 57205 28319 57239
rect 28261 57199 28319 57205
rect 29914 57196 29920 57248
rect 29972 57196 29978 57248
rect 30834 57196 30840 57248
rect 30892 57196 30898 57248
rect 31202 57196 31208 57248
rect 31260 57236 31266 57248
rect 32493 57239 32551 57245
rect 32493 57236 32505 57239
rect 31260 57208 32505 57236
rect 31260 57196 31266 57208
rect 32493 57205 32505 57208
rect 32539 57205 32551 57239
rect 32493 57199 32551 57205
rect 33410 57196 33416 57248
rect 33468 57196 33474 57248
rect 34790 57196 34796 57248
rect 34848 57236 34854 57248
rect 35069 57239 35127 57245
rect 35069 57236 35081 57239
rect 34848 57208 35081 57236
rect 34848 57196 34854 57208
rect 35069 57205 35081 57208
rect 35115 57205 35127 57239
rect 35069 57199 35127 57205
rect 35618 57196 35624 57248
rect 35676 57236 35682 57248
rect 35989 57239 36047 57245
rect 35989 57236 36001 57239
rect 35676 57208 36001 57236
rect 35676 57196 35682 57208
rect 35989 57205 36001 57208
rect 36035 57205 36047 57239
rect 35989 57199 36047 57205
rect 37090 57196 37096 57248
rect 37148 57236 37154 57248
rect 37645 57239 37703 57245
rect 37645 57236 37657 57239
rect 37148 57208 37657 57236
rect 37148 57196 37154 57208
rect 37645 57205 37657 57208
rect 37691 57205 37703 57239
rect 37645 57199 37703 57205
rect 37918 57196 37924 57248
rect 37976 57236 37982 57248
rect 38565 57239 38623 57245
rect 38565 57236 38577 57239
rect 37976 57208 38577 57236
rect 37976 57196 37982 57208
rect 38565 57205 38577 57208
rect 38611 57205 38623 57239
rect 38565 57199 38623 57205
rect 39298 57196 39304 57248
rect 39356 57236 39362 57248
rect 40221 57239 40279 57245
rect 40221 57236 40233 57239
rect 39356 57208 40233 57236
rect 39356 57196 39362 57208
rect 40221 57205 40233 57208
rect 40267 57205 40279 57239
rect 40221 57199 40279 57205
rect 40310 57196 40316 57248
rect 40368 57236 40374 57248
rect 41141 57239 41199 57245
rect 41141 57236 41153 57239
rect 40368 57208 41153 57236
rect 40368 57196 40374 57208
rect 41141 57205 41153 57208
rect 41187 57205 41199 57239
rect 41141 57199 41199 57205
rect 41690 57196 41696 57248
rect 41748 57236 41754 57248
rect 42797 57239 42855 57245
rect 42797 57236 42809 57239
rect 41748 57208 42809 57236
rect 41748 57196 41754 57208
rect 42797 57205 42809 57208
rect 42843 57205 42855 57239
rect 42797 57199 42855 57205
rect 43622 57196 43628 57248
rect 43680 57236 43686 57248
rect 43717 57239 43775 57245
rect 43717 57236 43729 57239
rect 43680 57208 43729 57236
rect 43680 57196 43686 57208
rect 43717 57205 43729 57208
rect 43763 57205 43775 57239
rect 43717 57199 43775 57205
rect 45370 57196 45376 57248
rect 45428 57196 45434 57248
rect 46290 57196 46296 57248
rect 46348 57196 46354 57248
rect 46382 57196 46388 57248
rect 46440 57236 46446 57248
rect 47949 57239 48007 57245
rect 47949 57236 47961 57239
rect 46440 57208 47961 57236
rect 46440 57196 46446 57208
rect 47949 57205 47961 57208
rect 47995 57205 48007 57239
rect 47949 57199 48007 57205
rect 48866 57196 48872 57248
rect 48924 57196 48930 57248
rect 49050 57196 49056 57248
rect 49108 57236 49114 57248
rect 50525 57239 50583 57245
rect 50525 57236 50537 57239
rect 49108 57208 50537 57236
rect 49108 57196 49114 57208
rect 50525 57205 50537 57208
rect 50571 57205 50583 57239
rect 50525 57199 50583 57205
rect 51442 57196 51448 57248
rect 51500 57196 51506 57248
rect 51718 57196 51724 57248
rect 51776 57236 51782 57248
rect 53101 57239 53159 57245
rect 53101 57236 53113 57239
rect 51776 57208 53113 57236
rect 51776 57196 51782 57208
rect 53101 57205 53113 57208
rect 53147 57205 53159 57239
rect 53101 57199 53159 57205
rect 53926 57196 53932 57248
rect 53984 57236 53990 57248
rect 54021 57239 54079 57245
rect 54021 57236 54033 57239
rect 53984 57208 54033 57236
rect 53984 57196 53990 57208
rect 54021 57205 54033 57208
rect 54067 57205 54079 57239
rect 54021 57199 54079 57205
rect 54110 57196 54116 57248
rect 54168 57236 54174 57248
rect 55677 57239 55735 57245
rect 55677 57236 55689 57239
rect 54168 57208 55689 57236
rect 54168 57196 54174 57208
rect 55677 57205 55689 57208
rect 55723 57205 55735 57239
rect 55677 57199 55735 57205
rect 57238 57196 57244 57248
rect 57296 57196 57302 57248
rect 58250 57196 58256 57248
rect 58308 57196 58314 57248
rect 1104 57146 58880 57168
rect 1104 57094 4214 57146
rect 4266 57094 4278 57146
rect 4330 57094 4342 57146
rect 4394 57094 4406 57146
rect 4458 57094 4470 57146
rect 4522 57094 34934 57146
rect 34986 57094 34998 57146
rect 35050 57094 35062 57146
rect 35114 57094 35126 57146
rect 35178 57094 35190 57146
rect 35242 57094 58880 57146
rect 1104 57072 58880 57094
rect 22186 56992 22192 57044
rect 22244 57032 22250 57044
rect 31570 57032 31576 57044
rect 22244 57004 31576 57032
rect 22244 56992 22250 57004
rect 31570 56992 31576 57004
rect 31628 56992 31634 57044
rect 57422 56992 57428 57044
rect 57480 57032 57486 57044
rect 58986 57032 58992 57044
rect 57480 57004 58992 57032
rect 57480 56992 57486 57004
rect 58986 56992 58992 57004
rect 59044 56992 59050 57044
rect 53558 56924 53564 56976
rect 53616 56964 53622 56976
rect 58250 56964 58256 56976
rect 53616 56936 58256 56964
rect 53616 56924 53622 56936
rect 58250 56924 58256 56936
rect 58308 56924 58314 56976
rect 17954 56856 17960 56908
rect 18012 56896 18018 56908
rect 30466 56896 30472 56908
rect 18012 56868 30472 56896
rect 18012 56856 18018 56868
rect 30466 56856 30472 56868
rect 30524 56856 30530 56908
rect 58986 56896 58992 56908
rect 56060 56868 58992 56896
rect 56060 56837 56088 56868
rect 58986 56856 58992 56868
rect 59044 56856 59050 56908
rect 56045 56831 56103 56837
rect 56045 56797 56057 56831
rect 56091 56797 56103 56831
rect 56045 56791 56103 56797
rect 56778 56788 56784 56840
rect 56836 56788 56842 56840
rect 57606 56788 57612 56840
rect 57664 56828 57670 56840
rect 57793 56831 57851 56837
rect 57793 56828 57805 56831
rect 57664 56800 57805 56828
rect 57664 56788 57670 56800
rect 57793 56797 57805 56800
rect 57839 56797 57851 56831
rect 57793 56791 57851 56797
rect 52454 56720 52460 56772
rect 52512 56760 52518 56772
rect 57057 56763 57115 56769
rect 57057 56760 57069 56763
rect 52512 56732 57069 56760
rect 52512 56720 52518 56732
rect 57057 56729 57069 56732
rect 57103 56729 57115 56763
rect 57057 56723 57115 56729
rect 58161 56763 58219 56769
rect 58161 56729 58173 56763
rect 58207 56760 58219 56763
rect 59446 56760 59452 56772
rect 58207 56732 59452 56760
rect 58207 56729 58219 56732
rect 58161 56723 58219 56729
rect 59446 56720 59452 56732
rect 59504 56720 59510 56772
rect 56226 56652 56232 56704
rect 56284 56652 56290 56704
rect 1104 56602 58880 56624
rect 1104 56550 19574 56602
rect 19626 56550 19638 56602
rect 19690 56550 19702 56602
rect 19754 56550 19766 56602
rect 19818 56550 19830 56602
rect 19882 56550 50294 56602
rect 50346 56550 50358 56602
rect 50410 56550 50422 56602
rect 50474 56550 50486 56602
rect 50538 56550 50550 56602
rect 50602 56550 58880 56602
rect 1104 56528 58880 56550
rect 58710 56488 58716 56500
rect 55876 56460 58716 56488
rect 55876 56429 55904 56460
rect 58710 56448 58716 56460
rect 58768 56448 58774 56500
rect 55861 56423 55919 56429
rect 55861 56389 55873 56423
rect 55907 56389 55919 56423
rect 55861 56383 55919 56389
rect 56597 56423 56655 56429
rect 56597 56389 56609 56423
rect 56643 56420 56655 56423
rect 56686 56420 56692 56432
rect 56643 56392 56692 56420
rect 56643 56389 56655 56392
rect 56597 56383 56655 56389
rect 56686 56380 56692 56392
rect 56744 56380 56750 56432
rect 57333 56423 57391 56429
rect 57333 56389 57345 56423
rect 57379 56420 57391 56423
rect 58986 56420 58992 56432
rect 57379 56392 58992 56420
rect 57379 56389 57391 56392
rect 57333 56383 57391 56389
rect 58986 56380 58992 56392
rect 59044 56380 59050 56432
rect 934 56312 940 56364
rect 992 56352 998 56364
rect 1581 56355 1639 56361
rect 1581 56352 1593 56355
rect 992 56324 1593 56352
rect 992 56312 998 56324
rect 1581 56321 1593 56324
rect 1627 56321 1639 56355
rect 1581 56315 1639 56321
rect 58158 56312 58164 56364
rect 58216 56312 58222 56364
rect 1857 56287 1915 56293
rect 1857 56253 1869 56287
rect 1903 56284 1915 56287
rect 18598 56284 18604 56296
rect 1903 56256 18604 56284
rect 1903 56253 1915 56256
rect 1857 56247 1915 56253
rect 18598 56244 18604 56256
rect 18656 56244 18662 56296
rect 55214 56244 55220 56296
rect 55272 56284 55278 56296
rect 58345 56287 58403 56293
rect 58345 56284 58357 56287
rect 55272 56256 58357 56284
rect 55272 56244 55278 56256
rect 58345 56253 58357 56256
rect 58391 56253 58403 56287
rect 58345 56247 58403 56253
rect 53834 56176 53840 56228
rect 53892 56216 53898 56228
rect 57517 56219 57575 56225
rect 57517 56216 57529 56219
rect 53892 56188 57529 56216
rect 53892 56176 53898 56188
rect 57517 56185 57529 56188
rect 57563 56185 57575 56219
rect 57517 56179 57575 56185
rect 52546 56108 52552 56160
rect 52604 56148 52610 56160
rect 55953 56151 56011 56157
rect 55953 56148 55965 56151
rect 52604 56120 55965 56148
rect 52604 56108 52610 56120
rect 55953 56117 55965 56120
rect 55999 56117 56011 56151
rect 55953 56111 56011 56117
rect 56042 56108 56048 56160
rect 56100 56148 56106 56160
rect 56689 56151 56747 56157
rect 56689 56148 56701 56151
rect 56100 56120 56701 56148
rect 56100 56108 56106 56120
rect 56689 56117 56701 56120
rect 56735 56117 56747 56151
rect 56689 56111 56747 56117
rect 1104 56058 58880 56080
rect 1104 56006 4214 56058
rect 4266 56006 4278 56058
rect 4330 56006 4342 56058
rect 4394 56006 4406 56058
rect 4458 56006 4470 56058
rect 4522 56006 34934 56058
rect 34986 56006 34998 56058
rect 35050 56006 35062 56058
rect 35114 56006 35126 56058
rect 35178 56006 35190 56058
rect 35242 56006 58880 56058
rect 1104 55984 58880 56006
rect 26786 55836 26792 55888
rect 26844 55876 26850 55888
rect 52454 55876 52460 55888
rect 26844 55848 52460 55876
rect 26844 55836 26850 55848
rect 52454 55836 52460 55848
rect 52512 55836 52518 55888
rect 53190 55836 53196 55888
rect 53248 55876 53254 55888
rect 58253 55879 58311 55885
rect 58253 55876 58265 55879
rect 53248 55848 58265 55876
rect 53248 55836 53254 55848
rect 58253 55845 58265 55848
rect 58299 55845 58311 55879
rect 58253 55839 58311 55845
rect 934 55700 940 55752
rect 992 55740 998 55752
rect 1581 55743 1639 55749
rect 1581 55740 1593 55743
rect 992 55712 1593 55740
rect 992 55700 998 55712
rect 1581 55709 1593 55712
rect 1627 55709 1639 55743
rect 1581 55703 1639 55709
rect 57422 55700 57428 55752
rect 57480 55700 57486 55752
rect 58069 55743 58127 55749
rect 58069 55709 58081 55743
rect 58115 55740 58127 55743
rect 58986 55740 58992 55752
rect 58115 55712 58992 55740
rect 58115 55709 58127 55712
rect 58069 55703 58127 55709
rect 58986 55700 58992 55712
rect 59044 55700 59050 55752
rect 1857 55675 1915 55681
rect 1857 55641 1869 55675
rect 1903 55672 1915 55675
rect 21358 55672 21364 55684
rect 1903 55644 21364 55672
rect 1903 55641 1915 55644
rect 1857 55635 1915 55641
rect 21358 55632 21364 55644
rect 21416 55632 21422 55684
rect 57514 55564 57520 55616
rect 57572 55564 57578 55616
rect 1104 55514 58880 55536
rect 1104 55462 19574 55514
rect 19626 55462 19638 55514
rect 19690 55462 19702 55514
rect 19754 55462 19766 55514
rect 19818 55462 19830 55514
rect 19882 55462 50294 55514
rect 50346 55462 50358 55514
rect 50410 55462 50422 55514
rect 50474 55462 50486 55514
rect 50538 55462 50550 55514
rect 50602 55462 58880 55514
rect 1104 55440 58880 55462
rect 58253 55403 58311 55409
rect 58253 55369 58265 55403
rect 58299 55400 58311 55403
rect 59078 55400 59084 55412
rect 58299 55372 59084 55400
rect 58299 55369 58311 55372
rect 58253 55363 58311 55369
rect 59078 55360 59084 55372
rect 59136 55360 59142 55412
rect 1026 55224 1032 55276
rect 1084 55264 1090 55276
rect 1673 55267 1731 55273
rect 1673 55264 1685 55267
rect 1084 55236 1685 55264
rect 1084 55224 1090 55236
rect 1673 55233 1685 55236
rect 1719 55233 1731 55267
rect 1673 55227 1731 55233
rect 58069 55267 58127 55273
rect 58069 55233 58081 55267
rect 58115 55264 58127 55267
rect 58802 55264 58808 55276
rect 58115 55236 58808 55264
rect 58115 55233 58127 55236
rect 58069 55227 58127 55233
rect 58802 55224 58808 55236
rect 58860 55224 58866 55276
rect 1946 55020 1952 55072
rect 2004 55020 2010 55072
rect 1104 54970 58880 54992
rect 1104 54918 4214 54970
rect 4266 54918 4278 54970
rect 4330 54918 4342 54970
rect 4394 54918 4406 54970
rect 4458 54918 4470 54970
rect 4522 54918 34934 54970
rect 34986 54918 34998 54970
rect 35050 54918 35062 54970
rect 35114 54918 35126 54970
rect 35178 54918 35190 54970
rect 35242 54918 58880 54970
rect 1104 54896 58880 54918
rect 57425 54655 57483 54661
rect 57425 54621 57437 54655
rect 57471 54652 57483 54655
rect 58986 54652 58992 54664
rect 57471 54624 58992 54652
rect 57471 54621 57483 54624
rect 57425 54615 57483 54621
rect 58986 54612 58992 54624
rect 59044 54612 59050 54664
rect 934 54544 940 54596
rect 992 54584 998 54596
rect 1673 54587 1731 54593
rect 1673 54584 1685 54587
rect 992 54556 1685 54584
rect 992 54544 998 54556
rect 1673 54553 1685 54556
rect 1719 54553 1731 54587
rect 1673 54547 1731 54553
rect 2041 54587 2099 54593
rect 2041 54553 2053 54587
rect 2087 54584 2099 54587
rect 2682 54584 2688 54596
rect 2087 54556 2688 54584
rect 2087 54553 2099 54556
rect 2041 54547 2099 54553
rect 2682 54544 2688 54556
rect 2740 54544 2746 54596
rect 58161 54587 58219 54593
rect 58161 54553 58173 54587
rect 58207 54584 58219 54587
rect 58894 54584 58900 54596
rect 58207 54556 58900 54584
rect 58207 54553 58219 54556
rect 58161 54547 58219 54553
rect 58894 54544 58900 54556
rect 58952 54544 58958 54596
rect 56594 54476 56600 54528
rect 56652 54516 56658 54528
rect 57517 54519 57575 54525
rect 57517 54516 57529 54519
rect 56652 54488 57529 54516
rect 56652 54476 56658 54488
rect 57517 54485 57529 54488
rect 57563 54485 57575 54519
rect 57517 54479 57575 54485
rect 58250 54476 58256 54528
rect 58308 54476 58314 54528
rect 1104 54426 58880 54448
rect 1104 54374 19574 54426
rect 19626 54374 19638 54426
rect 19690 54374 19702 54426
rect 19754 54374 19766 54426
rect 19818 54374 19830 54426
rect 19882 54374 50294 54426
rect 50346 54374 50358 54426
rect 50410 54374 50422 54426
rect 50474 54374 50486 54426
rect 50538 54374 50550 54426
rect 50602 54374 58880 54426
rect 1104 54352 58880 54374
rect 1026 54136 1032 54188
rect 1084 54176 1090 54188
rect 1673 54179 1731 54185
rect 1673 54176 1685 54179
rect 1084 54148 1685 54176
rect 1084 54136 1090 54148
rect 1673 54145 1685 54148
rect 1719 54145 1731 54179
rect 1673 54139 1731 54145
rect 58069 54179 58127 54185
rect 58069 54145 58081 54179
rect 58115 54176 58127 54179
rect 58986 54176 58992 54188
rect 58115 54148 58992 54176
rect 58115 54145 58127 54148
rect 58069 54139 58127 54145
rect 58986 54136 58992 54148
rect 59044 54136 59050 54188
rect 1949 53975 2007 53981
rect 1949 53941 1961 53975
rect 1995 53972 2007 53975
rect 2590 53972 2596 53984
rect 1995 53944 2596 53972
rect 1995 53941 2007 53944
rect 1949 53935 2007 53941
rect 2590 53932 2596 53944
rect 2648 53932 2654 53984
rect 58253 53975 58311 53981
rect 58253 53941 58265 53975
rect 58299 53972 58311 53975
rect 58526 53972 58532 53984
rect 58299 53944 58532 53972
rect 58299 53941 58311 53944
rect 58253 53935 58311 53941
rect 58526 53932 58532 53944
rect 58584 53932 58590 53984
rect 1104 53882 58880 53904
rect 1104 53830 4214 53882
rect 4266 53830 4278 53882
rect 4330 53830 4342 53882
rect 4394 53830 4406 53882
rect 4458 53830 4470 53882
rect 4522 53830 34934 53882
rect 34986 53830 34998 53882
rect 35050 53830 35062 53882
rect 35114 53830 35126 53882
rect 35178 53830 35190 53882
rect 35242 53830 58880 53882
rect 1104 53808 58880 53830
rect 934 53456 940 53508
rect 992 53496 998 53508
rect 1673 53499 1731 53505
rect 1673 53496 1685 53499
rect 992 53468 1685 53496
rect 992 53456 998 53468
rect 1673 53465 1685 53468
rect 1719 53465 1731 53499
rect 1673 53459 1731 53465
rect 58158 53456 58164 53508
rect 58216 53456 58222 53508
rect 58345 53499 58403 53505
rect 58345 53465 58357 53499
rect 58391 53496 58403 53499
rect 58434 53496 58440 53508
rect 58391 53468 58440 53496
rect 58391 53465 58403 53468
rect 58345 53459 58403 53465
rect 58434 53456 58440 53468
rect 58492 53456 58498 53508
rect 1949 53431 2007 53437
rect 1949 53397 1961 53431
rect 1995 53428 2007 53431
rect 47854 53428 47860 53440
rect 1995 53400 47860 53428
rect 1995 53397 2007 53400
rect 1949 53391 2007 53397
rect 47854 53388 47860 53400
rect 47912 53388 47918 53440
rect 1104 53338 58880 53360
rect 1104 53286 19574 53338
rect 19626 53286 19638 53338
rect 19690 53286 19702 53338
rect 19754 53286 19766 53338
rect 19818 53286 19830 53338
rect 19882 53286 50294 53338
rect 50346 53286 50358 53338
rect 50410 53286 50422 53338
rect 50474 53286 50486 53338
rect 50538 53286 50550 53338
rect 50602 53286 58880 53338
rect 1104 53264 58880 53286
rect 1946 53184 1952 53236
rect 2004 53224 2010 53236
rect 2004 53196 45554 53224
rect 2004 53184 2010 53196
rect 1026 53048 1032 53100
rect 1084 53088 1090 53100
rect 1673 53091 1731 53097
rect 1673 53088 1685 53091
rect 1084 53060 1685 53088
rect 1084 53048 1090 53060
rect 1673 53057 1685 53060
rect 1719 53057 1731 53091
rect 45526 53088 45554 53196
rect 48225 53091 48283 53097
rect 48225 53088 48237 53091
rect 45526 53060 48237 53088
rect 1673 53051 1731 53057
rect 48225 53057 48237 53060
rect 48271 53057 48283 53091
rect 48225 53051 48283 53057
rect 48409 53091 48467 53097
rect 48409 53057 48421 53091
rect 48455 53057 48467 53091
rect 48409 53051 48467 53057
rect 48777 53091 48835 53097
rect 48777 53057 48789 53091
rect 48823 53088 48835 53091
rect 52454 53088 52460 53100
rect 48823 53060 52460 53088
rect 48823 53057 48835 53060
rect 48777 53051 48835 53057
rect 48130 52980 48136 53032
rect 48188 53020 48194 53032
rect 48424 53020 48452 53051
rect 52454 53048 52460 53060
rect 52512 53048 52518 53100
rect 58069 53091 58127 53097
rect 58069 53057 58081 53091
rect 58115 53088 58127 53091
rect 58894 53088 58900 53100
rect 58115 53060 58900 53088
rect 58115 53057 58127 53060
rect 58069 53051 58127 53057
rect 58894 53048 58900 53060
rect 58952 53048 58958 53100
rect 48188 52992 48452 53020
rect 48188 52980 48194 52992
rect 48498 52980 48504 53032
rect 48556 53020 48562 53032
rect 48685 53023 48743 53029
rect 48685 53020 48697 53023
rect 48556 52992 48697 53020
rect 48556 52980 48562 52992
rect 48685 52989 48697 52992
rect 48731 52989 48743 53023
rect 48685 52983 48743 52989
rect 1949 52887 2007 52893
rect 1949 52853 1961 52887
rect 1995 52884 2007 52887
rect 11698 52884 11704 52896
rect 1995 52856 11704 52884
rect 1995 52853 2007 52856
rect 1949 52847 2007 52853
rect 11698 52844 11704 52856
rect 11756 52844 11762 52896
rect 48038 52844 48044 52896
rect 48096 52844 48102 52896
rect 58066 52844 58072 52896
rect 58124 52884 58130 52896
rect 58253 52887 58311 52893
rect 58253 52884 58265 52887
rect 58124 52856 58265 52884
rect 58124 52844 58130 52856
rect 58253 52853 58265 52856
rect 58299 52853 58311 52887
rect 58253 52847 58311 52853
rect 1104 52794 58880 52816
rect 1104 52742 4214 52794
rect 4266 52742 4278 52794
rect 4330 52742 4342 52794
rect 4394 52742 4406 52794
rect 4458 52742 4470 52794
rect 4522 52742 34934 52794
rect 34986 52742 34998 52794
rect 35050 52742 35062 52794
rect 35114 52742 35126 52794
rect 35178 52742 35190 52794
rect 35242 52742 58880 52794
rect 1104 52720 58880 52742
rect 47670 52640 47676 52692
rect 47728 52640 47734 52692
rect 55950 52572 55956 52624
rect 56008 52612 56014 52624
rect 58158 52612 58164 52624
rect 56008 52584 58164 52612
rect 56008 52572 56014 52584
rect 58158 52572 58164 52584
rect 58216 52572 58222 52624
rect 58250 52544 58256 52556
rect 42444 52516 58256 52544
rect 11882 52436 11888 52488
rect 11940 52476 11946 52488
rect 41785 52479 41843 52485
rect 41785 52476 41797 52479
rect 11940 52448 41797 52476
rect 11940 52436 11946 52448
rect 41785 52445 41797 52448
rect 41831 52476 41843 52479
rect 42153 52479 42211 52485
rect 42153 52476 42165 52479
rect 41831 52448 42165 52476
rect 41831 52445 41843 52448
rect 41785 52439 41843 52445
rect 42153 52445 42165 52448
rect 42199 52445 42211 52479
rect 42153 52439 42211 52445
rect 42334 52436 42340 52488
rect 42392 52436 42398 52488
rect 42444 52485 42472 52516
rect 58250 52504 58256 52516
rect 58308 52504 58314 52556
rect 42429 52479 42487 52485
rect 42429 52445 42441 52479
rect 42475 52445 42487 52479
rect 42429 52439 42487 52445
rect 42518 52436 42524 52488
rect 42576 52436 42582 52488
rect 47854 52436 47860 52488
rect 47912 52436 47918 52488
rect 48041 52479 48099 52485
rect 48041 52445 48053 52479
rect 48087 52476 48099 52479
rect 48130 52476 48136 52488
rect 48087 52448 48136 52476
rect 48087 52445 48099 52448
rect 48041 52439 48099 52445
rect 48130 52436 48136 52448
rect 48188 52436 48194 52488
rect 48409 52479 48467 52485
rect 48409 52445 48421 52479
rect 48455 52445 48467 52479
rect 48409 52439 48467 52445
rect 934 52368 940 52420
rect 992 52408 998 52420
rect 1673 52411 1731 52417
rect 1673 52408 1685 52411
rect 992 52380 1685 52408
rect 992 52368 998 52380
rect 1673 52377 1685 52380
rect 1719 52377 1731 52411
rect 1673 52371 1731 52377
rect 2038 52368 2044 52420
rect 2096 52368 2102 52420
rect 48424 52408 48452 52439
rect 48498 52436 48504 52488
rect 48556 52436 48562 52488
rect 57514 52476 57520 52488
rect 48608 52448 57520 52476
rect 48608 52408 48636 52448
rect 57514 52436 57520 52448
rect 57572 52436 57578 52488
rect 57885 52479 57943 52485
rect 57885 52445 57897 52479
rect 57931 52476 57943 52479
rect 58986 52476 58992 52488
rect 57931 52448 58992 52476
rect 57931 52445 57943 52448
rect 57885 52439 57943 52445
rect 58986 52436 58992 52448
rect 59044 52436 59050 52488
rect 48424 52380 48636 52408
rect 58158 52368 58164 52420
rect 58216 52368 58222 52420
rect 42702 52300 42708 52352
rect 42760 52300 42766 52352
rect 1104 52250 58880 52272
rect 1104 52198 19574 52250
rect 19626 52198 19638 52250
rect 19690 52198 19702 52250
rect 19754 52198 19766 52250
rect 19818 52198 19830 52250
rect 19882 52198 50294 52250
rect 50346 52198 50358 52250
rect 50410 52198 50422 52250
rect 50474 52198 50486 52250
rect 50538 52198 50550 52250
rect 50602 52198 58880 52250
rect 1104 52176 58880 52198
rect 57333 52071 57391 52077
rect 57333 52037 57345 52071
rect 57379 52068 57391 52071
rect 58986 52068 58992 52080
rect 57379 52040 58992 52068
rect 57379 52037 57391 52040
rect 57333 52031 57391 52037
rect 58986 52028 58992 52040
rect 59044 52028 59050 52080
rect 1026 51960 1032 52012
rect 1084 52000 1090 52012
rect 1581 52003 1639 52009
rect 1581 52000 1593 52003
rect 1084 51972 1593 52000
rect 1084 51960 1090 51972
rect 1581 51969 1593 51972
rect 1627 51969 1639 52003
rect 48225 52003 48283 52009
rect 48225 52000 48237 52003
rect 1581 51963 1639 51969
rect 26206 51972 48237 52000
rect 2038 51892 2044 51944
rect 2096 51932 2102 51944
rect 26206 51932 26234 51972
rect 48225 51969 48237 51972
rect 48271 51969 48283 52003
rect 48225 51963 48283 51969
rect 48409 52003 48467 52009
rect 48409 51969 48421 52003
rect 48455 51969 48467 52003
rect 48409 51963 48467 51969
rect 48777 52003 48835 52009
rect 48777 51969 48789 52003
rect 48823 52000 48835 52003
rect 53558 52000 53564 52012
rect 48823 51972 53564 52000
rect 48823 51969 48835 51972
rect 48777 51963 48835 51969
rect 2096 51904 26234 51932
rect 2096 51892 2102 51904
rect 47762 51892 47768 51944
rect 47820 51892 47826 51944
rect 48130 51892 48136 51944
rect 48188 51932 48194 51944
rect 48424 51932 48452 51963
rect 53558 51960 53564 51972
rect 53616 51960 53622 52012
rect 58069 52003 58127 52009
rect 58069 51969 58081 52003
rect 58115 52000 58127 52003
rect 58802 52000 58808 52012
rect 58115 51972 58808 52000
rect 58115 51969 58127 51972
rect 58069 51963 58127 51969
rect 58802 51960 58808 51972
rect 58860 51960 58866 52012
rect 48188 51904 48452 51932
rect 48188 51892 48194 51904
rect 48498 51892 48504 51944
rect 48556 51932 48562 51944
rect 48685 51935 48743 51941
rect 48685 51932 48697 51935
rect 48556 51904 48697 51932
rect 48556 51892 48562 51904
rect 48685 51901 48697 51904
rect 48731 51901 48743 51935
rect 48685 51895 48743 51901
rect 37274 51824 37280 51876
rect 37332 51864 37338 51876
rect 57517 51867 57575 51873
rect 57517 51864 57529 51867
rect 37332 51836 57529 51864
rect 37332 51824 37338 51836
rect 57517 51833 57529 51836
rect 57563 51833 57575 51867
rect 57517 51827 57575 51833
rect 1765 51799 1823 51805
rect 1765 51765 1777 51799
rect 1811 51796 1823 51799
rect 46842 51796 46848 51808
rect 1811 51768 46848 51796
rect 1811 51765 1823 51768
rect 1765 51759 1823 51765
rect 46842 51756 46848 51768
rect 46900 51756 46906 51808
rect 57974 51756 57980 51808
rect 58032 51796 58038 51808
rect 58253 51799 58311 51805
rect 58253 51796 58265 51799
rect 58032 51768 58265 51796
rect 58032 51756 58038 51768
rect 58253 51765 58265 51768
rect 58299 51765 58311 51799
rect 58253 51759 58311 51765
rect 1104 51706 58880 51728
rect 1104 51654 4214 51706
rect 4266 51654 4278 51706
rect 4330 51654 4342 51706
rect 4394 51654 4406 51706
rect 4458 51654 4470 51706
rect 4522 51654 34934 51706
rect 34986 51654 34998 51706
rect 35050 51654 35062 51706
rect 35114 51654 35126 51706
rect 35178 51654 35190 51706
rect 35242 51654 58880 51706
rect 1104 51632 58880 51654
rect 2682 51552 2688 51604
rect 2740 51592 2746 51604
rect 2740 51564 49280 51592
rect 2740 51552 2746 51564
rect 47397 51527 47455 51533
rect 47397 51493 47409 51527
rect 47443 51524 47455 51527
rect 47946 51524 47952 51536
rect 47443 51496 47952 51524
rect 47443 51493 47455 51496
rect 47397 51487 47455 51493
rect 47946 51484 47952 51496
rect 48004 51484 48010 51536
rect 48130 51484 48136 51536
rect 48188 51524 48194 51536
rect 48188 51496 49096 51524
rect 48188 51484 48194 51496
rect 48590 51456 48596 51468
rect 48424 51428 48596 51456
rect 36906 51348 36912 51400
rect 36964 51348 36970 51400
rect 37090 51397 37096 51400
rect 37057 51391 37096 51397
rect 37057 51357 37069 51391
rect 37057 51351 37096 51357
rect 37090 51348 37096 51351
rect 37148 51348 37154 51400
rect 37274 51348 37280 51400
rect 37332 51348 37338 51400
rect 37415 51391 37473 51397
rect 37415 51357 37427 51391
rect 37461 51388 37473 51391
rect 42518 51388 42524 51400
rect 37461 51360 42524 51388
rect 37461 51357 37473 51360
rect 37415 51351 37473 51357
rect 42518 51348 42524 51360
rect 42576 51348 42582 51400
rect 46842 51348 46848 51400
rect 46900 51348 46906 51400
rect 47265 51391 47323 51397
rect 47265 51357 47277 51391
rect 47311 51388 47323 51391
rect 48222 51388 48228 51400
rect 47311 51360 48228 51388
rect 47311 51357 47323 51360
rect 47265 51351 47323 51357
rect 48222 51348 48228 51360
rect 48280 51348 48286 51400
rect 48424 51397 48452 51428
rect 48590 51416 48596 51428
rect 48648 51416 48654 51468
rect 48409 51391 48467 51397
rect 48409 51357 48421 51391
rect 48455 51357 48467 51391
rect 48409 51351 48467 51357
rect 48685 51391 48743 51397
rect 48685 51357 48697 51391
rect 48731 51357 48743 51391
rect 48685 51351 48743 51357
rect 48777 51391 48835 51397
rect 48777 51357 48789 51391
rect 48823 51388 48835 51391
rect 48866 51388 48872 51400
rect 48823 51360 48872 51388
rect 48823 51357 48835 51360
rect 48777 51351 48835 51357
rect 934 51280 940 51332
rect 992 51320 998 51332
rect 1673 51323 1731 51329
rect 1673 51320 1685 51323
rect 992 51292 1685 51320
rect 992 51280 998 51292
rect 1673 51289 1685 51292
rect 1719 51289 1731 51323
rect 1673 51283 1731 51289
rect 2038 51280 2044 51332
rect 2096 51280 2102 51332
rect 37182 51280 37188 51332
rect 37240 51280 37246 51332
rect 47026 51280 47032 51332
rect 47084 51280 47090 51332
rect 47121 51323 47179 51329
rect 47121 51289 47133 51323
rect 47167 51289 47179 51323
rect 47121 51283 47179 51289
rect 37550 51212 37556 51264
rect 37608 51212 37614 51264
rect 47136 51252 47164 51283
rect 47486 51280 47492 51332
rect 47544 51320 47550 51332
rect 47949 51323 48007 51329
rect 47949 51320 47961 51323
rect 47544 51292 47961 51320
rect 47544 51280 47550 51292
rect 47949 51289 47961 51292
rect 47995 51289 48007 51323
rect 48700 51320 48728 51351
rect 48866 51348 48872 51360
rect 48924 51348 48930 51400
rect 49068 51397 49096 51496
rect 49252 51397 49280 51564
rect 49053 51391 49111 51397
rect 49053 51357 49065 51391
rect 49099 51357 49111 51391
rect 49053 51351 49111 51357
rect 49237 51391 49295 51397
rect 49237 51357 49249 51391
rect 49283 51357 49295 51391
rect 49237 51351 49295 51357
rect 57333 51391 57391 51397
rect 57333 51357 57345 51391
rect 57379 51388 57391 51391
rect 58986 51388 58992 51400
rect 57379 51360 58992 51388
rect 57379 51357 57391 51360
rect 57333 51351 57391 51357
rect 58986 51348 58992 51360
rect 59044 51348 59050 51400
rect 52638 51320 52644 51332
rect 48700 51292 52644 51320
rect 47949 51283 48007 51289
rect 52638 51280 52644 51292
rect 52696 51280 52702 51332
rect 58161 51323 58219 51329
rect 58161 51289 58173 51323
rect 58207 51320 58219 51323
rect 58894 51320 58900 51332
rect 58207 51292 58900 51320
rect 58207 51289 58219 51292
rect 58161 51283 58219 51289
rect 58894 51280 58900 51292
rect 58952 51280 58958 51332
rect 53834 51252 53840 51264
rect 47136 51224 53840 51252
rect 53834 51212 53840 51224
rect 53892 51212 53898 51264
rect 57514 51212 57520 51264
rect 57572 51212 57578 51264
rect 58253 51255 58311 51261
rect 58253 51221 58265 51255
rect 58299 51252 58311 51255
rect 58710 51252 58716 51264
rect 58299 51224 58716 51252
rect 58299 51221 58311 51224
rect 58253 51215 58311 51221
rect 58710 51212 58716 51224
rect 58768 51212 58774 51264
rect 1104 51162 58880 51184
rect 1104 51110 19574 51162
rect 19626 51110 19638 51162
rect 19690 51110 19702 51162
rect 19754 51110 19766 51162
rect 19818 51110 19830 51162
rect 19882 51110 50294 51162
rect 50346 51110 50358 51162
rect 50410 51110 50422 51162
rect 50474 51110 50486 51162
rect 50538 51110 50550 51162
rect 50602 51110 58880 51162
rect 1104 51088 58880 51110
rect 55214 51048 55220 51060
rect 48608 51020 55220 51048
rect 47026 50940 47032 50992
rect 47084 50980 47090 50992
rect 48130 50980 48136 50992
rect 47084 50952 48136 50980
rect 47084 50940 47090 50952
rect 48130 50940 48136 50952
rect 48188 50980 48194 50992
rect 48188 50952 48268 50980
rect 48188 50940 48194 50952
rect 1026 50872 1032 50924
rect 1084 50912 1090 50924
rect 48240 50921 48268 50952
rect 48608 50921 48636 51020
rect 55214 51008 55220 51020
rect 55272 51008 55278 51060
rect 48682 50940 48688 50992
rect 48740 50980 48746 50992
rect 49697 50983 49755 50989
rect 49697 50980 49709 50983
rect 48740 50952 49709 50980
rect 48740 50940 48746 50952
rect 49697 50949 49709 50952
rect 49743 50949 49755 50983
rect 49697 50943 49755 50949
rect 49789 50983 49847 50989
rect 49789 50949 49801 50983
rect 49835 50980 49847 50983
rect 54110 50980 54116 50992
rect 49835 50952 54116 50980
rect 49835 50949 49847 50952
rect 49789 50943 49847 50949
rect 54110 50940 54116 50952
rect 54168 50940 54174 50992
rect 1673 50915 1731 50921
rect 1673 50912 1685 50915
rect 1084 50884 1685 50912
rect 1084 50872 1090 50884
rect 1673 50881 1685 50884
rect 1719 50881 1731 50915
rect 48041 50915 48099 50921
rect 48041 50912 48053 50915
rect 1673 50875 1731 50881
rect 22066 50884 48053 50912
rect 2038 50804 2044 50856
rect 2096 50844 2102 50856
rect 22066 50844 22094 50884
rect 48041 50881 48053 50884
rect 48087 50881 48099 50915
rect 48041 50875 48099 50881
rect 48225 50915 48283 50921
rect 48225 50881 48237 50915
rect 48271 50881 48283 50915
rect 48225 50875 48283 50881
rect 48593 50915 48651 50921
rect 48593 50881 48605 50915
rect 48639 50881 48651 50915
rect 48593 50875 48651 50881
rect 48866 50872 48872 50924
rect 48924 50912 48930 50924
rect 49421 50915 49479 50921
rect 49421 50912 49433 50915
rect 48924 50884 49433 50912
rect 48924 50872 48930 50884
rect 49421 50881 49433 50884
rect 49467 50881 49479 50915
rect 49421 50875 49479 50881
rect 49514 50915 49572 50921
rect 49514 50881 49526 50915
rect 49560 50881 49572 50915
rect 49886 50915 49944 50921
rect 49886 50912 49898 50915
rect 49514 50875 49572 50881
rect 49620 50884 49898 50912
rect 2096 50816 22094 50844
rect 2096 50804 2102 50816
rect 47302 50804 47308 50856
rect 47360 50844 47366 50856
rect 47581 50847 47639 50853
rect 47581 50844 47593 50847
rect 47360 50816 47593 50844
rect 47360 50804 47366 50816
rect 47581 50813 47593 50816
rect 47627 50813 47639 50847
rect 47581 50807 47639 50813
rect 48498 50804 48504 50856
rect 48556 50804 48562 50856
rect 49528 50844 49556 50875
rect 49068 50816 49556 50844
rect 1949 50711 2007 50717
rect 1949 50677 1961 50711
rect 1995 50708 2007 50711
rect 2406 50708 2412 50720
rect 1995 50680 2412 50708
rect 1995 50677 2007 50680
rect 1949 50671 2007 50677
rect 2406 50668 2412 50680
rect 2464 50668 2470 50720
rect 2590 50668 2596 50720
rect 2648 50708 2654 50720
rect 49068 50717 49096 50816
rect 49234 50736 49240 50788
rect 49292 50776 49298 50788
rect 49620 50776 49648 50884
rect 49886 50881 49898 50884
rect 49932 50881 49944 50915
rect 49886 50875 49944 50881
rect 58161 50915 58219 50921
rect 58161 50881 58173 50915
rect 58207 50912 58219 50915
rect 58250 50912 58256 50924
rect 58207 50884 58256 50912
rect 58207 50881 58219 50884
rect 58161 50875 58219 50881
rect 58250 50872 58256 50884
rect 58308 50872 58314 50924
rect 55858 50804 55864 50856
rect 55916 50844 55922 50856
rect 58066 50844 58072 50856
rect 55916 50816 58072 50844
rect 55916 50804 55922 50816
rect 58066 50804 58072 50816
rect 58124 50804 58130 50856
rect 49292 50748 49648 50776
rect 49292 50736 49298 50748
rect 49053 50711 49111 50717
rect 49053 50708 49065 50711
rect 2648 50680 49065 50708
rect 2648 50668 2654 50680
rect 49053 50677 49065 50680
rect 49099 50677 49111 50711
rect 49053 50671 49111 50677
rect 49142 50668 49148 50720
rect 49200 50708 49206 50720
rect 50065 50711 50123 50717
rect 50065 50708 50077 50711
rect 49200 50680 50077 50708
rect 49200 50668 49206 50680
rect 50065 50677 50077 50680
rect 50111 50677 50123 50711
rect 50065 50671 50123 50677
rect 58066 50668 58072 50720
rect 58124 50708 58130 50720
rect 58253 50711 58311 50717
rect 58253 50708 58265 50711
rect 58124 50680 58265 50708
rect 58124 50668 58130 50680
rect 58253 50677 58265 50680
rect 58299 50677 58311 50711
rect 58253 50671 58311 50677
rect 1104 50618 58880 50640
rect 1104 50566 4214 50618
rect 4266 50566 4278 50618
rect 4330 50566 4342 50618
rect 4394 50566 4406 50618
rect 4458 50566 4470 50618
rect 4522 50566 34934 50618
rect 34986 50566 34998 50618
rect 35050 50566 35062 50618
rect 35114 50566 35126 50618
rect 35178 50566 35190 50618
rect 35242 50566 58880 50618
rect 1104 50544 58880 50566
rect 48498 50464 48504 50516
rect 48556 50504 48562 50516
rect 49418 50504 49424 50516
rect 48556 50476 49424 50504
rect 48556 50464 48562 50476
rect 49418 50464 49424 50476
rect 49476 50464 49482 50516
rect 48590 50396 48596 50448
rect 48648 50436 48654 50448
rect 49234 50436 49240 50448
rect 48648 50408 49240 50436
rect 48648 50396 48654 50408
rect 49234 50396 49240 50408
rect 49292 50396 49298 50448
rect 56042 50436 56048 50448
rect 49344 50408 56048 50436
rect 49053 50371 49111 50377
rect 49053 50337 49065 50371
rect 49099 50368 49111 50371
rect 49142 50368 49148 50380
rect 49099 50340 49148 50368
rect 49099 50337 49111 50340
rect 49053 50331 49111 50337
rect 49142 50328 49148 50340
rect 49200 50328 49206 50380
rect 49344 50309 49372 50408
rect 56042 50396 56048 50408
rect 56100 50396 56106 50448
rect 49418 50328 49424 50380
rect 49476 50328 49482 50380
rect 58342 50328 58348 50380
rect 58400 50368 58406 50380
rect 59078 50368 59084 50380
rect 58400 50340 59084 50368
rect 58400 50328 58406 50340
rect 59078 50328 59084 50340
rect 59136 50328 59142 50380
rect 48961 50303 49019 50309
rect 48961 50269 48973 50303
rect 49007 50269 49019 50303
rect 48961 50263 49019 50269
rect 49329 50303 49387 50309
rect 49329 50269 49341 50303
rect 49375 50269 49387 50303
rect 49329 50263 49387 50269
rect 934 50192 940 50244
rect 992 50232 998 50244
rect 1673 50235 1731 50241
rect 1673 50232 1685 50235
rect 992 50204 1685 50232
rect 992 50192 998 50204
rect 1673 50201 1685 50204
rect 1719 50201 1731 50235
rect 1673 50195 1731 50201
rect 48317 50235 48375 50241
rect 48317 50201 48329 50235
rect 48363 50232 48375 50235
rect 48774 50232 48780 50244
rect 48363 50204 48780 50232
rect 48363 50201 48375 50204
rect 48317 50195 48375 50201
rect 48774 50192 48780 50204
rect 48832 50192 48838 50244
rect 48976 50232 49004 50263
rect 49602 50232 49608 50244
rect 48976 50204 49608 50232
rect 49602 50192 49608 50204
rect 49660 50192 49666 50244
rect 58158 50192 58164 50244
rect 58216 50192 58222 50244
rect 1949 50167 2007 50173
rect 1949 50133 1961 50167
rect 1995 50164 2007 50167
rect 43070 50164 43076 50176
rect 1995 50136 43076 50164
rect 1995 50133 2007 50136
rect 1949 50127 2007 50133
rect 43070 50124 43076 50136
rect 43128 50124 43134 50176
rect 56134 50124 56140 50176
rect 56192 50164 56198 50176
rect 58253 50167 58311 50173
rect 58253 50164 58265 50167
rect 56192 50136 58265 50164
rect 56192 50124 56198 50136
rect 58253 50133 58265 50136
rect 58299 50133 58311 50167
rect 58253 50127 58311 50133
rect 1104 50074 58880 50096
rect 1104 50022 19574 50074
rect 19626 50022 19638 50074
rect 19690 50022 19702 50074
rect 19754 50022 19766 50074
rect 19818 50022 19830 50074
rect 19882 50022 50294 50074
rect 50346 50022 50358 50074
rect 50410 50022 50422 50074
rect 50474 50022 50486 50074
rect 50538 50022 50550 50074
rect 50602 50022 58880 50074
rect 1104 50000 58880 50022
rect 47026 49892 47032 49904
rect 43272 49864 47032 49892
rect 43272 49836 43300 49864
rect 47026 49852 47032 49864
rect 47084 49852 47090 49904
rect 1026 49784 1032 49836
rect 1084 49824 1090 49836
rect 1673 49827 1731 49833
rect 1673 49824 1685 49827
rect 1084 49796 1685 49824
rect 1084 49784 1090 49796
rect 1673 49793 1685 49796
rect 1719 49793 1731 49827
rect 1673 49787 1731 49793
rect 42518 49784 42524 49836
rect 42576 49824 42582 49836
rect 42576 49796 42748 49824
rect 42576 49784 42582 49796
rect 1854 49716 1860 49768
rect 1912 49756 1918 49768
rect 1949 49759 2007 49765
rect 1949 49756 1961 49759
rect 1912 49728 1961 49756
rect 1912 49716 1918 49728
rect 1949 49725 1961 49728
rect 1995 49725 2007 49759
rect 1949 49719 2007 49725
rect 42610 49716 42616 49768
rect 42668 49716 42674 49768
rect 42720 49756 42748 49796
rect 43070 49784 43076 49836
rect 43128 49784 43134 49836
rect 43254 49784 43260 49836
rect 43312 49784 43318 49836
rect 43625 49827 43683 49833
rect 43625 49793 43637 49827
rect 43671 49824 43683 49827
rect 56594 49824 56600 49836
rect 43671 49796 56600 49824
rect 43671 49793 43683 49796
rect 43625 49787 43683 49793
rect 56594 49784 56600 49796
rect 56652 49784 56658 49836
rect 58161 49827 58219 49833
rect 58161 49793 58173 49827
rect 58207 49824 58219 49827
rect 58986 49824 58992 49836
rect 58207 49796 58992 49824
rect 58207 49793 58219 49796
rect 58161 49787 58219 49793
rect 58986 49784 58992 49796
rect 59044 49784 59050 49836
rect 43533 49759 43591 49765
rect 43533 49756 43545 49759
rect 42720 49728 43545 49756
rect 43533 49725 43545 49728
rect 43579 49756 43591 49759
rect 48498 49756 48504 49768
rect 43579 49728 48504 49756
rect 43579 49725 43591 49728
rect 43533 49719 43591 49725
rect 48498 49716 48504 49728
rect 48556 49716 48562 49768
rect 58345 49759 58403 49765
rect 58345 49725 58357 49759
rect 58391 49756 58403 49759
rect 58618 49756 58624 49768
rect 58391 49728 58624 49756
rect 58391 49725 58403 49728
rect 58345 49719 58403 49725
rect 58618 49716 58624 49728
rect 58676 49716 58682 49768
rect 1104 49530 58880 49552
rect 1104 49478 4214 49530
rect 4266 49478 4278 49530
rect 4330 49478 4342 49530
rect 4394 49478 4406 49530
rect 4458 49478 4470 49530
rect 4522 49478 34934 49530
rect 34986 49478 34998 49530
rect 35050 49478 35062 49530
rect 35114 49478 35126 49530
rect 35178 49478 35190 49530
rect 35242 49478 58880 49530
rect 1104 49456 58880 49478
rect 30834 49280 30840 49292
rect 30208 49252 30840 49280
rect 30208 49221 30236 49252
rect 30834 49240 30840 49252
rect 30892 49240 30898 49292
rect 30193 49215 30251 49221
rect 30193 49181 30205 49215
rect 30239 49181 30251 49215
rect 30193 49175 30251 49181
rect 30466 49172 30472 49224
rect 30524 49172 30530 49224
rect 30561 49215 30619 49221
rect 30561 49181 30573 49215
rect 30607 49181 30619 49215
rect 30561 49175 30619 49181
rect 934 49104 940 49156
rect 992 49144 998 49156
rect 1673 49147 1731 49153
rect 1673 49144 1685 49147
rect 992 49116 1685 49144
rect 992 49104 998 49116
rect 1673 49113 1685 49116
rect 1719 49113 1731 49147
rect 1673 49107 1731 49113
rect 30374 49104 30380 49156
rect 30432 49104 30438 49156
rect 30576 49144 30604 49175
rect 31386 49144 31392 49156
rect 30576 49116 31392 49144
rect 1946 49036 1952 49088
rect 2004 49036 2010 49088
rect 28350 49036 28356 49088
rect 28408 49076 28414 49088
rect 30576 49076 30604 49116
rect 31386 49104 31392 49116
rect 31444 49104 31450 49156
rect 57974 49104 57980 49156
rect 58032 49104 58038 49156
rect 28408 49048 30604 49076
rect 30745 49079 30803 49085
rect 28408 49036 28414 49048
rect 30745 49045 30757 49079
rect 30791 49076 30803 49079
rect 30926 49076 30932 49088
rect 30791 49048 30932 49076
rect 30791 49045 30803 49048
rect 30745 49039 30803 49045
rect 30926 49036 30932 49048
rect 30984 49036 30990 49088
rect 58066 49036 58072 49088
rect 58124 49036 58130 49088
rect 1104 48986 58880 49008
rect 1104 48934 19574 48986
rect 19626 48934 19638 48986
rect 19690 48934 19702 48986
rect 19754 48934 19766 48986
rect 19818 48934 19830 48986
rect 19882 48934 50294 48986
rect 50346 48934 50358 48986
rect 50410 48934 50422 48986
rect 50474 48934 50486 48986
rect 50538 48934 50550 48986
rect 50602 48934 58880 48986
rect 1104 48912 58880 48934
rect 10229 48807 10287 48813
rect 10229 48773 10241 48807
rect 10275 48804 10287 48807
rect 57882 48804 57888 48816
rect 10275 48776 10456 48804
rect 10275 48773 10287 48776
rect 10229 48767 10287 48773
rect 1026 48696 1032 48748
rect 1084 48736 1090 48748
rect 1673 48739 1731 48745
rect 1673 48736 1685 48739
rect 1084 48708 1685 48736
rect 1084 48696 1090 48708
rect 1673 48705 1685 48708
rect 1719 48705 1731 48739
rect 1673 48699 1731 48705
rect 9950 48696 9956 48748
rect 10008 48696 10014 48748
rect 10134 48696 10140 48748
rect 10192 48696 10198 48748
rect 10326 48739 10384 48745
rect 10326 48705 10338 48739
rect 10372 48705 10384 48739
rect 10326 48699 10384 48705
rect 2222 48628 2228 48680
rect 2280 48668 2286 48680
rect 10336 48668 10364 48699
rect 2280 48640 10364 48668
rect 2280 48628 2286 48640
rect 1765 48535 1823 48541
rect 1765 48501 1777 48535
rect 1811 48532 1823 48535
rect 10428 48532 10456 48776
rect 31036 48776 57888 48804
rect 31036 48745 31064 48776
rect 57882 48764 57888 48776
rect 57940 48764 57946 48816
rect 30745 48739 30803 48745
rect 30745 48705 30757 48739
rect 30791 48705 30803 48739
rect 30745 48699 30803 48705
rect 31021 48739 31079 48745
rect 31021 48705 31033 48739
rect 31067 48705 31079 48739
rect 31021 48699 31079 48705
rect 31113 48739 31171 48745
rect 31113 48705 31125 48739
rect 31159 48705 31171 48739
rect 31113 48699 31171 48705
rect 30760 48600 30788 48699
rect 31128 48668 31156 48699
rect 31386 48696 31392 48748
rect 31444 48696 31450 48748
rect 31570 48696 31576 48748
rect 31628 48696 31634 48748
rect 58069 48739 58127 48745
rect 58069 48705 58081 48739
rect 58115 48736 58127 48739
rect 58802 48736 58808 48748
rect 58115 48708 58808 48736
rect 58115 48705 58127 48708
rect 58069 48699 58127 48705
rect 58802 48696 58808 48708
rect 58860 48696 58866 48748
rect 33042 48668 33048 48680
rect 31128 48640 33048 48668
rect 33042 48628 33048 48640
rect 33100 48628 33106 48680
rect 31478 48600 31484 48612
rect 30760 48572 31484 48600
rect 31478 48560 31484 48572
rect 31536 48560 31542 48612
rect 1811 48504 10456 48532
rect 1811 48501 1823 48504
rect 1765 48495 1823 48501
rect 10502 48492 10508 48544
rect 10560 48492 10566 48544
rect 30377 48535 30435 48541
rect 30377 48501 30389 48535
rect 30423 48532 30435 48535
rect 30650 48532 30656 48544
rect 30423 48504 30656 48532
rect 30423 48501 30435 48504
rect 30377 48495 30435 48501
rect 30650 48492 30656 48504
rect 30708 48492 30714 48544
rect 56042 48492 56048 48544
rect 56100 48532 56106 48544
rect 58253 48535 58311 48541
rect 58253 48532 58265 48535
rect 56100 48504 58265 48532
rect 56100 48492 56106 48504
rect 58253 48501 58265 48504
rect 58299 48501 58311 48535
rect 58253 48495 58311 48501
rect 1104 48442 58880 48464
rect 1104 48390 4214 48442
rect 4266 48390 4278 48442
rect 4330 48390 4342 48442
rect 4394 48390 4406 48442
rect 4458 48390 4470 48442
rect 4522 48390 34934 48442
rect 34986 48390 34998 48442
rect 35050 48390 35062 48442
rect 35114 48390 35126 48442
rect 35178 48390 35190 48442
rect 35242 48390 58880 48442
rect 1104 48368 58880 48390
rect 35710 48288 35716 48340
rect 35768 48328 35774 48340
rect 35894 48328 35900 48340
rect 35768 48300 35900 48328
rect 35768 48288 35774 48300
rect 35894 48288 35900 48300
rect 35952 48288 35958 48340
rect 57882 48288 57888 48340
rect 57940 48328 57946 48340
rect 58986 48328 58992 48340
rect 57940 48300 58992 48328
rect 57940 48288 57946 48300
rect 58986 48288 58992 48300
rect 59044 48288 59050 48340
rect 31386 48220 31392 48272
rect 31444 48260 31450 48272
rect 58158 48260 58164 48272
rect 31444 48232 58164 48260
rect 31444 48220 31450 48232
rect 58158 48220 58164 48232
rect 58216 48220 58222 48272
rect 10502 48152 10508 48204
rect 10560 48192 10566 48204
rect 40954 48192 40960 48204
rect 10560 48164 40960 48192
rect 10560 48152 10566 48164
rect 40954 48152 40960 48164
rect 41012 48152 41018 48204
rect 30374 48084 30380 48136
rect 30432 48124 30438 48136
rect 31202 48133 31208 48136
rect 31021 48127 31079 48133
rect 31021 48124 31033 48127
rect 30432 48096 31033 48124
rect 30432 48084 30438 48096
rect 31021 48093 31033 48096
rect 31067 48093 31079 48127
rect 31021 48087 31079 48093
rect 31169 48127 31208 48133
rect 31169 48093 31181 48127
rect 31169 48087 31208 48093
rect 31202 48084 31208 48087
rect 31260 48084 31266 48136
rect 31386 48084 31392 48136
rect 31444 48084 31450 48136
rect 31478 48084 31484 48136
rect 31536 48133 31542 48136
rect 31536 48124 31544 48133
rect 31536 48096 31581 48124
rect 31536 48087 31544 48096
rect 31536 48084 31542 48087
rect 34882 48084 34888 48136
rect 34940 48084 34946 48136
rect 35161 48127 35219 48133
rect 35161 48124 35173 48127
rect 34992 48096 35173 48124
rect 934 48016 940 48068
rect 992 48056 998 48068
rect 1673 48059 1731 48065
rect 1673 48056 1685 48059
rect 992 48028 1685 48056
rect 992 48016 998 48028
rect 1673 48025 1685 48028
rect 1719 48025 1731 48059
rect 1673 48019 1731 48025
rect 31294 48016 31300 48068
rect 31352 48016 31358 48068
rect 34790 48016 34796 48068
rect 34848 48056 34854 48068
rect 34992 48056 35020 48096
rect 35161 48093 35173 48096
rect 35207 48093 35219 48127
rect 35161 48087 35219 48093
rect 35253 48127 35311 48133
rect 35253 48093 35265 48127
rect 35299 48124 35311 48127
rect 35894 48124 35900 48136
rect 35299 48096 35900 48124
rect 35299 48093 35311 48096
rect 35253 48087 35311 48093
rect 35894 48084 35900 48096
rect 35952 48124 35958 48136
rect 37182 48124 37188 48136
rect 35952 48096 37188 48124
rect 35952 48084 35958 48096
rect 37182 48084 37188 48096
rect 37240 48124 37246 48136
rect 41782 48124 41788 48136
rect 37240 48096 41788 48124
rect 37240 48084 37246 48096
rect 41782 48084 41788 48096
rect 41840 48084 41846 48136
rect 57149 48127 57207 48133
rect 57149 48093 57161 48127
rect 57195 48093 57207 48127
rect 57149 48087 57207 48093
rect 34848 48028 35020 48056
rect 35069 48059 35127 48065
rect 34848 48016 34854 48028
rect 35069 48025 35081 48059
rect 35115 48025 35127 48059
rect 41598 48056 41604 48068
rect 35069 48019 35127 48025
rect 35360 48028 41604 48056
rect 1765 47991 1823 47997
rect 1765 47957 1777 47991
rect 1811 47988 1823 47991
rect 30834 47988 30840 48000
rect 1811 47960 30840 47988
rect 1811 47957 1823 47960
rect 1765 47951 1823 47957
rect 30834 47948 30840 47960
rect 30892 47948 30898 48000
rect 31662 47948 31668 48000
rect 31720 47948 31726 48000
rect 35084 47988 35112 48019
rect 35360 47988 35388 48028
rect 35912 48000 35940 48028
rect 41598 48016 41604 48028
rect 41656 48016 41662 48068
rect 57164 48056 57192 48087
rect 57882 48084 57888 48136
rect 57940 48084 57946 48136
rect 58986 48124 58992 48136
rect 57992 48096 58992 48124
rect 57992 48056 58020 48096
rect 58986 48084 58992 48096
rect 59044 48084 59050 48136
rect 57164 48028 58020 48056
rect 58161 48059 58219 48065
rect 58161 48025 58173 48059
rect 58207 48056 58219 48059
rect 59078 48056 59084 48068
rect 58207 48028 59084 48056
rect 58207 48025 58219 48028
rect 58161 48019 58219 48025
rect 59078 48016 59084 48028
rect 59136 48016 59142 48068
rect 35084 47960 35388 47988
rect 35434 47948 35440 48000
rect 35492 47948 35498 48000
rect 35894 47948 35900 48000
rect 35952 47948 35958 48000
rect 57330 47948 57336 48000
rect 57388 47948 57394 48000
rect 1104 47898 58880 47920
rect 1104 47846 19574 47898
rect 19626 47846 19638 47898
rect 19690 47846 19702 47898
rect 19754 47846 19766 47898
rect 19818 47846 19830 47898
rect 19882 47846 50294 47898
rect 50346 47846 50358 47898
rect 50410 47846 50422 47898
rect 50474 47846 50486 47898
rect 50538 47846 50550 47898
rect 50602 47846 58880 47898
rect 1104 47824 58880 47846
rect 34882 47744 34888 47796
rect 34940 47784 34946 47796
rect 35342 47784 35348 47796
rect 34940 47756 35348 47784
rect 34940 47744 34946 47756
rect 35342 47744 35348 47756
rect 35400 47744 35406 47796
rect 35866 47756 45554 47784
rect 31113 47719 31171 47725
rect 31113 47685 31125 47719
rect 31159 47716 31171 47719
rect 35866 47716 35894 47756
rect 31159 47688 35894 47716
rect 31159 47685 31171 47688
rect 31113 47679 31171 47685
rect 40954 47676 40960 47728
rect 41012 47676 41018 47728
rect 41598 47676 41604 47728
rect 41656 47676 41662 47728
rect 41690 47676 41696 47728
rect 41748 47676 41754 47728
rect 45526 47716 45554 47756
rect 58434 47716 58440 47728
rect 45526 47688 58440 47716
rect 58434 47676 58440 47688
rect 58492 47676 58498 47728
rect 1026 47608 1032 47660
rect 1084 47648 1090 47660
rect 1581 47651 1639 47657
rect 1581 47648 1593 47651
rect 1084 47620 1593 47648
rect 1084 47608 1090 47620
rect 1581 47617 1593 47620
rect 1627 47617 1639 47651
rect 1581 47611 1639 47617
rect 30374 47608 30380 47660
rect 30432 47648 30438 47660
rect 30745 47651 30803 47657
rect 30745 47648 30757 47651
rect 30432 47620 30757 47648
rect 30432 47608 30438 47620
rect 30745 47617 30757 47620
rect 30791 47617 30803 47651
rect 30745 47611 30803 47617
rect 30834 47608 30840 47660
rect 30892 47608 30898 47660
rect 31018 47608 31024 47660
rect 31076 47608 31082 47660
rect 31251 47651 31309 47657
rect 31251 47617 31263 47651
rect 31297 47648 31309 47651
rect 31478 47648 31484 47660
rect 31297 47620 31484 47648
rect 31297 47617 31309 47620
rect 31251 47611 31309 47617
rect 31478 47608 31484 47620
rect 31536 47648 31542 47660
rect 32950 47648 32956 47660
rect 31536 47620 32956 47648
rect 31536 47608 31542 47620
rect 32950 47608 32956 47620
rect 33008 47608 33014 47660
rect 33042 47608 33048 47660
rect 33100 47648 33106 47660
rect 35434 47648 35440 47660
rect 33100 47620 35440 47648
rect 33100 47608 33106 47620
rect 35434 47608 35440 47620
rect 35492 47608 35498 47660
rect 40972 47648 41000 47676
rect 41325 47651 41383 47657
rect 41325 47648 41337 47651
rect 40972 47620 41337 47648
rect 41325 47617 41337 47620
rect 41371 47617 41383 47651
rect 41325 47611 41383 47617
rect 41473 47651 41531 47657
rect 41473 47617 41485 47651
rect 41519 47648 41531 47651
rect 41519 47617 41552 47648
rect 41473 47611 41552 47617
rect 41524 47580 41552 47611
rect 41782 47608 41788 47660
rect 41840 47657 41846 47660
rect 41840 47611 41848 47657
rect 57241 47651 57299 47657
rect 57241 47617 57253 47651
rect 57287 47617 57299 47651
rect 57241 47611 57299 47617
rect 58069 47651 58127 47657
rect 58069 47617 58081 47651
rect 58115 47648 58127 47651
rect 58894 47648 58900 47660
rect 58115 47620 58900 47648
rect 58115 47617 58127 47620
rect 58069 47611 58127 47617
rect 41840 47608 41846 47611
rect 43070 47580 43076 47592
rect 41524 47552 43076 47580
rect 43070 47540 43076 47552
rect 43128 47540 43134 47592
rect 57256 47580 57284 47611
rect 58894 47608 58900 47620
rect 58952 47608 58958 47660
rect 58986 47580 58992 47592
rect 57256 47552 58992 47580
rect 58986 47540 58992 47552
rect 59044 47540 59050 47592
rect 1765 47447 1823 47453
rect 1765 47413 1777 47447
rect 1811 47444 1823 47447
rect 14458 47444 14464 47456
rect 1811 47416 14464 47444
rect 1811 47413 1823 47416
rect 1765 47407 1823 47413
rect 14458 47404 14464 47416
rect 14516 47404 14522 47456
rect 31386 47404 31392 47456
rect 31444 47404 31450 47456
rect 41969 47447 42027 47453
rect 41969 47413 41981 47447
rect 42015 47444 42027 47447
rect 42150 47444 42156 47456
rect 42015 47416 42156 47444
rect 42015 47413 42027 47416
rect 41969 47407 42027 47413
rect 42150 47404 42156 47416
rect 42208 47404 42214 47456
rect 57422 47404 57428 47456
rect 57480 47404 57486 47456
rect 58253 47447 58311 47453
rect 58253 47413 58265 47447
rect 58299 47444 58311 47447
rect 58434 47444 58440 47456
rect 58299 47416 58440 47444
rect 58299 47413 58311 47416
rect 58253 47407 58311 47413
rect 58434 47404 58440 47416
rect 58492 47404 58498 47456
rect 1104 47354 58880 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 58880 47354
rect 1104 47280 58880 47302
rect 58253 47175 58311 47181
rect 58253 47141 58265 47175
rect 58299 47172 58311 47175
rect 58802 47172 58808 47184
rect 58299 47144 58808 47172
rect 58299 47141 58311 47144
rect 58253 47135 58311 47141
rect 58802 47132 58808 47144
rect 58860 47132 58866 47184
rect 30466 46996 30472 47048
rect 30524 47036 30530 47048
rect 31294 47036 31300 47048
rect 30524 47008 31300 47036
rect 30524 46996 30530 47008
rect 31294 46996 31300 47008
rect 31352 47036 31358 47048
rect 32674 47036 32680 47048
rect 31352 47008 32680 47036
rect 31352 46996 31358 47008
rect 32674 46996 32680 47008
rect 32732 47036 32738 47048
rect 35710 47036 35716 47048
rect 32732 47008 35716 47036
rect 32732 46996 32738 47008
rect 35710 46996 35716 47008
rect 35768 46996 35774 47048
rect 58069 47039 58127 47045
rect 58069 47005 58081 47039
rect 58115 47036 58127 47039
rect 58986 47036 58992 47048
rect 58115 47008 58992 47036
rect 58115 47005 58127 47008
rect 58069 46999 58127 47005
rect 58986 46996 58992 47008
rect 59044 46996 59050 47048
rect 934 46928 940 46980
rect 992 46968 998 46980
rect 1673 46971 1731 46977
rect 1673 46968 1685 46971
rect 992 46940 1685 46968
rect 992 46928 998 46940
rect 1673 46937 1685 46940
rect 1719 46937 1731 46971
rect 1673 46931 1731 46937
rect 1857 46971 1915 46977
rect 1857 46937 1869 46971
rect 1903 46968 1915 46971
rect 32306 46968 32312 46980
rect 1903 46940 32312 46968
rect 1903 46937 1915 46940
rect 1857 46931 1915 46937
rect 32306 46928 32312 46940
rect 32364 46928 32370 46980
rect 1104 46810 58880 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 50294 46810
rect 50346 46758 50358 46810
rect 50410 46758 50422 46810
rect 50474 46758 50486 46810
rect 50538 46758 50550 46810
rect 50602 46758 58880 46810
rect 1104 46736 58880 46758
rect 33137 46631 33195 46637
rect 33137 46628 33149 46631
rect 32324 46600 33149 46628
rect 32324 46572 32352 46600
rect 33137 46597 33149 46600
rect 33183 46597 33195 46631
rect 33137 46591 33195 46597
rect 1026 46520 1032 46572
rect 1084 46560 1090 46572
rect 1581 46563 1639 46569
rect 1581 46560 1593 46563
rect 1084 46532 1593 46560
rect 1084 46520 1090 46532
rect 1581 46529 1593 46532
rect 1627 46529 1639 46563
rect 1581 46523 1639 46529
rect 32306 46520 32312 46572
rect 32364 46520 32370 46572
rect 32493 46563 32551 46569
rect 32493 46529 32505 46563
rect 32539 46529 32551 46563
rect 32493 46523 32551 46529
rect 32585 46563 32643 46569
rect 32585 46529 32597 46563
rect 32631 46529 32643 46563
rect 32585 46523 32643 46529
rect 31018 46452 31024 46504
rect 31076 46492 31082 46504
rect 32508 46492 32536 46523
rect 31076 46464 32536 46492
rect 32600 46492 32628 46523
rect 32674 46520 32680 46572
rect 32732 46520 32738 46572
rect 58158 46520 58164 46572
rect 58216 46520 58222 46572
rect 37918 46492 37924 46504
rect 32600 46464 37924 46492
rect 31076 46452 31082 46464
rect 32508 46424 32536 46464
rect 37918 46452 37924 46464
rect 37976 46452 37982 46504
rect 50706 46452 50712 46504
rect 50764 46492 50770 46504
rect 58526 46492 58532 46504
rect 50764 46464 58532 46492
rect 50764 46452 50770 46464
rect 58526 46452 58532 46464
rect 58584 46452 58590 46504
rect 35526 46424 35532 46436
rect 32508 46396 35532 46424
rect 35526 46384 35532 46396
rect 35584 46384 35590 46436
rect 1765 46359 1823 46365
rect 1765 46325 1777 46359
rect 1811 46356 1823 46359
rect 26970 46356 26976 46368
rect 1811 46328 26976 46356
rect 1811 46325 1823 46328
rect 1765 46319 1823 46325
rect 26970 46316 26976 46328
rect 27028 46316 27034 46368
rect 32306 46316 32312 46368
rect 32364 46356 32370 46368
rect 32861 46359 32919 46365
rect 32861 46356 32873 46359
rect 32364 46328 32873 46356
rect 32364 46316 32370 46328
rect 32861 46325 32873 46328
rect 32907 46325 32919 46359
rect 32861 46319 32919 46325
rect 58250 46316 58256 46368
rect 58308 46316 58314 46368
rect 1104 46266 58880 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 58880 46266
rect 1104 46192 58880 46214
rect 36906 46112 36912 46164
rect 36964 46152 36970 46164
rect 37001 46155 37059 46161
rect 37001 46152 37013 46155
rect 36964 46124 37013 46152
rect 36964 46112 36970 46124
rect 37001 46121 37013 46124
rect 37047 46121 37059 46155
rect 37001 46115 37059 46121
rect 934 45908 940 45960
rect 992 45948 998 45960
rect 1581 45951 1639 45957
rect 1581 45948 1593 45951
rect 992 45920 1593 45948
rect 992 45908 998 45920
rect 1581 45917 1593 45920
rect 1627 45917 1639 45951
rect 1581 45911 1639 45917
rect 26970 45908 26976 45960
rect 27028 45948 27034 45960
rect 36449 45951 36507 45957
rect 36449 45948 36461 45951
rect 27028 45920 36461 45948
rect 27028 45908 27034 45920
rect 36449 45917 36461 45920
rect 36495 45917 36507 45951
rect 36449 45911 36507 45917
rect 36814 45908 36820 45960
rect 36872 45908 36878 45960
rect 57885 45951 57943 45957
rect 57885 45917 57897 45951
rect 57931 45948 57943 45951
rect 58986 45948 58992 45960
rect 57931 45920 58992 45948
rect 57931 45917 57943 45920
rect 57885 45911 57943 45917
rect 58986 45908 58992 45920
rect 59044 45908 59050 45960
rect 35526 45840 35532 45892
rect 35584 45880 35590 45892
rect 36633 45883 36691 45889
rect 36633 45880 36645 45883
rect 35584 45852 36645 45880
rect 35584 45840 35590 45852
rect 36633 45849 36645 45852
rect 36679 45849 36691 45883
rect 36633 45843 36691 45849
rect 36725 45883 36783 45889
rect 36725 45849 36737 45883
rect 36771 45880 36783 45883
rect 38286 45880 38292 45892
rect 36771 45852 38292 45880
rect 36771 45849 36783 45852
rect 36725 45843 36783 45849
rect 1762 45772 1768 45824
rect 1820 45772 1826 45824
rect 36648 45812 36676 45843
rect 38286 45840 38292 45852
rect 38344 45840 38350 45892
rect 58066 45840 58072 45892
rect 58124 45880 58130 45892
rect 58161 45883 58219 45889
rect 58161 45880 58173 45883
rect 58124 45852 58173 45880
rect 58124 45840 58130 45852
rect 58161 45849 58173 45852
rect 58207 45849 58219 45883
rect 58161 45843 58219 45849
rect 48682 45812 48688 45824
rect 36648 45784 48688 45812
rect 48682 45772 48688 45784
rect 48740 45772 48746 45824
rect 1104 45722 58880 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 50294 45722
rect 50346 45670 50358 45722
rect 50410 45670 50422 45722
rect 50474 45670 50486 45722
rect 50538 45670 50550 45722
rect 50602 45670 58880 45722
rect 1104 45648 58880 45670
rect 35526 45568 35532 45620
rect 35584 45568 35590 45620
rect 29730 45500 29736 45552
rect 29788 45540 29794 45552
rect 29788 45512 35480 45540
rect 29788 45500 29794 45512
rect 1026 45432 1032 45484
rect 1084 45472 1090 45484
rect 1581 45475 1639 45481
rect 1581 45472 1593 45475
rect 1084 45444 1593 45472
rect 1084 45432 1090 45444
rect 1581 45441 1593 45444
rect 1627 45441 1639 45475
rect 1581 45435 1639 45441
rect 32306 45432 32312 45484
rect 32364 45432 32370 45484
rect 32398 45432 32404 45484
rect 32456 45432 32462 45484
rect 32582 45432 32588 45484
rect 32640 45432 32646 45484
rect 32674 45432 32680 45484
rect 32732 45432 32738 45484
rect 32784 45481 32812 45512
rect 32774 45475 32832 45481
rect 32774 45441 32786 45475
rect 32820 45441 32832 45475
rect 32774 45435 32832 45441
rect 35345 45475 35403 45481
rect 35345 45441 35357 45475
rect 35391 45441 35403 45475
rect 35345 45435 35403 45441
rect 1762 45364 1768 45416
rect 1820 45404 1826 45416
rect 34977 45407 35035 45413
rect 34977 45404 34989 45407
rect 1820 45376 34989 45404
rect 1820 45364 1826 45376
rect 34977 45373 34989 45376
rect 35023 45404 35035 45407
rect 35360 45404 35388 45435
rect 35023 45376 35388 45404
rect 35452 45404 35480 45512
rect 35544 45481 35572 45568
rect 35618 45500 35624 45552
rect 35676 45500 35682 45552
rect 35894 45540 35900 45552
rect 35866 45500 35900 45540
rect 35952 45540 35958 45552
rect 36814 45540 36820 45552
rect 35952 45512 36820 45540
rect 35952 45500 35958 45512
rect 36814 45500 36820 45512
rect 36872 45500 36878 45552
rect 35529 45475 35587 45481
rect 35529 45441 35541 45475
rect 35575 45441 35587 45475
rect 35529 45435 35587 45441
rect 35710 45432 35716 45484
rect 35768 45432 35774 45484
rect 35866 45404 35894 45500
rect 58158 45432 58164 45484
rect 58216 45432 58222 45484
rect 58342 45432 58348 45484
rect 58400 45472 58406 45484
rect 58526 45472 58532 45484
rect 58400 45444 58532 45472
rect 58400 45432 58406 45444
rect 58526 45432 58532 45444
rect 58584 45432 58590 45484
rect 35452 45376 35894 45404
rect 35023 45373 35035 45376
rect 34977 45367 35035 45373
rect 32582 45296 32588 45348
rect 32640 45336 32646 45348
rect 42334 45336 42340 45348
rect 32640 45308 42340 45336
rect 32640 45296 32646 45308
rect 42334 45296 42340 45308
rect 42392 45296 42398 45348
rect 1765 45271 1823 45277
rect 1765 45237 1777 45271
rect 1811 45268 1823 45271
rect 7190 45268 7196 45280
rect 1811 45240 7196 45268
rect 1811 45237 1823 45240
rect 1765 45231 1823 45237
rect 7190 45228 7196 45240
rect 7248 45228 7254 45280
rect 32766 45228 32772 45280
rect 32824 45268 32830 45280
rect 32953 45271 33011 45277
rect 32953 45268 32965 45271
rect 32824 45240 32965 45268
rect 32824 45228 32830 45240
rect 32953 45237 32965 45240
rect 32999 45237 33011 45271
rect 32953 45231 33011 45237
rect 35897 45271 35955 45277
rect 35897 45237 35909 45271
rect 35943 45268 35955 45271
rect 36446 45268 36452 45280
rect 35943 45240 36452 45268
rect 35943 45237 35955 45240
rect 35897 45231 35955 45237
rect 36446 45228 36452 45240
rect 36504 45228 36510 45280
rect 58250 45228 58256 45280
rect 58308 45228 58314 45280
rect 1104 45178 58880 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 58880 45178
rect 1104 45104 58880 45126
rect 6730 45024 6736 45076
rect 6788 45064 6794 45076
rect 32398 45064 32404 45076
rect 6788 45036 32404 45064
rect 6788 45024 6794 45036
rect 32398 45024 32404 45036
rect 32456 45024 32462 45076
rect 58342 45064 58348 45076
rect 49160 45036 58348 45064
rect 39390 44956 39396 45008
rect 39448 44996 39454 45008
rect 39448 44968 45554 44996
rect 39448 44956 39454 44968
rect 934 44752 940 44804
rect 992 44792 998 44804
rect 1673 44795 1731 44801
rect 1673 44792 1685 44795
rect 992 44764 1685 44792
rect 992 44752 998 44764
rect 1673 44761 1685 44764
rect 1719 44761 1731 44795
rect 1673 44755 1731 44761
rect 1857 44795 1915 44801
rect 1857 44761 1869 44795
rect 1903 44792 1915 44795
rect 2130 44792 2136 44804
rect 1903 44764 2136 44792
rect 1903 44761 1915 44764
rect 1857 44755 1915 44761
rect 2130 44752 2136 44764
rect 2188 44752 2194 44804
rect 45526 44792 45554 44968
rect 49160 44937 49188 45036
rect 58342 45024 58348 45036
rect 58400 45024 58406 45076
rect 57330 44996 57336 45008
rect 49252 44968 57336 44996
rect 49145 44931 49203 44937
rect 49145 44897 49157 44931
rect 49191 44897 49203 44931
rect 49145 44891 49203 44897
rect 47210 44820 47216 44872
rect 47268 44860 47274 44872
rect 49053 44863 49111 44869
rect 49053 44860 49065 44863
rect 47268 44832 49065 44860
rect 47268 44820 47274 44832
rect 49053 44829 49065 44832
rect 49099 44829 49111 44863
rect 49053 44823 49111 44829
rect 49252 44792 49280 44968
rect 57330 44956 57336 44968
rect 57388 44956 57394 45008
rect 49326 44888 49332 44940
rect 49384 44888 49390 44940
rect 58894 44928 58900 44940
rect 57256 44900 58900 44928
rect 57256 44869 57284 44900
rect 58894 44888 58900 44900
rect 58952 44888 58958 44940
rect 49421 44863 49479 44869
rect 49421 44829 49433 44863
rect 49467 44829 49479 44863
rect 49421 44823 49479 44829
rect 57241 44863 57299 44869
rect 57241 44829 57253 44863
rect 57287 44829 57299 44863
rect 57241 44823 57299 44829
rect 57885 44863 57943 44869
rect 57885 44829 57897 44863
rect 57931 44860 57943 44863
rect 58986 44860 58992 44872
rect 57931 44832 58992 44860
rect 57931 44829 57943 44832
rect 57885 44823 57943 44829
rect 45526 44764 49280 44792
rect 49436 44792 49464 44823
rect 58986 44820 58992 44832
rect 59044 44820 59050 44872
rect 58161 44795 58219 44801
rect 49436 44764 57468 44792
rect 48682 44684 48688 44736
rect 48740 44684 48746 44736
rect 57330 44684 57336 44736
rect 57388 44684 57394 44736
rect 57440 44724 57468 44764
rect 58161 44761 58173 44795
rect 58207 44792 58219 44795
rect 59262 44792 59268 44804
rect 58207 44764 59268 44792
rect 58207 44761 58219 44764
rect 58161 44755 58219 44761
rect 59262 44752 59268 44764
rect 59320 44752 59326 44804
rect 58710 44724 58716 44736
rect 57440 44696 58716 44724
rect 58710 44684 58716 44696
rect 58768 44684 58774 44736
rect 1104 44634 58880 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 50294 44634
rect 50346 44582 50358 44634
rect 50410 44582 50422 44634
rect 50474 44582 50486 44634
rect 50538 44582 50550 44634
rect 50602 44582 58880 44634
rect 1104 44560 58880 44582
rect 41690 44412 41696 44464
rect 41748 44452 41754 44464
rect 41969 44455 42027 44461
rect 41969 44452 41981 44455
rect 41748 44424 41981 44452
rect 41748 44412 41754 44424
rect 41969 44421 41981 44424
rect 42015 44452 42027 44455
rect 42610 44452 42616 44464
rect 42015 44424 42616 44452
rect 42015 44421 42027 44424
rect 41969 44415 42027 44421
rect 42610 44412 42616 44424
rect 42668 44412 42674 44464
rect 1026 44344 1032 44396
rect 1084 44384 1090 44396
rect 1581 44387 1639 44393
rect 1581 44384 1593 44387
rect 1084 44356 1593 44384
rect 1084 44344 1090 44356
rect 1581 44353 1593 44356
rect 1627 44353 1639 44387
rect 1581 44347 1639 44353
rect 41414 44344 41420 44396
rect 41472 44384 41478 44396
rect 49326 44384 49332 44396
rect 41472 44356 49332 44384
rect 41472 44344 41478 44356
rect 49326 44344 49332 44356
rect 49384 44344 49390 44396
rect 58069 44387 58127 44393
rect 58069 44353 58081 44387
rect 58115 44384 58127 44387
rect 58986 44384 58992 44396
rect 58115 44356 58992 44384
rect 58115 44353 58127 44356
rect 58069 44347 58127 44353
rect 58986 44344 58992 44356
rect 59044 44344 59050 44396
rect 1765 44183 1823 44189
rect 1765 44149 1777 44183
rect 1811 44180 1823 44183
rect 26970 44180 26976 44192
rect 1811 44152 26976 44180
rect 1811 44149 1823 44152
rect 1765 44143 1823 44149
rect 26970 44140 26976 44152
rect 27028 44140 27034 44192
rect 58250 44140 58256 44192
rect 58308 44140 58314 44192
rect 1104 44090 58880 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 58880 44090
rect 1104 44016 58880 44038
rect 41616 43812 45554 43840
rect 41322 43732 41328 43784
rect 41380 43732 41386 43784
rect 41616 43781 41644 43812
rect 41601 43775 41659 43781
rect 41601 43741 41613 43775
rect 41647 43741 41659 43775
rect 41601 43735 41659 43741
rect 41690 43732 41696 43784
rect 41748 43732 41754 43784
rect 42613 43775 42671 43781
rect 42613 43741 42625 43775
rect 42659 43741 42671 43775
rect 45526 43772 45554 43812
rect 56134 43772 56140 43784
rect 45526 43744 56140 43772
rect 42613 43735 42671 43741
rect 934 43664 940 43716
rect 992 43704 998 43716
rect 1673 43707 1731 43713
rect 1673 43704 1685 43707
rect 992 43676 1685 43704
rect 992 43664 998 43676
rect 1673 43673 1685 43676
rect 1719 43673 1731 43707
rect 1673 43667 1731 43673
rect 1857 43707 1915 43713
rect 1857 43673 1869 43707
rect 1903 43704 1915 43707
rect 2314 43704 2320 43716
rect 1903 43676 2320 43704
rect 1903 43673 1915 43676
rect 1857 43667 1915 43673
rect 2314 43664 2320 43676
rect 2372 43664 2378 43716
rect 36998 43664 37004 43716
rect 37056 43704 37062 43716
rect 41509 43707 41567 43713
rect 41509 43704 41521 43707
rect 37056 43676 41521 43704
rect 37056 43664 37062 43676
rect 41509 43673 41521 43676
rect 41555 43673 41567 43707
rect 42429 43707 42487 43713
rect 42429 43704 42441 43707
rect 41509 43667 41567 43673
rect 41616 43676 42441 43704
rect 37918 43596 37924 43648
rect 37976 43636 37982 43648
rect 41616 43636 41644 43676
rect 42429 43673 42441 43676
rect 42475 43673 42487 43707
rect 42429 43667 42487 43673
rect 37976 43608 41644 43636
rect 41877 43639 41935 43645
rect 37976 43596 37982 43608
rect 41877 43605 41889 43639
rect 41923 43636 41935 43639
rect 42628 43636 42656 43735
rect 56134 43732 56140 43744
rect 56192 43732 56198 43784
rect 58066 43732 58072 43784
rect 58124 43732 58130 43784
rect 42886 43664 42892 43716
rect 42944 43704 42950 43716
rect 47210 43704 47216 43716
rect 42944 43676 47216 43704
rect 42944 43664 42950 43676
rect 47210 43664 47216 43676
rect 47268 43664 47274 43716
rect 41923 43608 42656 43636
rect 42797 43639 42855 43645
rect 41923 43605 41935 43608
rect 41877 43599 41935 43605
rect 42797 43605 42809 43639
rect 42843 43636 42855 43639
rect 57330 43636 57336 43648
rect 42843 43608 57336 43636
rect 42843 43605 42855 43608
rect 42797 43599 42855 43605
rect 57330 43596 57336 43608
rect 57388 43596 57394 43648
rect 58253 43639 58311 43645
rect 58253 43605 58265 43639
rect 58299 43636 58311 43639
rect 58710 43636 58716 43648
rect 58299 43608 58716 43636
rect 58299 43605 58311 43608
rect 58253 43599 58311 43605
rect 58710 43596 58716 43608
rect 58768 43596 58774 43648
rect 1104 43546 58880 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 50294 43546
rect 50346 43494 50358 43546
rect 50410 43494 50422 43546
rect 50474 43494 50486 43546
rect 50538 43494 50550 43546
rect 50602 43494 58880 43546
rect 1104 43472 58880 43494
rect 11698 43392 11704 43444
rect 11756 43432 11762 43444
rect 26142 43432 26148 43444
rect 11756 43404 26148 43432
rect 11756 43392 11762 43404
rect 26142 43392 26148 43404
rect 26200 43392 26206 43444
rect 33778 43392 33784 43444
rect 33836 43432 33842 43444
rect 42886 43432 42892 43444
rect 33836 43404 42892 43432
rect 33836 43392 33842 43404
rect 42886 43392 42892 43404
rect 42944 43392 42950 43444
rect 57882 43392 57888 43444
rect 57940 43432 57946 43444
rect 58066 43432 58072 43444
rect 57940 43404 58072 43432
rect 57940 43392 57946 43404
rect 58066 43392 58072 43404
rect 58124 43392 58130 43444
rect 1026 43256 1032 43308
rect 1084 43296 1090 43308
rect 1581 43299 1639 43305
rect 1581 43296 1593 43299
rect 1084 43268 1593 43296
rect 1084 43256 1090 43268
rect 1581 43265 1593 43268
rect 1627 43265 1639 43299
rect 1581 43259 1639 43265
rect 58069 43299 58127 43305
rect 58069 43265 58081 43299
rect 58115 43296 58127 43299
rect 58986 43296 58992 43308
rect 58115 43268 58992 43296
rect 58115 43265 58127 43268
rect 58069 43259 58127 43265
rect 58986 43256 58992 43268
rect 59044 43256 59050 43308
rect 1765 43095 1823 43101
rect 1765 43061 1777 43095
rect 1811 43092 1823 43095
rect 11698 43092 11704 43104
rect 1811 43064 11704 43092
rect 1811 43061 1823 43064
rect 1765 43055 1823 43061
rect 11698 43052 11704 43064
rect 11756 43052 11762 43104
rect 58253 43095 58311 43101
rect 58253 43061 58265 43095
rect 58299 43092 58311 43095
rect 59170 43092 59176 43104
rect 58299 43064 59176 43092
rect 58299 43061 58311 43064
rect 58253 43055 58311 43061
rect 59170 43052 59176 43064
rect 59228 43052 59234 43104
rect 1104 43002 58880 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 58880 43002
rect 1104 42928 58880 42950
rect 57977 42687 58035 42693
rect 57977 42653 57989 42687
rect 58023 42684 58035 42687
rect 58894 42684 58900 42696
rect 58023 42656 58900 42684
rect 58023 42653 58035 42656
rect 57977 42647 58035 42653
rect 58894 42644 58900 42656
rect 58952 42644 58958 42696
rect 934 42576 940 42628
rect 992 42616 998 42628
rect 1673 42619 1731 42625
rect 1673 42616 1685 42619
rect 992 42588 1685 42616
rect 992 42576 998 42588
rect 1673 42585 1685 42588
rect 1719 42585 1731 42619
rect 1673 42579 1731 42585
rect 1765 42551 1823 42557
rect 1765 42517 1777 42551
rect 1811 42548 1823 42551
rect 27890 42548 27896 42560
rect 1811 42520 27896 42548
rect 1811 42517 1823 42520
rect 1765 42511 1823 42517
rect 27890 42508 27896 42520
rect 27948 42508 27954 42560
rect 58253 42551 58311 42557
rect 58253 42517 58265 42551
rect 58299 42548 58311 42551
rect 58894 42548 58900 42560
rect 58299 42520 58900 42548
rect 58299 42517 58311 42520
rect 58253 42511 58311 42517
rect 58894 42508 58900 42520
rect 58952 42508 58958 42560
rect 1104 42458 58880 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 50294 42458
rect 50346 42406 50358 42458
rect 50410 42406 50422 42458
rect 50474 42406 50486 42458
rect 50538 42406 50550 42458
rect 50602 42406 58880 42458
rect 1104 42384 58880 42406
rect 31018 42344 31024 42356
rect 28092 42316 31024 42344
rect 28092 42288 28120 42316
rect 31018 42304 31024 42316
rect 31076 42304 31082 42356
rect 28074 42236 28080 42288
rect 28132 42236 28138 42288
rect 28166 42236 28172 42288
rect 28224 42236 28230 42288
rect 50890 42236 50896 42288
rect 50948 42276 50954 42288
rect 58526 42276 58532 42288
rect 50948 42248 58532 42276
rect 50948 42236 50954 42248
rect 58526 42236 58532 42248
rect 58584 42236 58590 42288
rect 1026 42168 1032 42220
rect 1084 42208 1090 42220
rect 1673 42211 1731 42217
rect 1673 42208 1685 42211
rect 1084 42180 1685 42208
rect 1084 42168 1090 42180
rect 1673 42177 1685 42180
rect 1719 42177 1731 42211
rect 1673 42171 1731 42177
rect 27890 42168 27896 42220
rect 27948 42168 27954 42220
rect 28258 42168 28264 42220
rect 28316 42208 28322 42220
rect 30466 42208 30472 42220
rect 28316 42180 30472 42208
rect 28316 42168 28322 42180
rect 30466 42168 30472 42180
rect 30524 42168 30530 42220
rect 58342 42168 58348 42220
rect 58400 42168 58406 42220
rect 37734 42100 37740 42152
rect 37792 42140 37798 42152
rect 56042 42140 56048 42152
rect 37792 42112 56048 42140
rect 37792 42100 37798 42112
rect 56042 42100 56048 42112
rect 56100 42100 56106 42152
rect 14458 42032 14464 42084
rect 14516 42072 14522 42084
rect 22738 42072 22744 42084
rect 14516 42044 22744 42072
rect 14516 42032 14522 42044
rect 22738 42032 22744 42044
rect 22796 42032 22802 42084
rect 33502 42032 33508 42084
rect 33560 42072 33566 42084
rect 55950 42072 55956 42084
rect 33560 42044 55956 42072
rect 33560 42032 33566 42044
rect 55950 42032 55956 42044
rect 56008 42032 56014 42084
rect 1765 42007 1823 42013
rect 1765 41973 1777 42007
rect 1811 42004 1823 42007
rect 26418 42004 26424 42016
rect 1811 41976 26424 42004
rect 1811 41973 1823 41976
rect 1765 41967 1823 41973
rect 26418 41964 26424 41976
rect 26476 41964 26482 42016
rect 28445 42007 28503 42013
rect 28445 41973 28457 42007
rect 28491 42004 28503 42007
rect 28534 42004 28540 42016
rect 28491 41976 28540 42004
rect 28491 41973 28503 41976
rect 28445 41967 28503 41973
rect 28534 41964 28540 41976
rect 28592 41964 28598 42016
rect 1104 41914 58880 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 58880 41914
rect 1104 41840 58880 41862
rect 26973 41735 27031 41741
rect 26973 41701 26985 41735
rect 27019 41732 27031 41735
rect 31846 41732 31852 41744
rect 27019 41704 31852 41732
rect 27019 41701 27031 41704
rect 26973 41695 27031 41701
rect 31846 41692 31852 41704
rect 31904 41692 31910 41744
rect 934 41556 940 41608
rect 992 41596 998 41608
rect 1581 41599 1639 41605
rect 1581 41596 1593 41599
rect 992 41568 1593 41596
rect 992 41556 998 41568
rect 1581 41565 1593 41568
rect 1627 41565 1639 41599
rect 1581 41559 1639 41565
rect 26418 41556 26424 41608
rect 26476 41556 26482 41608
rect 26694 41556 26700 41608
rect 26752 41556 26758 41608
rect 26841 41599 26899 41605
rect 26841 41565 26853 41599
rect 26887 41596 26899 41599
rect 28258 41596 28264 41608
rect 26887 41568 28264 41596
rect 26887 41565 26899 41568
rect 26841 41559 26899 41565
rect 28258 41556 28264 41568
rect 28316 41596 28322 41608
rect 28718 41596 28724 41608
rect 28316 41568 28724 41596
rect 28316 41556 28322 41568
rect 28718 41556 28724 41568
rect 28776 41556 28782 41608
rect 58345 41599 58403 41605
rect 58345 41565 58357 41599
rect 58391 41596 58403 41599
rect 58986 41596 58992 41608
rect 58391 41568 58992 41596
rect 58391 41565 58403 41568
rect 58345 41559 58403 41565
rect 58986 41556 58992 41568
rect 59044 41556 59050 41608
rect 26605 41531 26663 41537
rect 26605 41497 26617 41531
rect 26651 41528 26663 41531
rect 28074 41528 28080 41540
rect 26651 41500 28080 41528
rect 26651 41497 26663 41500
rect 26605 41491 26663 41497
rect 28074 41488 28080 41500
rect 28132 41488 28138 41540
rect 1765 41463 1823 41469
rect 1765 41429 1777 41463
rect 1811 41460 1823 41463
rect 21266 41460 21272 41472
rect 1811 41432 21272 41460
rect 1811 41429 1823 41432
rect 1765 41423 1823 41429
rect 21266 41420 21272 41432
rect 21324 41420 21330 41472
rect 1104 41370 58880 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 50294 41370
rect 50346 41318 50358 41370
rect 50410 41318 50422 41370
rect 50474 41318 50486 41370
rect 50538 41318 50550 41370
rect 50602 41318 58880 41370
rect 1104 41296 58880 41318
rect 1026 41080 1032 41132
rect 1084 41120 1090 41132
rect 1581 41123 1639 41129
rect 1581 41120 1593 41123
rect 1084 41092 1593 41120
rect 1084 41080 1090 41092
rect 1581 41089 1593 41092
rect 1627 41089 1639 41123
rect 1581 41083 1639 41089
rect 1765 40919 1823 40925
rect 1765 40885 1777 40919
rect 1811 40916 1823 40919
rect 9214 40916 9220 40928
rect 1811 40888 9220 40916
rect 1811 40885 1823 40888
rect 1765 40879 1823 40885
rect 9214 40876 9220 40888
rect 9272 40876 9278 40928
rect 58526 40876 58532 40928
rect 58584 40916 58590 40928
rect 58802 40916 58808 40928
rect 58584 40888 58808 40916
rect 58584 40876 58590 40888
rect 58802 40876 58808 40888
rect 58860 40876 58866 40928
rect 1104 40826 58880 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 58880 40826
rect 1104 40752 58880 40774
rect 58802 40672 58808 40724
rect 58860 40712 58866 40724
rect 59078 40712 59084 40724
rect 58860 40684 59084 40712
rect 58860 40672 58866 40684
rect 59078 40672 59084 40684
rect 59136 40672 59142 40724
rect 9677 40647 9735 40653
rect 9677 40613 9689 40647
rect 9723 40644 9735 40647
rect 9723 40616 40540 40644
rect 9723 40613 9735 40616
rect 9677 40607 9735 40613
rect 1857 40579 1915 40585
rect 1857 40545 1869 40579
rect 1903 40576 1915 40579
rect 1903 40548 9444 40576
rect 1903 40545 1915 40548
rect 1857 40539 1915 40545
rect 9122 40468 9128 40520
rect 9180 40468 9186 40520
rect 9416 40517 9444 40548
rect 9582 40517 9588 40520
rect 9401 40511 9459 40517
rect 9401 40477 9413 40511
rect 9447 40477 9459 40511
rect 9401 40471 9459 40477
rect 9545 40511 9588 40517
rect 9545 40477 9557 40511
rect 9545 40471 9588 40477
rect 9582 40468 9588 40471
rect 9640 40468 9646 40520
rect 31386 40468 31392 40520
rect 31444 40468 31450 40520
rect 40221 40511 40279 40517
rect 40221 40477 40233 40511
rect 40267 40477 40279 40511
rect 40221 40471 40279 40477
rect 934 40400 940 40452
rect 992 40440 998 40452
rect 1673 40443 1731 40449
rect 1673 40440 1685 40443
rect 992 40412 1685 40440
rect 992 40400 998 40412
rect 1673 40409 1685 40412
rect 1719 40409 1731 40443
rect 1673 40403 1731 40409
rect 9306 40400 9312 40452
rect 9364 40440 9370 40452
rect 10134 40440 10140 40452
rect 9364 40412 10140 40440
rect 9364 40400 9370 40412
rect 10134 40400 10140 40412
rect 10192 40400 10198 40452
rect 31205 40443 31263 40449
rect 31205 40409 31217 40443
rect 31251 40440 31263 40443
rect 40037 40443 40095 40449
rect 40037 40440 40049 40443
rect 31251 40412 40049 40440
rect 31251 40409 31263 40412
rect 31205 40403 31263 40409
rect 40037 40409 40049 40412
rect 40083 40409 40095 40443
rect 40236 40440 40264 40471
rect 40310 40468 40316 40520
rect 40368 40468 40374 40520
rect 40512 40517 40540 40616
rect 40497 40511 40555 40517
rect 40497 40477 40509 40511
rect 40543 40477 40555 40511
rect 40497 40471 40555 40477
rect 40586 40468 40592 40520
rect 40644 40468 40650 40520
rect 43714 40440 43720 40452
rect 40236 40412 43720 40440
rect 40037 40403 40095 40409
rect 43714 40400 43720 40412
rect 43772 40440 43778 40452
rect 49142 40440 49148 40452
rect 43772 40412 49148 40440
rect 43772 40400 43778 40412
rect 49142 40400 49148 40412
rect 49200 40400 49206 40452
rect 31478 40332 31484 40384
rect 31536 40332 31542 40384
rect 1104 40282 58880 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 50294 40282
rect 50346 40230 50358 40282
rect 50410 40230 50422 40282
rect 50474 40230 50486 40282
rect 50538 40230 50550 40282
rect 50602 40230 58880 40282
rect 1104 40208 58880 40230
rect 1026 40060 1032 40112
rect 1084 40100 1090 40112
rect 1673 40103 1731 40109
rect 1673 40100 1685 40103
rect 1084 40072 1685 40100
rect 1084 40060 1090 40072
rect 1673 40069 1685 40072
rect 1719 40069 1731 40103
rect 1673 40063 1731 40069
rect 58342 39856 58348 39908
rect 58400 39856 58406 39908
rect 1765 39831 1823 39837
rect 1765 39797 1777 39831
rect 1811 39828 1823 39831
rect 7650 39828 7656 39840
rect 1811 39800 7656 39828
rect 1811 39797 1823 39800
rect 1765 39791 1823 39797
rect 7650 39788 7656 39800
rect 7708 39788 7714 39840
rect 1104 39738 58880 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 58880 39738
rect 1104 39664 58880 39686
rect 7926 39516 7932 39568
rect 7984 39516 7990 39568
rect 7374 39380 7380 39432
rect 7432 39380 7438 39432
rect 7650 39380 7656 39432
rect 7708 39380 7714 39432
rect 7834 39429 7840 39432
rect 7797 39423 7840 39429
rect 7797 39389 7809 39423
rect 7797 39383 7840 39389
rect 7834 39380 7840 39383
rect 7892 39380 7898 39432
rect 9214 39380 9220 39432
rect 9272 39420 9278 39432
rect 29546 39420 29552 39432
rect 9272 39392 29552 39420
rect 9272 39380 9278 39392
rect 29546 39380 29552 39392
rect 29604 39380 29610 39432
rect 934 39312 940 39364
rect 992 39352 998 39364
rect 1673 39355 1731 39361
rect 1673 39352 1685 39355
rect 992 39324 1685 39352
rect 992 39312 998 39324
rect 1673 39321 1685 39324
rect 1719 39321 1731 39355
rect 1673 39315 1731 39321
rect 4890 39312 4896 39364
rect 4948 39352 4954 39364
rect 7561 39355 7619 39361
rect 7561 39352 7573 39355
rect 4948 39324 7573 39352
rect 4948 39312 4954 39324
rect 7561 39321 7573 39324
rect 7607 39352 7619 39355
rect 9306 39352 9312 39364
rect 7607 39324 9312 39352
rect 7607 39321 7619 39324
rect 7561 39315 7619 39321
rect 9306 39312 9312 39324
rect 9364 39312 9370 39364
rect 11698 39312 11704 39364
rect 11756 39352 11762 39364
rect 29362 39352 29368 39364
rect 11756 39324 29368 39352
rect 11756 39312 11762 39324
rect 29362 39312 29368 39324
rect 29420 39312 29426 39364
rect 1765 39287 1823 39293
rect 1765 39253 1777 39287
rect 1811 39284 1823 39287
rect 32674 39284 32680 39296
rect 1811 39256 32680 39284
rect 1811 39253 1823 39256
rect 1765 39247 1823 39253
rect 32674 39244 32680 39256
rect 32732 39244 32738 39296
rect 1104 39194 58880 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 50294 39194
rect 50346 39142 50358 39194
rect 50410 39142 50422 39194
rect 50474 39142 50486 39194
rect 50538 39142 50550 39194
rect 50602 39142 58880 39194
rect 1104 39120 58880 39142
rect 32953 39015 33011 39021
rect 32953 38981 32965 39015
rect 32999 39012 33011 39015
rect 55858 39012 55864 39024
rect 32999 38984 55864 39012
rect 32999 38981 33011 38984
rect 32953 38975 33011 38981
rect 55858 38972 55864 38984
rect 55916 38972 55922 39024
rect 1026 38904 1032 38956
rect 1084 38944 1090 38956
rect 1673 38947 1731 38953
rect 1673 38944 1685 38947
rect 1084 38916 1685 38944
rect 1084 38904 1090 38916
rect 1673 38913 1685 38916
rect 1719 38913 1731 38947
rect 1673 38907 1731 38913
rect 32674 38904 32680 38956
rect 32732 38904 32738 38956
rect 32858 38904 32864 38956
rect 32916 38904 32922 38956
rect 33042 38904 33048 38956
rect 33100 38904 33106 38956
rect 1857 38811 1915 38817
rect 1857 38777 1869 38811
rect 1903 38808 1915 38811
rect 4982 38808 4988 38820
rect 1903 38780 4988 38808
rect 1903 38777 1915 38780
rect 1857 38771 1915 38777
rect 4982 38768 4988 38780
rect 5040 38768 5046 38820
rect 29454 38700 29460 38752
rect 29512 38740 29518 38752
rect 31478 38740 31484 38752
rect 29512 38712 31484 38740
rect 29512 38700 29518 38712
rect 31478 38700 31484 38712
rect 31536 38700 31542 38752
rect 33229 38743 33287 38749
rect 33229 38709 33241 38743
rect 33275 38740 33287 38743
rect 33686 38740 33692 38752
rect 33275 38712 33692 38740
rect 33275 38709 33287 38712
rect 33229 38703 33287 38709
rect 33686 38700 33692 38712
rect 33744 38700 33750 38752
rect 58342 38700 58348 38752
rect 58400 38700 58406 38752
rect 1104 38650 58880 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 58880 38650
rect 1104 38576 58880 38598
rect 7834 38496 7840 38548
rect 7892 38536 7898 38548
rect 9582 38536 9588 38548
rect 7892 38508 9588 38536
rect 7892 38496 7898 38508
rect 9582 38496 9588 38508
rect 9640 38536 9646 38548
rect 11422 38536 11428 38548
rect 9640 38508 11428 38536
rect 9640 38496 9646 38508
rect 11422 38496 11428 38508
rect 11480 38496 11486 38548
rect 5258 38428 5264 38480
rect 5316 38428 5322 38480
rect 58158 38428 58164 38480
rect 58216 38468 58222 38480
rect 58434 38468 58440 38480
rect 58216 38440 58440 38468
rect 58216 38428 58222 38440
rect 58434 38428 58440 38440
rect 58492 38428 58498 38480
rect 33042 38360 33048 38412
rect 33100 38400 33106 38412
rect 33413 38403 33471 38409
rect 33413 38400 33425 38403
rect 33100 38372 33425 38400
rect 33100 38360 33106 38372
rect 33413 38369 33425 38372
rect 33459 38400 33471 38403
rect 33459 38372 35894 38400
rect 33459 38369 33471 38372
rect 33413 38363 33471 38369
rect 4706 38292 4712 38344
rect 4764 38292 4770 38344
rect 4890 38292 4896 38344
rect 4948 38292 4954 38344
rect 4982 38292 4988 38344
rect 5040 38292 5046 38344
rect 5082 38335 5140 38341
rect 5082 38301 5094 38335
rect 5128 38332 5140 38335
rect 7834 38332 7840 38344
rect 5128 38304 7840 38332
rect 5128 38301 5140 38304
rect 5082 38295 5140 38301
rect 934 38224 940 38276
rect 992 38264 998 38276
rect 1673 38267 1731 38273
rect 1673 38264 1685 38267
rect 992 38236 1685 38264
rect 992 38224 998 38236
rect 1673 38233 1685 38236
rect 1719 38233 1731 38267
rect 1673 38227 1731 38233
rect 3602 38224 3608 38276
rect 3660 38264 3666 38276
rect 5092 38264 5120 38295
rect 7834 38292 7840 38304
rect 7892 38292 7898 38344
rect 21266 38292 21272 38344
rect 21324 38332 21330 38344
rect 27154 38332 27160 38344
rect 21324 38304 27160 38332
rect 21324 38292 21330 38304
rect 27154 38292 27160 38304
rect 27212 38292 27218 38344
rect 33137 38335 33195 38341
rect 33137 38301 33149 38335
rect 33183 38332 33195 38335
rect 33226 38332 33232 38344
rect 33183 38304 33232 38332
rect 33183 38301 33195 38304
rect 33137 38295 33195 38301
rect 33226 38292 33232 38304
rect 33284 38292 33290 38344
rect 3660 38236 5120 38264
rect 35866 38264 35894 38372
rect 41414 38264 41420 38276
rect 35866 38236 41420 38264
rect 3660 38224 3666 38236
rect 41414 38224 41420 38236
rect 41472 38224 41478 38276
rect 1765 38199 1823 38205
rect 1765 38165 1777 38199
rect 1811 38196 1823 38199
rect 32674 38196 32680 38208
rect 1811 38168 32680 38196
rect 1811 38165 1823 38168
rect 1765 38159 1823 38165
rect 32674 38156 32680 38168
rect 32732 38156 32738 38208
rect 1104 38106 58880 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 50294 38106
rect 50346 38054 50358 38106
rect 50410 38054 50422 38106
rect 50474 38054 50486 38106
rect 50538 38054 50550 38106
rect 50602 38054 58880 38106
rect 1104 38032 58880 38054
rect 7190 37884 7196 37936
rect 7248 37924 7254 37936
rect 30558 37924 30564 37936
rect 7248 37896 30564 37924
rect 7248 37884 7254 37896
rect 30558 37884 30564 37896
rect 30616 37884 30622 37936
rect 32953 37927 33011 37933
rect 32953 37893 32965 37927
rect 32999 37924 33011 37927
rect 32999 37896 35894 37924
rect 32999 37893 33011 37896
rect 32953 37887 33011 37893
rect 1026 37816 1032 37868
rect 1084 37856 1090 37868
rect 1673 37859 1731 37865
rect 1673 37856 1685 37859
rect 1084 37828 1685 37856
rect 1084 37816 1090 37828
rect 1673 37825 1685 37828
rect 1719 37825 1731 37859
rect 1673 37819 1731 37825
rect 32674 37816 32680 37868
rect 32732 37816 32738 37868
rect 32858 37816 32864 37868
rect 32916 37816 32922 37868
rect 33042 37816 33048 37868
rect 33100 37865 33106 37868
rect 33100 37856 33108 37865
rect 35866 37856 35894 37896
rect 53282 37884 53288 37936
rect 53340 37924 53346 37936
rect 58066 37924 58072 37936
rect 53340 37896 58072 37924
rect 53340 37884 53346 37896
rect 58066 37884 58072 37896
rect 58124 37884 58130 37936
rect 57514 37856 57520 37868
rect 33100 37828 33145 37856
rect 35866 37828 57520 37856
rect 33100 37819 33108 37828
rect 33100 37816 33106 37819
rect 57514 37816 57520 37828
rect 57572 37816 57578 37868
rect 1857 37723 1915 37729
rect 1857 37689 1869 37723
rect 1903 37720 1915 37723
rect 3694 37720 3700 37732
rect 1903 37692 3700 37720
rect 1903 37689 1915 37692
rect 1857 37683 1915 37689
rect 3694 37680 3700 37692
rect 3752 37680 3758 37732
rect 33229 37655 33287 37661
rect 33229 37621 33241 37655
rect 33275 37652 33287 37655
rect 33594 37652 33600 37664
rect 33275 37624 33600 37652
rect 33275 37621 33287 37624
rect 33229 37615 33287 37621
rect 33594 37612 33600 37624
rect 33652 37612 33658 37664
rect 1104 37562 58880 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 58880 37562
rect 1104 37488 58880 37510
rect 1857 37315 1915 37321
rect 1857 37281 1869 37315
rect 1903 37312 1915 37315
rect 19426 37312 19432 37324
rect 1903 37284 19432 37312
rect 1903 37281 1915 37284
rect 1857 37275 1915 37281
rect 19426 37272 19432 37284
rect 19484 37272 19490 37324
rect 57514 37204 57520 37256
rect 57572 37244 57578 37256
rect 57885 37247 57943 37253
rect 57885 37244 57897 37247
rect 57572 37216 57897 37244
rect 57572 37204 57578 37216
rect 57885 37213 57897 37216
rect 57931 37213 57943 37247
rect 57885 37207 57943 37213
rect 58161 37247 58219 37253
rect 58161 37213 58173 37247
rect 58207 37244 58219 37247
rect 58986 37244 58992 37256
rect 58207 37216 58992 37244
rect 58207 37213 58219 37216
rect 58161 37207 58219 37213
rect 58986 37204 58992 37216
rect 59044 37204 59050 37256
rect 934 37136 940 37188
rect 992 37176 998 37188
rect 1673 37179 1731 37185
rect 1673 37176 1685 37179
rect 992 37148 1685 37176
rect 992 37136 998 37148
rect 1673 37145 1685 37148
rect 1719 37145 1731 37179
rect 1673 37139 1731 37145
rect 1104 37018 58880 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 50294 37018
rect 50346 36966 50358 37018
rect 50410 36966 50422 37018
rect 50474 36966 50486 37018
rect 50538 36966 50550 37018
rect 50602 36966 58880 37018
rect 1104 36944 58880 36966
rect 3418 36864 3424 36916
rect 3476 36904 3482 36916
rect 3476 36876 4476 36904
rect 3476 36864 3482 36876
rect 1026 36728 1032 36780
rect 1084 36768 1090 36780
rect 1673 36771 1731 36777
rect 1673 36768 1685 36771
rect 1084 36740 1685 36768
rect 1084 36728 1090 36740
rect 1673 36737 1685 36740
rect 1719 36737 1731 36771
rect 1673 36731 1731 36737
rect 3142 36728 3148 36780
rect 3200 36768 3206 36780
rect 3602 36768 3608 36780
rect 3200 36740 3608 36768
rect 3200 36728 3206 36740
rect 3602 36728 3608 36740
rect 3660 36728 3666 36780
rect 3694 36728 3700 36780
rect 3752 36728 3758 36780
rect 3878 36728 3884 36780
rect 3936 36768 3942 36780
rect 4448 36777 4476 36876
rect 3973 36771 4031 36777
rect 3973 36768 3985 36771
rect 3936 36740 3985 36768
rect 3936 36728 3942 36740
rect 3973 36737 3985 36740
rect 4019 36737 4031 36771
rect 3973 36731 4031 36737
rect 4249 36771 4307 36777
rect 4249 36737 4261 36771
rect 4295 36737 4307 36771
rect 4249 36731 4307 36737
rect 4433 36771 4491 36777
rect 4433 36737 4445 36771
rect 4479 36737 4491 36771
rect 4433 36731 4491 36737
rect 4264 36700 4292 36731
rect 19334 36728 19340 36780
rect 19392 36768 19398 36780
rect 19705 36771 19763 36777
rect 19705 36768 19717 36771
rect 19392 36740 19717 36768
rect 19392 36728 19398 36740
rect 19705 36737 19717 36740
rect 19751 36737 19763 36771
rect 19705 36731 19763 36737
rect 58066 36728 58072 36780
rect 58124 36728 58130 36780
rect 4614 36700 4620 36712
rect 4264 36672 4620 36700
rect 4614 36660 4620 36672
rect 4672 36700 4678 36712
rect 4890 36700 4896 36712
rect 4672 36672 4896 36700
rect 4672 36660 4678 36672
rect 4890 36660 4896 36672
rect 4948 36660 4954 36712
rect 11422 36660 11428 36712
rect 11480 36700 11486 36712
rect 21450 36700 21456 36712
rect 11480 36672 21456 36700
rect 11480 36660 11486 36672
rect 21450 36660 21456 36672
rect 21508 36660 21514 36712
rect 1857 36635 1915 36641
rect 1857 36601 1869 36635
rect 1903 36632 1915 36635
rect 2038 36632 2044 36644
rect 1903 36604 2044 36632
rect 1903 36601 1915 36604
rect 1857 36595 1915 36601
rect 2038 36592 2044 36604
rect 2096 36592 2102 36644
rect 31018 36632 31024 36644
rect 19628 36604 31024 36632
rect 3237 36567 3295 36573
rect 3237 36533 3249 36567
rect 3283 36564 3295 36567
rect 19628 36564 19656 36604
rect 31018 36592 31024 36604
rect 31076 36592 31082 36644
rect 3283 36536 19656 36564
rect 58253 36567 58311 36573
rect 3283 36533 3295 36536
rect 3237 36527 3295 36533
rect 58253 36533 58265 36567
rect 58299 36564 58311 36567
rect 59538 36564 59544 36576
rect 58299 36536 59544 36564
rect 58299 36533 58311 36536
rect 58253 36527 58311 36533
rect 59538 36524 59544 36536
rect 59596 36524 59602 36576
rect 1104 36474 58880 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 58880 36474
rect 1104 36400 58880 36422
rect 58158 36184 58164 36236
rect 58216 36184 58222 36236
rect 934 36116 940 36168
rect 992 36156 998 36168
rect 1581 36159 1639 36165
rect 1581 36156 1593 36159
rect 992 36128 1593 36156
rect 992 36116 998 36128
rect 1581 36125 1593 36128
rect 1627 36125 1639 36159
rect 1581 36119 1639 36125
rect 19426 36116 19432 36168
rect 19484 36156 19490 36168
rect 19889 36159 19947 36165
rect 19889 36156 19901 36159
rect 19484 36128 19901 36156
rect 19484 36116 19490 36128
rect 19889 36125 19901 36128
rect 19935 36125 19947 36159
rect 19889 36119 19947 36125
rect 20162 36116 20168 36168
rect 20220 36116 20226 36168
rect 20257 36159 20315 36165
rect 20257 36125 20269 36159
rect 20303 36156 20315 36159
rect 27798 36156 27804 36168
rect 20303 36128 27804 36156
rect 20303 36125 20315 36128
rect 20257 36119 20315 36125
rect 27798 36116 27804 36128
rect 27856 36156 27862 36168
rect 28350 36156 28356 36168
rect 27856 36128 28356 36156
rect 27856 36116 27862 36128
rect 28350 36116 28356 36128
rect 28408 36116 28414 36168
rect 30374 36116 30380 36168
rect 30432 36116 30438 36168
rect 30650 36116 30656 36168
rect 30708 36116 30714 36168
rect 31018 36116 31024 36168
rect 31076 36116 31082 36168
rect 31386 36116 31392 36168
rect 31444 36116 31450 36168
rect 55950 36116 55956 36168
rect 56008 36156 56014 36168
rect 57885 36159 57943 36165
rect 57885 36156 57897 36159
rect 56008 36128 57897 36156
rect 56008 36116 56014 36128
rect 57885 36125 57897 36128
rect 57931 36125 57943 36159
rect 57885 36119 57943 36125
rect 20073 36091 20131 36097
rect 20073 36057 20085 36091
rect 20119 36088 20131 36091
rect 21450 36088 21456 36100
rect 20119 36060 21456 36088
rect 20119 36057 20131 36060
rect 20073 36051 20131 36057
rect 21450 36048 21456 36060
rect 21508 36088 21514 36100
rect 31294 36088 31300 36100
rect 21508 36060 31300 36088
rect 21508 36048 21514 36060
rect 31294 36048 31300 36060
rect 31352 36088 31358 36100
rect 32858 36088 32864 36100
rect 31352 36060 32864 36088
rect 31352 36048 31358 36060
rect 32858 36048 32864 36060
rect 32916 36048 32922 36100
rect 1765 36023 1823 36029
rect 1765 35989 1777 36023
rect 1811 36020 1823 36023
rect 3418 36020 3424 36032
rect 1811 35992 3424 36020
rect 1811 35989 1823 35992
rect 1765 35983 1823 35989
rect 3418 35980 3424 35992
rect 3476 35980 3482 36032
rect 20441 36023 20499 36029
rect 20441 35989 20453 36023
rect 20487 36020 20499 36023
rect 28626 36020 28632 36032
rect 20487 35992 28632 36020
rect 20487 35989 20499 35992
rect 20441 35983 20499 35989
rect 28626 35980 28632 35992
rect 28684 35980 28690 36032
rect 30466 35980 30472 36032
rect 30524 35980 30530 36032
rect 45002 35980 45008 36032
rect 45060 36020 45066 36032
rect 46290 36020 46296 36032
rect 45060 35992 46296 36020
rect 45060 35980 45066 35992
rect 46290 35980 46296 35992
rect 46348 35980 46354 36032
rect 1104 35930 58880 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 50294 35930
rect 50346 35878 50358 35930
rect 50410 35878 50422 35930
rect 50474 35878 50486 35930
rect 50538 35878 50550 35930
rect 50602 35878 58880 35930
rect 1104 35856 58880 35878
rect 3237 35819 3295 35825
rect 3237 35785 3249 35819
rect 3283 35816 3295 35819
rect 3878 35816 3884 35828
rect 3283 35788 3884 35816
rect 3283 35785 3295 35788
rect 3237 35779 3295 35785
rect 3878 35776 3884 35788
rect 3936 35776 3942 35828
rect 28258 35776 28264 35828
rect 28316 35816 28322 35828
rect 33410 35816 33416 35828
rect 28316 35788 33416 35816
rect 28316 35776 28322 35788
rect 33410 35776 33416 35788
rect 33468 35776 33474 35828
rect 57974 35748 57980 35760
rect 2700 35720 57980 35748
rect 1026 35640 1032 35692
rect 1084 35680 1090 35692
rect 2700 35689 2728 35720
rect 57974 35708 57980 35720
rect 58032 35708 58038 35760
rect 58158 35708 58164 35760
rect 58216 35708 58222 35760
rect 1673 35683 1731 35689
rect 1673 35680 1685 35683
rect 1084 35652 1685 35680
rect 1084 35640 1090 35652
rect 1673 35649 1685 35652
rect 1719 35649 1731 35683
rect 1673 35643 1731 35649
rect 2409 35683 2467 35689
rect 2409 35649 2421 35683
rect 2455 35680 2467 35683
rect 2685 35683 2743 35689
rect 2685 35680 2697 35683
rect 2455 35652 2697 35680
rect 2455 35649 2467 35652
rect 2409 35643 2467 35649
rect 2685 35649 2697 35652
rect 2731 35649 2743 35683
rect 2685 35643 2743 35649
rect 2866 35640 2872 35692
rect 2924 35640 2930 35692
rect 2958 35640 2964 35692
rect 3016 35640 3022 35692
rect 3053 35683 3111 35689
rect 3053 35649 3065 35683
rect 3099 35680 3111 35683
rect 4062 35680 4068 35692
rect 3099 35652 4068 35680
rect 3099 35649 3111 35652
rect 3053 35643 3111 35649
rect 4062 35640 4068 35652
rect 4120 35640 4126 35692
rect 28169 35683 28227 35689
rect 28169 35649 28181 35683
rect 28215 35649 28227 35683
rect 28169 35643 28227 35649
rect 1946 35572 1952 35624
rect 2004 35612 2010 35624
rect 28184 35612 28212 35643
rect 28258 35640 28264 35692
rect 28316 35640 28322 35692
rect 28442 35640 28448 35692
rect 28500 35640 28506 35692
rect 28537 35683 28595 35689
rect 28537 35649 28549 35683
rect 28583 35680 28595 35683
rect 28626 35680 28632 35692
rect 28583 35652 28632 35680
rect 28583 35649 28595 35652
rect 28537 35643 28595 35649
rect 28626 35640 28632 35652
rect 28684 35640 28690 35692
rect 29086 35640 29092 35692
rect 29144 35640 29150 35692
rect 30834 35640 30840 35692
rect 30892 35680 30898 35692
rect 33229 35683 33287 35689
rect 33229 35680 33241 35683
rect 30892 35652 33241 35680
rect 30892 35640 30898 35652
rect 33229 35649 33241 35652
rect 33275 35649 33287 35683
rect 33229 35643 33287 35649
rect 28718 35612 28724 35624
rect 2004 35584 16574 35612
rect 28184 35584 28724 35612
rect 2004 35572 2010 35584
rect 1857 35547 1915 35553
rect 1857 35513 1869 35547
rect 1903 35544 1915 35547
rect 16546 35544 16574 35584
rect 28718 35572 28724 35584
rect 28776 35612 28782 35624
rect 29365 35615 29423 35621
rect 29365 35612 29377 35615
rect 28776 35584 29377 35612
rect 28776 35572 28782 35584
rect 29365 35581 29377 35584
rect 29411 35581 29423 35615
rect 33244 35612 33272 35643
rect 33318 35640 33324 35692
rect 33376 35640 33382 35692
rect 33410 35640 33416 35692
rect 33468 35680 33474 35692
rect 33505 35683 33563 35689
rect 33505 35680 33517 35683
rect 33468 35652 33517 35680
rect 33468 35640 33474 35652
rect 33505 35649 33517 35652
rect 33551 35649 33563 35683
rect 33505 35643 33563 35649
rect 33597 35683 33655 35689
rect 33597 35649 33609 35683
rect 33643 35680 33655 35683
rect 33686 35680 33692 35692
rect 33643 35652 33692 35680
rect 33643 35649 33655 35652
rect 33597 35643 33655 35649
rect 33686 35640 33692 35652
rect 33744 35640 33750 35692
rect 34790 35680 34796 35692
rect 33796 35652 34796 35680
rect 33796 35612 33824 35652
rect 34790 35640 34796 35652
rect 34848 35640 34854 35692
rect 33244 35584 33824 35612
rect 29365 35575 29423 35581
rect 33870 35572 33876 35624
rect 33928 35612 33934 35624
rect 43714 35612 43720 35624
rect 33928 35584 43720 35612
rect 33928 35572 33934 35584
rect 43714 35572 43720 35584
rect 43772 35572 43778 35624
rect 41138 35544 41144 35556
rect 1903 35516 6914 35544
rect 16546 35516 41144 35544
rect 1903 35513 1915 35516
rect 1857 35507 1915 35513
rect 6886 35476 6914 35516
rect 41138 35504 41144 35516
rect 41196 35504 41202 35556
rect 58345 35547 58403 35553
rect 58345 35513 58357 35547
rect 58391 35544 58403 35547
rect 59722 35544 59728 35556
rect 58391 35516 59728 35544
rect 58391 35513 58403 35516
rect 58345 35507 58403 35513
rect 59722 35504 59728 35516
rect 59780 35504 59786 35556
rect 23198 35476 23204 35488
rect 6886 35448 23204 35476
rect 23198 35436 23204 35448
rect 23256 35436 23262 35488
rect 27982 35436 27988 35488
rect 28040 35436 28046 35488
rect 28442 35436 28448 35488
rect 28500 35476 28506 35488
rect 30098 35476 30104 35488
rect 28500 35448 30104 35476
rect 28500 35436 28506 35448
rect 30098 35436 30104 35448
rect 30156 35436 30162 35488
rect 33045 35479 33103 35485
rect 33045 35445 33057 35479
rect 33091 35476 33103 35479
rect 33134 35476 33140 35488
rect 33091 35448 33140 35476
rect 33091 35445 33103 35448
rect 33045 35439 33103 35445
rect 33134 35436 33140 35448
rect 33192 35436 33198 35488
rect 1104 35386 58880 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 58880 35386
rect 1104 35312 58880 35334
rect 1762 35232 1768 35284
rect 1820 35272 1826 35284
rect 26694 35272 26700 35284
rect 1820 35244 26700 35272
rect 1820 35232 1826 35244
rect 26694 35232 26700 35244
rect 26752 35232 26758 35284
rect 31021 35275 31079 35281
rect 31021 35241 31033 35275
rect 31067 35272 31079 35275
rect 31386 35272 31392 35284
rect 31067 35244 31392 35272
rect 31067 35241 31079 35244
rect 31021 35235 31079 35241
rect 31386 35232 31392 35244
rect 31444 35232 31450 35284
rect 33870 35272 33876 35284
rect 31726 35244 33876 35272
rect 29086 35164 29092 35216
rect 29144 35204 29150 35216
rect 31726 35204 31754 35244
rect 33870 35232 33876 35244
rect 33928 35232 33934 35284
rect 29144 35176 31754 35204
rect 32401 35207 32459 35213
rect 29144 35164 29150 35176
rect 32401 35173 32413 35207
rect 32447 35204 32459 35207
rect 32953 35207 33011 35213
rect 32953 35204 32965 35207
rect 32447 35176 32965 35204
rect 32447 35173 32459 35176
rect 32401 35167 32459 35173
rect 32953 35173 32965 35176
rect 32999 35173 33011 35207
rect 57422 35204 57428 35216
rect 32953 35167 33011 35173
rect 33060 35176 57428 35204
rect 33060 35136 33088 35176
rect 57422 35164 57428 35176
rect 57480 35164 57486 35216
rect 31864 35108 33088 35136
rect 30469 35071 30527 35077
rect 30469 35037 30481 35071
rect 30515 35068 30527 35071
rect 30558 35068 30564 35080
rect 30515 35040 30564 35068
rect 30515 35037 30527 35040
rect 30469 35031 30527 35037
rect 30558 35028 30564 35040
rect 30616 35028 30622 35080
rect 30834 35028 30840 35080
rect 30892 35028 30898 35080
rect 31864 35077 31892 35108
rect 33226 35096 33232 35148
rect 33284 35136 33290 35148
rect 33410 35136 33416 35148
rect 33284 35108 33416 35136
rect 33284 35096 33290 35108
rect 33410 35096 33416 35108
rect 33468 35096 33474 35148
rect 33686 35096 33692 35148
rect 33744 35136 33750 35148
rect 58342 35136 58348 35148
rect 33744 35108 58348 35136
rect 33744 35096 33750 35108
rect 58342 35096 58348 35108
rect 58400 35096 58406 35148
rect 31849 35071 31907 35077
rect 31849 35037 31861 35071
rect 31895 35037 31907 35071
rect 32217 35071 32275 35077
rect 32217 35068 32229 35071
rect 31849 35031 31907 35037
rect 31956 35040 32229 35068
rect 934 34960 940 35012
rect 992 35000 998 35012
rect 1673 35003 1731 35009
rect 1673 35000 1685 35003
rect 992 34972 1685 35000
rect 992 34960 998 34972
rect 1673 34969 1685 34972
rect 1719 34969 1731 35003
rect 1673 34963 1731 34969
rect 28074 34960 28080 35012
rect 28132 35000 28138 35012
rect 30653 35003 30711 35009
rect 30653 35000 30665 35003
rect 28132 34972 30665 35000
rect 28132 34960 28138 34972
rect 30653 34969 30665 34972
rect 30699 34969 30711 35003
rect 30653 34963 30711 34969
rect 30742 34960 30748 35012
rect 30800 34960 30806 35012
rect 30852 34972 31156 35000
rect 1765 34935 1823 34941
rect 1765 34901 1777 34935
rect 1811 34932 1823 34935
rect 30852 34932 30880 34972
rect 1811 34904 30880 34932
rect 31128 34932 31156 34972
rect 31570 34960 31576 35012
rect 31628 35000 31634 35012
rect 31956 35000 31984 35040
rect 32217 35037 32229 35040
rect 32263 35037 32275 35071
rect 32217 35031 32275 35037
rect 31628 34972 31984 35000
rect 31628 34960 31634 34972
rect 32030 34960 32036 35012
rect 32088 34960 32094 35012
rect 32125 35003 32183 35009
rect 32125 34969 32137 35003
rect 32171 34969 32183 35003
rect 32232 35000 32260 35031
rect 32766 35028 32772 35080
rect 32824 35068 32830 35080
rect 32861 35071 32919 35077
rect 32861 35068 32873 35071
rect 32824 35040 32873 35068
rect 32824 35028 32830 35040
rect 32861 35037 32873 35040
rect 32907 35037 32919 35071
rect 32861 35031 32919 35037
rect 33134 35028 33140 35080
rect 33192 35028 33198 35080
rect 42242 35028 42248 35080
rect 42300 35028 42306 35080
rect 42705 35071 42763 35077
rect 42705 35037 42717 35071
rect 42751 35068 42763 35071
rect 42794 35068 42800 35080
rect 42751 35040 42800 35068
rect 42751 35037 42763 35040
rect 42705 35031 42763 35037
rect 42794 35028 42800 35040
rect 42852 35068 42858 35080
rect 43254 35068 43260 35080
rect 42852 35040 43260 35068
rect 42852 35028 42858 35040
rect 43254 35028 43260 35040
rect 43312 35028 43318 35080
rect 57606 35028 57612 35080
rect 57664 35068 57670 35080
rect 57885 35071 57943 35077
rect 57885 35068 57897 35071
rect 57664 35040 57897 35068
rect 57664 35028 57670 35040
rect 57885 35037 57897 35040
rect 57931 35037 57943 35071
rect 57885 35031 57943 35037
rect 32950 35000 32956 35012
rect 32232 34972 32956 35000
rect 32125 34963 32183 34969
rect 32140 34932 32168 34963
rect 32950 34960 32956 34972
rect 33008 34960 33014 35012
rect 58158 34960 58164 35012
rect 58216 34960 58222 35012
rect 59078 34960 59084 35012
rect 59136 35000 59142 35012
rect 59354 35000 59360 35012
rect 59136 34972 59360 35000
rect 59136 34960 59142 34972
rect 59354 34960 59360 34972
rect 59412 34960 59418 35012
rect 31128 34904 32168 34932
rect 1811 34901 1823 34904
rect 1765 34895 1823 34901
rect 32214 34892 32220 34944
rect 32272 34932 32278 34944
rect 32766 34932 32772 34944
rect 32272 34904 32772 34932
rect 32272 34892 32278 34904
rect 32766 34892 32772 34904
rect 32824 34892 32830 34944
rect 33321 34935 33379 34941
rect 33321 34901 33333 34935
rect 33367 34932 33379 34935
rect 33410 34932 33416 34944
rect 33367 34904 33416 34932
rect 33367 34901 33379 34904
rect 33321 34895 33379 34901
rect 33410 34892 33416 34904
rect 33468 34892 33474 34944
rect 1104 34842 58880 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 50294 34842
rect 50346 34790 50358 34842
rect 50410 34790 50422 34842
rect 50474 34790 50486 34842
rect 50538 34790 50550 34842
rect 50602 34790 58880 34842
rect 1104 34768 58880 34790
rect 1762 34688 1768 34740
rect 1820 34688 1826 34740
rect 10134 34688 10140 34740
rect 10192 34728 10198 34740
rect 24394 34728 24400 34740
rect 10192 34700 24400 34728
rect 10192 34688 10198 34700
rect 24394 34688 24400 34700
rect 24452 34688 24458 34740
rect 33413 34731 33471 34737
rect 33413 34728 33425 34731
rect 24504 34700 33425 34728
rect 5258 34620 5264 34672
rect 5316 34660 5322 34672
rect 24504 34660 24532 34700
rect 33413 34697 33425 34700
rect 33459 34728 33471 34731
rect 34054 34728 34060 34740
rect 33459 34700 34060 34728
rect 33459 34697 33471 34700
rect 33413 34691 33471 34697
rect 34054 34688 34060 34700
rect 34112 34688 34118 34740
rect 41138 34688 41144 34740
rect 41196 34688 41202 34740
rect 42794 34728 42800 34740
rect 41708 34700 42800 34728
rect 33686 34660 33692 34672
rect 5316 34632 24532 34660
rect 32692 34632 33692 34660
rect 5316 34620 5322 34632
rect 1026 34552 1032 34604
rect 1084 34592 1090 34604
rect 1673 34595 1731 34601
rect 1673 34592 1685 34595
rect 1084 34564 1685 34592
rect 1084 34552 1090 34564
rect 1673 34561 1685 34564
rect 1719 34561 1731 34595
rect 1673 34555 1731 34561
rect 24302 34552 24308 34604
rect 24360 34592 24366 34604
rect 24360 34564 24532 34592
rect 24360 34552 24366 34564
rect 24504 34524 24532 34564
rect 24578 34552 24584 34604
rect 24636 34592 24642 34604
rect 24673 34595 24731 34601
rect 24673 34592 24685 34595
rect 24636 34564 24685 34592
rect 24636 34552 24642 34564
rect 24673 34561 24685 34564
rect 24719 34561 24731 34595
rect 32398 34592 32404 34604
rect 24673 34555 24731 34561
rect 25424 34564 32404 34592
rect 25424 34524 25452 34564
rect 32398 34552 32404 34564
rect 32456 34552 32462 34604
rect 32490 34552 32496 34604
rect 32548 34552 32554 34604
rect 32692 34601 32720 34632
rect 33686 34620 33692 34632
rect 33744 34620 33750 34672
rect 33781 34663 33839 34669
rect 33781 34629 33793 34663
rect 33827 34660 33839 34663
rect 37550 34660 37556 34672
rect 33827 34632 37556 34660
rect 33827 34629 33839 34632
rect 33781 34623 33839 34629
rect 37550 34620 37556 34632
rect 37608 34620 37614 34672
rect 32641 34595 32720 34601
rect 32641 34561 32653 34595
rect 32687 34564 32720 34595
rect 32687 34561 32699 34564
rect 32641 34555 32699 34561
rect 32766 34552 32772 34604
rect 32824 34552 32830 34604
rect 32861 34595 32919 34601
rect 32861 34561 32873 34595
rect 32907 34561 32919 34595
rect 32861 34555 32919 34561
rect 24504 34496 25452 34524
rect 26694 34484 26700 34536
rect 26752 34524 26758 34536
rect 32876 34524 32904 34555
rect 32950 34552 32956 34604
rect 33008 34601 33014 34604
rect 33008 34592 33016 34601
rect 34698 34592 34704 34604
rect 33008 34564 33053 34592
rect 34164 34564 34704 34592
rect 33008 34555 33016 34564
rect 33008 34552 33014 34555
rect 34164 34533 34192 34564
rect 34698 34552 34704 34564
rect 34756 34552 34762 34604
rect 41156 34592 41184 34688
rect 41708 34669 41736 34700
rect 42794 34688 42800 34700
rect 42852 34688 42858 34740
rect 58253 34731 58311 34737
rect 58253 34697 58265 34731
rect 58299 34728 58311 34731
rect 59078 34728 59084 34740
rect 58299 34700 59084 34728
rect 58299 34697 58311 34700
rect 58253 34691 58311 34697
rect 59078 34688 59084 34700
rect 59136 34688 59142 34740
rect 41693 34663 41751 34669
rect 41693 34629 41705 34663
rect 41739 34629 41751 34663
rect 41693 34623 41751 34629
rect 41785 34663 41843 34669
rect 41785 34629 41797 34663
rect 41831 34660 41843 34663
rect 42426 34660 42432 34672
rect 41831 34632 42432 34660
rect 41831 34629 41843 34632
rect 41785 34623 41843 34629
rect 42426 34620 42432 34632
rect 42484 34620 42490 34672
rect 41509 34595 41567 34601
rect 41509 34592 41521 34595
rect 41156 34564 41521 34592
rect 41509 34561 41521 34564
rect 41555 34561 41567 34595
rect 41877 34595 41935 34601
rect 41877 34592 41889 34595
rect 41509 34555 41567 34561
rect 41708 34564 41889 34592
rect 41708 34536 41736 34564
rect 41877 34561 41889 34564
rect 41923 34561 41935 34595
rect 41877 34555 41935 34561
rect 42794 34552 42800 34604
rect 42852 34592 42858 34604
rect 43257 34595 43315 34601
rect 43257 34592 43269 34595
rect 42852 34564 43269 34592
rect 42852 34552 42858 34564
rect 43257 34561 43269 34564
rect 43303 34561 43315 34595
rect 43257 34555 43315 34561
rect 43622 34552 43628 34604
rect 43680 34552 43686 34604
rect 43714 34552 43720 34604
rect 43772 34552 43778 34604
rect 58066 34552 58072 34604
rect 58124 34552 58130 34604
rect 26752 34496 32904 34524
rect 34149 34527 34207 34533
rect 26752 34484 26758 34496
rect 34149 34493 34161 34527
rect 34195 34493 34207 34527
rect 34149 34487 34207 34493
rect 34330 34484 34336 34536
rect 34388 34484 34394 34536
rect 41690 34484 41696 34536
rect 41748 34484 41754 34536
rect 43165 34527 43223 34533
rect 43165 34524 43177 34527
rect 42076 34496 43177 34524
rect 33137 34459 33195 34465
rect 33137 34425 33149 34459
rect 33183 34456 33195 34459
rect 33919 34459 33977 34465
rect 33919 34456 33931 34459
rect 33183 34428 33931 34456
rect 33183 34425 33195 34428
rect 33137 34419 33195 34425
rect 33919 34425 33931 34428
rect 33965 34425 33977 34459
rect 33919 34419 33977 34425
rect 34054 34416 34060 34468
rect 34112 34416 34118 34468
rect 42076 34465 42104 34496
rect 43165 34493 43177 34496
rect 43211 34493 43223 34527
rect 43165 34487 43223 34493
rect 42061 34459 42119 34465
rect 42061 34425 42073 34459
rect 42107 34425 42119 34459
rect 42061 34419 42119 34425
rect 42705 34391 42763 34397
rect 42705 34357 42717 34391
rect 42751 34388 42763 34391
rect 42978 34388 42984 34400
rect 42751 34360 42984 34388
rect 42751 34357 42763 34360
rect 42705 34351 42763 34357
rect 42978 34348 42984 34360
rect 43036 34348 43042 34400
rect 1104 34298 58880 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 58880 34298
rect 1104 34224 58880 34246
rect 34698 34144 34704 34196
rect 34756 34184 34762 34196
rect 35253 34187 35311 34193
rect 35253 34184 35265 34187
rect 34756 34156 35265 34184
rect 34756 34144 34762 34156
rect 35253 34153 35265 34156
rect 35299 34153 35311 34187
rect 58526 34184 58532 34196
rect 35253 34147 35311 34153
rect 35866 34156 58532 34184
rect 4062 34076 4068 34128
rect 4120 34116 4126 34128
rect 4525 34119 4583 34125
rect 4120 34088 4384 34116
rect 4120 34076 4126 34088
rect 1857 34051 1915 34057
rect 1857 34017 1869 34051
rect 1903 34048 1915 34051
rect 1903 34020 4292 34048
rect 1903 34017 1915 34020
rect 1857 34011 1915 34017
rect 3970 33940 3976 33992
rect 4028 33940 4034 33992
rect 4264 33989 4292 34020
rect 4356 33989 4384 34088
rect 4525 34085 4537 34119
rect 4571 34116 4583 34119
rect 35866 34116 35894 34156
rect 58526 34144 58532 34156
rect 58584 34144 58590 34196
rect 4571 34088 6914 34116
rect 4571 34085 4583 34088
rect 4525 34079 4583 34085
rect 6886 34048 6914 34088
rect 34164 34088 35894 34116
rect 34164 34048 34192 34088
rect 42794 34076 42800 34128
rect 42852 34076 42858 34128
rect 6886 34020 22094 34048
rect 4249 33983 4307 33989
rect 4249 33949 4261 33983
rect 4295 33949 4307 33983
rect 4249 33943 4307 33949
rect 4346 33983 4404 33989
rect 4346 33949 4358 33983
rect 4392 33949 4404 33983
rect 22066 33980 22094 34020
rect 34072 34020 34192 34048
rect 34885 34051 34943 34057
rect 34072 33989 34100 34020
rect 34885 34017 34897 34051
rect 34931 34048 34943 34051
rect 39942 34048 39948 34060
rect 34931 34020 39948 34048
rect 34931 34017 34943 34020
rect 34885 34011 34943 34017
rect 39942 34008 39948 34020
rect 40000 34008 40006 34060
rect 42702 34008 42708 34060
rect 42760 34048 42766 34060
rect 42760 34020 43392 34048
rect 42760 34008 42766 34020
rect 33873 33983 33931 33989
rect 33873 33980 33885 33983
rect 22066 33952 33885 33980
rect 4346 33943 4404 33949
rect 33873 33949 33885 33952
rect 33919 33949 33931 33983
rect 33873 33943 33931 33949
rect 34057 33983 34115 33989
rect 34057 33949 34069 33983
rect 34103 33949 34115 33983
rect 34057 33943 34115 33949
rect 34149 33983 34207 33989
rect 34149 33949 34161 33983
rect 34195 33949 34207 33983
rect 34149 33943 34207 33949
rect 934 33872 940 33924
rect 992 33912 998 33924
rect 1673 33915 1731 33921
rect 1673 33912 1685 33915
rect 992 33884 1685 33912
rect 992 33872 998 33884
rect 1673 33881 1685 33884
rect 1719 33881 1731 33915
rect 1673 33875 1731 33881
rect 4157 33915 4215 33921
rect 4157 33881 4169 33915
rect 4203 33912 4215 33915
rect 4614 33912 4620 33924
rect 4203 33884 4620 33912
rect 4203 33881 4215 33884
rect 4157 33875 4215 33881
rect 4614 33872 4620 33884
rect 4672 33872 4678 33924
rect 32766 33872 32772 33924
rect 32824 33912 32830 33924
rect 33778 33912 33784 33924
rect 32824 33884 33784 33912
rect 32824 33872 32830 33884
rect 33778 33872 33784 33884
rect 33836 33912 33842 33924
rect 34164 33912 34192 33943
rect 34790 33940 34796 33992
rect 34848 33980 34854 33992
rect 35069 33983 35127 33989
rect 35069 33980 35081 33983
rect 34848 33952 35081 33980
rect 34848 33940 34854 33952
rect 35069 33949 35081 33952
rect 35115 33980 35127 33983
rect 42981 33983 43039 33989
rect 42981 33980 42993 33983
rect 35115 33952 42993 33980
rect 35115 33949 35127 33952
rect 35069 33943 35127 33949
rect 42981 33949 42993 33952
rect 43027 33949 43039 33983
rect 42981 33943 43039 33949
rect 43070 33940 43076 33992
rect 43128 33940 43134 33992
rect 43162 33940 43168 33992
rect 43220 33980 43226 33992
rect 43364 33989 43392 34020
rect 47946 34008 47952 34060
rect 48004 34008 48010 34060
rect 49050 34048 49056 34060
rect 48240 34020 49056 34048
rect 43257 33983 43315 33989
rect 43257 33980 43269 33983
rect 43220 33952 43269 33980
rect 43220 33940 43226 33952
rect 43257 33949 43269 33952
rect 43303 33949 43315 33983
rect 43257 33943 43315 33949
rect 43349 33983 43407 33989
rect 43349 33949 43361 33983
rect 43395 33949 43407 33983
rect 43349 33943 43407 33949
rect 47670 33940 47676 33992
rect 47728 33980 47734 33992
rect 48240 33989 48268 34020
rect 49050 34008 49056 34020
rect 49108 34008 49114 34060
rect 47857 33983 47915 33989
rect 47857 33980 47869 33983
rect 47728 33952 47869 33980
rect 47728 33940 47734 33952
rect 47857 33949 47869 33952
rect 47903 33949 47915 33983
rect 47857 33943 47915 33949
rect 48225 33983 48283 33989
rect 48225 33949 48237 33983
rect 48271 33949 48283 33983
rect 48225 33943 48283 33949
rect 48317 33983 48375 33989
rect 48317 33949 48329 33983
rect 48363 33949 48375 33983
rect 48317 33943 48375 33949
rect 33836 33884 34192 33912
rect 33836 33872 33842 33884
rect 46014 33872 46020 33924
rect 46072 33912 46078 33924
rect 47213 33915 47271 33921
rect 47213 33912 47225 33915
rect 46072 33884 47225 33912
rect 46072 33872 46078 33884
rect 47213 33881 47225 33884
rect 47259 33881 47271 33915
rect 48332 33912 48360 33943
rect 56686 33940 56692 33992
rect 56744 33980 56750 33992
rect 57885 33983 57943 33989
rect 57885 33980 57897 33983
rect 56744 33952 57897 33980
rect 56744 33940 56750 33952
rect 57885 33949 57897 33952
rect 57931 33949 57943 33983
rect 57885 33943 57943 33949
rect 47213 33875 47271 33881
rect 47872 33884 48360 33912
rect 47872 33856 47900 33884
rect 58158 33872 58164 33924
rect 58216 33872 58222 33924
rect 33962 33844 33968 33856
rect 34020 33853 34026 33856
rect 33929 33816 33968 33844
rect 33962 33804 33968 33816
rect 34020 33807 34029 33853
rect 34020 33804 34026 33807
rect 47854 33804 47860 33856
rect 47912 33804 47918 33856
rect 1104 33754 58880 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 50294 33754
rect 50346 33702 50358 33754
rect 50410 33702 50422 33754
rect 50474 33702 50486 33754
rect 50538 33702 50550 33754
rect 50602 33702 58880 33754
rect 1104 33680 58880 33702
rect 33226 33600 33232 33652
rect 33284 33600 33290 33652
rect 1857 33575 1915 33581
rect 1857 33541 1869 33575
rect 1903 33572 1915 33575
rect 2958 33572 2964 33584
rect 1903 33544 2964 33572
rect 1903 33541 1915 33544
rect 1857 33535 1915 33541
rect 2958 33532 2964 33544
rect 3016 33532 3022 33584
rect 33962 33532 33968 33584
rect 34020 33572 34026 33584
rect 34020 33544 34744 33572
rect 34020 33532 34026 33544
rect 1026 33464 1032 33516
rect 1084 33504 1090 33516
rect 1673 33507 1731 33513
rect 1673 33504 1685 33507
rect 1084 33476 1685 33504
rect 1084 33464 1090 33476
rect 1673 33473 1685 33476
rect 1719 33473 1731 33507
rect 1673 33467 1731 33473
rect 30098 33464 30104 33516
rect 30156 33504 30162 33516
rect 33134 33504 33140 33516
rect 30156 33476 33140 33504
rect 30156 33464 30162 33476
rect 33134 33464 33140 33476
rect 33192 33504 33198 33516
rect 33229 33507 33287 33513
rect 33229 33504 33241 33507
rect 33192 33476 33241 33504
rect 33192 33464 33198 33476
rect 33229 33473 33241 33476
rect 33275 33473 33287 33507
rect 33229 33467 33287 33473
rect 33594 33464 33600 33516
rect 33652 33464 33658 33516
rect 34716 33513 34744 33544
rect 34149 33507 34207 33513
rect 34149 33473 34161 33507
rect 34195 33473 34207 33507
rect 34149 33467 34207 33473
rect 34701 33507 34759 33513
rect 34701 33473 34713 33507
rect 34747 33473 34759 33507
rect 34701 33467 34759 33473
rect 34164 33436 34192 33467
rect 58066 33464 58072 33516
rect 58124 33464 58130 33516
rect 37090 33436 37096 33448
rect 34164 33408 37096 33436
rect 37090 33396 37096 33408
rect 37148 33396 37154 33448
rect 50982 33260 50988 33312
rect 51040 33300 51046 33312
rect 51442 33300 51448 33312
rect 51040 33272 51448 33300
rect 51040 33260 51046 33272
rect 51442 33260 51448 33272
rect 51500 33260 51506 33312
rect 58253 33303 58311 33309
rect 58253 33269 58265 33303
rect 58299 33300 58311 33303
rect 59630 33300 59636 33312
rect 58299 33272 59636 33300
rect 58299 33269 58311 33272
rect 58253 33263 58311 33269
rect 59630 33260 59636 33272
rect 59688 33260 59694 33312
rect 1104 33210 58880 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 58880 33210
rect 1104 33136 58880 33158
rect 1946 33056 1952 33108
rect 2004 33096 2010 33108
rect 2406 33096 2412 33108
rect 2004 33068 2412 33096
rect 2004 33056 2010 33068
rect 2406 33056 2412 33068
rect 2464 33056 2470 33108
rect 29730 33056 29736 33108
rect 29788 33096 29794 33108
rect 30190 33096 30196 33108
rect 29788 33068 30196 33096
rect 29788 33056 29794 33068
rect 30190 33056 30196 33068
rect 30248 33056 30254 33108
rect 50798 33056 50804 33108
rect 50856 33096 50862 33108
rect 57238 33096 57244 33108
rect 50856 33068 57244 33096
rect 50856 33056 50862 33068
rect 57238 33056 57244 33068
rect 57296 33056 57302 33108
rect 2222 32920 2228 32972
rect 2280 32960 2286 32972
rect 2406 32960 2412 32972
rect 2280 32932 2412 32960
rect 2280 32920 2286 32932
rect 2406 32920 2412 32932
rect 2464 32920 2470 32972
rect 23014 32920 23020 32972
rect 23072 32960 23078 32972
rect 29822 32960 29828 32972
rect 23072 32932 29828 32960
rect 23072 32920 23078 32932
rect 29822 32920 29828 32932
rect 29880 32920 29886 32972
rect 27893 32895 27951 32901
rect 27893 32861 27905 32895
rect 27939 32892 27951 32895
rect 28258 32892 28264 32904
rect 27939 32864 28264 32892
rect 27939 32861 27951 32864
rect 27893 32855 27951 32861
rect 28258 32852 28264 32864
rect 28316 32892 28322 32904
rect 42242 32892 42248 32904
rect 28316 32864 42248 32892
rect 28316 32852 28322 32864
rect 42242 32852 42248 32864
rect 42300 32852 42306 32904
rect 49878 32852 49884 32904
rect 49936 32892 49942 32904
rect 57885 32895 57943 32901
rect 57885 32892 57897 32895
rect 49936 32864 57897 32892
rect 49936 32852 49942 32864
rect 57885 32861 57897 32864
rect 57931 32861 57943 32895
rect 57885 32855 57943 32861
rect 934 32784 940 32836
rect 992 32824 998 32836
rect 1673 32827 1731 32833
rect 1673 32824 1685 32827
rect 992 32796 1685 32824
rect 992 32784 998 32796
rect 1673 32793 1685 32796
rect 1719 32793 1731 32827
rect 1673 32787 1731 32793
rect 27706 32784 27712 32836
rect 27764 32824 27770 32836
rect 28074 32824 28080 32836
rect 27764 32796 28080 32824
rect 27764 32784 27770 32796
rect 28074 32784 28080 32796
rect 28132 32824 28138 32836
rect 28353 32827 28411 32833
rect 28353 32824 28365 32827
rect 28132 32796 28365 32824
rect 28132 32784 28138 32796
rect 28353 32793 28365 32796
rect 28399 32793 28411 32827
rect 28353 32787 28411 32793
rect 58158 32784 58164 32836
rect 58216 32784 58222 32836
rect 1765 32759 1823 32765
rect 1765 32725 1777 32759
rect 1811 32756 1823 32759
rect 2314 32756 2320 32768
rect 1811 32728 2320 32756
rect 1811 32725 1823 32728
rect 1765 32719 1823 32725
rect 2314 32716 2320 32728
rect 2372 32716 2378 32768
rect 3418 32716 3424 32768
rect 3476 32756 3482 32768
rect 59262 32756 59268 32768
rect 3476 32728 59268 32756
rect 3476 32716 3482 32728
rect 59262 32716 59268 32728
rect 59320 32716 59326 32768
rect 1104 32666 58880 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 50294 32666
rect 50346 32614 50358 32666
rect 50410 32614 50422 32666
rect 50474 32614 50486 32666
rect 50538 32614 50550 32666
rect 50602 32614 58880 32666
rect 1104 32592 58880 32614
rect 2406 32552 2412 32564
rect 2240 32524 2412 32552
rect 2240 32493 2268 32524
rect 2406 32512 2412 32524
rect 2464 32512 2470 32564
rect 2866 32512 2872 32564
rect 2924 32552 2930 32564
rect 3234 32552 3240 32564
rect 2924 32524 3240 32552
rect 2924 32512 2930 32524
rect 3234 32512 3240 32524
rect 3292 32552 3298 32564
rect 3292 32524 3648 32552
rect 3292 32512 3298 32524
rect 2225 32487 2283 32493
rect 2225 32453 2237 32487
rect 2271 32453 2283 32487
rect 2225 32447 2283 32453
rect 2314 32444 2320 32496
rect 2372 32444 2378 32496
rect 3620 32493 3648 32524
rect 28166 32512 28172 32564
rect 28224 32552 28230 32564
rect 46474 32552 46480 32564
rect 28224 32524 46480 32552
rect 28224 32512 28230 32524
rect 46474 32512 46480 32524
rect 46532 32512 46538 32564
rect 3053 32487 3111 32493
rect 3053 32453 3065 32487
rect 3099 32484 3111 32487
rect 3605 32487 3663 32493
rect 3099 32456 3464 32484
rect 3099 32453 3111 32456
rect 3053 32447 3111 32453
rect 3436 32428 3464 32456
rect 3605 32453 3617 32487
rect 3651 32453 3663 32487
rect 3605 32447 3663 32453
rect 19978 32444 19984 32496
rect 20036 32484 20042 32496
rect 28261 32487 28319 32493
rect 28261 32484 28273 32487
rect 20036 32456 28273 32484
rect 20036 32444 20042 32456
rect 28261 32453 28273 32456
rect 28307 32453 28319 32487
rect 31478 32484 31484 32496
rect 28261 32447 28319 32453
rect 29012 32456 31484 32484
rect 2041 32419 2099 32425
rect 2041 32385 2053 32419
rect 2087 32416 2099 32419
rect 2130 32416 2136 32428
rect 2087 32388 2136 32416
rect 2087 32385 2099 32388
rect 2041 32379 2099 32385
rect 2130 32376 2136 32388
rect 2188 32376 2194 32428
rect 2409 32419 2467 32425
rect 2409 32385 2421 32419
rect 2455 32416 2467 32419
rect 2498 32416 2504 32428
rect 2455 32388 2504 32416
rect 2455 32385 2467 32388
rect 2409 32379 2467 32385
rect 2498 32376 2504 32388
rect 2556 32376 2562 32428
rect 3326 32376 3332 32428
rect 3384 32376 3390 32428
rect 3418 32376 3424 32428
rect 3476 32416 3482 32428
rect 3476 32388 3521 32416
rect 3476 32376 3482 32388
rect 3694 32376 3700 32428
rect 3752 32376 3758 32428
rect 3794 32419 3852 32425
rect 3794 32385 3806 32419
rect 3840 32416 3852 32419
rect 4062 32416 4068 32428
rect 3840 32388 4068 32416
rect 3840 32385 3852 32388
rect 3794 32379 3852 32385
rect 2516 32348 2544 32376
rect 3804 32348 3832 32379
rect 4062 32376 4068 32388
rect 4120 32416 4126 32428
rect 11790 32416 11796 32428
rect 4120 32388 11796 32416
rect 4120 32376 4126 32388
rect 11790 32376 11796 32388
rect 11848 32376 11854 32428
rect 27890 32376 27896 32428
rect 27948 32376 27954 32428
rect 28442 32425 28448 32428
rect 27986 32419 28044 32425
rect 27986 32385 27998 32419
rect 28032 32385 28044 32419
rect 28169 32419 28227 32425
rect 28169 32416 28181 32419
rect 27986 32379 28044 32385
rect 28092 32388 28181 32416
rect 2516 32320 3832 32348
rect 27614 32308 27620 32360
rect 27672 32348 27678 32360
rect 28000 32348 28028 32379
rect 27672 32320 28028 32348
rect 27672 32308 27678 32320
rect 28092 32292 28120 32388
rect 28169 32385 28181 32388
rect 28215 32385 28227 32419
rect 28169 32379 28227 32385
rect 28399 32419 28448 32425
rect 28399 32385 28411 32419
rect 28445 32385 28448 32419
rect 28399 32379 28448 32385
rect 28442 32376 28448 32379
rect 28500 32376 28506 32428
rect 29012 32425 29040 32456
rect 31478 32444 31484 32456
rect 31536 32444 31542 32496
rect 37553 32487 37611 32493
rect 37553 32484 37565 32487
rect 31726 32456 37565 32484
rect 28997 32419 29055 32425
rect 28997 32385 29009 32419
rect 29043 32385 29055 32419
rect 28997 32379 29055 32385
rect 29273 32419 29331 32425
rect 29273 32385 29285 32419
rect 29319 32385 29331 32419
rect 29273 32379 29331 32385
rect 29288 32348 29316 32379
rect 28424 32320 29316 32348
rect 3973 32283 4031 32289
rect 3973 32249 3985 32283
rect 4019 32280 4031 32283
rect 4019 32252 19334 32280
rect 4019 32249 4031 32252
rect 3973 32243 4031 32249
rect 2590 32172 2596 32224
rect 2648 32172 2654 32224
rect 19306 32212 19334 32252
rect 28074 32240 28080 32292
rect 28132 32240 28138 32292
rect 28424 32212 28452 32320
rect 29546 32308 29552 32360
rect 29604 32308 29610 32360
rect 29822 32308 29828 32360
rect 29880 32348 29886 32360
rect 31726 32348 31754 32456
rect 37553 32453 37565 32456
rect 37599 32453 37611 32487
rect 37553 32447 37611 32453
rect 43070 32444 43076 32496
rect 43128 32484 43134 32496
rect 54570 32484 54576 32496
rect 43128 32456 54576 32484
rect 43128 32444 43134 32456
rect 54570 32444 54576 32456
rect 54628 32444 54634 32496
rect 39942 32376 39948 32428
rect 40000 32416 40006 32428
rect 52822 32416 52828 32428
rect 40000 32388 52828 32416
rect 40000 32376 40006 32388
rect 52822 32376 52828 32388
rect 52880 32376 52886 32428
rect 58066 32376 58072 32428
rect 58124 32376 58130 32428
rect 29880 32320 31754 32348
rect 29880 32308 29886 32320
rect 28537 32283 28595 32289
rect 28537 32249 28549 32283
rect 28583 32280 28595 32283
rect 29089 32283 29147 32289
rect 29089 32280 29101 32283
rect 28583 32252 29101 32280
rect 28583 32249 28595 32252
rect 28537 32243 28595 32249
rect 29089 32249 29101 32252
rect 29135 32249 29147 32283
rect 29089 32243 29147 32249
rect 19306 32184 28452 32212
rect 28626 32172 28632 32224
rect 28684 32212 28690 32224
rect 30190 32212 30196 32224
rect 28684 32184 30196 32212
rect 28684 32172 28690 32184
rect 30190 32172 30196 32184
rect 30248 32172 30254 32224
rect 37826 32172 37832 32224
rect 37884 32172 37890 32224
rect 57974 32172 57980 32224
rect 58032 32212 58038 32224
rect 58253 32215 58311 32221
rect 58253 32212 58265 32215
rect 58032 32184 58265 32212
rect 58032 32172 58038 32184
rect 58253 32181 58265 32184
rect 58299 32181 58311 32215
rect 58253 32175 58311 32181
rect 1104 32122 58880 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 58880 32122
rect 1104 32048 58880 32070
rect 2501 32011 2559 32017
rect 2501 31977 2513 32011
rect 2547 32008 2559 32011
rect 27614 32008 27620 32020
rect 2547 31980 27620 32008
rect 2547 31977 2559 31980
rect 2501 31971 2559 31977
rect 27614 31968 27620 31980
rect 27672 31968 27678 32020
rect 27890 31968 27896 32020
rect 27948 32008 27954 32020
rect 28169 32011 28227 32017
rect 28169 32008 28181 32011
rect 27948 31980 28181 32008
rect 27948 31968 27954 31980
rect 28169 31977 28181 31980
rect 28215 31977 28227 32011
rect 28169 31971 28227 31977
rect 37090 31968 37096 32020
rect 37148 31968 37154 32020
rect 37826 31968 37832 32020
rect 37884 32008 37890 32020
rect 47762 32008 47768 32020
rect 37884 31980 47768 32008
rect 37884 31968 37890 31980
rect 47762 31968 47768 31980
rect 47820 31968 47826 32020
rect 1857 31943 1915 31949
rect 1857 31909 1869 31943
rect 1903 31940 1915 31943
rect 3694 31940 3700 31952
rect 1903 31912 3700 31940
rect 1903 31909 1915 31912
rect 1857 31903 1915 31909
rect 3694 31900 3700 31912
rect 3752 31900 3758 31952
rect 27341 31943 27399 31949
rect 27341 31909 27353 31943
rect 27387 31940 27399 31943
rect 27387 31912 27936 31940
rect 27387 31909 27399 31912
rect 27341 31903 27399 31909
rect 1026 31832 1032 31884
rect 1084 31872 1090 31884
rect 1084 31844 2452 31872
rect 1084 31832 1090 31844
rect 934 31764 940 31816
rect 992 31804 998 31816
rect 2424 31813 2452 31844
rect 26970 31832 26976 31884
rect 27028 31872 27034 31884
rect 27908 31872 27936 31912
rect 28166 31872 28172 31884
rect 27028 31844 27660 31872
rect 27028 31832 27034 31844
rect 27632 31813 27660 31844
rect 27908 31844 28172 31872
rect 1673 31807 1731 31813
rect 1673 31804 1685 31807
rect 992 31776 1685 31804
rect 992 31764 998 31776
rect 1673 31773 1685 31776
rect 1719 31773 1731 31807
rect 1673 31767 1731 31773
rect 2409 31807 2467 31813
rect 2409 31773 2421 31807
rect 2455 31773 2467 31807
rect 2409 31767 2467 31773
rect 27617 31807 27675 31813
rect 27617 31773 27629 31807
rect 27663 31773 27675 31807
rect 27617 31767 27675 31773
rect 27706 31764 27712 31816
rect 27764 31804 27770 31816
rect 27908 31813 27936 31844
rect 28166 31832 28172 31844
rect 28224 31832 28230 31884
rect 37844 31872 37872 31968
rect 54478 31900 54484 31952
rect 54536 31940 54542 31952
rect 54536 31912 57192 31940
rect 54536 31900 54542 31912
rect 36740 31844 37872 31872
rect 27801 31807 27859 31813
rect 27801 31804 27813 31807
rect 27764 31776 27813 31804
rect 27764 31764 27770 31776
rect 27801 31773 27813 31776
rect 27847 31773 27859 31807
rect 27801 31767 27859 31773
rect 27893 31807 27951 31813
rect 27893 31773 27905 31807
rect 27939 31773 27951 31807
rect 27893 31767 27951 31773
rect 27985 31807 28043 31813
rect 27985 31773 27997 31807
rect 28031 31804 28043 31807
rect 28074 31804 28080 31816
rect 28031 31776 28080 31804
rect 28031 31773 28043 31776
rect 27985 31767 28043 31773
rect 28074 31764 28080 31776
rect 28132 31804 28138 31816
rect 30834 31804 30840 31816
rect 28132 31776 30840 31804
rect 28132 31764 28138 31776
rect 30834 31764 30840 31776
rect 30892 31764 30898 31816
rect 36446 31764 36452 31816
rect 36504 31764 36510 31816
rect 36630 31813 36636 31816
rect 36597 31807 36636 31813
rect 36597 31773 36609 31807
rect 36597 31767 36636 31773
rect 36630 31764 36636 31767
rect 36688 31764 36694 31816
rect 36740 31813 36768 31844
rect 36725 31807 36783 31813
rect 36725 31773 36737 31807
rect 36771 31773 36783 31807
rect 36725 31767 36783 31773
rect 36814 31764 36820 31816
rect 36872 31764 36878 31816
rect 36998 31813 37004 31816
rect 36955 31807 37004 31813
rect 36955 31773 36967 31807
rect 37001 31773 37004 31807
rect 36955 31767 37004 31773
rect 36998 31764 37004 31767
rect 37056 31764 37062 31816
rect 56965 31807 57023 31813
rect 56965 31773 56977 31807
rect 57011 31804 57023 31807
rect 57054 31804 57060 31816
rect 57011 31776 57060 31804
rect 57011 31773 57023 31776
rect 56965 31767 57023 31773
rect 57054 31764 57060 31776
rect 57112 31764 57118 31816
rect 57164 31804 57192 31912
rect 57241 31875 57299 31881
rect 57241 31841 57253 31875
rect 57287 31872 57299 31875
rect 58894 31872 58900 31884
rect 57287 31844 58900 31872
rect 57287 31841 57299 31844
rect 57241 31835 57299 31841
rect 58894 31832 58900 31844
rect 58952 31832 58958 31884
rect 57885 31807 57943 31813
rect 57164 31776 57836 31804
rect 57808 31736 57836 31776
rect 57885 31773 57897 31807
rect 57931 31804 57943 31807
rect 58986 31804 58992 31816
rect 57931 31776 58992 31804
rect 57931 31773 57943 31776
rect 57885 31767 57943 31773
rect 58986 31764 58992 31776
rect 59044 31764 59050 31816
rect 58161 31739 58219 31745
rect 58161 31736 58173 31739
rect 57808 31708 58173 31736
rect 58161 31705 58173 31708
rect 58207 31705 58219 31739
rect 58161 31699 58219 31705
rect 1104 31578 58880 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 50294 31578
rect 50346 31526 50358 31578
rect 50410 31526 50422 31578
rect 50474 31526 50486 31578
rect 50538 31526 50550 31578
rect 50602 31526 58880 31578
rect 1104 31504 58880 31526
rect 2593 31467 2651 31473
rect 2593 31433 2605 31467
rect 2639 31464 2651 31467
rect 3326 31464 3332 31476
rect 2639 31436 3332 31464
rect 2639 31433 2651 31436
rect 2593 31427 2651 31433
rect 3326 31424 3332 31436
rect 3384 31424 3390 31476
rect 48225 31399 48283 31405
rect 48225 31365 48237 31399
rect 48271 31396 48283 31399
rect 58434 31396 58440 31408
rect 48271 31368 58440 31396
rect 48271 31365 48283 31368
rect 48225 31359 48283 31365
rect 58434 31356 58440 31368
rect 58492 31356 58498 31408
rect 2038 31288 2044 31340
rect 2096 31288 2102 31340
rect 2225 31331 2283 31337
rect 2225 31297 2237 31331
rect 2271 31297 2283 31331
rect 2225 31291 2283 31297
rect 2240 31260 2268 31291
rect 2314 31288 2320 31340
rect 2372 31288 2378 31340
rect 2409 31331 2467 31337
rect 2409 31297 2421 31331
rect 2455 31328 2467 31331
rect 2682 31328 2688 31340
rect 2455 31300 2688 31328
rect 2455 31297 2467 31300
rect 2409 31291 2467 31297
rect 2682 31288 2688 31300
rect 2740 31288 2746 31340
rect 48041 31331 48099 31337
rect 48041 31297 48053 31331
rect 48087 31328 48099 31331
rect 48130 31328 48136 31340
rect 48087 31300 48136 31328
rect 48087 31297 48099 31300
rect 48041 31291 48099 31297
rect 48130 31288 48136 31300
rect 48188 31288 48194 31340
rect 48314 31288 48320 31340
rect 48372 31288 48378 31340
rect 58066 31288 58072 31340
rect 58124 31288 58130 31340
rect 19426 31260 19432 31272
rect 2240 31232 19432 31260
rect 19426 31220 19432 31232
rect 19484 31220 19490 31272
rect 45554 31084 45560 31136
rect 45612 31124 45618 31136
rect 47857 31127 47915 31133
rect 47857 31124 47869 31127
rect 45612 31096 47869 31124
rect 45612 31084 45618 31096
rect 47857 31093 47869 31096
rect 47903 31093 47915 31127
rect 47857 31087 47915 31093
rect 58250 31084 58256 31136
rect 58308 31084 58314 31136
rect 1104 31034 58880 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 58880 31034
rect 1104 30960 58880 30982
rect 27614 30880 27620 30932
rect 27672 30920 27678 30932
rect 30742 30920 30748 30932
rect 27672 30892 30748 30920
rect 27672 30880 27678 30892
rect 30742 30880 30748 30892
rect 30800 30880 30806 30932
rect 48130 30880 48136 30932
rect 48188 30880 48194 30932
rect 58250 30920 58256 30932
rect 51046 30892 58256 30920
rect 29914 30852 29920 30864
rect 28373 30824 29920 30852
rect 934 30676 940 30728
rect 992 30716 998 30728
rect 1673 30719 1731 30725
rect 1673 30716 1685 30719
rect 992 30688 1685 30716
rect 992 30676 998 30688
rect 1673 30685 1685 30688
rect 1719 30685 1731 30719
rect 1673 30679 1731 30685
rect 26234 30676 26240 30728
rect 26292 30716 26298 30728
rect 28373 30725 28401 30824
rect 29914 30812 29920 30824
rect 29972 30812 29978 30864
rect 43898 30812 43904 30864
rect 43956 30852 43962 30864
rect 51046 30852 51074 30892
rect 58250 30880 58256 30892
rect 58308 30880 58314 30932
rect 43956 30824 51074 30852
rect 43956 30812 43962 30824
rect 29362 30744 29368 30796
rect 29420 30784 29426 30796
rect 29420 30756 29868 30784
rect 29420 30744 29426 30756
rect 28261 30719 28319 30725
rect 28261 30716 28273 30719
rect 26292 30688 28273 30716
rect 26292 30676 26298 30688
rect 28261 30685 28273 30688
rect 28307 30685 28319 30719
rect 28261 30679 28319 30685
rect 28354 30719 28412 30725
rect 28354 30685 28366 30719
rect 28400 30685 28412 30719
rect 28354 30679 28412 30685
rect 28718 30676 28724 30728
rect 28776 30725 28782 30728
rect 28776 30679 28784 30725
rect 28776 30676 28782 30679
rect 29638 30676 29644 30728
rect 29696 30716 29702 30728
rect 29840 30725 29868 30756
rect 41414 30744 41420 30796
rect 41472 30784 41478 30796
rect 41472 30756 47992 30784
rect 41472 30744 41478 30756
rect 30282 30725 30288 30728
rect 29733 30719 29791 30725
rect 29733 30716 29745 30719
rect 29696 30688 29745 30716
rect 29696 30676 29702 30688
rect 29733 30685 29745 30688
rect 29779 30685 29791 30719
rect 29733 30679 29791 30685
rect 29826 30719 29884 30725
rect 29826 30685 29838 30719
rect 29872 30685 29884 30719
rect 29826 30679 29884 30685
rect 30239 30719 30288 30725
rect 30239 30685 30251 30719
rect 30285 30685 30288 30719
rect 30239 30679 30288 30685
rect 30282 30676 30288 30679
rect 30340 30676 30346 30728
rect 31573 30719 31631 30725
rect 31573 30685 31585 30719
rect 31619 30716 31631 30719
rect 46566 30716 46572 30728
rect 31619 30688 46572 30716
rect 31619 30685 31631 30688
rect 31573 30679 31631 30685
rect 46566 30676 46572 30688
rect 46624 30676 46630 30728
rect 47578 30676 47584 30728
rect 47636 30676 47642 30728
rect 47762 30676 47768 30728
rect 47820 30676 47826 30728
rect 47964 30725 47992 30756
rect 47949 30719 48007 30725
rect 47949 30685 47961 30719
rect 47995 30685 48007 30719
rect 58618 30716 58624 30728
rect 47949 30679 48007 30685
rect 51046 30688 58624 30716
rect 28166 30608 28172 30660
rect 28224 30648 28230 30660
rect 28537 30651 28595 30657
rect 28537 30648 28549 30651
rect 28224 30620 28549 30648
rect 28224 30608 28230 30620
rect 28537 30617 28549 30620
rect 28583 30617 28595 30651
rect 28537 30611 28595 30617
rect 28626 30608 28632 30660
rect 28684 30608 28690 30660
rect 30009 30651 30067 30657
rect 30009 30648 30021 30651
rect 28828 30620 30021 30648
rect 1762 30540 1768 30592
rect 1820 30540 1826 30592
rect 27706 30540 27712 30592
rect 27764 30580 27770 30592
rect 28828 30580 28856 30620
rect 30009 30617 30021 30620
rect 30055 30617 30067 30651
rect 30009 30611 30067 30617
rect 30101 30651 30159 30657
rect 30101 30617 30113 30651
rect 30147 30648 30159 30651
rect 30147 30620 31754 30648
rect 30147 30617 30159 30620
rect 30101 30611 30159 30617
rect 27764 30552 28856 30580
rect 28905 30583 28963 30589
rect 27764 30540 27770 30552
rect 28905 30549 28917 30583
rect 28951 30580 28963 30583
rect 29730 30580 29736 30592
rect 28951 30552 29736 30580
rect 28951 30549 28963 30552
rect 28905 30543 28963 30549
rect 29730 30540 29736 30552
rect 29788 30540 29794 30592
rect 30374 30540 30380 30592
rect 30432 30540 30438 30592
rect 31726 30580 31754 30620
rect 32122 30608 32128 30660
rect 32180 30608 32186 30660
rect 36538 30580 36544 30592
rect 31726 30552 36544 30580
rect 36538 30540 36544 30552
rect 36596 30540 36602 30592
rect 47780 30580 47808 30676
rect 47857 30651 47915 30657
rect 47857 30617 47869 30651
rect 47903 30648 47915 30651
rect 51046 30648 51074 30688
rect 58618 30676 58624 30688
rect 58676 30676 58682 30728
rect 47903 30620 51074 30648
rect 47903 30617 47915 30620
rect 47857 30611 47915 30617
rect 58158 30608 58164 30660
rect 58216 30608 58222 30660
rect 48682 30580 48688 30592
rect 47780 30552 48688 30580
rect 48682 30540 48688 30552
rect 48740 30540 48746 30592
rect 56318 30540 56324 30592
rect 56376 30580 56382 30592
rect 58253 30583 58311 30589
rect 58253 30580 58265 30583
rect 56376 30552 58265 30580
rect 56376 30540 56382 30552
rect 58253 30549 58265 30552
rect 58299 30549 58311 30583
rect 58253 30543 58311 30549
rect 1104 30490 58880 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 50294 30490
rect 50346 30438 50358 30490
rect 50410 30438 50422 30490
rect 50474 30438 50486 30490
rect 50538 30438 50550 30490
rect 50602 30438 58880 30490
rect 1104 30416 58880 30438
rect 1762 30336 1768 30388
rect 1820 30376 1826 30388
rect 28626 30376 28632 30388
rect 1820 30348 28632 30376
rect 1820 30336 1826 30348
rect 28626 30336 28632 30348
rect 28684 30336 28690 30388
rect 29638 30336 29644 30388
rect 29696 30376 29702 30388
rect 30098 30376 30104 30388
rect 29696 30348 30104 30376
rect 29696 30336 29702 30348
rect 30098 30336 30104 30348
rect 30156 30376 30162 30388
rect 30834 30376 30840 30388
rect 30156 30348 30840 30376
rect 30156 30336 30162 30348
rect 30834 30336 30840 30348
rect 30892 30336 30898 30388
rect 934 30268 940 30320
rect 992 30308 998 30320
rect 1673 30311 1731 30317
rect 1673 30308 1685 30311
rect 992 30280 1685 30308
rect 992 30268 998 30280
rect 1673 30277 1685 30280
rect 1719 30277 1731 30311
rect 1673 30271 1731 30277
rect 1857 30311 1915 30317
rect 1857 30277 1869 30311
rect 1903 30308 1915 30311
rect 2777 30311 2835 30317
rect 2777 30308 2789 30311
rect 1903 30280 2789 30308
rect 1903 30277 1915 30280
rect 1857 30271 1915 30277
rect 2777 30277 2789 30280
rect 2823 30277 2835 30311
rect 2777 30271 2835 30277
rect 6886 30280 17080 30308
rect 2590 30200 2596 30252
rect 2648 30200 2654 30252
rect 2682 30200 2688 30252
rect 2740 30240 2746 30252
rect 2869 30243 2927 30249
rect 2869 30240 2881 30243
rect 2740 30212 2881 30240
rect 2740 30200 2746 30212
rect 2869 30209 2881 30212
rect 2915 30240 2927 30243
rect 6886 30240 6914 30280
rect 2915 30212 6914 30240
rect 2915 30209 2927 30212
rect 2869 30203 2927 30209
rect 13814 30200 13820 30252
rect 13872 30240 13878 30252
rect 17052 30249 17080 30280
rect 17126 30268 17132 30320
rect 17184 30268 17190 30320
rect 22830 30268 22836 30320
rect 22888 30268 22894 30320
rect 29730 30268 29736 30320
rect 29788 30308 29794 30320
rect 29788 30280 30788 30308
rect 29788 30268 29794 30280
rect 16853 30243 16911 30249
rect 16853 30240 16865 30243
rect 13872 30212 16865 30240
rect 13872 30200 13878 30212
rect 16853 30209 16865 30212
rect 16899 30209 16911 30243
rect 16853 30203 16911 30209
rect 17037 30243 17095 30249
rect 17037 30209 17049 30243
rect 17083 30209 17095 30243
rect 17037 30203 17095 30209
rect 17052 30172 17080 30203
rect 17218 30200 17224 30252
rect 17276 30200 17282 30252
rect 22462 30200 22468 30252
rect 22520 30240 22526 30252
rect 22741 30243 22799 30249
rect 22741 30240 22753 30243
rect 22520 30212 22753 30240
rect 22520 30200 22526 30212
rect 22741 30209 22753 30212
rect 22787 30209 22799 30243
rect 22741 30203 22799 30209
rect 22922 30200 22928 30252
rect 22980 30200 22986 30252
rect 23106 30249 23112 30252
rect 23063 30243 23112 30249
rect 23063 30209 23075 30243
rect 23109 30209 23112 30243
rect 23063 30203 23112 30209
rect 23106 30200 23112 30203
rect 23164 30200 23170 30252
rect 23198 30200 23204 30252
rect 23256 30200 23262 30252
rect 23290 30200 23296 30252
rect 23348 30240 23354 30252
rect 24210 30240 24216 30252
rect 23348 30212 24216 30240
rect 23348 30200 23354 30212
rect 24210 30200 24216 30212
rect 24268 30240 24274 30252
rect 28718 30240 28724 30252
rect 24268 30212 28724 30240
rect 24268 30200 24274 30212
rect 28718 30200 28724 30212
rect 28776 30200 28782 30252
rect 30285 30243 30343 30249
rect 30285 30209 30297 30243
rect 30331 30209 30343 30243
rect 30285 30203 30343 30209
rect 22370 30172 22376 30184
rect 17052 30144 22376 30172
rect 22370 30132 22376 30144
rect 22428 30132 22434 30184
rect 26234 30172 26240 30184
rect 22480 30144 26240 30172
rect 17405 30107 17463 30113
rect 17405 30073 17417 30107
rect 17451 30104 17463 30107
rect 22480 30104 22508 30144
rect 26234 30132 26240 30144
rect 26292 30132 26298 30184
rect 30006 30132 30012 30184
rect 30064 30172 30070 30184
rect 30300 30172 30328 30203
rect 30374 30200 30380 30252
rect 30432 30200 30438 30252
rect 30760 30249 30788 30280
rect 48222 30268 48228 30320
rect 48280 30308 48286 30320
rect 53190 30308 53196 30320
rect 48280 30280 53196 30308
rect 48280 30268 48286 30280
rect 53190 30268 53196 30280
rect 53248 30268 53254 30320
rect 30745 30243 30803 30249
rect 30745 30209 30757 30243
rect 30791 30209 30803 30243
rect 30745 30203 30803 30209
rect 31202 30200 31208 30252
rect 31260 30200 31266 30252
rect 31481 30243 31539 30249
rect 31481 30209 31493 30243
rect 31527 30240 31539 30243
rect 32122 30240 32128 30252
rect 31527 30212 32128 30240
rect 31527 30209 31539 30212
rect 31481 30203 31539 30209
rect 32122 30200 32128 30212
rect 32180 30240 32186 30252
rect 36814 30240 36820 30252
rect 32180 30212 36820 30240
rect 32180 30200 32186 30212
rect 36814 30200 36820 30212
rect 36872 30200 36878 30252
rect 47578 30200 47584 30252
rect 47636 30240 47642 30252
rect 52730 30240 52736 30252
rect 47636 30212 52736 30240
rect 47636 30200 47642 30212
rect 52730 30200 52736 30212
rect 52788 30200 52794 30252
rect 58066 30200 58072 30252
rect 58124 30200 58130 30252
rect 30064 30144 31754 30172
rect 30064 30132 30070 30144
rect 17451 30076 22508 30104
rect 22557 30107 22615 30113
rect 17451 30073 17463 30076
rect 17405 30067 17463 30073
rect 22557 30073 22569 30107
rect 22603 30104 22615 30107
rect 31726 30104 31754 30144
rect 45554 30104 45560 30116
rect 22603 30076 31616 30104
rect 31726 30076 45560 30104
rect 22603 30073 22615 30076
rect 22557 30067 22615 30073
rect 2409 30039 2467 30045
rect 2409 30005 2421 30039
rect 2455 30036 2467 30039
rect 22278 30036 22284 30048
rect 2455 30008 22284 30036
rect 2455 30005 2467 30008
rect 2409 29999 2467 30005
rect 22278 29996 22284 30008
rect 22336 29996 22342 30048
rect 22830 29996 22836 30048
rect 22888 30036 22894 30048
rect 23750 30036 23756 30048
rect 22888 30008 23756 30036
rect 22888 29996 22894 30008
rect 23750 29996 23756 30008
rect 23808 29996 23814 30048
rect 28166 29996 28172 30048
rect 28224 30036 28230 30048
rect 28350 30036 28356 30048
rect 28224 30008 28356 30036
rect 28224 29996 28230 30008
rect 28350 29996 28356 30008
rect 28408 30036 28414 30048
rect 30558 30036 30564 30048
rect 28408 30008 30564 30036
rect 28408 29996 28414 30008
rect 30558 29996 30564 30008
rect 30616 29996 30622 30048
rect 31588 30036 31616 30076
rect 45554 30064 45560 30076
rect 45612 30064 45618 30116
rect 32582 30036 32588 30048
rect 31588 30008 32588 30036
rect 32582 29996 32588 30008
rect 32640 29996 32646 30048
rect 41874 29996 41880 30048
rect 41932 30036 41938 30048
rect 58253 30039 58311 30045
rect 58253 30036 58265 30039
rect 41932 30008 58265 30036
rect 41932 29996 41938 30008
rect 58253 30005 58265 30008
rect 58299 30005 58311 30039
rect 58253 29999 58311 30005
rect 1104 29946 58880 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 58880 29946
rect 1104 29872 58880 29894
rect 32677 29835 32735 29841
rect 32677 29832 32689 29835
rect 22066 29804 32689 29832
rect 1857 29767 1915 29773
rect 1857 29733 1869 29767
rect 1903 29764 1915 29767
rect 2314 29764 2320 29776
rect 1903 29736 2320 29764
rect 1903 29733 1915 29736
rect 1857 29727 1915 29733
rect 2314 29724 2320 29736
rect 2372 29724 2378 29776
rect 7926 29724 7932 29776
rect 7984 29764 7990 29776
rect 22066 29764 22094 29804
rect 32677 29801 32689 29804
rect 32723 29801 32735 29835
rect 32677 29795 32735 29801
rect 7984 29736 22094 29764
rect 7984 29724 7990 29736
rect 27982 29724 27988 29776
rect 28040 29764 28046 29776
rect 28537 29767 28595 29773
rect 28537 29764 28549 29767
rect 28040 29736 28549 29764
rect 28040 29724 28046 29736
rect 28537 29733 28549 29736
rect 28583 29733 28595 29767
rect 28537 29727 28595 29733
rect 29825 29767 29883 29773
rect 29825 29733 29837 29767
rect 29871 29764 29883 29767
rect 30374 29764 30380 29776
rect 29871 29736 30380 29764
rect 29871 29733 29883 29736
rect 29825 29727 29883 29733
rect 30374 29724 30380 29736
rect 30432 29724 30438 29776
rect 32582 29724 32588 29776
rect 32640 29724 32646 29776
rect 33318 29724 33324 29776
rect 33376 29764 33382 29776
rect 33376 29736 34100 29764
rect 33376 29724 33382 29736
rect 23106 29696 23112 29708
rect 19306 29668 23112 29696
rect 934 29588 940 29640
rect 992 29628 998 29640
rect 1673 29631 1731 29637
rect 1673 29628 1685 29631
rect 992 29600 1685 29628
rect 992 29588 998 29600
rect 1673 29597 1685 29600
rect 1719 29597 1731 29631
rect 1673 29591 1731 29597
rect 1026 29520 1032 29572
rect 1084 29560 1090 29572
rect 2409 29563 2467 29569
rect 2409 29560 2421 29563
rect 1084 29532 2421 29560
rect 1084 29520 1090 29532
rect 2409 29529 2421 29532
rect 2455 29529 2467 29563
rect 2409 29523 2467 29529
rect 11790 29520 11796 29572
rect 11848 29560 11854 29572
rect 19306 29560 19334 29668
rect 23106 29656 23112 29668
rect 23164 29696 23170 29708
rect 31386 29696 31392 29708
rect 23164 29668 23888 29696
rect 23164 29656 23170 29668
rect 23201 29631 23259 29637
rect 23201 29597 23213 29631
rect 23247 29628 23259 29631
rect 23290 29628 23296 29640
rect 23247 29600 23296 29628
rect 23247 29597 23259 29600
rect 23201 29591 23259 29597
rect 23290 29588 23296 29600
rect 23348 29588 23354 29640
rect 23860 29637 23888 29668
rect 28368 29668 31392 29696
rect 23845 29631 23903 29637
rect 23845 29597 23857 29631
rect 23891 29628 23903 29631
rect 28368 29628 28396 29668
rect 31386 29656 31392 29668
rect 31444 29656 31450 29708
rect 32309 29699 32367 29705
rect 32309 29665 32321 29699
rect 32355 29696 32367 29699
rect 33962 29696 33968 29708
rect 32355 29668 33968 29696
rect 32355 29665 32367 29668
rect 32309 29659 32367 29665
rect 33962 29656 33968 29668
rect 34020 29656 34026 29708
rect 34072 29696 34100 29736
rect 36630 29724 36636 29776
rect 36688 29764 36694 29776
rect 51534 29764 51540 29776
rect 36688 29736 51540 29764
rect 36688 29724 36694 29736
rect 51534 29724 51540 29736
rect 51592 29724 51598 29776
rect 49694 29696 49700 29708
rect 34072 29668 49700 29696
rect 49694 29656 49700 29668
rect 49752 29656 49758 29708
rect 58158 29656 58164 29708
rect 58216 29656 58222 29708
rect 23891 29600 28396 29628
rect 23891 29597 23903 29600
rect 23845 29591 23903 29597
rect 28442 29588 28448 29640
rect 28500 29588 28506 29640
rect 28718 29588 28724 29640
rect 28776 29588 28782 29640
rect 29730 29588 29736 29640
rect 29788 29588 29794 29640
rect 30006 29588 30012 29640
rect 30064 29588 30070 29640
rect 32582 29588 32588 29640
rect 32640 29628 32646 29640
rect 32769 29631 32827 29637
rect 32769 29628 32781 29631
rect 32640 29600 32781 29628
rect 32640 29588 32646 29600
rect 32769 29597 32781 29600
rect 32815 29597 32827 29631
rect 32769 29591 32827 29597
rect 33045 29631 33103 29637
rect 33045 29597 33057 29631
rect 33091 29597 33103 29631
rect 33045 29591 33103 29597
rect 11848 29532 19334 29560
rect 28169 29563 28227 29569
rect 11848 29520 11854 29532
rect 28169 29529 28181 29563
rect 28215 29560 28227 29563
rect 28736 29560 28764 29588
rect 28215 29532 28764 29560
rect 28215 29529 28227 29532
rect 28169 29523 28227 29529
rect 29178 29520 29184 29572
rect 29236 29520 29242 29572
rect 30116 29532 30328 29560
rect 2314 29452 2320 29504
rect 2372 29492 2378 29504
rect 2501 29495 2559 29501
rect 2501 29492 2513 29495
rect 2372 29464 2513 29492
rect 2372 29452 2378 29464
rect 2501 29461 2513 29464
rect 2547 29461 2559 29495
rect 2501 29455 2559 29461
rect 13906 29452 13912 29504
rect 13964 29492 13970 29504
rect 15010 29492 15016 29504
rect 13964 29464 15016 29492
rect 13964 29452 13970 29464
rect 15010 29452 15016 29464
rect 15068 29492 15074 29504
rect 28626 29492 28632 29504
rect 15068 29464 28632 29492
rect 15068 29452 15074 29464
rect 28626 29452 28632 29464
rect 28684 29492 28690 29504
rect 30116 29492 30144 29532
rect 28684 29464 30144 29492
rect 28684 29452 28690 29464
rect 30190 29452 30196 29504
rect 30248 29452 30254 29504
rect 30300 29492 30328 29532
rect 30558 29520 30564 29572
rect 30616 29560 30622 29572
rect 33060 29560 33088 29591
rect 57698 29588 57704 29640
rect 57756 29628 57762 29640
rect 57885 29631 57943 29637
rect 57885 29628 57897 29631
rect 57756 29600 57897 29628
rect 57756 29588 57762 29600
rect 57885 29597 57897 29600
rect 57931 29597 57943 29631
rect 57885 29591 57943 29597
rect 30616 29532 33088 29560
rect 30616 29520 30622 29532
rect 32030 29492 32036 29504
rect 30300 29464 32036 29492
rect 32030 29452 32036 29464
rect 32088 29452 32094 29504
rect 32953 29495 33011 29501
rect 32953 29461 32965 29495
rect 32999 29492 33011 29495
rect 39298 29492 39304 29504
rect 32999 29464 39304 29492
rect 32999 29461 33011 29464
rect 32953 29455 33011 29461
rect 39298 29452 39304 29464
rect 39356 29452 39362 29504
rect 1104 29402 58880 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 50294 29402
rect 50346 29350 50358 29402
rect 50410 29350 50422 29402
rect 50474 29350 50486 29402
rect 50538 29350 50550 29402
rect 50602 29350 58880 29402
rect 1104 29328 58880 29350
rect 2406 29288 2412 29300
rect 2240 29260 2412 29288
rect 2240 29229 2268 29260
rect 2406 29248 2412 29260
rect 2464 29248 2470 29300
rect 2610 29291 2668 29297
rect 2610 29257 2622 29291
rect 2656 29288 2668 29291
rect 22278 29288 22284 29300
rect 2656 29260 22284 29288
rect 2656 29257 2668 29260
rect 2610 29251 2668 29257
rect 22278 29248 22284 29260
rect 22336 29248 22342 29300
rect 22462 29248 22468 29300
rect 22520 29248 22526 29300
rect 22738 29248 22744 29300
rect 22796 29248 22802 29300
rect 22922 29248 22928 29300
rect 22980 29288 22986 29300
rect 23382 29288 23388 29300
rect 22980 29260 23388 29288
rect 22980 29248 22986 29260
rect 23382 29248 23388 29260
rect 23440 29288 23446 29300
rect 24305 29291 24363 29297
rect 23440 29260 23520 29288
rect 23440 29248 23446 29260
rect 2225 29223 2283 29229
rect 2225 29189 2237 29223
rect 2271 29189 2283 29223
rect 2225 29183 2283 29189
rect 2314 29180 2320 29232
rect 2372 29180 2378 29232
rect 2041 29155 2099 29161
rect 2041 29121 2053 29155
rect 2087 29152 2099 29155
rect 2130 29152 2136 29164
rect 2087 29124 2136 29152
rect 2087 29121 2099 29124
rect 2041 29115 2099 29121
rect 2130 29112 2136 29124
rect 2188 29112 2194 29164
rect 2414 29155 2472 29161
rect 2414 29121 2426 29155
rect 2460 29152 2472 29155
rect 2682 29152 2688 29164
rect 2460 29124 2688 29152
rect 2460 29121 2472 29124
rect 2414 29115 2472 29121
rect 2424 29084 2452 29115
rect 2682 29112 2688 29124
rect 2740 29112 2746 29164
rect 22097 29155 22155 29161
rect 22097 29121 22109 29155
rect 22143 29152 22155 29155
rect 22738 29152 22744 29164
rect 22143 29124 22744 29152
rect 22143 29121 22155 29124
rect 22097 29115 22155 29121
rect 22738 29112 22744 29124
rect 22796 29112 22802 29164
rect 23198 29112 23204 29164
rect 23256 29112 23262 29164
rect 23492 29161 23520 29260
rect 24305 29257 24317 29291
rect 24351 29288 24363 29291
rect 28902 29288 28908 29300
rect 24351 29260 28908 29288
rect 24351 29257 24363 29260
rect 24305 29251 24363 29257
rect 28902 29248 28908 29260
rect 28960 29248 28966 29300
rect 23566 29180 23572 29232
rect 23624 29220 23630 29232
rect 58342 29220 58348 29232
rect 23624 29192 31616 29220
rect 23624 29180 23630 29192
rect 23477 29155 23535 29161
rect 23477 29121 23489 29155
rect 23523 29121 23535 29155
rect 23477 29115 23535 29121
rect 23750 29112 23756 29164
rect 23808 29112 23814 29164
rect 24489 29155 24547 29161
rect 24489 29121 24501 29155
rect 24535 29121 24547 29155
rect 24489 29115 24547 29121
rect 28445 29155 28503 29161
rect 28445 29121 28457 29155
rect 28491 29121 28503 29155
rect 28445 29115 28503 29121
rect 2148 29056 2452 29084
rect 2148 29028 2176 29056
rect 3234 29044 3240 29096
rect 3292 29084 3298 29096
rect 13906 29084 13912 29096
rect 3292 29056 13912 29084
rect 3292 29044 3298 29056
rect 13906 29044 13912 29056
rect 13964 29044 13970 29096
rect 22189 29087 22247 29093
rect 22189 29053 22201 29087
rect 22235 29053 22247 29087
rect 24504 29084 24532 29115
rect 24946 29084 24952 29096
rect 22189 29047 22247 29053
rect 23400 29056 24952 29084
rect 2130 28976 2136 29028
rect 2188 28976 2194 29028
rect 22204 29016 22232 29047
rect 23400 29016 23428 29056
rect 24946 29044 24952 29056
rect 25004 29044 25010 29096
rect 22204 28988 23428 29016
rect 28169 29019 28227 29025
rect 28169 28985 28181 29019
rect 28215 29016 28227 29019
rect 28460 29016 28488 29115
rect 28626 29112 28632 29164
rect 28684 29112 28690 29164
rect 28718 29112 28724 29164
rect 28776 29112 28782 29164
rect 28810 29112 28816 29164
rect 28868 29112 28874 29164
rect 29638 29112 29644 29164
rect 29696 29112 29702 29164
rect 31018 29112 31024 29164
rect 31076 29152 31082 29164
rect 31588 29161 31616 29192
rect 41386 29192 58348 29220
rect 31297 29155 31355 29161
rect 31297 29152 31309 29155
rect 31076 29124 31309 29152
rect 31076 29112 31082 29124
rect 31297 29121 31309 29124
rect 31343 29121 31355 29155
rect 31297 29115 31355 29121
rect 31573 29155 31631 29161
rect 31573 29121 31585 29155
rect 31619 29121 31631 29155
rect 31573 29115 31631 29121
rect 28644 29084 28672 29112
rect 29917 29087 29975 29093
rect 29917 29084 29929 29087
rect 28644 29056 29929 29084
rect 29917 29053 29929 29056
rect 29963 29053 29975 29087
rect 29917 29047 29975 29053
rect 31481 29087 31539 29093
rect 31481 29053 31493 29087
rect 31527 29084 31539 29087
rect 31662 29084 31668 29096
rect 31527 29056 31668 29084
rect 31527 29053 31539 29056
rect 31481 29047 31539 29053
rect 31662 29044 31668 29056
rect 31720 29044 31726 29096
rect 41386 29016 41414 29192
rect 58342 29180 58348 29192
rect 58400 29180 58406 29232
rect 58066 29112 58072 29164
rect 58124 29112 58130 29164
rect 28215 28988 41414 29016
rect 58253 29019 58311 29025
rect 28215 28985 28227 28988
rect 28169 28979 28227 28985
rect 58253 28985 58265 29019
rect 58299 29016 58311 29019
rect 58434 29016 58440 29028
rect 58299 28988 58440 29016
rect 58299 28985 58311 28988
rect 58253 28979 58311 28985
rect 58434 28976 58440 28988
rect 58492 28976 58498 29028
rect 22281 28951 22339 28957
rect 22281 28917 22293 28951
rect 22327 28948 22339 28951
rect 24486 28948 24492 28960
rect 22327 28920 24492 28948
rect 22327 28917 22339 28920
rect 22281 28911 22339 28917
rect 24486 28908 24492 28920
rect 24544 28908 24550 28960
rect 28994 28908 29000 28960
rect 29052 28908 29058 28960
rect 30926 28908 30932 28960
rect 30984 28948 30990 28960
rect 31297 28951 31355 28957
rect 31297 28948 31309 28951
rect 30984 28920 31309 28948
rect 30984 28908 30990 28920
rect 31297 28917 31309 28920
rect 31343 28917 31355 28951
rect 31297 28911 31355 28917
rect 31754 28908 31760 28960
rect 31812 28908 31818 28960
rect 1104 28858 58880 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 58880 28858
rect 1104 28784 58880 28806
rect 28442 28704 28448 28756
rect 28500 28744 28506 28756
rect 28810 28744 28816 28756
rect 28500 28716 28816 28744
rect 28500 28704 28506 28716
rect 28810 28704 28816 28716
rect 28868 28704 28874 28756
rect 28905 28747 28963 28753
rect 28905 28713 28917 28747
rect 28951 28744 28963 28747
rect 28994 28744 29000 28756
rect 28951 28716 29000 28744
rect 28951 28713 28963 28716
rect 28905 28707 28963 28713
rect 28994 28704 29000 28716
rect 29052 28704 29058 28756
rect 36998 28744 37004 28756
rect 30576 28716 37004 28744
rect 24302 28636 24308 28688
rect 24360 28676 24366 28688
rect 30374 28676 30380 28688
rect 24360 28648 30380 28676
rect 24360 28636 24366 28648
rect 30374 28636 30380 28648
rect 30432 28636 30438 28688
rect 19426 28568 19432 28620
rect 19484 28608 19490 28620
rect 23109 28611 23167 28617
rect 23109 28608 23121 28611
rect 19484 28580 23121 28608
rect 19484 28568 19490 28580
rect 23109 28577 23121 28580
rect 23155 28577 23167 28611
rect 23109 28571 23167 28577
rect 23658 28568 23664 28620
rect 23716 28608 23722 28620
rect 24029 28611 24087 28617
rect 24029 28608 24041 28611
rect 23716 28580 24041 28608
rect 23716 28568 23722 28580
rect 24029 28577 24041 28580
rect 24075 28608 24087 28611
rect 25498 28608 25504 28620
rect 24075 28580 25504 28608
rect 24075 28577 24087 28580
rect 24029 28571 24087 28577
rect 25498 28568 25504 28580
rect 25556 28608 25562 28620
rect 25710 28611 25768 28617
rect 25710 28608 25722 28611
rect 25556 28580 25722 28608
rect 25556 28568 25562 28580
rect 25710 28577 25722 28580
rect 25756 28577 25768 28611
rect 30466 28608 30472 28620
rect 25710 28571 25768 28577
rect 28920 28580 30472 28608
rect 934 28500 940 28552
rect 992 28540 998 28552
rect 1673 28543 1731 28549
rect 1673 28540 1685 28543
rect 992 28512 1685 28540
rect 992 28500 998 28512
rect 1673 28509 1685 28512
rect 1719 28509 1731 28543
rect 1673 28503 1731 28509
rect 23290 28500 23296 28552
rect 23348 28540 23354 28552
rect 23477 28543 23535 28549
rect 23477 28540 23489 28543
rect 23348 28512 23489 28540
rect 23348 28500 23354 28512
rect 23477 28509 23489 28512
rect 23523 28509 23535 28543
rect 23477 28503 23535 28509
rect 23569 28543 23627 28549
rect 23569 28509 23581 28543
rect 23615 28540 23627 28543
rect 23750 28540 23756 28552
rect 23615 28512 23756 28540
rect 23615 28509 23627 28512
rect 23569 28503 23627 28509
rect 23017 28475 23075 28481
rect 23017 28441 23029 28475
rect 23063 28472 23075 28475
rect 23382 28472 23388 28484
rect 23063 28444 23388 28472
rect 23063 28441 23075 28444
rect 23017 28435 23075 28441
rect 23382 28432 23388 28444
rect 23440 28432 23446 28484
rect 23492 28472 23520 28503
rect 23750 28500 23756 28512
rect 23808 28500 23814 28552
rect 24578 28500 24584 28552
rect 24636 28540 24642 28552
rect 25225 28543 25283 28549
rect 25225 28540 25237 28543
rect 24636 28512 25237 28540
rect 24636 28500 24642 28512
rect 25225 28509 25237 28512
rect 25271 28540 25283 28543
rect 25866 28540 25872 28552
rect 25271 28512 25872 28540
rect 25271 28509 25283 28512
rect 25225 28503 25283 28509
rect 25866 28500 25872 28512
rect 25924 28500 25930 28552
rect 28534 28500 28540 28552
rect 28592 28540 28598 28552
rect 28629 28543 28687 28549
rect 28629 28540 28641 28543
rect 28592 28512 28641 28540
rect 28592 28500 28598 28512
rect 28629 28509 28641 28512
rect 28675 28509 28687 28543
rect 28629 28503 28687 28509
rect 28810 28500 28816 28552
rect 28868 28500 28874 28552
rect 28920 28549 28948 28580
rect 30466 28568 30472 28580
rect 30524 28568 30530 28620
rect 28905 28543 28963 28549
rect 28905 28509 28917 28543
rect 28951 28509 28963 28543
rect 28905 28503 28963 28509
rect 29825 28543 29883 28549
rect 29825 28509 29837 28543
rect 29871 28509 29883 28543
rect 30576 28540 30604 28716
rect 36998 28704 37004 28716
rect 37056 28704 37062 28756
rect 31754 28676 31760 28688
rect 31588 28648 31760 28676
rect 31588 28549 31616 28648
rect 31754 28636 31760 28648
rect 31812 28636 31818 28688
rect 49053 28679 49111 28685
rect 49053 28676 49065 28679
rect 42444 28648 49065 28676
rect 29825 28503 29883 28509
rect 30208 28512 30604 28540
rect 31573 28543 31631 28549
rect 25593 28475 25651 28481
rect 25593 28472 25605 28475
rect 23492 28444 25605 28472
rect 25593 28441 25605 28444
rect 25639 28441 25651 28475
rect 25593 28435 25651 28441
rect 28718 28432 28724 28484
rect 28776 28472 28782 28484
rect 29840 28472 29868 28503
rect 28776 28444 29868 28472
rect 28776 28432 28782 28444
rect 30006 28432 30012 28484
rect 30064 28472 30070 28484
rect 30208 28481 30236 28512
rect 31573 28509 31585 28543
rect 31619 28509 31631 28543
rect 31573 28503 31631 28509
rect 31757 28543 31815 28549
rect 31757 28509 31769 28543
rect 31803 28540 31815 28543
rect 37918 28540 37924 28552
rect 31803 28512 37924 28540
rect 31803 28509 31815 28512
rect 31757 28503 31815 28509
rect 37918 28500 37924 28512
rect 37976 28500 37982 28552
rect 42150 28500 42156 28552
rect 42208 28540 42214 28552
rect 42444 28549 42472 28648
rect 49053 28645 49065 28648
rect 49099 28645 49111 28679
rect 49053 28639 49111 28645
rect 52178 28608 52184 28620
rect 48792 28580 52184 28608
rect 42245 28543 42303 28549
rect 42245 28540 42257 28543
rect 42208 28512 42257 28540
rect 42208 28500 42214 28512
rect 42245 28509 42257 28512
rect 42291 28509 42303 28543
rect 42245 28503 42303 28509
rect 42429 28543 42487 28549
rect 42429 28509 42441 28543
rect 42475 28509 42487 28543
rect 42429 28503 42487 28509
rect 48409 28543 48467 28549
rect 48409 28509 48421 28543
rect 48455 28509 48467 28543
rect 48409 28503 48467 28509
rect 48557 28543 48615 28549
rect 48557 28509 48569 28543
rect 48603 28540 48615 28543
rect 48792 28540 48820 28580
rect 52178 28568 52184 28580
rect 52236 28568 52242 28620
rect 58158 28568 58164 28620
rect 58216 28568 58222 28620
rect 48603 28512 48820 28540
rect 48915 28543 48973 28549
rect 48603 28509 48615 28512
rect 48557 28503 48615 28509
rect 48915 28509 48927 28543
rect 48961 28540 48973 28543
rect 49234 28540 49240 28552
rect 48961 28512 49240 28540
rect 48961 28509 48973 28512
rect 48915 28503 48973 28509
rect 30193 28475 30251 28481
rect 30193 28472 30205 28475
rect 30064 28444 30205 28472
rect 30064 28432 30070 28444
rect 30193 28441 30205 28444
rect 30239 28441 30251 28475
rect 30193 28435 30251 28441
rect 30282 28432 30288 28484
rect 30340 28472 30346 28484
rect 41690 28472 41696 28484
rect 30340 28444 41696 28472
rect 30340 28432 30346 28444
rect 41690 28432 41696 28444
rect 41748 28472 41754 28484
rect 42058 28472 42064 28484
rect 41748 28444 42064 28472
rect 41748 28432 41754 28444
rect 42058 28432 42064 28444
rect 42116 28432 42122 28484
rect 1765 28407 1823 28413
rect 1765 28373 1777 28407
rect 1811 28404 1823 28407
rect 13814 28404 13820 28416
rect 1811 28376 13820 28404
rect 1811 28373 1823 28376
rect 1765 28367 1823 28373
rect 13814 28364 13820 28376
rect 13872 28364 13878 28416
rect 25406 28364 25412 28416
rect 25464 28404 25470 28416
rect 25501 28407 25559 28413
rect 25501 28404 25513 28407
rect 25464 28376 25513 28404
rect 25464 28364 25470 28376
rect 25501 28373 25513 28376
rect 25547 28373 25559 28407
rect 25501 28367 25559 28373
rect 25869 28407 25927 28413
rect 25869 28373 25881 28407
rect 25915 28404 25927 28407
rect 27982 28404 27988 28416
rect 25915 28376 27988 28404
rect 25915 28373 25927 28376
rect 25869 28367 25927 28373
rect 27982 28364 27988 28376
rect 28040 28364 28046 28416
rect 29089 28407 29147 28413
rect 29089 28373 29101 28407
rect 29135 28404 29147 28407
rect 31570 28404 31576 28416
rect 29135 28376 31576 28404
rect 29135 28373 29147 28376
rect 29089 28367 29147 28373
rect 31570 28364 31576 28376
rect 31628 28364 31634 28416
rect 31849 28407 31907 28413
rect 31849 28373 31861 28407
rect 31895 28404 31907 28407
rect 31938 28404 31944 28416
rect 31895 28376 31944 28404
rect 31895 28373 31907 28376
rect 31849 28367 31907 28373
rect 31938 28364 31944 28376
rect 31996 28364 32002 28416
rect 41230 28364 41236 28416
rect 41288 28404 41294 28416
rect 42521 28407 42579 28413
rect 42521 28404 42533 28407
rect 41288 28376 42533 28404
rect 41288 28364 41294 28376
rect 42521 28373 42533 28376
rect 42567 28373 42579 28407
rect 48424 28404 48452 28503
rect 49234 28500 49240 28512
rect 49292 28500 49298 28552
rect 56594 28500 56600 28552
rect 56652 28540 56658 28552
rect 57885 28543 57943 28549
rect 57885 28540 57897 28543
rect 56652 28512 57897 28540
rect 56652 28500 56658 28512
rect 57885 28509 57897 28512
rect 57931 28509 57943 28543
rect 57885 28503 57943 28509
rect 48682 28432 48688 28484
rect 48740 28432 48746 28484
rect 48777 28475 48835 28481
rect 48777 28441 48789 28475
rect 48823 28472 48835 28475
rect 50706 28472 50712 28484
rect 48823 28444 50712 28472
rect 48823 28441 48835 28444
rect 48777 28435 48835 28441
rect 50706 28432 50712 28444
rect 50764 28432 50770 28484
rect 48866 28404 48872 28416
rect 48424 28376 48872 28404
rect 42521 28367 42579 28373
rect 48866 28364 48872 28376
rect 48924 28364 48930 28416
rect 1104 28314 58880 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 50294 28314
rect 50346 28262 50358 28314
rect 50410 28262 50422 28314
rect 50474 28262 50486 28314
rect 50538 28262 50550 28314
rect 50602 28262 58880 28314
rect 1104 28240 58880 28262
rect 18966 28160 18972 28212
rect 19024 28200 19030 28212
rect 22278 28200 22284 28212
rect 19024 28172 22284 28200
rect 19024 28160 19030 28172
rect 22278 28160 22284 28172
rect 22336 28160 22342 28212
rect 22462 28160 22468 28212
rect 22520 28200 22526 28212
rect 24302 28200 24308 28212
rect 22520 28172 24308 28200
rect 22520 28160 22526 28172
rect 24302 28160 24308 28172
rect 24360 28160 24366 28212
rect 25593 28203 25651 28209
rect 25593 28169 25605 28203
rect 25639 28200 25651 28203
rect 28718 28200 28724 28212
rect 25639 28172 28724 28200
rect 25639 28169 25651 28172
rect 25593 28163 25651 28169
rect 28718 28160 28724 28172
rect 28776 28160 28782 28212
rect 28810 28160 28816 28212
rect 28868 28200 28874 28212
rect 29089 28203 29147 28209
rect 29089 28200 29101 28203
rect 28868 28172 29101 28200
rect 28868 28160 28874 28172
rect 29089 28169 29101 28172
rect 29135 28169 29147 28203
rect 29089 28163 29147 28169
rect 30098 28160 30104 28212
rect 30156 28200 30162 28212
rect 31389 28203 31447 28209
rect 30156 28172 31248 28200
rect 30156 28160 30162 28172
rect 934 28092 940 28144
rect 992 28132 998 28144
rect 1673 28135 1731 28141
rect 1673 28132 1685 28135
rect 992 28104 1685 28132
rect 992 28092 998 28104
rect 1673 28101 1685 28104
rect 1719 28101 1731 28135
rect 1673 28095 1731 28101
rect 15378 28092 15384 28144
rect 15436 28132 15442 28144
rect 31113 28135 31171 28141
rect 31113 28132 31125 28135
rect 15436 28104 19334 28132
rect 15436 28092 15442 28104
rect 19306 28064 19334 28104
rect 22112 28104 28856 28132
rect 22112 28064 22140 28104
rect 19306 28036 22140 28064
rect 23201 28067 23259 28073
rect 23201 28033 23213 28067
rect 23247 28064 23259 28067
rect 23290 28064 23296 28076
rect 23247 28036 23296 28064
rect 23247 28033 23259 28036
rect 23201 28027 23259 28033
rect 23290 28024 23296 28036
rect 23348 28024 23354 28076
rect 23382 28024 23388 28076
rect 23440 28024 23446 28076
rect 23750 28024 23756 28076
rect 23808 28024 23814 28076
rect 24486 28024 24492 28076
rect 24544 28024 24550 28076
rect 24946 28024 24952 28076
rect 25004 28064 25010 28076
rect 25041 28067 25099 28073
rect 25041 28064 25053 28067
rect 25004 28036 25053 28064
rect 25004 28024 25010 28036
rect 25041 28033 25053 28036
rect 25087 28033 25099 28067
rect 25041 28027 25099 28033
rect 25498 28024 25504 28076
rect 25556 28024 25562 28076
rect 25590 28024 25596 28076
rect 25648 28024 25654 28076
rect 25866 28024 25872 28076
rect 25924 28064 25930 28076
rect 27157 28067 27215 28073
rect 27157 28064 27169 28067
rect 25924 28036 27169 28064
rect 25924 28024 25930 28036
rect 27157 28033 27169 28036
rect 27203 28033 27215 28067
rect 27157 28027 27215 28033
rect 28534 28024 28540 28076
rect 28592 28024 28598 28076
rect 28828 28073 28856 28104
rect 29196 28104 31125 28132
rect 28721 28067 28779 28073
rect 28721 28033 28733 28067
rect 28767 28033 28779 28067
rect 28721 28027 28779 28033
rect 28813 28067 28871 28073
rect 28813 28033 28825 28067
rect 28859 28033 28871 28067
rect 28813 28027 28871 28033
rect 22278 27956 22284 28008
rect 22336 27996 22342 28008
rect 22336 27968 26188 27996
rect 22336 27956 22342 27968
rect 25038 27888 25044 27940
rect 25096 27928 25102 27940
rect 26050 27928 26056 27940
rect 25096 27900 26056 27928
rect 25096 27888 25102 27900
rect 26050 27888 26056 27900
rect 26108 27888 26114 27940
rect 26160 27928 26188 27968
rect 27338 27956 27344 28008
rect 27396 27956 27402 28008
rect 27522 27956 27528 28008
rect 27580 27996 27586 28008
rect 28736 27996 28764 28027
rect 28902 28024 28908 28076
rect 28960 28024 28966 28076
rect 28994 27996 29000 28008
rect 27580 27968 29000 27996
rect 27580 27956 27586 27968
rect 28994 27956 29000 27968
rect 29052 27956 29058 28008
rect 29196 27928 29224 28104
rect 31113 28101 31125 28104
rect 31159 28101 31171 28135
rect 31113 28095 31171 28101
rect 29362 28024 29368 28076
rect 29420 28064 29426 28076
rect 29641 28067 29699 28073
rect 29641 28064 29653 28067
rect 29420 28036 29653 28064
rect 29420 28024 29426 28036
rect 29641 28033 29653 28036
rect 29687 28064 29699 28067
rect 30006 28064 30012 28076
rect 29687 28036 30012 28064
rect 29687 28033 29699 28036
rect 29641 28027 29699 28033
rect 30006 28024 30012 28036
rect 30064 28024 30070 28076
rect 30466 28024 30472 28076
rect 30524 28064 30530 28076
rect 31220 28073 31248 28172
rect 31389 28169 31401 28203
rect 31435 28200 31447 28203
rect 31478 28200 31484 28212
rect 31435 28172 31484 28200
rect 31435 28169 31447 28172
rect 31389 28163 31447 28169
rect 31478 28160 31484 28172
rect 31536 28160 31542 28212
rect 48314 28132 48320 28144
rect 31588 28104 48320 28132
rect 30745 28067 30803 28073
rect 30745 28064 30757 28067
rect 30524 28036 30757 28064
rect 30524 28024 30530 28036
rect 30745 28033 30757 28036
rect 30791 28033 30803 28067
rect 30745 28027 30803 28033
rect 30838 28067 30896 28073
rect 30838 28033 30850 28067
rect 30884 28033 30896 28067
rect 30838 28027 30896 28033
rect 31021 28067 31079 28073
rect 31021 28033 31033 28067
rect 31067 28033 31079 28067
rect 31021 28027 31079 28033
rect 31210 28067 31268 28073
rect 31210 28033 31222 28067
rect 31256 28033 31268 28067
rect 31210 28027 31268 28033
rect 29917 27999 29975 28005
rect 29917 27996 29929 27999
rect 26160 27900 29224 27928
rect 29564 27968 29929 27996
rect 1765 27863 1823 27869
rect 1765 27829 1777 27863
rect 1811 27860 1823 27863
rect 28626 27860 28632 27872
rect 1811 27832 28632 27860
rect 1811 27829 1823 27832
rect 1765 27823 1823 27829
rect 28626 27820 28632 27832
rect 28684 27820 28690 27872
rect 28994 27820 29000 27872
rect 29052 27860 29058 27872
rect 29564 27860 29592 27968
rect 29917 27965 29929 27968
rect 29963 27996 29975 27999
rect 30282 27996 30288 28008
rect 29963 27968 30288 27996
rect 29963 27965 29975 27968
rect 29917 27959 29975 27965
rect 30282 27956 30288 27968
rect 30340 27956 30346 28008
rect 30852 27928 30880 28027
rect 31036 27996 31064 28027
rect 31110 27996 31116 28008
rect 31036 27968 31116 27996
rect 31110 27956 31116 27968
rect 31168 27996 31174 28008
rect 31588 27996 31616 28104
rect 48314 28092 48320 28104
rect 48372 28092 48378 28144
rect 58710 28132 58716 28144
rect 51046 28104 58716 28132
rect 51046 28064 51074 28104
rect 58710 28092 58716 28104
rect 58768 28092 58774 28144
rect 31168 27968 31616 27996
rect 38626 28036 51074 28064
rect 31168 27956 31174 27968
rect 38626 27928 38654 28036
rect 58066 28024 58072 28076
rect 58124 28024 58130 28076
rect 30852 27900 38654 27928
rect 29052 27832 29592 27860
rect 29052 27820 29058 27832
rect 42610 27820 42616 27872
rect 42668 27860 42674 27872
rect 58253 27863 58311 27869
rect 58253 27860 58265 27863
rect 42668 27832 58265 27860
rect 42668 27820 42674 27832
rect 58253 27829 58265 27832
rect 58299 27829 58311 27863
rect 58253 27823 58311 27829
rect 1104 27770 58880 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 58880 27770
rect 1104 27696 58880 27718
rect 22370 27616 22376 27668
rect 22428 27656 22434 27668
rect 28442 27656 28448 27668
rect 22428 27628 28448 27656
rect 22428 27616 22434 27628
rect 23658 27548 23664 27600
rect 23716 27548 23722 27600
rect 26326 27548 26332 27600
rect 26384 27588 26390 27600
rect 27338 27588 27344 27600
rect 26384 27560 27344 27588
rect 26384 27548 26390 27560
rect 23014 27480 23020 27532
rect 23072 27480 23078 27532
rect 23676 27520 23704 27548
rect 23492 27492 23704 27520
rect 934 27412 940 27464
rect 992 27452 998 27464
rect 1673 27455 1731 27461
rect 1673 27452 1685 27455
rect 992 27424 1685 27452
rect 992 27412 998 27424
rect 1673 27421 1685 27424
rect 1719 27421 1731 27455
rect 1673 27415 1731 27421
rect 22094 27412 22100 27464
rect 22152 27452 22158 27464
rect 23032 27452 23060 27480
rect 23109 27455 23167 27461
rect 23109 27452 23121 27455
rect 22152 27424 23121 27452
rect 22152 27412 22158 27424
rect 23109 27421 23121 27424
rect 23155 27421 23167 27455
rect 23109 27415 23167 27421
rect 23290 27412 23296 27464
rect 23348 27452 23354 27464
rect 23492 27461 23520 27492
rect 23477 27455 23535 27461
rect 23477 27452 23489 27455
rect 23348 27424 23489 27452
rect 23348 27412 23354 27424
rect 23477 27421 23489 27424
rect 23523 27421 23535 27455
rect 23477 27415 23535 27421
rect 23566 27412 23572 27464
rect 23624 27412 23630 27464
rect 23658 27412 23664 27464
rect 23716 27452 23722 27464
rect 24029 27455 24087 27461
rect 24029 27452 24041 27455
rect 23716 27424 24041 27452
rect 23716 27412 23722 27424
rect 24029 27421 24041 27424
rect 24075 27452 24087 27455
rect 24946 27452 24952 27464
rect 24075 27424 24952 27452
rect 24075 27421 24087 27424
rect 24029 27415 24087 27421
rect 24946 27412 24952 27424
rect 25004 27452 25010 27464
rect 25222 27452 25228 27464
rect 25004 27424 25228 27452
rect 25004 27412 25010 27424
rect 25222 27412 25228 27424
rect 25280 27412 25286 27464
rect 25406 27412 25412 27464
rect 25464 27412 25470 27464
rect 25498 27412 25504 27464
rect 25556 27452 25562 27464
rect 26605 27455 26663 27461
rect 26605 27452 26617 27455
rect 25556 27424 26617 27452
rect 25556 27412 25562 27424
rect 26605 27421 26617 27424
rect 26651 27421 26663 27455
rect 26712 27452 26740 27560
rect 27338 27548 27344 27560
rect 27396 27548 27402 27600
rect 26789 27455 26847 27461
rect 26789 27452 26801 27455
rect 26712 27424 26801 27452
rect 26605 27415 26663 27421
rect 26789 27421 26801 27424
rect 26835 27421 26847 27455
rect 26789 27415 26847 27421
rect 26970 27412 26976 27464
rect 27028 27412 27034 27464
rect 27062 27412 27068 27464
rect 27120 27412 27126 27464
rect 27433 27455 27491 27461
rect 27433 27421 27445 27455
rect 27479 27452 27491 27455
rect 27706 27452 27712 27464
rect 27479 27424 27712 27452
rect 27479 27421 27491 27424
rect 27433 27415 27491 27421
rect 27706 27412 27712 27424
rect 27764 27412 27770 27464
rect 28175 27461 28203 27628
rect 28442 27616 28448 27628
rect 28500 27656 28506 27668
rect 30466 27656 30472 27668
rect 28500 27628 28994 27656
rect 28500 27616 28506 27628
rect 28966 27588 28994 27628
rect 30300 27628 30472 27656
rect 30098 27588 30104 27600
rect 28966 27560 30104 27588
rect 30098 27548 30104 27560
rect 30156 27548 30162 27600
rect 30300 27597 30328 27628
rect 30466 27616 30472 27628
rect 30524 27616 30530 27668
rect 33134 27656 33140 27668
rect 30576 27628 33140 27656
rect 30285 27591 30343 27597
rect 30285 27557 30297 27591
rect 30331 27557 30343 27591
rect 30285 27551 30343 27557
rect 30374 27548 30380 27600
rect 30432 27588 30438 27600
rect 30576 27588 30604 27628
rect 33134 27616 33140 27628
rect 33192 27656 33198 27668
rect 34146 27656 34152 27668
rect 33192 27628 34152 27656
rect 33192 27616 33198 27628
rect 34146 27616 34152 27628
rect 34204 27616 34210 27668
rect 34256 27628 34468 27656
rect 30432 27560 30604 27588
rect 30432 27548 30438 27560
rect 31662 27548 31668 27600
rect 31720 27588 31726 27600
rect 32493 27591 32551 27597
rect 32493 27588 32505 27591
rect 31720 27560 32505 27588
rect 31720 27548 31726 27560
rect 32493 27557 32505 27560
rect 32539 27557 32551 27591
rect 34256 27588 34284 27628
rect 32493 27551 32551 27557
rect 33612 27560 34284 27588
rect 34440 27588 34468 27628
rect 34440 27560 41414 27588
rect 28626 27480 28632 27532
rect 28684 27520 28690 27532
rect 33612 27520 33640 27560
rect 28684 27492 33640 27520
rect 28684 27480 28690 27492
rect 33778 27480 33784 27532
rect 33836 27480 33842 27532
rect 41386 27520 41414 27560
rect 45462 27548 45468 27600
rect 45520 27588 45526 27600
rect 49605 27591 49663 27597
rect 49605 27588 49617 27591
rect 45520 27560 49617 27588
rect 45520 27548 45526 27560
rect 49605 27557 49617 27560
rect 49651 27557 49663 27591
rect 49605 27551 49663 27557
rect 48958 27520 48964 27532
rect 41386 27492 48964 27520
rect 48958 27480 48964 27492
rect 49016 27480 49022 27532
rect 51350 27520 51356 27532
rect 49068 27492 51356 27520
rect 27985 27455 28043 27461
rect 27985 27452 27997 27455
rect 27816 27424 27997 27452
rect 23017 27387 23075 27393
rect 23017 27353 23029 27387
rect 23063 27353 23075 27387
rect 25590 27384 25596 27396
rect 23017 27347 23075 27353
rect 24872 27356 25596 27384
rect 1765 27319 1823 27325
rect 1765 27285 1777 27319
rect 1811 27316 1823 27319
rect 18966 27316 18972 27328
rect 1811 27288 18972 27316
rect 1811 27285 1823 27288
rect 1765 27279 1823 27285
rect 18966 27276 18972 27288
rect 19024 27276 19030 27328
rect 23032 27316 23060 27347
rect 24872 27328 24900 27356
rect 25590 27344 25596 27356
rect 25648 27384 25654 27396
rect 25777 27387 25835 27393
rect 25777 27384 25789 27387
rect 25648 27356 25789 27384
rect 25648 27344 25654 27356
rect 25777 27353 25789 27356
rect 25823 27384 25835 27387
rect 26234 27384 26240 27396
rect 25823 27356 26240 27384
rect 25823 27353 25835 27356
rect 25777 27347 25835 27353
rect 26234 27344 26240 27356
rect 26292 27384 26298 27396
rect 26697 27387 26755 27393
rect 26697 27384 26709 27387
rect 26292 27356 26709 27384
rect 26292 27344 26298 27356
rect 26697 27353 26709 27356
rect 26743 27353 26755 27387
rect 26697 27347 26755 27353
rect 23750 27316 23756 27328
rect 23032 27288 23756 27316
rect 23750 27276 23756 27288
rect 23808 27316 23814 27328
rect 24854 27316 24860 27328
rect 23808 27288 24860 27316
rect 23808 27276 23814 27288
rect 24854 27276 24860 27288
rect 24912 27276 24918 27328
rect 26050 27276 26056 27328
rect 26108 27316 26114 27328
rect 26326 27316 26332 27328
rect 26108 27288 26332 27316
rect 26108 27276 26114 27288
rect 26326 27276 26332 27288
rect 26384 27276 26390 27328
rect 26421 27319 26479 27325
rect 26421 27285 26433 27319
rect 26467 27316 26479 27319
rect 26510 27316 26516 27328
rect 26467 27288 26516 27316
rect 26467 27285 26479 27288
rect 26421 27279 26479 27285
rect 26510 27276 26516 27288
rect 26568 27276 26574 27328
rect 26602 27276 26608 27328
rect 26660 27316 26666 27328
rect 27816 27316 27844 27424
rect 27985 27421 27997 27424
rect 28031 27421 28043 27455
rect 27985 27415 28043 27421
rect 28123 27455 28203 27461
rect 28123 27421 28135 27455
rect 28169 27424 28203 27455
rect 28169 27421 28181 27424
rect 28123 27415 28181 27421
rect 28442 27412 28448 27464
rect 28500 27452 28506 27464
rect 30469 27455 30527 27461
rect 30469 27452 30481 27455
rect 28500 27424 30481 27452
rect 28500 27412 28506 27424
rect 30469 27421 30481 27424
rect 30515 27421 30527 27455
rect 30469 27415 30527 27421
rect 30650 27412 30656 27464
rect 30708 27412 30714 27464
rect 30837 27455 30895 27461
rect 30837 27421 30849 27455
rect 30883 27452 30895 27455
rect 30926 27452 30932 27464
rect 30883 27424 30932 27452
rect 30883 27421 30895 27424
rect 30837 27415 30895 27421
rect 30926 27412 30932 27424
rect 30984 27412 30990 27464
rect 32214 27412 32220 27464
rect 32272 27412 32278 27464
rect 32306 27412 32312 27464
rect 32364 27412 32370 27464
rect 32953 27455 33011 27461
rect 32953 27421 32965 27455
rect 32999 27421 33011 27455
rect 32953 27415 33011 27421
rect 27890 27344 27896 27396
rect 27948 27344 27954 27396
rect 32968 27384 32996 27415
rect 33502 27412 33508 27464
rect 33560 27412 33566 27464
rect 33962 27412 33968 27464
rect 34020 27412 34026 27464
rect 49068 27461 49096 27492
rect 51350 27480 51356 27492
rect 51408 27480 51414 27532
rect 58161 27523 58219 27529
rect 58161 27489 58173 27523
rect 58207 27520 58219 27523
rect 58986 27520 58992 27532
rect 58207 27492 58992 27520
rect 58207 27489 58219 27492
rect 58161 27483 58219 27489
rect 58986 27480 58992 27492
rect 59044 27480 59050 27532
rect 49053 27455 49111 27461
rect 49053 27421 49065 27455
rect 49099 27421 49111 27455
rect 49053 27415 49111 27421
rect 49418 27412 49424 27464
rect 49476 27461 49482 27464
rect 49476 27452 49484 27461
rect 49476 27424 49521 27452
rect 49476 27415 49484 27424
rect 49476 27412 49482 27415
rect 56870 27412 56876 27464
rect 56928 27452 56934 27464
rect 57885 27455 57943 27461
rect 57885 27452 57897 27455
rect 56928 27424 57897 27452
rect 56928 27412 56934 27424
rect 57885 27421 57897 27424
rect 57931 27421 57943 27455
rect 57885 27415 57943 27421
rect 35342 27384 35348 27396
rect 28184 27356 35348 27384
rect 28184 27328 28212 27356
rect 35342 27344 35348 27356
rect 35400 27344 35406 27396
rect 48682 27344 48688 27396
rect 48740 27384 48746 27396
rect 49237 27387 49295 27393
rect 49237 27384 49249 27387
rect 48740 27356 49249 27384
rect 48740 27344 48746 27356
rect 49237 27353 49249 27356
rect 49283 27353 49295 27387
rect 49237 27347 49295 27353
rect 49329 27387 49387 27393
rect 49329 27353 49341 27387
rect 49375 27384 49387 27387
rect 50890 27384 50896 27396
rect 49375 27356 50896 27384
rect 49375 27353 49387 27356
rect 49329 27347 49387 27353
rect 50890 27344 50896 27356
rect 50948 27344 50954 27396
rect 26660 27288 27844 27316
rect 26660 27276 26666 27288
rect 28166 27276 28172 27328
rect 28224 27276 28230 27328
rect 28261 27319 28319 27325
rect 28261 27285 28273 27319
rect 28307 27316 28319 27319
rect 28442 27316 28448 27328
rect 28307 27288 28448 27316
rect 28307 27285 28319 27288
rect 28261 27279 28319 27285
rect 28442 27276 28448 27288
rect 28500 27276 28506 27328
rect 33594 27276 33600 27328
rect 33652 27316 33658 27328
rect 33714 27319 33772 27325
rect 33714 27316 33726 27319
rect 33652 27288 33726 27316
rect 33652 27276 33658 27288
rect 33714 27285 33726 27288
rect 33760 27285 33772 27319
rect 33714 27279 33772 27285
rect 1104 27226 58880 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 50294 27226
rect 50346 27174 50358 27226
rect 50410 27174 50422 27226
rect 50474 27174 50486 27226
rect 50538 27174 50550 27226
rect 50602 27174 58880 27226
rect 1104 27152 58880 27174
rect 23566 27072 23572 27124
rect 23624 27112 23630 27124
rect 25038 27112 25044 27124
rect 23624 27084 25044 27112
rect 23624 27072 23630 27084
rect 25038 27072 25044 27084
rect 25096 27112 25102 27124
rect 25314 27112 25320 27124
rect 25096 27084 25320 27112
rect 25096 27072 25102 27084
rect 25314 27072 25320 27084
rect 25372 27072 25378 27124
rect 26050 27072 26056 27124
rect 26108 27072 26114 27124
rect 26234 27072 26240 27124
rect 26292 27072 26298 27124
rect 26326 27072 26332 27124
rect 26384 27072 26390 27124
rect 26418 27072 26424 27124
rect 26476 27112 26482 27124
rect 30650 27112 30656 27124
rect 26476 27084 30656 27112
rect 26476 27072 26482 27084
rect 30650 27072 30656 27084
rect 30708 27072 30714 27124
rect 31018 27072 31024 27124
rect 31076 27072 31082 27124
rect 59170 27112 59176 27124
rect 41386 27084 59176 27112
rect 934 27004 940 27056
rect 992 27044 998 27056
rect 1673 27047 1731 27053
rect 1673 27044 1685 27047
rect 992 27016 1685 27044
rect 992 27004 998 27016
rect 1673 27013 1685 27016
rect 1719 27013 1731 27047
rect 1673 27007 1731 27013
rect 1854 27004 1860 27056
rect 1912 27044 1918 27056
rect 25498 27044 25504 27056
rect 1912 27016 25504 27044
rect 1912 27004 1918 27016
rect 25498 27004 25504 27016
rect 25556 27004 25562 27056
rect 26142 27004 26148 27056
rect 26200 27004 26206 27056
rect 26513 27047 26571 27053
rect 26513 27013 26525 27047
rect 26559 27044 26571 27047
rect 26970 27044 26976 27056
rect 26559 27016 26976 27044
rect 26559 27013 26571 27016
rect 26513 27007 26571 27013
rect 1026 26936 1032 26988
rect 1084 26976 1090 26988
rect 2409 26979 2467 26985
rect 2409 26976 2421 26979
rect 1084 26948 2421 26976
rect 1084 26936 1090 26948
rect 2409 26945 2421 26948
rect 2455 26945 2467 26979
rect 2409 26939 2467 26945
rect 23014 26936 23020 26988
rect 23072 26936 23078 26988
rect 23382 26936 23388 26988
rect 23440 26936 23446 26988
rect 23477 26979 23535 26985
rect 23477 26945 23489 26979
rect 23523 26976 23535 26979
rect 24578 26976 24584 26988
rect 23523 26948 24584 26976
rect 23523 26945 23535 26948
rect 23477 26939 23535 26945
rect 24578 26936 24584 26948
rect 24636 26936 24642 26988
rect 24854 26936 24860 26988
rect 24912 26936 24918 26988
rect 25038 26936 25044 26988
rect 25096 26936 25102 26988
rect 25130 26936 25136 26988
rect 25188 26936 25194 26988
rect 25222 26936 25228 26988
rect 25280 26976 25286 26988
rect 25280 26948 25325 26976
rect 25280 26936 25286 26948
rect 22922 26868 22928 26920
rect 22980 26868 22986 26920
rect 23937 26911 23995 26917
rect 23937 26877 23949 26911
rect 23983 26908 23995 26911
rect 24486 26908 24492 26920
rect 23983 26880 24492 26908
rect 23983 26877 23995 26880
rect 23937 26871 23995 26877
rect 24486 26868 24492 26880
rect 24544 26908 24550 26920
rect 24946 26908 24952 26920
rect 24544 26880 24952 26908
rect 24544 26868 24550 26880
rect 24946 26868 24952 26880
rect 25004 26868 25010 26920
rect 26602 26908 26608 26920
rect 25056 26880 26608 26908
rect 1857 26843 1915 26849
rect 1857 26809 1869 26843
rect 1903 26840 1915 26843
rect 25056 26840 25084 26880
rect 26602 26868 26608 26880
rect 26660 26868 26666 26920
rect 1903 26812 25084 26840
rect 25501 26843 25559 26849
rect 1903 26809 1915 26812
rect 1857 26803 1915 26809
rect 25501 26809 25513 26843
rect 25547 26840 25559 26843
rect 25590 26840 25596 26852
rect 25547 26812 25596 26840
rect 25547 26809 25559 26812
rect 25501 26803 25559 26809
rect 25590 26800 25596 26812
rect 25648 26840 25654 26852
rect 26712 26840 26740 27016
rect 26970 27004 26976 27016
rect 27028 27004 27034 27056
rect 27706 27004 27712 27056
rect 27764 27044 27770 27056
rect 30558 27044 30564 27056
rect 27764 27016 30564 27044
rect 27764 27004 27770 27016
rect 30558 27004 30564 27016
rect 30616 27004 30622 27056
rect 32030 27004 32036 27056
rect 32088 27044 32094 27056
rect 41386 27044 41414 27084
rect 59170 27072 59176 27084
rect 59228 27072 59234 27124
rect 32088 27016 41414 27044
rect 32088 27004 32094 27016
rect 58158 27004 58164 27056
rect 58216 27004 58222 27056
rect 27982 26936 27988 26988
rect 28040 26936 28046 26988
rect 28537 26979 28595 26985
rect 28537 26945 28549 26979
rect 28583 26976 28595 26979
rect 29086 26976 29092 26988
rect 28583 26948 29092 26976
rect 28583 26945 28595 26948
rect 28537 26939 28595 26945
rect 29086 26936 29092 26948
rect 29144 26936 29150 26988
rect 30469 26979 30527 26985
rect 30469 26945 30481 26979
rect 30515 26945 30527 26979
rect 30469 26939 30527 26945
rect 30484 26908 30512 26939
rect 30650 26936 30656 26988
rect 30708 26936 30714 26988
rect 30742 26936 30748 26988
rect 30800 26936 30806 26988
rect 30837 26979 30895 26985
rect 30837 26945 30849 26979
rect 30883 26976 30895 26979
rect 31386 26976 31392 26988
rect 30883 26948 31392 26976
rect 30883 26945 30895 26948
rect 30837 26939 30895 26945
rect 31386 26936 31392 26948
rect 31444 26936 31450 26988
rect 32766 26936 32772 26988
rect 32824 26936 32830 26988
rect 32950 26936 32956 26988
rect 33008 26936 33014 26988
rect 33134 26936 33140 26988
rect 33192 26936 33198 26988
rect 42794 26936 42800 26988
rect 42852 26976 42858 26988
rect 43162 26976 43168 26988
rect 42852 26948 43168 26976
rect 42852 26936 42858 26948
rect 43162 26936 43168 26948
rect 43220 26936 43226 26988
rect 30926 26908 30932 26920
rect 30484 26880 30932 26908
rect 30926 26868 30932 26880
rect 30984 26908 30990 26920
rect 31662 26908 31668 26920
rect 30984 26880 31668 26908
rect 30984 26868 30990 26880
rect 31662 26868 31668 26880
rect 31720 26868 31726 26920
rect 34146 26868 34152 26920
rect 34204 26908 34210 26920
rect 47210 26908 47216 26920
rect 34204 26880 47216 26908
rect 34204 26868 34210 26880
rect 47210 26868 47216 26880
rect 47268 26908 47274 26920
rect 49418 26908 49424 26920
rect 47268 26880 49424 26908
rect 47268 26868 47274 26880
rect 49418 26868 49424 26880
rect 49476 26868 49482 26920
rect 25648 26812 26740 26840
rect 25648 26800 25654 26812
rect 27062 26800 27068 26852
rect 27120 26840 27126 26852
rect 27120 26812 31754 26840
rect 27120 26800 27126 26812
rect 2501 26775 2559 26781
rect 2501 26741 2513 26775
rect 2547 26772 2559 26775
rect 30006 26772 30012 26784
rect 2547 26744 30012 26772
rect 2547 26741 2559 26744
rect 2501 26735 2559 26741
rect 30006 26732 30012 26744
rect 30064 26732 30070 26784
rect 31726 26772 31754 26812
rect 32582 26800 32588 26852
rect 32640 26800 32646 26852
rect 43714 26800 43720 26852
rect 43772 26840 43778 26852
rect 43772 26812 51074 26840
rect 43772 26800 43778 26812
rect 45462 26772 45468 26784
rect 31726 26744 45468 26772
rect 45462 26732 45468 26744
rect 45520 26732 45526 26784
rect 51046 26772 51074 26812
rect 58253 26775 58311 26781
rect 58253 26772 58265 26775
rect 51046 26744 58265 26772
rect 58253 26741 58265 26744
rect 58299 26741 58311 26775
rect 58253 26735 58311 26741
rect 1104 26682 58880 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 58880 26682
rect 1104 26608 58880 26630
rect 22922 26528 22928 26580
rect 22980 26568 22986 26580
rect 23477 26571 23535 26577
rect 23477 26568 23489 26571
rect 22980 26540 23489 26568
rect 22980 26528 22986 26540
rect 23477 26537 23489 26540
rect 23523 26568 23535 26571
rect 25406 26568 25412 26580
rect 23523 26540 25412 26568
rect 23523 26537 23535 26540
rect 23477 26531 23535 26537
rect 25406 26528 25412 26540
rect 25464 26528 25470 26580
rect 27890 26528 27896 26580
rect 27948 26568 27954 26580
rect 29914 26568 29920 26580
rect 27948 26540 29920 26568
rect 27948 26528 27954 26540
rect 29914 26528 29920 26540
rect 29972 26528 29978 26580
rect 30653 26571 30711 26577
rect 30653 26568 30665 26571
rect 30024 26540 30665 26568
rect 25041 26503 25099 26509
rect 25041 26469 25053 26503
rect 25087 26500 25099 26503
rect 25087 26472 25452 26500
rect 25087 26469 25099 26472
rect 25041 26463 25099 26469
rect 25424 26432 25452 26472
rect 25608 26472 29684 26500
rect 25608 26432 25636 26472
rect 28166 26432 28172 26444
rect 25424 26404 25636 26432
rect 25700 26404 28172 26432
rect 1581 26367 1639 26373
rect 1581 26333 1593 26367
rect 1627 26364 1639 26367
rect 20162 26364 20168 26376
rect 1627 26336 20168 26364
rect 1627 26333 1639 26336
rect 1581 26327 1639 26333
rect 20162 26324 20168 26336
rect 20220 26324 20226 26376
rect 25225 26367 25283 26373
rect 25225 26364 25237 26367
rect 20916 26336 25237 26364
rect 934 26256 940 26308
rect 992 26296 998 26308
rect 1857 26299 1915 26305
rect 1857 26296 1869 26299
rect 992 26268 1869 26296
rect 992 26256 998 26268
rect 1857 26265 1869 26268
rect 1903 26265 1915 26299
rect 1857 26259 1915 26265
rect 1946 26256 1952 26308
rect 2004 26296 2010 26308
rect 20916 26296 20944 26336
rect 25225 26333 25237 26336
rect 25271 26333 25283 26367
rect 25225 26327 25283 26333
rect 25406 26324 25412 26376
rect 25464 26373 25470 26376
rect 25464 26367 25507 26373
rect 25495 26333 25507 26367
rect 25464 26327 25507 26333
rect 25464 26324 25470 26327
rect 25590 26324 25596 26376
rect 25648 26324 25654 26376
rect 2004 26268 20944 26296
rect 2004 26256 2010 26268
rect 23198 26256 23204 26308
rect 23256 26296 23262 26308
rect 23385 26299 23443 26305
rect 23385 26296 23397 26299
rect 23256 26268 23397 26296
rect 23256 26256 23262 26268
rect 23385 26265 23397 26268
rect 23431 26265 23443 26299
rect 23385 26259 23443 26265
rect 24854 26256 24860 26308
rect 24912 26296 24918 26308
rect 25327 26299 25385 26305
rect 25327 26296 25339 26299
rect 24912 26268 25339 26296
rect 24912 26256 24918 26268
rect 25327 26265 25339 26268
rect 25373 26265 25385 26299
rect 25700 26296 25728 26404
rect 28166 26392 28172 26404
rect 28224 26392 28230 26444
rect 28350 26392 28356 26444
rect 28408 26392 28414 26444
rect 26510 26324 26516 26376
rect 26568 26324 26574 26376
rect 27893 26367 27951 26373
rect 27893 26333 27905 26367
rect 27939 26364 27951 26367
rect 29086 26364 29092 26376
rect 27939 26336 29092 26364
rect 27939 26333 27951 26336
rect 27893 26327 27951 26333
rect 29086 26324 29092 26336
rect 29144 26324 29150 26376
rect 25327 26259 25385 26265
rect 25424 26268 25728 26296
rect 24762 26188 24768 26240
rect 24820 26228 24826 26240
rect 25424 26228 25452 26268
rect 26326 26256 26332 26308
rect 26384 26256 26390 26308
rect 26694 26256 26700 26308
rect 26752 26296 26758 26308
rect 26881 26299 26939 26305
rect 26881 26296 26893 26299
rect 26752 26268 26893 26296
rect 26752 26256 26758 26268
rect 26881 26265 26893 26268
rect 26927 26265 26939 26299
rect 29656 26296 29684 26472
rect 30024 26432 30052 26540
rect 30653 26537 30665 26540
rect 30699 26568 30711 26571
rect 59354 26568 59360 26580
rect 30699 26540 59360 26568
rect 30699 26537 30711 26540
rect 30653 26531 30711 26537
rect 59354 26528 59360 26540
rect 59412 26528 59418 26580
rect 43254 26500 43260 26512
rect 30760 26472 43260 26500
rect 30760 26432 30788 26472
rect 43254 26460 43260 26472
rect 43312 26460 43318 26512
rect 47946 26460 47952 26512
rect 48004 26500 48010 26512
rect 49605 26503 49663 26509
rect 49605 26500 49617 26503
rect 48004 26472 49617 26500
rect 48004 26460 48010 26472
rect 49605 26469 49617 26472
rect 49651 26469 49663 26503
rect 49605 26463 49663 26469
rect 29748 26404 30052 26432
rect 30576 26404 30788 26432
rect 31481 26435 31539 26441
rect 29748 26373 29776 26404
rect 29733 26367 29791 26373
rect 29733 26333 29745 26367
rect 29779 26333 29791 26367
rect 29733 26327 29791 26333
rect 29914 26324 29920 26376
rect 29972 26324 29978 26376
rect 30006 26324 30012 26376
rect 30064 26324 30070 26376
rect 30098 26324 30104 26376
rect 30156 26324 30162 26376
rect 30576 26296 30604 26404
rect 31481 26401 31493 26435
rect 31527 26432 31539 26435
rect 31662 26432 31668 26444
rect 31527 26404 31668 26432
rect 31527 26401 31539 26404
rect 31481 26395 31539 26401
rect 31662 26392 31668 26404
rect 31720 26392 31726 26444
rect 32950 26432 32956 26444
rect 31772 26404 32956 26432
rect 30650 26324 30656 26376
rect 30708 26364 30714 26376
rect 31573 26367 31631 26373
rect 31573 26364 31585 26367
rect 30708 26336 31585 26364
rect 30708 26324 30714 26336
rect 31573 26333 31585 26336
rect 31619 26364 31631 26367
rect 31772 26364 31800 26404
rect 32950 26392 32956 26404
rect 33008 26392 33014 26444
rect 35342 26392 35348 26444
rect 35400 26432 35406 26444
rect 37826 26432 37832 26444
rect 35400 26404 37832 26432
rect 35400 26392 35406 26404
rect 37826 26392 37832 26404
rect 37884 26432 37890 26444
rect 48774 26432 48780 26444
rect 37884 26404 48780 26432
rect 37884 26392 37890 26404
rect 31619 26336 31800 26364
rect 32033 26367 32091 26373
rect 31619 26333 31631 26336
rect 31573 26327 31631 26333
rect 32033 26333 32045 26367
rect 32079 26364 32091 26367
rect 42794 26364 42800 26376
rect 32079 26336 42800 26364
rect 32079 26333 32091 26336
rect 32033 26327 32091 26333
rect 29656 26268 30604 26296
rect 26881 26259 26939 26265
rect 30742 26256 30748 26308
rect 30800 26296 30806 26308
rect 32048 26296 32076 26327
rect 42794 26324 42800 26336
rect 42852 26364 42858 26376
rect 43070 26364 43076 26376
rect 42852 26336 43076 26364
rect 42852 26324 42858 26336
rect 43070 26324 43076 26336
rect 43128 26324 43134 26376
rect 43254 26324 43260 26376
rect 43312 26364 43318 26376
rect 47857 26367 47915 26373
rect 47857 26364 47869 26367
rect 43312 26336 47869 26364
rect 43312 26324 43318 26336
rect 47857 26333 47869 26336
rect 47903 26333 47915 26367
rect 47857 26327 47915 26333
rect 47950 26367 48008 26373
rect 47950 26333 47962 26367
rect 47996 26333 48008 26367
rect 47950 26327 48008 26333
rect 30800 26268 32076 26296
rect 30800 26256 30806 26268
rect 43162 26256 43168 26308
rect 43220 26296 43226 26308
rect 43714 26296 43720 26308
rect 43220 26268 43720 26296
rect 43220 26256 43226 26268
rect 43714 26256 43720 26268
rect 43772 26256 43778 26308
rect 24820 26200 25452 26228
rect 24820 26188 24826 26200
rect 30282 26188 30288 26240
rect 30340 26188 30346 26240
rect 47964 26228 47992 26327
rect 48222 26324 48228 26376
rect 48280 26324 48286 26376
rect 48332 26373 48360 26404
rect 48774 26392 48780 26404
rect 48832 26432 48838 26444
rect 49234 26432 49240 26444
rect 48832 26404 49240 26432
rect 48832 26392 48838 26404
rect 49234 26392 49240 26404
rect 49292 26392 49298 26444
rect 52914 26432 52920 26444
rect 49344 26404 52920 26432
rect 48322 26367 48380 26373
rect 48322 26333 48334 26367
rect 48368 26333 48380 26367
rect 48322 26327 48380 26333
rect 48958 26324 48964 26376
rect 49016 26324 49022 26376
rect 49109 26367 49167 26373
rect 49109 26333 49121 26367
rect 49155 26364 49167 26367
rect 49344 26364 49372 26404
rect 52914 26392 52920 26404
rect 52972 26392 52978 26444
rect 58158 26392 58164 26444
rect 58216 26392 58222 26444
rect 49155 26336 49372 26364
rect 49155 26333 49167 26336
rect 49109 26327 49167 26333
rect 49418 26324 49424 26376
rect 49476 26373 49482 26376
rect 49476 26364 49484 26373
rect 49476 26336 49521 26364
rect 49476 26327 49484 26336
rect 49476 26324 49482 26327
rect 53098 26324 53104 26376
rect 53156 26364 53162 26376
rect 57885 26367 57943 26373
rect 57885 26364 57897 26367
rect 53156 26336 57897 26364
rect 53156 26324 53162 26336
rect 57885 26333 57897 26336
rect 57931 26333 57943 26367
rect 57885 26327 57943 26333
rect 48133 26299 48191 26305
rect 48133 26265 48145 26299
rect 48179 26296 48191 26299
rect 48682 26296 48688 26308
rect 48179 26268 48688 26296
rect 48179 26265 48191 26268
rect 48133 26259 48191 26265
rect 48682 26256 48688 26268
rect 48740 26296 48746 26308
rect 49237 26299 49295 26305
rect 49237 26296 49249 26299
rect 48740 26268 49249 26296
rect 48740 26256 48746 26268
rect 49237 26265 49249 26268
rect 49283 26265 49295 26299
rect 49237 26259 49295 26265
rect 49329 26299 49387 26305
rect 49329 26265 49341 26299
rect 49375 26265 49387 26299
rect 49329 26259 49387 26265
rect 48222 26228 48228 26240
rect 47964 26200 48228 26228
rect 48222 26188 48228 26200
rect 48280 26188 48286 26240
rect 48406 26188 48412 26240
rect 48464 26228 48470 26240
rect 48501 26231 48559 26237
rect 48501 26228 48513 26231
rect 48464 26200 48513 26228
rect 48464 26188 48470 26200
rect 48501 26197 48513 26200
rect 48547 26197 48559 26231
rect 49344 26228 49372 26259
rect 56226 26228 56232 26240
rect 49344 26200 56232 26228
rect 48501 26191 48559 26197
rect 56226 26188 56232 26200
rect 56284 26188 56290 26240
rect 1104 26138 58880 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 50294 26138
rect 50346 26086 50358 26138
rect 50410 26086 50422 26138
rect 50474 26086 50486 26138
rect 50538 26086 50550 26138
rect 50602 26086 58880 26138
rect 1104 26064 58880 26086
rect 23014 26024 23020 26036
rect 22296 25996 23020 26024
rect 20162 25916 20168 25968
rect 20220 25956 20226 25968
rect 21177 25959 21235 25965
rect 21177 25956 21189 25959
rect 20220 25928 21189 25956
rect 20220 25916 20226 25928
rect 21177 25925 21189 25928
rect 21223 25925 21235 25959
rect 21177 25919 21235 25925
rect 1578 25848 1584 25900
rect 1636 25848 1642 25900
rect 20990 25848 20996 25900
rect 21048 25848 21054 25900
rect 21453 25891 21511 25897
rect 21453 25857 21465 25891
rect 21499 25888 21511 25891
rect 22296 25888 22324 25996
rect 23014 25984 23020 25996
rect 23072 25984 23078 26036
rect 24578 25984 24584 26036
rect 24636 25984 24642 26036
rect 32582 25984 32588 26036
rect 32640 26024 32646 26036
rect 41782 26024 41788 26036
rect 32640 25996 41788 26024
rect 32640 25984 32646 25996
rect 41782 25984 41788 25996
rect 41840 25984 41846 26036
rect 22922 25916 22928 25968
rect 22980 25916 22986 25968
rect 23477 25959 23535 25965
rect 23477 25925 23489 25959
rect 23523 25956 23535 25959
rect 23658 25956 23664 25968
rect 23523 25928 23664 25956
rect 23523 25925 23535 25928
rect 23477 25919 23535 25925
rect 23658 25916 23664 25928
rect 23716 25916 23722 25968
rect 23934 25916 23940 25968
rect 23992 25956 23998 25968
rect 28537 25959 28595 25965
rect 28537 25956 28549 25959
rect 23992 25928 28549 25956
rect 23992 25916 23998 25928
rect 21499 25860 22324 25888
rect 21499 25857 21511 25860
rect 21453 25851 21511 25857
rect 22370 25848 22376 25900
rect 22428 25888 22434 25900
rect 23017 25891 23075 25897
rect 23017 25888 23029 25891
rect 22428 25860 23029 25888
rect 22428 25848 22434 25860
rect 23017 25857 23029 25860
rect 23063 25857 23075 25891
rect 23017 25851 23075 25857
rect 23290 25848 23296 25900
rect 23348 25888 23354 25900
rect 23385 25891 23443 25897
rect 23385 25888 23397 25891
rect 23348 25860 23397 25888
rect 23348 25848 23354 25860
rect 23385 25857 23397 25860
rect 23431 25857 23443 25891
rect 23385 25851 23443 25857
rect 24026 25848 24032 25900
rect 24084 25888 24090 25900
rect 27172 25897 27200 25928
rect 28537 25925 28549 25928
rect 28583 25925 28595 25959
rect 28537 25919 28595 25925
rect 29086 25916 29092 25968
rect 29144 25956 29150 25968
rect 29144 25928 38608 25956
rect 29144 25916 29150 25928
rect 24489 25891 24547 25897
rect 24489 25888 24501 25891
rect 24084 25860 24501 25888
rect 24084 25848 24090 25860
rect 24489 25857 24501 25860
rect 24535 25857 24547 25891
rect 24489 25851 24547 25857
rect 27157 25891 27215 25897
rect 27157 25857 27169 25891
rect 27203 25857 27215 25891
rect 27157 25851 27215 25857
rect 28166 25848 28172 25900
rect 28224 25848 28230 25900
rect 30098 25848 30104 25900
rect 30156 25848 30162 25900
rect 30193 25891 30251 25897
rect 30193 25857 30205 25891
rect 30239 25888 30251 25891
rect 30282 25888 30288 25900
rect 30239 25860 30288 25888
rect 30239 25857 30251 25860
rect 30193 25851 30251 25857
rect 30282 25848 30288 25860
rect 30340 25848 30346 25900
rect 30374 25848 30380 25900
rect 30432 25848 30438 25900
rect 36998 25848 37004 25900
rect 37056 25888 37062 25900
rect 38580 25897 38608 25928
rect 42058 25916 42064 25968
rect 42116 25956 42122 25968
rect 43533 25959 43591 25965
rect 43533 25956 43545 25959
rect 42116 25928 43545 25956
rect 42116 25916 42122 25928
rect 43533 25925 43545 25928
rect 43579 25925 43591 25959
rect 43533 25919 43591 25925
rect 43625 25959 43683 25965
rect 43625 25925 43637 25959
rect 43671 25956 43683 25959
rect 45370 25956 45376 25968
rect 43671 25928 45376 25956
rect 43671 25925 43683 25928
rect 43625 25919 43683 25925
rect 45370 25916 45376 25928
rect 45428 25916 45434 25968
rect 58158 25916 58164 25968
rect 58216 25916 58222 25968
rect 37645 25891 37703 25897
rect 37645 25888 37657 25891
rect 37056 25860 37657 25888
rect 37056 25848 37062 25860
rect 37645 25857 37657 25860
rect 37691 25857 37703 25891
rect 37645 25851 37703 25857
rect 38565 25891 38623 25897
rect 38565 25857 38577 25891
rect 38611 25857 38623 25891
rect 38565 25851 38623 25857
rect 41782 25848 41788 25900
rect 41840 25888 41846 25900
rect 43254 25888 43260 25900
rect 41840 25860 43260 25888
rect 41840 25848 41846 25860
rect 43254 25848 43260 25860
rect 43312 25848 43318 25900
rect 43438 25897 43444 25900
rect 43405 25891 43444 25897
rect 43405 25857 43417 25891
rect 43405 25851 43444 25857
rect 43438 25848 43444 25851
rect 43496 25848 43502 25900
rect 43806 25897 43812 25900
rect 43763 25891 43812 25897
rect 43763 25857 43775 25891
rect 43809 25857 43812 25891
rect 43763 25851 43812 25857
rect 43778 25848 43812 25851
rect 43864 25848 43870 25900
rect 934 25780 940 25832
rect 992 25820 998 25832
rect 1765 25823 1823 25829
rect 1765 25820 1777 25823
rect 992 25792 1777 25820
rect 992 25780 998 25792
rect 1765 25789 1777 25792
rect 1811 25789 1823 25823
rect 1765 25783 1823 25789
rect 23566 25780 23572 25832
rect 23624 25820 23630 25832
rect 23937 25823 23995 25829
rect 23937 25820 23949 25823
rect 23624 25792 23949 25820
rect 23624 25780 23630 25792
rect 23937 25789 23949 25792
rect 23983 25820 23995 25823
rect 24578 25820 24584 25832
rect 23983 25792 24584 25820
rect 23983 25789 23995 25792
rect 23937 25783 23995 25789
rect 24578 25780 24584 25792
rect 24636 25780 24642 25832
rect 27433 25823 27491 25829
rect 27433 25789 27445 25823
rect 27479 25820 27491 25823
rect 27706 25820 27712 25832
rect 27479 25792 27712 25820
rect 27479 25789 27491 25792
rect 27433 25783 27491 25789
rect 27706 25780 27712 25792
rect 27764 25820 27770 25832
rect 28258 25820 28264 25832
rect 27764 25792 28264 25820
rect 27764 25780 27770 25792
rect 28258 25780 28264 25792
rect 28316 25780 28322 25832
rect 30558 25780 30564 25832
rect 30616 25780 30622 25832
rect 37550 25780 37556 25832
rect 37608 25820 37614 25832
rect 37829 25823 37887 25829
rect 37829 25820 37841 25823
rect 37608 25792 37841 25820
rect 37608 25780 37614 25792
rect 37829 25789 37841 25792
rect 37875 25820 37887 25823
rect 38470 25820 38476 25832
rect 37875 25792 38476 25820
rect 37875 25789 37887 25792
rect 37829 25783 37887 25789
rect 38470 25780 38476 25792
rect 38528 25780 38534 25832
rect 38838 25780 38844 25832
rect 38896 25820 38902 25832
rect 43778 25820 43806 25848
rect 38896 25792 43806 25820
rect 38896 25780 38902 25792
rect 47118 25780 47124 25832
rect 47176 25820 47182 25832
rect 48866 25820 48872 25832
rect 47176 25792 48872 25820
rect 47176 25780 47182 25792
rect 48866 25780 48872 25792
rect 48924 25780 48930 25832
rect 23106 25712 23112 25764
rect 23164 25752 23170 25764
rect 27890 25752 27896 25764
rect 23164 25724 27896 25752
rect 23164 25712 23170 25724
rect 27890 25712 27896 25724
rect 27948 25712 27954 25764
rect 32214 25712 32220 25764
rect 32272 25752 32278 25764
rect 50062 25752 50068 25764
rect 32272 25724 50068 25752
rect 32272 25712 32278 25724
rect 50062 25712 50068 25724
rect 50120 25712 50126 25764
rect 26326 25644 26332 25696
rect 26384 25684 26390 25696
rect 43901 25687 43959 25693
rect 43901 25684 43913 25687
rect 26384 25656 43913 25684
rect 26384 25644 26390 25656
rect 43901 25653 43913 25656
rect 43947 25653 43959 25687
rect 43901 25647 43959 25653
rect 46750 25644 46756 25696
rect 46808 25684 46814 25696
rect 58253 25687 58311 25693
rect 58253 25684 58265 25687
rect 46808 25656 58265 25684
rect 46808 25644 46814 25656
rect 58253 25653 58265 25656
rect 58299 25653 58311 25687
rect 58253 25647 58311 25653
rect 1104 25594 58880 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 58880 25594
rect 1104 25520 58880 25542
rect 1578 25440 1584 25492
rect 1636 25480 1642 25492
rect 2685 25483 2743 25489
rect 2685 25480 2697 25483
rect 1636 25452 2697 25480
rect 1636 25440 1642 25452
rect 2685 25449 2697 25452
rect 2731 25449 2743 25483
rect 2685 25443 2743 25449
rect 23477 25483 23535 25489
rect 23477 25449 23489 25483
rect 23523 25480 23535 25483
rect 28166 25480 28172 25492
rect 23523 25452 28172 25480
rect 23523 25449 23535 25452
rect 23477 25443 23535 25449
rect 28166 25440 28172 25452
rect 28224 25440 28230 25492
rect 30098 25440 30104 25492
rect 30156 25480 30162 25492
rect 37921 25483 37979 25489
rect 37921 25480 37933 25483
rect 30156 25452 37933 25480
rect 30156 25440 30162 25452
rect 37921 25449 37933 25452
rect 37967 25449 37979 25483
rect 47854 25480 47860 25492
rect 37921 25443 37979 25449
rect 46584 25452 47860 25480
rect 22741 25415 22799 25421
rect 22741 25381 22753 25415
rect 22787 25412 22799 25415
rect 23658 25412 23664 25424
rect 22787 25384 23664 25412
rect 22787 25381 22799 25384
rect 22741 25375 22799 25381
rect 23658 25372 23664 25384
rect 23716 25412 23722 25424
rect 37642 25412 37648 25424
rect 23716 25384 24992 25412
rect 23716 25372 23722 25384
rect 22922 25304 22928 25356
rect 22980 25344 22986 25356
rect 23293 25347 23351 25353
rect 23293 25344 23305 25347
rect 22980 25316 23305 25344
rect 22980 25304 22986 25316
rect 23293 25313 23305 25316
rect 23339 25313 23351 25347
rect 23293 25307 23351 25313
rect 23474 25304 23480 25356
rect 23532 25344 23538 25356
rect 23532 25316 24532 25344
rect 23532 25304 23538 25316
rect 24504 25288 24532 25316
rect 24578 25304 24584 25356
rect 24636 25344 24642 25356
rect 24964 25353 24992 25384
rect 25056 25384 37648 25412
rect 24949 25347 25007 25353
rect 24636 25316 24808 25344
rect 24636 25304 24642 25316
rect 1581 25279 1639 25285
rect 1581 25245 1593 25279
rect 1627 25276 1639 25279
rect 1627 25248 2452 25276
rect 1627 25245 1639 25248
rect 1581 25239 1639 25245
rect 934 25168 940 25220
rect 992 25208 998 25220
rect 1857 25211 1915 25217
rect 1857 25208 1869 25211
rect 992 25180 1869 25208
rect 992 25168 998 25180
rect 1857 25177 1869 25180
rect 1903 25177 1915 25211
rect 2424 25208 2452 25248
rect 2498 25236 2504 25288
rect 2556 25236 2562 25288
rect 2655 25279 2713 25285
rect 2655 25245 2667 25279
rect 2701 25276 2713 25279
rect 3142 25276 3148 25288
rect 2701 25248 3148 25276
rect 2701 25245 2713 25248
rect 2655 25239 2713 25245
rect 3142 25236 3148 25248
rect 3200 25236 3206 25288
rect 23201 25279 23259 25285
rect 23201 25245 23213 25279
rect 23247 25276 23259 25279
rect 23566 25276 23572 25288
rect 23247 25248 23572 25276
rect 23247 25245 23259 25248
rect 23201 25239 23259 25245
rect 23566 25236 23572 25248
rect 23624 25236 23630 25288
rect 24486 25236 24492 25288
rect 24544 25276 24550 25288
rect 24673 25279 24731 25285
rect 24673 25276 24685 25279
rect 24544 25248 24685 25276
rect 24544 25236 24550 25248
rect 24673 25245 24685 25248
rect 24719 25245 24731 25279
rect 24780 25276 24808 25316
rect 24949 25313 24961 25347
rect 24995 25313 25007 25347
rect 24949 25307 25007 25313
rect 25056 25276 25084 25384
rect 37642 25372 37648 25384
rect 37700 25372 37706 25424
rect 43806 25372 43812 25424
rect 43864 25412 43870 25424
rect 45094 25412 45100 25424
rect 43864 25384 45100 25412
rect 43864 25372 43870 25384
rect 45094 25372 45100 25384
rect 45152 25412 45158 25424
rect 46584 25412 46612 25452
rect 47854 25440 47860 25452
rect 47912 25440 47918 25492
rect 45152 25384 46612 25412
rect 47044 25384 47348 25412
rect 45152 25372 45158 25384
rect 27706 25344 27712 25356
rect 27356 25316 27712 25344
rect 24780 25248 25084 25276
rect 24673 25239 24731 25245
rect 27154 25236 27160 25288
rect 27212 25236 27218 25288
rect 27356 25285 27384 25316
rect 27706 25304 27712 25316
rect 27764 25304 27770 25356
rect 27890 25304 27896 25356
rect 27948 25344 27954 25356
rect 28629 25347 28687 25353
rect 28629 25344 28641 25347
rect 27948 25316 28641 25344
rect 27948 25304 27954 25316
rect 28629 25313 28641 25316
rect 28675 25313 28687 25347
rect 39482 25344 39488 25356
rect 28629 25307 28687 25313
rect 37568 25316 39488 25344
rect 27341 25279 27399 25285
rect 27341 25245 27353 25279
rect 27387 25245 27399 25279
rect 27341 25239 27399 25245
rect 27522 25236 27528 25288
rect 27580 25236 27586 25288
rect 27614 25236 27620 25288
rect 27672 25276 27678 25288
rect 28169 25279 28227 25285
rect 28169 25276 28181 25279
rect 27672 25248 28181 25276
rect 27672 25236 27678 25248
rect 28169 25245 28181 25248
rect 28215 25245 28227 25279
rect 28169 25239 28227 25245
rect 28258 25236 28264 25288
rect 28316 25236 28322 25288
rect 28442 25236 28448 25288
rect 28500 25236 28506 25288
rect 29733 25279 29791 25285
rect 29733 25245 29745 25279
rect 29779 25276 29791 25279
rect 30742 25276 30748 25288
rect 29779 25248 30748 25276
rect 29779 25245 29791 25248
rect 29733 25239 29791 25245
rect 30742 25236 30748 25248
rect 30800 25236 30806 25288
rect 37274 25236 37280 25288
rect 37332 25236 37338 25288
rect 37425 25279 37483 25285
rect 37425 25245 37437 25279
rect 37471 25276 37483 25279
rect 37568 25276 37596 25316
rect 39482 25304 39488 25316
rect 39540 25304 39546 25356
rect 37471 25248 37596 25276
rect 37471 25245 37483 25248
rect 37425 25239 37483 25245
rect 37642 25236 37648 25288
rect 37700 25236 37706 25288
rect 37783 25279 37841 25285
rect 37783 25245 37795 25279
rect 37829 25276 37841 25279
rect 38838 25276 38844 25288
rect 37829 25248 38844 25276
rect 37829 25245 37841 25248
rect 37783 25239 37841 25245
rect 38838 25236 38844 25248
rect 38896 25236 38902 25288
rect 43254 25236 43260 25288
rect 43312 25276 43318 25288
rect 45922 25276 45928 25288
rect 43312 25248 45928 25276
rect 43312 25236 43318 25248
rect 45922 25236 45928 25248
rect 45980 25276 45986 25288
rect 46198 25285 46204 25288
rect 46017 25279 46075 25285
rect 46017 25276 46029 25279
rect 45980 25248 46029 25276
rect 45980 25236 45986 25248
rect 46017 25245 46029 25248
rect 46063 25245 46075 25279
rect 46017 25239 46075 25245
rect 46165 25279 46204 25285
rect 46165 25245 46177 25279
rect 46165 25239 46204 25245
rect 46198 25236 46204 25239
rect 46256 25236 46262 25288
rect 46382 25236 46388 25288
rect 46440 25236 46446 25288
rect 46497 25285 46525 25384
rect 47044 25344 47072 25384
rect 46584 25316 47072 25344
rect 46482 25279 46540 25285
rect 46482 25245 46494 25279
rect 46528 25245 46540 25279
rect 46482 25239 46540 25245
rect 22741 25211 22799 25217
rect 2424 25180 6914 25208
rect 1857 25171 1915 25177
rect 6886 25140 6914 25180
rect 22741 25177 22753 25211
rect 22787 25208 22799 25211
rect 23290 25208 23296 25220
rect 22787 25180 23296 25208
rect 22787 25177 22799 25180
rect 22741 25171 22799 25177
rect 23290 25168 23296 25180
rect 23348 25168 23354 25220
rect 27430 25168 27436 25220
rect 27488 25168 27494 25220
rect 28350 25168 28356 25220
rect 28408 25208 28414 25220
rect 28408 25180 31754 25208
rect 28408 25168 28414 25180
rect 22278 25140 22284 25152
rect 6886 25112 22284 25140
rect 22278 25100 22284 25112
rect 22336 25100 22342 25152
rect 27709 25143 27767 25149
rect 27709 25109 27721 25143
rect 27755 25140 27767 25143
rect 28074 25140 28080 25152
rect 27755 25112 28080 25140
rect 27755 25109 27767 25112
rect 27709 25103 27767 25109
rect 28074 25100 28080 25112
rect 28132 25100 28138 25152
rect 31018 25100 31024 25152
rect 31076 25100 31082 25152
rect 31726 25140 31754 25180
rect 37550 25168 37556 25220
rect 37608 25168 37614 25220
rect 37752 25180 38056 25208
rect 37752 25140 37780 25180
rect 31726 25112 37780 25140
rect 38028 25140 38056 25180
rect 38470 25168 38476 25220
rect 38528 25208 38534 25220
rect 46290 25208 46296 25220
rect 38528 25180 46296 25208
rect 38528 25168 38534 25180
rect 46290 25168 46296 25180
rect 46348 25168 46354 25220
rect 46584 25140 46612 25316
rect 47118 25236 47124 25288
rect 47176 25236 47182 25288
rect 47214 25279 47272 25285
rect 47214 25245 47226 25279
rect 47260 25245 47272 25279
rect 47214 25239 47272 25245
rect 47026 25168 47032 25220
rect 47084 25208 47090 25220
rect 47228 25208 47256 25239
rect 47084 25180 47256 25208
rect 47320 25208 47348 25384
rect 51718 25344 51724 25356
rect 47504 25316 51724 25344
rect 47394 25236 47400 25288
rect 47452 25236 47458 25288
rect 47504 25285 47532 25316
rect 51718 25304 51724 25316
rect 51776 25304 51782 25356
rect 47489 25279 47547 25285
rect 47489 25245 47501 25279
rect 47535 25245 47547 25279
rect 47489 25239 47547 25245
rect 47586 25279 47644 25285
rect 47586 25245 47598 25279
rect 47632 25276 47644 25279
rect 47632 25248 48360 25276
rect 47632 25245 47644 25248
rect 47586 25239 47644 25245
rect 47596 25208 47624 25239
rect 48225 25211 48283 25217
rect 48225 25208 48237 25211
rect 47320 25180 47624 25208
rect 47688 25180 48237 25208
rect 47084 25168 47090 25180
rect 38028 25112 46612 25140
rect 46661 25143 46719 25149
rect 46661 25109 46673 25143
rect 46707 25140 46719 25143
rect 47688 25140 47716 25180
rect 48225 25177 48237 25180
rect 48271 25177 48283 25211
rect 48332 25208 48360 25248
rect 48406 25236 48412 25288
rect 48464 25236 48470 25288
rect 57882 25236 57888 25288
rect 57940 25236 57946 25288
rect 49050 25208 49056 25220
rect 48332 25180 49056 25208
rect 48225 25171 48283 25177
rect 49050 25168 49056 25180
rect 49108 25168 49114 25220
rect 58158 25168 58164 25220
rect 58216 25168 58222 25220
rect 46707 25112 47716 25140
rect 46707 25109 46719 25112
rect 46661 25103 46719 25109
rect 47762 25100 47768 25152
rect 47820 25100 47826 25152
rect 47854 25100 47860 25152
rect 47912 25140 47918 25152
rect 48501 25143 48559 25149
rect 48501 25140 48513 25143
rect 47912 25112 48513 25140
rect 47912 25100 47918 25112
rect 48501 25109 48513 25112
rect 48547 25109 48559 25143
rect 48501 25103 48559 25109
rect 1104 25050 58880 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 50294 25050
rect 50346 24998 50358 25050
rect 50410 24998 50422 25050
rect 50474 24998 50486 25050
rect 50538 24998 50550 25050
rect 50602 24998 58880 25050
rect 1104 24976 58880 24998
rect 2498 24896 2504 24948
rect 2556 24936 2562 24948
rect 2556 24908 2728 24936
rect 2556 24896 2562 24908
rect 1578 24760 1584 24812
rect 1636 24760 1642 24812
rect 2406 24760 2412 24812
rect 2464 24800 2470 24812
rect 2501 24803 2559 24809
rect 2501 24800 2513 24803
rect 2464 24772 2513 24800
rect 2464 24760 2470 24772
rect 2501 24769 2513 24772
rect 2547 24769 2559 24803
rect 2501 24763 2559 24769
rect 2594 24803 2652 24809
rect 2594 24769 2606 24803
rect 2640 24769 2652 24803
rect 2700 24800 2728 24908
rect 23290 24896 23296 24948
rect 23348 24936 23354 24948
rect 23348 24908 24072 24936
rect 23348 24896 23354 24908
rect 22278 24828 22284 24880
rect 22336 24828 22342 24880
rect 23658 24868 23664 24880
rect 23308 24840 23664 24868
rect 15746 24800 15752 24812
rect 2700 24772 15752 24800
rect 2594 24763 2652 24769
rect 934 24692 940 24744
rect 992 24732 998 24744
rect 1765 24735 1823 24741
rect 1765 24732 1777 24735
rect 992 24704 1777 24732
rect 992 24692 998 24704
rect 1765 24701 1777 24704
rect 1811 24701 1823 24735
rect 1765 24695 1823 24701
rect 2130 24692 2136 24744
rect 2188 24732 2194 24744
rect 2608 24732 2636 24763
rect 15746 24760 15752 24772
rect 15804 24760 15810 24812
rect 20990 24760 20996 24812
rect 21048 24800 21054 24812
rect 22097 24803 22155 24809
rect 22097 24800 22109 24803
rect 21048 24772 22109 24800
rect 21048 24760 21054 24772
rect 22097 24769 22109 24772
rect 22143 24800 22155 24803
rect 22186 24800 22192 24812
rect 22143 24772 22192 24800
rect 22143 24769 22155 24772
rect 22097 24763 22155 24769
rect 22186 24760 22192 24772
rect 22244 24760 22250 24812
rect 23308 24809 23336 24840
rect 23658 24828 23664 24840
rect 23716 24828 23722 24880
rect 23293 24803 23351 24809
rect 23293 24769 23305 24803
rect 23339 24769 23351 24803
rect 23293 24763 23351 24769
rect 23569 24803 23627 24809
rect 23569 24769 23581 24803
rect 23615 24800 23627 24803
rect 23768 24800 23796 24908
rect 24044 24868 24072 24908
rect 24210 24896 24216 24948
rect 24268 24896 24274 24948
rect 37274 24896 37280 24948
rect 37332 24936 37338 24948
rect 38013 24939 38071 24945
rect 38013 24936 38025 24939
rect 37332 24908 38025 24936
rect 37332 24896 37338 24908
rect 38013 24905 38025 24908
rect 38059 24905 38071 24939
rect 38013 24899 38071 24905
rect 46290 24896 46296 24948
rect 46348 24936 46354 24948
rect 47394 24936 47400 24948
rect 46348 24908 47400 24936
rect 46348 24896 46354 24908
rect 47394 24896 47400 24908
rect 47452 24936 47458 24948
rect 47578 24936 47584 24948
rect 47452 24908 47584 24936
rect 47452 24896 47458 24908
rect 47578 24896 47584 24908
rect 47636 24896 47642 24948
rect 25593 24871 25651 24877
rect 25593 24868 25605 24871
rect 24044 24840 25605 24868
rect 25593 24837 25605 24840
rect 25639 24837 25651 24871
rect 28350 24868 28356 24880
rect 25593 24831 25651 24837
rect 27724 24840 28356 24868
rect 23615 24772 23796 24800
rect 23615 24769 23627 24772
rect 23569 24763 23627 24769
rect 24026 24760 24032 24812
rect 24084 24760 24090 24812
rect 24581 24803 24639 24809
rect 24581 24800 24593 24803
rect 24136 24772 24593 24800
rect 2188 24704 2636 24732
rect 22373 24735 22431 24741
rect 2188 24692 2194 24704
rect 22373 24701 22385 24735
rect 22419 24732 22431 24735
rect 22419 24704 23520 24732
rect 22419 24701 22431 24704
rect 22373 24695 22431 24701
rect 23492 24676 23520 24704
rect 2869 24667 2927 24673
rect 2869 24633 2881 24667
rect 2915 24664 2927 24667
rect 2958 24664 2964 24676
rect 2915 24636 2964 24664
rect 2915 24633 2927 24636
rect 2869 24627 2927 24633
rect 2958 24624 2964 24636
rect 3016 24624 3022 24676
rect 23474 24624 23480 24676
rect 23532 24624 23538 24676
rect 23198 24556 23204 24608
rect 23256 24596 23262 24608
rect 24136 24596 24164 24772
rect 24581 24769 24593 24772
rect 24627 24769 24639 24803
rect 24581 24763 24639 24769
rect 24854 24760 24860 24812
rect 24912 24800 24918 24812
rect 25130 24800 25136 24812
rect 24912 24772 25136 24800
rect 24912 24760 24918 24772
rect 25130 24760 25136 24772
rect 25188 24800 25194 24812
rect 25225 24803 25283 24809
rect 25225 24800 25237 24803
rect 25188 24772 25237 24800
rect 25188 24760 25194 24772
rect 25225 24769 25237 24772
rect 25271 24769 25283 24803
rect 25225 24763 25283 24769
rect 25682 24760 25688 24812
rect 25740 24800 25746 24812
rect 27525 24803 27583 24809
rect 25740 24772 25912 24800
rect 25740 24760 25746 24772
rect 25884 24732 25912 24772
rect 27525 24769 27537 24803
rect 27571 24800 27583 24803
rect 27614 24800 27620 24812
rect 27571 24772 27620 24800
rect 27571 24769 27583 24772
rect 27525 24763 27583 24769
rect 27614 24760 27620 24772
rect 27672 24760 27678 24812
rect 27724 24809 27752 24840
rect 28350 24828 28356 24840
rect 28408 24828 28414 24880
rect 30469 24871 30527 24877
rect 30469 24868 30481 24871
rect 29012 24840 30481 24868
rect 27709 24803 27767 24809
rect 27709 24769 27721 24803
rect 27755 24769 27767 24803
rect 27709 24763 27767 24769
rect 27801 24803 27859 24809
rect 27801 24769 27813 24803
rect 27847 24769 27859 24803
rect 27985 24803 28043 24809
rect 27985 24800 27997 24803
rect 27801 24763 27859 24769
rect 27908 24772 27997 24800
rect 27816 24732 27844 24763
rect 25884 24704 27844 24732
rect 24302 24624 24308 24676
rect 24360 24664 24366 24676
rect 27908 24664 27936 24772
rect 27985 24769 27997 24772
rect 28031 24769 28043 24803
rect 27985 24763 28043 24769
rect 28074 24760 28080 24812
rect 28132 24760 28138 24812
rect 28721 24803 28779 24809
rect 28721 24769 28733 24803
rect 28767 24800 28779 24803
rect 28902 24800 28908 24812
rect 28767 24772 28908 24800
rect 28767 24769 28779 24772
rect 28721 24763 28779 24769
rect 28902 24760 28908 24772
rect 28960 24760 28966 24812
rect 28626 24692 28632 24744
rect 28684 24732 28690 24744
rect 29012 24732 29040 24840
rect 30469 24837 30481 24840
rect 30515 24868 30527 24871
rect 30742 24868 30748 24880
rect 30515 24840 30748 24868
rect 30515 24837 30527 24840
rect 30469 24831 30527 24837
rect 30742 24828 30748 24840
rect 30800 24868 30806 24880
rect 32766 24868 32772 24880
rect 30800 24840 32772 24868
rect 30800 24828 30806 24840
rect 32766 24828 32772 24840
rect 32824 24828 32830 24880
rect 37568 24840 37964 24868
rect 37461 24803 37519 24809
rect 37461 24769 37473 24803
rect 37507 24800 37519 24803
rect 37568 24800 37596 24840
rect 37507 24772 37596 24800
rect 37645 24803 37703 24809
rect 37507 24769 37519 24772
rect 37461 24763 37519 24769
rect 37645 24769 37657 24803
rect 37691 24769 37703 24803
rect 37645 24763 37703 24769
rect 28684 24704 29040 24732
rect 28684 24692 28690 24704
rect 29730 24692 29736 24744
rect 29788 24732 29794 24744
rect 31018 24732 31024 24744
rect 29788 24704 31024 24732
rect 29788 24692 29794 24704
rect 31018 24692 31024 24704
rect 31076 24692 31082 24744
rect 37366 24732 37372 24744
rect 31726 24704 37372 24732
rect 24360 24636 27936 24664
rect 24360 24624 24366 24636
rect 23256 24568 24164 24596
rect 27908 24596 27936 24636
rect 28074 24624 28080 24676
rect 28132 24664 28138 24676
rect 31726 24664 31754 24704
rect 37366 24692 37372 24704
rect 37424 24732 37430 24744
rect 37660 24732 37688 24763
rect 37734 24760 37740 24812
rect 37792 24760 37798 24812
rect 37826 24760 37832 24812
rect 37884 24760 37890 24812
rect 37936 24800 37964 24840
rect 47762 24828 47768 24880
rect 47820 24828 47826 24880
rect 48222 24828 48228 24880
rect 48280 24868 48286 24880
rect 51442 24868 51448 24880
rect 48280 24840 51448 24868
rect 48280 24828 48286 24840
rect 51442 24828 51448 24840
rect 51500 24828 51506 24880
rect 40678 24800 40684 24812
rect 37936 24772 40684 24800
rect 40678 24760 40684 24772
rect 40736 24760 40742 24812
rect 47946 24760 47952 24812
rect 48004 24760 48010 24812
rect 58066 24760 58072 24812
rect 58124 24760 58130 24812
rect 37424 24704 37688 24732
rect 37424 24692 37430 24704
rect 39298 24692 39304 24744
rect 39356 24732 39362 24744
rect 39356 24704 51074 24732
rect 39356 24692 39362 24704
rect 42978 24664 42984 24676
rect 28132 24636 31754 24664
rect 36464 24636 42984 24664
rect 28132 24624 28138 24636
rect 29730 24596 29736 24608
rect 27908 24568 29736 24596
rect 23256 24556 23262 24568
rect 29730 24556 29736 24568
rect 29788 24556 29794 24608
rect 31018 24556 31024 24608
rect 31076 24596 31082 24608
rect 36464 24596 36492 24636
rect 42978 24624 42984 24636
rect 43036 24624 43042 24676
rect 51046 24664 51074 24704
rect 58253 24667 58311 24673
rect 58253 24664 58265 24667
rect 51046 24636 58265 24664
rect 58253 24633 58265 24636
rect 58299 24633 58311 24667
rect 58253 24627 58311 24633
rect 31076 24568 36492 24596
rect 31076 24556 31082 24568
rect 36538 24556 36544 24608
rect 36596 24596 36602 24608
rect 40770 24596 40776 24608
rect 36596 24568 40776 24596
rect 36596 24556 36602 24568
rect 40770 24556 40776 24568
rect 40828 24556 40834 24608
rect 48038 24556 48044 24608
rect 48096 24556 48102 24608
rect 1104 24506 58880 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 58880 24506
rect 1104 24432 58880 24454
rect 1578 24352 1584 24404
rect 1636 24392 1642 24404
rect 2685 24395 2743 24401
rect 2685 24392 2697 24395
rect 1636 24364 2697 24392
rect 1636 24352 1642 24364
rect 2685 24361 2697 24364
rect 2731 24361 2743 24395
rect 27798 24392 27804 24404
rect 2685 24355 2743 24361
rect 22066 24364 27804 24392
rect 12802 24284 12808 24336
rect 12860 24324 12866 24336
rect 12860 24296 16574 24324
rect 12860 24284 12866 24296
rect 16114 24256 16120 24268
rect 1596 24228 16120 24256
rect 1596 24197 1624 24228
rect 16114 24216 16120 24228
rect 16172 24216 16178 24268
rect 16546 24256 16574 24296
rect 17218 24284 17224 24336
rect 17276 24324 17282 24336
rect 17770 24324 17776 24336
rect 17276 24296 17776 24324
rect 17276 24284 17282 24296
rect 17770 24284 17776 24296
rect 17828 24324 17834 24336
rect 22066 24324 22094 24364
rect 27798 24352 27804 24364
rect 27856 24352 27862 24404
rect 28258 24352 28264 24404
rect 28316 24392 28322 24404
rect 28813 24395 28871 24401
rect 28813 24392 28825 24395
rect 28316 24364 28825 24392
rect 28316 24352 28322 24364
rect 28813 24361 28825 24364
rect 28859 24361 28871 24395
rect 28813 24355 28871 24361
rect 30374 24352 30380 24404
rect 30432 24352 30438 24404
rect 36538 24392 36544 24404
rect 31726 24364 36544 24392
rect 17828 24296 22094 24324
rect 17828 24284 17834 24296
rect 28166 24284 28172 24336
rect 28224 24324 28230 24336
rect 28442 24324 28448 24336
rect 28224 24296 28448 24324
rect 28224 24284 28230 24296
rect 28442 24284 28448 24296
rect 28500 24284 28506 24336
rect 28534 24284 28540 24336
rect 28592 24324 28598 24336
rect 31726 24324 31754 24364
rect 36538 24352 36544 24364
rect 36596 24352 36602 24404
rect 37090 24352 37096 24404
rect 37148 24392 37154 24404
rect 41322 24392 41328 24404
rect 37148 24364 41328 24392
rect 37148 24352 37154 24364
rect 41322 24352 41328 24364
rect 41380 24352 41386 24404
rect 47670 24352 47676 24404
rect 47728 24352 47734 24404
rect 28592 24296 31754 24324
rect 28592 24284 28598 24296
rect 33134 24284 33140 24336
rect 33192 24324 33198 24336
rect 33192 24296 51074 24324
rect 33192 24284 33198 24296
rect 45186 24256 45192 24268
rect 16546 24228 28580 24256
rect 1581 24191 1639 24197
rect 1581 24157 1593 24191
rect 1627 24157 1639 24191
rect 1581 24151 1639 24157
rect 2406 24148 2412 24200
rect 2464 24188 2470 24200
rect 2682 24197 2688 24200
rect 2501 24191 2559 24197
rect 2501 24188 2513 24191
rect 2464 24160 2513 24188
rect 2464 24148 2470 24160
rect 2501 24157 2513 24160
rect 2547 24157 2559 24191
rect 2501 24151 2559 24157
rect 2655 24191 2688 24197
rect 2655 24157 2667 24191
rect 2655 24151 2688 24157
rect 2682 24148 2688 24151
rect 2740 24148 2746 24200
rect 23106 24148 23112 24200
rect 23164 24148 23170 24200
rect 23290 24148 23296 24200
rect 23348 24188 23354 24200
rect 23477 24191 23535 24197
rect 23477 24188 23489 24191
rect 23348 24160 23489 24188
rect 23348 24148 23354 24160
rect 23477 24157 23489 24160
rect 23523 24157 23535 24191
rect 23477 24151 23535 24157
rect 23658 24148 23664 24200
rect 23716 24188 23722 24200
rect 24029 24191 24087 24197
rect 24029 24188 24041 24191
rect 23716 24160 24041 24188
rect 23716 24148 23722 24160
rect 24029 24157 24041 24160
rect 24075 24157 24087 24191
rect 24029 24151 24087 24157
rect 28166 24148 28172 24200
rect 28224 24148 28230 24200
rect 28262 24191 28320 24197
rect 28262 24157 28274 24191
rect 28308 24157 28320 24191
rect 28262 24151 28320 24157
rect 934 24080 940 24132
rect 992 24120 998 24132
rect 1857 24123 1915 24129
rect 1857 24120 1869 24123
rect 992 24092 1869 24120
rect 992 24080 998 24092
rect 1857 24089 1869 24092
rect 1903 24089 1915 24123
rect 1857 24083 1915 24089
rect 23017 24123 23075 24129
rect 23017 24089 23029 24123
rect 23063 24089 23075 24123
rect 23017 24083 23075 24089
rect 23032 24052 23060 24083
rect 23198 24080 23204 24132
rect 23256 24120 23262 24132
rect 23569 24123 23627 24129
rect 23569 24120 23581 24123
rect 23256 24092 23581 24120
rect 23256 24080 23262 24092
rect 23569 24089 23581 24092
rect 23615 24089 23627 24123
rect 23569 24083 23627 24089
rect 27982 24080 27988 24132
rect 28040 24120 28046 24132
rect 28276 24120 28304 24151
rect 28442 24148 28448 24200
rect 28500 24148 28506 24200
rect 28552 24197 28580 24228
rect 36556 24228 45192 24256
rect 28537 24191 28595 24197
rect 28537 24157 28549 24191
rect 28583 24157 28595 24191
rect 28537 24151 28595 24157
rect 28626 24148 28632 24200
rect 28684 24197 28690 24200
rect 28684 24188 28692 24197
rect 28684 24160 28729 24188
rect 28684 24151 28692 24160
rect 28684 24148 28690 24151
rect 29730 24148 29736 24200
rect 29788 24148 29794 24200
rect 29822 24148 29828 24200
rect 29880 24148 29886 24200
rect 30282 24197 30288 24200
rect 30239 24191 30288 24197
rect 30239 24157 30251 24191
rect 30285 24157 30288 24191
rect 30239 24151 30288 24157
rect 30282 24148 30288 24151
rect 30340 24148 30346 24200
rect 28040 24092 28304 24120
rect 28460 24120 28488 24148
rect 29086 24120 29092 24132
rect 28460 24092 29092 24120
rect 28040 24080 28046 24092
rect 29086 24080 29092 24092
rect 29144 24080 29150 24132
rect 30009 24123 30067 24129
rect 30009 24089 30021 24123
rect 30055 24089 30067 24123
rect 30009 24083 30067 24089
rect 30101 24123 30159 24129
rect 30101 24089 30113 24123
rect 30147 24120 30159 24123
rect 36556 24120 36584 24228
rect 45186 24216 45192 24228
rect 45244 24216 45250 24268
rect 51046 24256 51074 24296
rect 54294 24256 54300 24268
rect 47412 24228 49188 24256
rect 51046 24228 54300 24256
rect 37274 24148 37280 24200
rect 37332 24148 37338 24200
rect 37366 24148 37372 24200
rect 37424 24188 37430 24200
rect 37461 24191 37519 24197
rect 37461 24188 37473 24191
rect 37424 24160 37473 24188
rect 37424 24148 37430 24160
rect 37461 24157 37473 24160
rect 37507 24157 37519 24191
rect 37461 24151 37519 24157
rect 37642 24148 37648 24200
rect 37700 24148 37706 24200
rect 40773 24191 40831 24197
rect 37798 24160 38654 24188
rect 30147 24092 36584 24120
rect 30147 24089 30159 24092
rect 30101 24083 30159 24089
rect 24026 24052 24032 24064
rect 23032 24024 24032 24052
rect 24026 24012 24032 24024
rect 24084 24012 24090 24064
rect 27706 24012 27712 24064
rect 27764 24052 27770 24064
rect 30024 24052 30052 24083
rect 36630 24080 36636 24132
rect 36688 24120 36694 24132
rect 37553 24123 37611 24129
rect 36688 24092 37504 24120
rect 36688 24080 36694 24092
rect 32030 24052 32036 24064
rect 27764 24024 32036 24052
rect 27764 24012 27770 24024
rect 32030 24012 32036 24024
rect 32088 24012 32094 24064
rect 37476 24052 37504 24092
rect 37553 24089 37565 24123
rect 37599 24120 37611 24123
rect 37798 24120 37826 24160
rect 37599 24092 37826 24120
rect 38626 24120 38654 24160
rect 40773 24157 40785 24191
rect 40819 24188 40831 24191
rect 42794 24188 42800 24200
rect 40819 24160 42800 24188
rect 40819 24157 40831 24160
rect 40773 24151 40831 24157
rect 42794 24148 42800 24160
rect 42852 24148 42858 24200
rect 46934 24148 46940 24200
rect 46992 24188 46998 24200
rect 47029 24191 47087 24197
rect 47029 24188 47041 24191
rect 46992 24160 47041 24188
rect 46992 24148 46998 24160
rect 47029 24157 47041 24160
rect 47075 24157 47087 24191
rect 47029 24151 47087 24157
rect 47177 24191 47235 24197
rect 47177 24157 47189 24191
rect 47223 24188 47235 24191
rect 47412 24188 47440 24228
rect 47578 24197 47584 24200
rect 47223 24160 47440 24188
rect 47535 24191 47584 24197
rect 47223 24157 47235 24160
rect 47177 24151 47235 24157
rect 47535 24157 47547 24191
rect 47581 24157 47584 24191
rect 47535 24151 47584 24157
rect 47578 24148 47584 24151
rect 47636 24148 47642 24200
rect 39390 24120 39396 24132
rect 38626 24092 39396 24120
rect 37599 24089 37611 24092
rect 37553 24083 37611 24089
rect 39390 24080 39396 24092
rect 39448 24080 39454 24132
rect 47305 24123 47363 24129
rect 47305 24120 47317 24123
rect 39500 24092 47317 24120
rect 37829 24055 37887 24061
rect 37829 24052 37841 24055
rect 37476 24024 37841 24052
rect 37829 24021 37841 24024
rect 37875 24021 37887 24055
rect 37829 24015 37887 24021
rect 37918 24012 37924 24064
rect 37976 24052 37982 24064
rect 39500 24052 39528 24092
rect 47305 24089 47317 24092
rect 47351 24089 47363 24123
rect 47305 24083 47363 24089
rect 47394 24080 47400 24132
rect 47452 24080 47458 24132
rect 37976 24024 39528 24052
rect 37976 24012 37982 24024
rect 40218 24012 40224 24064
rect 40276 24052 40282 24064
rect 40957 24055 41015 24061
rect 40957 24052 40969 24055
rect 40276 24024 40969 24052
rect 40276 24012 40282 24024
rect 40957 24021 40969 24024
rect 41003 24021 41015 24055
rect 49160 24052 49188 24228
rect 54294 24216 54300 24228
rect 54352 24216 54358 24268
rect 55214 24148 55220 24200
rect 55272 24188 55278 24200
rect 57885 24191 57943 24197
rect 57885 24188 57897 24191
rect 55272 24160 57897 24188
rect 55272 24148 55278 24160
rect 57885 24157 57897 24160
rect 57931 24157 57943 24191
rect 57885 24151 57943 24157
rect 58158 24080 58164 24132
rect 58216 24080 58222 24132
rect 53374 24052 53380 24064
rect 49160 24024 53380 24052
rect 40957 24015 41015 24021
rect 53374 24012 53380 24024
rect 53432 24012 53438 24064
rect 1104 23962 58880 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 50294 23962
rect 50346 23910 50358 23962
rect 50410 23910 50422 23962
rect 50474 23910 50486 23962
rect 50538 23910 50550 23962
rect 50602 23910 58880 23962
rect 1104 23888 58880 23910
rect 16114 23808 16120 23860
rect 16172 23808 16178 23860
rect 23198 23808 23204 23860
rect 23256 23808 23262 23860
rect 24394 23808 24400 23860
rect 24452 23808 24458 23860
rect 28166 23808 28172 23860
rect 28224 23848 28230 23860
rect 36630 23848 36636 23860
rect 28224 23820 36636 23848
rect 28224 23808 28230 23820
rect 36630 23808 36636 23820
rect 36688 23808 36694 23860
rect 36817 23851 36875 23857
rect 36817 23817 36829 23851
rect 36863 23817 36875 23851
rect 42150 23848 42156 23860
rect 36817 23811 36875 23817
rect 38396 23820 42156 23848
rect 20990 23780 20996 23792
rect 15764 23752 20996 23780
rect 15764 23724 15792 23752
rect 20990 23740 20996 23752
rect 21048 23740 21054 23792
rect 23216 23780 23244 23808
rect 23216 23752 24440 23780
rect 1581 23715 1639 23721
rect 1581 23681 1593 23715
rect 1627 23712 1639 23715
rect 2866 23712 2872 23724
rect 1627 23684 2872 23712
rect 1627 23681 1639 23684
rect 1581 23675 1639 23681
rect 2866 23672 2872 23684
rect 2924 23672 2930 23724
rect 15746 23672 15752 23724
rect 15804 23672 15810 23724
rect 15903 23715 15961 23721
rect 15903 23681 15915 23715
rect 15949 23712 15961 23715
rect 17770 23712 17776 23724
rect 15949 23684 17776 23712
rect 15949 23681 15961 23684
rect 15903 23675 15961 23681
rect 17770 23672 17776 23684
rect 17828 23672 17834 23724
rect 23477 23715 23535 23721
rect 23477 23681 23489 23715
rect 23523 23712 23535 23715
rect 23658 23712 23664 23724
rect 23523 23684 23664 23712
rect 23523 23681 23535 23684
rect 23477 23675 23535 23681
rect 23658 23672 23664 23684
rect 23716 23672 23722 23724
rect 23753 23715 23811 23721
rect 23753 23681 23765 23715
rect 23799 23681 23811 23715
rect 23753 23675 23811 23681
rect 934 23604 940 23656
rect 992 23644 998 23656
rect 1765 23647 1823 23653
rect 1765 23644 1777 23647
rect 992 23616 1777 23644
rect 992 23604 998 23616
rect 1765 23613 1777 23616
rect 1811 23613 1823 23647
rect 1765 23607 1823 23613
rect 23290 23604 23296 23656
rect 23348 23644 23354 23656
rect 23768 23644 23796 23675
rect 24026 23672 24032 23724
rect 24084 23672 24090 23724
rect 24412 23721 24440 23752
rect 27798 23740 27804 23792
rect 27856 23780 27862 23792
rect 28626 23780 28632 23792
rect 27856 23752 28632 23780
rect 27856 23740 27862 23752
rect 28626 23740 28632 23752
rect 28684 23740 28690 23792
rect 36832 23780 36860 23811
rect 37366 23780 37372 23792
rect 36832 23752 37372 23780
rect 37366 23740 37372 23752
rect 37424 23740 37430 23792
rect 24397 23715 24455 23721
rect 24397 23681 24409 23715
rect 24443 23681 24455 23715
rect 24397 23675 24455 23681
rect 34149 23715 34207 23721
rect 34149 23681 34161 23715
rect 34195 23681 34207 23715
rect 34149 23675 34207 23681
rect 34333 23715 34391 23721
rect 34333 23681 34345 23715
rect 34379 23712 34391 23715
rect 34422 23712 34428 23724
rect 34379 23684 34428 23712
rect 34379 23681 34391 23684
rect 34333 23675 34391 23681
rect 23348 23616 23796 23644
rect 23348 23604 23354 23616
rect 34164 23576 34192 23675
rect 34422 23672 34428 23684
rect 34480 23672 34486 23724
rect 36633 23715 36691 23721
rect 36633 23681 36645 23715
rect 36679 23712 36691 23715
rect 36906 23712 36912 23724
rect 36679 23684 36912 23712
rect 36679 23681 36691 23684
rect 36633 23675 36691 23681
rect 36906 23672 36912 23684
rect 36964 23672 36970 23724
rect 38396 23721 38424 23820
rect 42150 23808 42156 23820
rect 42208 23808 42214 23860
rect 42702 23780 42708 23792
rect 39132 23752 42708 23780
rect 39132 23721 39160 23752
rect 42702 23740 42708 23752
rect 42760 23740 42766 23792
rect 38381 23715 38439 23721
rect 38381 23681 38393 23715
rect 38427 23681 38439 23715
rect 38381 23675 38439 23681
rect 39117 23715 39175 23721
rect 39117 23681 39129 23715
rect 39163 23681 39175 23715
rect 39117 23675 39175 23681
rect 40221 23715 40279 23721
rect 40221 23681 40233 23715
rect 40267 23712 40279 23715
rect 40862 23712 40868 23724
rect 40267 23684 40868 23712
rect 40267 23681 40279 23684
rect 40221 23675 40279 23681
rect 40862 23672 40868 23684
rect 40920 23672 40926 23724
rect 40957 23715 41015 23721
rect 40957 23681 40969 23715
rect 41003 23712 41015 23715
rect 41003 23684 41414 23712
rect 41003 23681 41015 23684
rect 40957 23675 41015 23681
rect 35894 23604 35900 23656
rect 35952 23644 35958 23656
rect 41386 23644 41414 23684
rect 41690 23672 41696 23724
rect 41748 23672 41754 23724
rect 41877 23715 41935 23721
rect 41877 23681 41889 23715
rect 41923 23712 41935 23715
rect 42150 23712 42156 23724
rect 41923 23684 42156 23712
rect 41923 23681 41935 23684
rect 41877 23675 41935 23681
rect 42150 23672 42156 23684
rect 42208 23672 42214 23724
rect 58066 23672 58072 23724
rect 58124 23672 58130 23724
rect 42886 23644 42892 23656
rect 35952 23616 41184 23644
rect 41386 23616 42892 23644
rect 35952 23604 35958 23616
rect 36722 23576 36728 23588
rect 34164 23548 36728 23576
rect 36722 23536 36728 23548
rect 36780 23536 36786 23588
rect 39301 23579 39359 23585
rect 39301 23576 39313 23579
rect 36832 23548 39313 23576
rect 34146 23468 34152 23520
rect 34204 23468 34210 23520
rect 36354 23468 36360 23520
rect 36412 23508 36418 23520
rect 36832 23508 36860 23548
rect 39301 23545 39313 23548
rect 39347 23545 39359 23579
rect 39301 23539 39359 23545
rect 40126 23536 40132 23588
rect 40184 23576 40190 23588
rect 41156 23585 41184 23616
rect 42886 23604 42892 23616
rect 42944 23604 42950 23656
rect 41141 23579 41199 23585
rect 40184 23548 41092 23576
rect 40184 23536 40190 23548
rect 36412 23480 36860 23508
rect 36412 23468 36418 23480
rect 37458 23468 37464 23520
rect 37516 23508 37522 23520
rect 38565 23511 38623 23517
rect 38565 23508 38577 23511
rect 37516 23480 38577 23508
rect 37516 23468 37522 23480
rect 38565 23477 38577 23480
rect 38611 23477 38623 23511
rect 38565 23471 38623 23477
rect 40034 23468 40040 23520
rect 40092 23508 40098 23520
rect 40405 23511 40463 23517
rect 40405 23508 40417 23511
rect 40092 23480 40417 23508
rect 40092 23468 40098 23480
rect 40405 23477 40417 23480
rect 40451 23477 40463 23511
rect 41064 23508 41092 23548
rect 41141 23545 41153 23579
rect 41187 23545 41199 23579
rect 41141 23539 41199 23545
rect 41322 23536 41328 23588
rect 41380 23576 41386 23588
rect 58253 23579 58311 23585
rect 58253 23576 58265 23579
rect 41380 23548 58265 23576
rect 41380 23536 41386 23548
rect 58253 23545 58265 23548
rect 58299 23545 58311 23579
rect 58253 23539 58311 23545
rect 41785 23511 41843 23517
rect 41785 23508 41797 23511
rect 41064 23480 41797 23508
rect 40405 23471 40463 23477
rect 41785 23477 41797 23480
rect 41831 23477 41843 23511
rect 41785 23471 41843 23477
rect 1104 23418 58880 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 58880 23418
rect 1104 23344 58880 23366
rect 21358 23264 21364 23316
rect 21416 23304 21422 23316
rect 24670 23304 24676 23316
rect 21416 23276 24676 23304
rect 21416 23264 21422 23276
rect 24670 23264 24676 23276
rect 24728 23264 24734 23316
rect 36446 23304 36452 23316
rect 28966 23276 36452 23304
rect 2866 23196 2872 23248
rect 2924 23196 2930 23248
rect 23842 23196 23848 23248
rect 23900 23236 23906 23248
rect 26694 23236 26700 23248
rect 23900 23208 26700 23236
rect 23900 23196 23906 23208
rect 26694 23196 26700 23208
rect 26752 23236 26758 23248
rect 28966 23236 28994 23276
rect 36446 23264 36452 23276
rect 36504 23264 36510 23316
rect 36633 23307 36691 23313
rect 36633 23273 36645 23307
rect 36679 23304 36691 23307
rect 39114 23304 39120 23316
rect 36679 23276 39120 23304
rect 36679 23273 36691 23276
rect 36633 23267 36691 23273
rect 39114 23264 39120 23276
rect 39172 23264 39178 23316
rect 40221 23307 40279 23313
rect 40221 23273 40233 23307
rect 40267 23304 40279 23307
rect 40267 23276 40816 23304
rect 40267 23273 40279 23276
rect 40221 23267 40279 23273
rect 38013 23239 38071 23245
rect 38013 23236 38025 23239
rect 26752 23208 28994 23236
rect 33980 23208 38025 23236
rect 26752 23196 26758 23208
rect 2406 23128 2412 23180
rect 2464 23168 2470 23180
rect 31386 23168 31392 23180
rect 2464 23140 2544 23168
rect 2464 23128 2470 23140
rect 2516 23109 2544 23140
rect 30484 23140 31392 23168
rect 1581 23103 1639 23109
rect 1581 23069 1593 23103
rect 1627 23100 1639 23103
rect 2501 23103 2559 23109
rect 1627 23072 2452 23100
rect 1627 23069 1639 23072
rect 1581 23063 1639 23069
rect 934 22992 940 23044
rect 992 23032 998 23044
rect 1857 23035 1915 23041
rect 1857 23032 1869 23035
rect 992 23004 1869 23032
rect 992 22992 998 23004
rect 1857 23001 1869 23004
rect 1903 23001 1915 23035
rect 2424 23032 2452 23072
rect 2501 23069 2513 23103
rect 2547 23069 2559 23103
rect 2501 23063 2559 23069
rect 2655 23103 2713 23109
rect 2655 23069 2667 23103
rect 2701 23100 2713 23103
rect 3418 23100 3424 23112
rect 2701 23072 3424 23100
rect 2701 23069 2713 23072
rect 2655 23063 2713 23069
rect 3418 23060 3424 23072
rect 3476 23060 3482 23112
rect 29730 23060 29736 23112
rect 29788 23060 29794 23112
rect 30484 23109 30512 23140
rect 31386 23128 31392 23140
rect 31444 23128 31450 23180
rect 30469 23103 30527 23109
rect 30469 23069 30481 23103
rect 30515 23069 30527 23103
rect 30469 23063 30527 23069
rect 30650 23060 30656 23112
rect 30708 23060 30714 23112
rect 33229 23103 33287 23109
rect 33229 23069 33241 23103
rect 33275 23100 33287 23103
rect 33778 23100 33784 23112
rect 33275 23072 33784 23100
rect 33275 23069 33287 23072
rect 33229 23063 33287 23069
rect 33778 23060 33784 23072
rect 33836 23060 33842 23112
rect 33980 23109 34008 23208
rect 38013 23205 38025 23208
rect 38059 23205 38071 23239
rect 38013 23199 38071 23205
rect 36446 23128 36452 23180
rect 36504 23168 36510 23180
rect 37093 23171 37151 23177
rect 37093 23168 37105 23171
rect 36504 23140 37105 23168
rect 36504 23128 36510 23140
rect 37093 23137 37105 23140
rect 37139 23137 37151 23171
rect 37093 23131 37151 23137
rect 37185 23171 37243 23177
rect 37185 23137 37197 23171
rect 37231 23137 37243 23171
rect 39942 23168 39948 23180
rect 37185 23131 37243 23137
rect 37844 23140 39948 23168
rect 33965 23103 34023 23109
rect 33965 23069 33977 23103
rect 34011 23069 34023 23103
rect 33965 23063 34023 23069
rect 34882 23060 34888 23112
rect 34940 23060 34946 23112
rect 35894 23060 35900 23112
rect 35952 23060 35958 23112
rect 36814 23060 36820 23112
rect 36872 23100 36878 23112
rect 37200 23100 37228 23131
rect 37844 23109 37872 23140
rect 39942 23128 39948 23140
rect 40000 23128 40006 23180
rect 36872 23072 37228 23100
rect 37829 23103 37887 23109
rect 36872 23060 36878 23072
rect 37829 23069 37841 23103
rect 37875 23069 37887 23103
rect 37829 23063 37887 23069
rect 39117 23103 39175 23109
rect 39117 23069 39129 23103
rect 39163 23069 39175 23103
rect 39117 23063 39175 23069
rect 2774 23032 2780 23044
rect 2424 23004 2780 23032
rect 1857 22995 1915 23001
rect 2774 22992 2780 23004
rect 2832 22992 2838 23044
rect 29822 22992 29828 23044
rect 29880 23032 29886 23044
rect 30561 23035 30619 23041
rect 30561 23032 30573 23035
rect 29880 23004 30573 23032
rect 29880 22992 29886 23004
rect 30561 23001 30573 23004
rect 30607 23001 30619 23035
rect 30561 22995 30619 23001
rect 32766 22992 32772 23044
rect 32824 23032 32830 23044
rect 32824 23004 35112 23032
rect 32824 22992 32830 23004
rect 29546 22924 29552 22976
rect 29604 22964 29610 22976
rect 29917 22967 29975 22973
rect 29917 22964 29929 22967
rect 29604 22936 29929 22964
rect 29604 22924 29610 22936
rect 29917 22933 29929 22936
rect 29963 22933 29975 22967
rect 29917 22927 29975 22933
rect 33413 22967 33471 22973
rect 33413 22933 33425 22967
rect 33459 22964 33471 22967
rect 33502 22964 33508 22976
rect 33459 22936 33508 22964
rect 33459 22933 33471 22936
rect 33413 22927 33471 22933
rect 33502 22924 33508 22936
rect 33560 22924 33566 22976
rect 33686 22924 33692 22976
rect 33744 22964 33750 22976
rect 35084 22973 35112 23004
rect 35250 22992 35256 23044
rect 35308 23032 35314 23044
rect 36170 23032 36176 23044
rect 35308 23004 36176 23032
rect 35308 22992 35314 23004
rect 36170 22992 36176 23004
rect 36228 23032 36234 23044
rect 36906 23032 36912 23044
rect 36228 23004 36912 23032
rect 36228 22992 36234 23004
rect 36906 22992 36912 23004
rect 36964 23032 36970 23044
rect 37001 23035 37059 23041
rect 37001 23032 37013 23035
rect 36964 23004 37013 23032
rect 36964 22992 36970 23004
rect 37001 23001 37013 23004
rect 37047 23001 37059 23035
rect 37001 22995 37059 23001
rect 34149 22967 34207 22973
rect 34149 22964 34161 22967
rect 33744 22936 34161 22964
rect 33744 22924 33750 22936
rect 34149 22933 34161 22936
rect 34195 22933 34207 22967
rect 34149 22927 34207 22933
rect 35069 22967 35127 22973
rect 35069 22933 35081 22967
rect 35115 22933 35127 22967
rect 35069 22927 35127 22933
rect 35158 22924 35164 22976
rect 35216 22964 35222 22976
rect 36081 22967 36139 22973
rect 36081 22964 36093 22967
rect 35216 22936 36093 22964
rect 35216 22924 35222 22936
rect 36081 22933 36093 22936
rect 36127 22933 36139 22967
rect 36081 22927 36139 22933
rect 38838 22924 38844 22976
rect 38896 22924 38902 22976
rect 39132 22964 39160 23063
rect 39206 23060 39212 23112
rect 39264 23060 39270 23112
rect 39301 23103 39359 23109
rect 39301 23069 39313 23103
rect 39347 23069 39359 23103
rect 39301 23063 39359 23069
rect 39485 23103 39543 23109
rect 39485 23069 39497 23103
rect 39531 23100 39543 23103
rect 39574 23100 39580 23112
rect 39531 23072 39580 23100
rect 39531 23069 39543 23072
rect 39485 23063 39543 23069
rect 39316 23032 39344 23063
rect 39574 23060 39580 23072
rect 39632 23060 39638 23112
rect 40034 23060 40040 23112
rect 40092 23060 40098 23112
rect 40788 23109 40816 23276
rect 42886 23264 42892 23316
rect 42944 23264 42950 23316
rect 45738 23264 45744 23316
rect 45796 23304 45802 23316
rect 45796 23276 51074 23304
rect 45796 23264 45802 23276
rect 41414 23128 41420 23180
rect 41472 23168 41478 23180
rect 43438 23168 43444 23180
rect 41472 23140 43444 23168
rect 41472 23128 41478 23140
rect 43438 23128 43444 23140
rect 43496 23128 43502 23180
rect 51046 23168 51074 23276
rect 56505 23239 56563 23245
rect 56505 23205 56517 23239
rect 56551 23236 56563 23239
rect 56962 23236 56968 23248
rect 56551 23208 56968 23236
rect 56551 23205 56563 23208
rect 56505 23199 56563 23205
rect 56962 23196 56968 23208
rect 57020 23196 57026 23248
rect 51537 23171 51595 23177
rect 51537 23168 51549 23171
rect 51046 23140 51549 23168
rect 51537 23137 51549 23140
rect 51583 23168 51595 23171
rect 51902 23168 51908 23180
rect 51583 23140 51908 23168
rect 51583 23137 51595 23140
rect 51537 23131 51595 23137
rect 51902 23128 51908 23140
rect 51960 23128 51966 23180
rect 58250 23168 58256 23180
rect 56336 23140 58256 23168
rect 40773 23103 40831 23109
rect 40773 23069 40785 23103
rect 40819 23069 40831 23103
rect 40773 23063 40831 23069
rect 41874 23060 41880 23112
rect 41932 23060 41938 23112
rect 41966 23060 41972 23112
rect 42024 23060 42030 23112
rect 42058 23060 42064 23112
rect 42116 23060 42122 23112
rect 42242 23060 42248 23112
rect 42300 23060 42306 23112
rect 42518 23060 42524 23112
rect 42576 23100 42582 23112
rect 42705 23103 42763 23109
rect 42705 23100 42717 23103
rect 42576 23072 42717 23100
rect 42576 23060 42582 23072
rect 42705 23069 42717 23072
rect 42751 23069 42763 23103
rect 42705 23063 42763 23069
rect 48222 23060 48228 23112
rect 48280 23060 48286 23112
rect 48593 23103 48651 23109
rect 48593 23069 48605 23103
rect 48639 23100 48651 23103
rect 49234 23100 49240 23112
rect 48639 23072 49240 23100
rect 48639 23069 48651 23072
rect 48593 23063 48651 23069
rect 49234 23060 49240 23072
rect 49292 23060 49298 23112
rect 51626 23060 51632 23112
rect 51684 23100 51690 23112
rect 51721 23103 51779 23109
rect 51721 23100 51733 23103
rect 51684 23072 51733 23100
rect 51684 23060 51690 23072
rect 51721 23069 51733 23072
rect 51767 23069 51779 23103
rect 51721 23063 51779 23069
rect 55398 23060 55404 23112
rect 55456 23100 55462 23112
rect 56336 23109 56364 23140
rect 58250 23128 58256 23140
rect 58308 23128 58314 23180
rect 56137 23103 56195 23109
rect 56137 23100 56149 23103
rect 55456 23072 56149 23100
rect 55456 23060 55462 23072
rect 56137 23069 56149 23072
rect 56183 23069 56195 23103
rect 56137 23063 56195 23069
rect 56321 23103 56379 23109
rect 56321 23069 56333 23103
rect 56367 23069 56379 23103
rect 56965 23103 57023 23109
rect 56965 23100 56977 23103
rect 56321 23063 56379 23069
rect 56428 23072 56977 23100
rect 40126 23032 40132 23044
rect 39316 23004 40132 23032
rect 40126 22992 40132 23004
rect 40184 22992 40190 23044
rect 41138 23032 41144 23044
rect 40880 23004 41144 23032
rect 40880 22964 40908 23004
rect 41138 22992 41144 23004
rect 41196 23032 41202 23044
rect 41322 23032 41328 23044
rect 41196 23004 41328 23032
rect 41196 22992 41202 23004
rect 41322 22992 41328 23004
rect 41380 22992 41386 23044
rect 48314 22992 48320 23044
rect 48372 23032 48378 23044
rect 48409 23035 48467 23041
rect 48409 23032 48421 23035
rect 48372 23004 48421 23032
rect 48372 22992 48378 23004
rect 48409 23001 48421 23004
rect 48455 23001 48467 23035
rect 48409 22995 48467 23001
rect 48498 22992 48504 23044
rect 48556 22992 48562 23044
rect 53742 23032 53748 23044
rect 48608 23004 53748 23032
rect 39132 22936 40908 22964
rect 40957 22967 41015 22973
rect 40957 22933 40969 22967
rect 41003 22964 41015 22967
rect 41506 22964 41512 22976
rect 41003 22936 41512 22964
rect 41003 22933 41015 22936
rect 40957 22927 41015 22933
rect 41506 22924 41512 22936
rect 41564 22924 41570 22976
rect 41601 22967 41659 22973
rect 41601 22933 41613 22967
rect 41647 22964 41659 22967
rect 42334 22964 42340 22976
rect 41647 22936 42340 22964
rect 41647 22933 41659 22936
rect 41601 22927 41659 22933
rect 42334 22924 42340 22936
rect 42392 22924 42398 22976
rect 43806 22924 43812 22976
rect 43864 22964 43870 22976
rect 48608 22964 48636 23004
rect 53742 22992 53748 23004
rect 53800 22992 53806 23044
rect 53834 22992 53840 23044
rect 53892 23032 53898 23044
rect 56428 23032 56456 23072
rect 56965 23069 56977 23072
rect 57011 23069 57023 23103
rect 57885 23103 57943 23109
rect 57885 23100 57897 23103
rect 56965 23063 57023 23069
rect 57164 23072 57897 23100
rect 57164 23032 57192 23072
rect 57885 23069 57897 23072
rect 57931 23069 57943 23103
rect 57885 23063 57943 23069
rect 53892 23004 56456 23032
rect 56520 23004 57192 23032
rect 57241 23035 57299 23041
rect 53892 22992 53898 23004
rect 43864 22936 48636 22964
rect 43864 22924 43870 22936
rect 48682 22924 48688 22976
rect 48740 22964 48746 22976
rect 48777 22967 48835 22973
rect 48777 22964 48789 22967
rect 48740 22936 48789 22964
rect 48740 22924 48746 22936
rect 48777 22933 48789 22936
rect 48823 22933 48835 22967
rect 48777 22927 48835 22933
rect 51905 22967 51963 22973
rect 51905 22933 51917 22967
rect 51951 22964 51963 22967
rect 51994 22964 52000 22976
rect 51951 22936 52000 22964
rect 51951 22933 51963 22936
rect 51905 22927 51963 22933
rect 51994 22924 52000 22936
rect 52052 22924 52058 22976
rect 56410 22924 56416 22976
rect 56468 22964 56474 22976
rect 56520 22964 56548 23004
rect 57241 23001 57253 23035
rect 57287 23001 57299 23035
rect 57241 22995 57299 23001
rect 56468 22936 56548 22964
rect 57256 22964 57284 22995
rect 58158 22992 58164 23044
rect 58216 22992 58222 23044
rect 58986 22964 58992 22976
rect 57256 22936 58992 22964
rect 56468 22924 56474 22936
rect 58986 22924 58992 22936
rect 59044 22924 59050 22976
rect 1104 22874 58880 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 50294 22874
rect 50346 22822 50358 22874
rect 50410 22822 50422 22874
rect 50474 22822 50486 22874
rect 50538 22822 50550 22874
rect 50602 22822 58880 22874
rect 1104 22800 58880 22822
rect 2406 22720 2412 22772
rect 2464 22760 2470 22772
rect 2501 22763 2559 22769
rect 2501 22760 2513 22763
rect 2464 22732 2513 22760
rect 2464 22720 2470 22732
rect 2501 22729 2513 22732
rect 2547 22729 2559 22763
rect 2501 22723 2559 22729
rect 18506 22720 18512 22772
rect 18564 22760 18570 22772
rect 30190 22760 30196 22772
rect 18564 22732 30196 22760
rect 18564 22720 18570 22732
rect 30190 22720 30196 22732
rect 30248 22720 30254 22772
rect 33137 22763 33195 22769
rect 31726 22732 33088 22760
rect 22373 22695 22431 22701
rect 22373 22661 22385 22695
rect 22419 22692 22431 22695
rect 22462 22692 22468 22704
rect 22419 22664 22468 22692
rect 22419 22661 22431 22664
rect 22373 22655 22431 22661
rect 22462 22652 22468 22664
rect 22520 22652 22526 22704
rect 24118 22652 24124 22704
rect 24176 22692 24182 22704
rect 24762 22692 24768 22704
rect 24176 22664 24768 22692
rect 24176 22652 24182 22664
rect 24762 22652 24768 22664
rect 24820 22652 24826 22704
rect 31726 22692 31754 22732
rect 29472 22664 31754 22692
rect 2225 22627 2283 22633
rect 2225 22593 2237 22627
rect 2271 22624 2283 22627
rect 10502 22624 10508 22636
rect 2271 22596 10508 22624
rect 2271 22593 2283 22596
rect 2225 22587 2283 22593
rect 10502 22584 10508 22596
rect 10560 22584 10566 22636
rect 24394 22584 24400 22636
rect 24452 22624 24458 22636
rect 29472 22624 29500 22664
rect 24452 22596 29500 22624
rect 24452 22584 24458 22596
rect 29546 22584 29552 22636
rect 29604 22584 29610 22636
rect 30282 22584 30288 22636
rect 30340 22584 30346 22636
rect 32766 22584 32772 22636
rect 32824 22584 32830 22636
rect 31021 22559 31079 22565
rect 31021 22525 31033 22559
rect 31067 22556 31079 22559
rect 31570 22556 31576 22568
rect 31067 22528 31576 22556
rect 31067 22525 31079 22528
rect 31021 22519 31079 22525
rect 31570 22516 31576 22528
rect 31628 22556 31634 22568
rect 32677 22559 32735 22565
rect 32677 22556 32689 22559
rect 31628 22528 32689 22556
rect 31628 22516 31634 22528
rect 32677 22525 32689 22528
rect 32723 22525 32735 22559
rect 33060 22556 33088 22732
rect 33137 22729 33149 22763
rect 33183 22729 33195 22763
rect 33137 22723 33195 22729
rect 33152 22624 33180 22723
rect 33778 22720 33784 22772
rect 33836 22720 33842 22772
rect 34882 22720 34888 22772
rect 34940 22760 34946 22772
rect 37645 22763 37703 22769
rect 37645 22760 37657 22763
rect 34940 22732 37657 22760
rect 34940 22720 34946 22732
rect 37645 22729 37657 22732
rect 37691 22729 37703 22763
rect 37645 22723 37703 22729
rect 37734 22720 37740 22772
rect 37792 22760 37798 22772
rect 39942 22760 39948 22772
rect 37792 22732 39948 22760
rect 37792 22720 37798 22732
rect 39942 22720 39948 22732
rect 40000 22720 40006 22772
rect 40034 22720 40040 22772
rect 40092 22760 40098 22772
rect 40497 22763 40555 22769
rect 40497 22760 40509 22763
rect 40092 22732 40509 22760
rect 40092 22720 40098 22732
rect 40497 22729 40509 22732
rect 40543 22729 40555 22763
rect 40497 22723 40555 22729
rect 41598 22720 41604 22772
rect 41656 22760 41662 22772
rect 42610 22760 42616 22772
rect 41656 22732 42616 22760
rect 41656 22720 41662 22732
rect 42610 22720 42616 22732
rect 42668 22720 42674 22772
rect 42702 22720 42708 22772
rect 42760 22760 42766 22772
rect 42797 22763 42855 22769
rect 42797 22760 42809 22763
rect 42760 22732 42809 22760
rect 42760 22720 42766 22732
rect 42797 22729 42809 22732
rect 42843 22729 42855 22763
rect 44266 22760 44272 22772
rect 42797 22723 42855 22729
rect 43364 22732 44272 22760
rect 34701 22695 34759 22701
rect 34701 22661 34713 22695
rect 34747 22692 34759 22695
rect 35434 22692 35440 22704
rect 34747 22664 35440 22692
rect 34747 22661 34759 22664
rect 34701 22655 34759 22661
rect 35434 22652 35440 22664
rect 35492 22652 35498 22704
rect 38194 22692 38200 22704
rect 35544 22664 38200 22692
rect 33597 22627 33655 22633
rect 33597 22624 33609 22627
rect 33152 22596 33609 22624
rect 33597 22593 33609 22596
rect 33643 22593 33655 22627
rect 33597 22587 33655 22593
rect 34885 22627 34943 22633
rect 34885 22593 34897 22627
rect 34931 22624 34943 22627
rect 35250 22624 35256 22636
rect 34931 22596 35256 22624
rect 34931 22593 34943 22596
rect 34885 22587 34943 22593
rect 35250 22584 35256 22596
rect 35308 22584 35314 22636
rect 35544 22633 35572 22664
rect 38194 22652 38200 22664
rect 38252 22692 38258 22704
rect 38740 22695 38798 22701
rect 38252 22664 38516 22692
rect 38252 22652 38258 22664
rect 35529 22627 35587 22633
rect 35529 22593 35541 22627
rect 35575 22593 35587 22627
rect 35785 22627 35843 22633
rect 35785 22624 35797 22627
rect 35529 22587 35587 22593
rect 35636 22596 35797 22624
rect 35342 22556 35348 22568
rect 33060 22528 35348 22556
rect 32677 22519 32735 22525
rect 35342 22516 35348 22528
rect 35400 22516 35406 22568
rect 35434 22516 35440 22568
rect 35492 22556 35498 22568
rect 35636 22556 35664 22596
rect 35785 22593 35797 22596
rect 35831 22593 35843 22627
rect 35785 22587 35843 22593
rect 36078 22584 36084 22636
rect 36136 22624 36142 22636
rect 36136 22596 37412 22624
rect 36136 22584 36142 22596
rect 35492 22528 35664 22556
rect 37384 22556 37412 22596
rect 37458 22584 37464 22636
rect 37516 22584 37522 22636
rect 38488 22633 38516 22664
rect 38740 22661 38752 22695
rect 38786 22692 38798 22695
rect 38838 22692 38844 22704
rect 38786 22664 38844 22692
rect 38786 22661 38798 22664
rect 38740 22655 38798 22661
rect 38838 22652 38844 22664
rect 38896 22652 38902 22704
rect 40954 22692 40960 22704
rect 39776 22664 40960 22692
rect 38473 22627 38531 22633
rect 38473 22593 38485 22627
rect 38519 22593 38531 22627
rect 39776 22624 39804 22664
rect 40954 22652 40960 22664
rect 41012 22652 41018 22704
rect 43364 22692 43392 22732
rect 44266 22720 44272 22732
rect 44324 22720 44330 22772
rect 44358 22720 44364 22772
rect 44416 22760 44422 22772
rect 45465 22763 45523 22769
rect 45465 22760 45477 22763
rect 44416 22732 45477 22760
rect 44416 22720 44422 22732
rect 45465 22729 45477 22732
rect 45511 22760 45523 22763
rect 46569 22763 46627 22769
rect 46569 22760 46581 22763
rect 45511 22732 46581 22760
rect 45511 22729 45523 22732
rect 45465 22723 45523 22729
rect 46569 22729 46581 22732
rect 46615 22729 46627 22763
rect 46569 22723 46627 22729
rect 46658 22720 46664 22772
rect 46716 22760 46722 22772
rect 48038 22760 48044 22772
rect 46716 22732 48044 22760
rect 46716 22720 46722 22732
rect 48038 22720 48044 22732
rect 48096 22720 48102 22772
rect 48498 22720 48504 22772
rect 48556 22760 48562 22772
rect 49786 22760 49792 22772
rect 48556 22732 49792 22760
rect 48556 22720 48562 22732
rect 49786 22720 49792 22732
rect 49844 22760 49850 22772
rect 49881 22763 49939 22769
rect 49881 22760 49893 22763
rect 49844 22732 49893 22760
rect 49844 22720 49850 22732
rect 49881 22729 49893 22732
rect 49927 22729 49939 22763
rect 49881 22723 49939 22729
rect 49988 22732 51580 22760
rect 41708 22664 41920 22692
rect 40313 22627 40371 22633
rect 40313 22624 40325 22627
rect 38473 22587 38531 22593
rect 38580 22596 39804 22624
rect 39868 22596 40325 22624
rect 38580 22556 38608 22596
rect 37384 22528 38608 22556
rect 35492 22516 35498 22528
rect 31389 22491 31447 22497
rect 31389 22457 31401 22491
rect 31435 22488 31447 22491
rect 32214 22488 32220 22500
rect 31435 22460 32220 22488
rect 31435 22457 31447 22460
rect 31389 22451 31447 22457
rect 32214 22448 32220 22460
rect 32272 22448 32278 22500
rect 36906 22448 36912 22500
rect 36964 22448 36970 22500
rect 29733 22423 29791 22429
rect 29733 22389 29745 22423
rect 29779 22420 29791 22423
rect 30006 22420 30012 22432
rect 29779 22392 30012 22420
rect 29779 22389 29791 22392
rect 29733 22383 29791 22389
rect 30006 22380 30012 22392
rect 30064 22380 30070 22432
rect 30374 22380 30380 22432
rect 30432 22420 30438 22432
rect 30469 22423 30527 22429
rect 30469 22420 30481 22423
rect 30432 22392 30481 22420
rect 30432 22380 30438 22392
rect 30469 22389 30481 22392
rect 30515 22389 30527 22423
rect 30469 22383 30527 22389
rect 31481 22423 31539 22429
rect 31481 22389 31493 22423
rect 31527 22420 31539 22423
rect 32766 22420 32772 22432
rect 31527 22392 32772 22420
rect 31527 22389 31539 22392
rect 31481 22383 31539 22389
rect 32766 22380 32772 22392
rect 32824 22380 32830 22432
rect 35069 22423 35127 22429
rect 35069 22389 35081 22423
rect 35115 22420 35127 22423
rect 35894 22420 35900 22432
rect 35115 22392 35900 22420
rect 35115 22389 35127 22392
rect 35069 22383 35127 22389
rect 35894 22380 35900 22392
rect 35952 22380 35958 22432
rect 38838 22380 38844 22432
rect 38896 22420 38902 22432
rect 39868 22429 39896 22596
rect 40313 22593 40325 22596
rect 40359 22593 40371 22627
rect 40313 22587 40371 22593
rect 41598 22584 41604 22636
rect 41656 22584 41662 22636
rect 41708 22633 41736 22664
rect 41693 22627 41751 22633
rect 41693 22593 41705 22627
rect 41739 22593 41751 22627
rect 41693 22587 41751 22593
rect 41785 22627 41843 22633
rect 41785 22593 41797 22627
rect 41831 22593 41843 22627
rect 41785 22587 41843 22593
rect 41322 22516 41328 22568
rect 41380 22556 41386 22568
rect 41800 22556 41828 22587
rect 41380 22528 41828 22556
rect 41892 22556 41920 22664
rect 42260 22664 43392 22692
rect 42260 22636 42288 22664
rect 43438 22652 43444 22704
rect 43496 22692 43502 22704
rect 49988 22692 50016 22732
rect 51552 22692 51580 22732
rect 51626 22720 51632 22772
rect 51684 22720 51690 22772
rect 53742 22720 53748 22772
rect 53800 22760 53806 22772
rect 58253 22763 58311 22769
rect 58253 22760 58265 22763
rect 53800 22732 58265 22760
rect 53800 22720 53806 22732
rect 58253 22729 58265 22732
rect 58299 22729 58311 22763
rect 58253 22723 58311 22729
rect 57974 22692 57980 22704
rect 43496 22664 50016 22692
rect 50080 22664 51488 22692
rect 51552 22664 57980 22692
rect 43496 22652 43502 22664
rect 41969 22627 42027 22633
rect 41969 22593 41981 22627
rect 42015 22624 42027 22627
rect 42242 22624 42248 22636
rect 42015 22596 42248 22624
rect 42015 22593 42027 22596
rect 41969 22587 42027 22593
rect 42242 22584 42248 22596
rect 42300 22584 42306 22636
rect 42613 22627 42671 22633
rect 42613 22593 42625 22627
rect 42659 22624 42671 22627
rect 42702 22624 42708 22636
rect 42659 22596 42708 22624
rect 42659 22593 42671 22596
rect 42613 22587 42671 22593
rect 42702 22584 42708 22596
rect 42760 22584 42766 22636
rect 43346 22584 43352 22636
rect 43404 22584 43410 22636
rect 44174 22584 44180 22636
rect 44232 22624 44238 22636
rect 48774 22633 48780 22636
rect 44341 22627 44399 22633
rect 44341 22624 44353 22627
rect 44232 22596 44353 22624
rect 44232 22584 44238 22596
rect 44341 22593 44353 22596
rect 44387 22593 44399 22627
rect 44341 22587 44399 22593
rect 48768 22587 48780 22633
rect 48774 22584 48780 22587
rect 48832 22584 48838 22636
rect 49234 22584 49240 22636
rect 49292 22624 49298 22636
rect 50080 22624 50108 22664
rect 49292 22596 50108 22624
rect 49292 22584 49298 22596
rect 51074 22584 51080 22636
rect 51132 22584 51138 22636
rect 51460 22633 51488 22664
rect 57974 22652 57980 22664
rect 58032 22652 58038 22704
rect 51261 22627 51319 22633
rect 51261 22593 51273 22627
rect 51307 22593 51319 22627
rect 51261 22587 51319 22593
rect 51353 22627 51411 22633
rect 51353 22593 51365 22627
rect 51399 22593 51411 22627
rect 51353 22587 51411 22593
rect 51445 22627 51503 22633
rect 51445 22593 51457 22627
rect 51491 22624 51503 22627
rect 51718 22624 51724 22636
rect 51491 22596 51724 22624
rect 51491 22593 51503 22596
rect 51445 22587 51503 22593
rect 41892 22528 44036 22556
rect 41380 22516 41386 22528
rect 41414 22448 41420 22500
rect 41472 22488 41478 22500
rect 42518 22488 42524 22500
rect 41472 22460 42524 22488
rect 41472 22448 41478 22460
rect 42518 22448 42524 22460
rect 42576 22448 42582 22500
rect 39853 22423 39911 22429
rect 39853 22420 39865 22423
rect 38896 22392 39865 22420
rect 38896 22380 38902 22392
rect 39853 22389 39865 22392
rect 39899 22389 39911 22423
rect 39853 22383 39911 22389
rect 41325 22423 41383 22429
rect 41325 22389 41337 22423
rect 41371 22420 41383 22423
rect 42702 22420 42708 22432
rect 41371 22392 42708 22420
rect 41371 22389 41383 22392
rect 41325 22383 41383 22389
rect 42702 22380 42708 22392
rect 42760 22380 42766 22432
rect 43530 22380 43536 22432
rect 43588 22380 43594 22432
rect 44008 22420 44036 22528
rect 44082 22516 44088 22568
rect 44140 22516 44146 22568
rect 46566 22516 46572 22568
rect 46624 22556 46630 22568
rect 46753 22559 46811 22565
rect 46753 22556 46765 22559
rect 46624 22528 46765 22556
rect 46624 22516 46630 22528
rect 46753 22525 46765 22528
rect 46799 22556 46811 22559
rect 46842 22556 46848 22568
rect 46799 22528 46848 22556
rect 46799 22525 46811 22528
rect 46753 22519 46811 22525
rect 46842 22516 46848 22528
rect 46900 22516 46906 22568
rect 48406 22516 48412 22568
rect 48464 22556 48470 22568
rect 48501 22559 48559 22565
rect 48501 22556 48513 22559
rect 48464 22528 48513 22556
rect 48464 22516 48470 22528
rect 48501 22525 48513 22528
rect 48547 22525 48559 22559
rect 48501 22519 48559 22525
rect 51276 22488 51304 22587
rect 51368 22556 51396 22587
rect 51718 22584 51724 22596
rect 51776 22584 51782 22636
rect 53006 22624 53012 22636
rect 51828 22596 53012 22624
rect 51828 22556 51856 22596
rect 53006 22584 53012 22596
rect 53064 22584 53070 22636
rect 53101 22627 53159 22633
rect 53101 22593 53113 22627
rect 53147 22624 53159 22627
rect 54110 22624 54116 22636
rect 53147 22596 54116 22624
rect 53147 22593 53159 22596
rect 53101 22587 53159 22593
rect 54110 22584 54116 22596
rect 54168 22584 54174 22636
rect 56229 22627 56287 22633
rect 56229 22593 56241 22627
rect 56275 22624 56287 22627
rect 56318 22624 56324 22636
rect 56275 22596 56324 22624
rect 56275 22593 56287 22596
rect 56229 22587 56287 22593
rect 56318 22584 56324 22596
rect 56376 22584 56382 22636
rect 58066 22584 58072 22636
rect 58124 22584 58130 22636
rect 51368 22528 51856 22556
rect 51902 22516 51908 22568
rect 51960 22556 51966 22568
rect 52917 22559 52975 22565
rect 52917 22556 52929 22559
rect 51960 22528 52929 22556
rect 51960 22516 51966 22528
rect 52917 22525 52929 22528
rect 52963 22556 52975 22559
rect 55398 22556 55404 22568
rect 52963 22528 55404 22556
rect 52963 22525 52975 22528
rect 52917 22519 52975 22525
rect 55398 22516 55404 22528
rect 55456 22516 55462 22568
rect 56410 22516 56416 22568
rect 56468 22556 56474 22568
rect 56505 22559 56563 22565
rect 56505 22556 56517 22559
rect 56468 22528 56517 22556
rect 56468 22516 56474 22528
rect 56505 22525 56517 22528
rect 56551 22525 56563 22559
rect 56505 22519 56563 22525
rect 53006 22488 53012 22500
rect 51276 22460 53012 22488
rect 53006 22448 53012 22460
rect 53064 22448 53070 22500
rect 55214 22488 55220 22500
rect 53116 22460 55220 22488
rect 45554 22420 45560 22432
rect 44008 22392 45560 22420
rect 45554 22380 45560 22392
rect 45612 22380 45618 22432
rect 46201 22423 46259 22429
rect 46201 22389 46213 22423
rect 46247 22420 46259 22423
rect 49142 22420 49148 22432
rect 46247 22392 49148 22420
rect 46247 22389 46259 22392
rect 46201 22383 46259 22389
rect 49142 22380 49148 22392
rect 49200 22380 49206 22432
rect 49786 22380 49792 22432
rect 49844 22420 49850 22432
rect 53116 22420 53144 22460
rect 55214 22448 55220 22460
rect 55272 22448 55278 22500
rect 49844 22392 53144 22420
rect 49844 22380 49850 22392
rect 53282 22380 53288 22432
rect 53340 22380 53346 22432
rect 1104 22330 58880 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 58880 22330
rect 1104 22256 58880 22278
rect 2685 22219 2743 22225
rect 2685 22185 2697 22219
rect 2731 22216 2743 22219
rect 2774 22216 2780 22228
rect 2731 22188 2780 22216
rect 2731 22185 2743 22188
rect 2685 22179 2743 22185
rect 2774 22176 2780 22188
rect 2832 22176 2838 22228
rect 29089 22219 29147 22225
rect 29089 22185 29101 22219
rect 29135 22216 29147 22219
rect 29730 22216 29736 22228
rect 29135 22188 29736 22216
rect 29135 22185 29147 22188
rect 29089 22179 29147 22185
rect 29730 22176 29736 22188
rect 29788 22176 29794 22228
rect 30834 22176 30840 22228
rect 30892 22216 30898 22228
rect 30892 22188 31524 22216
rect 30892 22176 30898 22188
rect 22189 22151 22247 22157
rect 22189 22148 22201 22151
rect 13832 22120 22201 22148
rect 934 22040 940 22092
rect 992 22080 998 22092
rect 1765 22083 1823 22089
rect 1765 22080 1777 22083
rect 992 22052 1777 22080
rect 992 22040 998 22052
rect 1765 22049 1777 22052
rect 1811 22049 1823 22083
rect 13832 22080 13860 22120
rect 22189 22117 22201 22120
rect 22235 22117 22247 22151
rect 22189 22111 22247 22117
rect 31110 22108 31116 22160
rect 31168 22148 31174 22160
rect 31386 22148 31392 22160
rect 31168 22120 31392 22148
rect 31168 22108 31174 22120
rect 31386 22108 31392 22120
rect 31444 22108 31450 22160
rect 1765 22043 1823 22049
rect 2424 22052 13860 22080
rect 1581 22015 1639 22021
rect 1581 21981 1593 22015
rect 1627 22012 1639 22015
rect 2424 22012 2452 22052
rect 23474 22040 23480 22092
rect 23532 22080 23538 22092
rect 28074 22080 28080 22092
rect 23532 22052 28080 22080
rect 23532 22040 23538 22052
rect 28074 22040 28080 22052
rect 28132 22040 28138 22092
rect 31496 22080 31524 22188
rect 31570 22176 31576 22228
rect 31628 22176 31634 22228
rect 32214 22176 32220 22228
rect 32272 22176 32278 22228
rect 35434 22176 35440 22228
rect 35492 22176 35498 22228
rect 37734 22216 37740 22228
rect 35728 22188 37740 22216
rect 32950 22108 32956 22160
rect 33008 22148 33014 22160
rect 35728 22148 35756 22188
rect 37734 22176 37740 22188
rect 37792 22176 37798 22228
rect 38102 22176 38108 22228
rect 38160 22216 38166 22228
rect 39850 22216 39856 22228
rect 38160 22188 39856 22216
rect 38160 22176 38166 22188
rect 39850 22176 39856 22188
rect 39908 22176 39914 22228
rect 48774 22176 48780 22228
rect 48832 22216 48838 22228
rect 48869 22219 48927 22225
rect 48869 22216 48881 22219
rect 48832 22188 48881 22216
rect 48832 22176 48838 22188
rect 48869 22185 48881 22188
rect 48915 22185 48927 22219
rect 48869 22179 48927 22185
rect 49142 22176 49148 22228
rect 49200 22216 49206 22228
rect 49200 22188 53052 22216
rect 49200 22176 49206 22188
rect 35802 22148 35808 22160
rect 33008 22120 35756 22148
rect 33008 22108 33014 22120
rect 35801 22108 35808 22148
rect 35860 22108 35866 22160
rect 38746 22108 38752 22160
rect 38804 22108 38810 22160
rect 38930 22108 38936 22160
rect 38988 22108 38994 22160
rect 39114 22108 39120 22160
rect 39172 22148 39178 22160
rect 47121 22151 47179 22157
rect 39172 22120 39344 22148
rect 39172 22108 39178 22120
rect 33686 22080 33692 22092
rect 31312 22052 33692 22080
rect 1627 21984 2452 22012
rect 1627 21981 1639 21984
rect 1581 21975 1639 21981
rect 2498 21972 2504 22024
rect 2556 21972 2562 22024
rect 2590 21972 2596 22024
rect 2648 22012 2654 22024
rect 2648 21984 6914 22012
rect 2648 21972 2654 21984
rect 6886 21876 6914 21984
rect 10134 21972 10140 22024
rect 10192 22012 10198 22024
rect 10502 22012 10508 22024
rect 10192 21984 10508 22012
rect 10192 21972 10198 21984
rect 10502 21972 10508 21984
rect 10560 22012 10566 22024
rect 22002 22012 22008 22024
rect 10560 21984 22008 22012
rect 10560 21972 10566 21984
rect 22002 21972 22008 21984
rect 22060 21972 22066 22024
rect 22465 22015 22523 22021
rect 22465 21981 22477 22015
rect 22511 22012 22523 22015
rect 24118 22012 24124 22024
rect 22511 21984 24124 22012
rect 22511 21981 22523 21984
rect 22465 21975 22523 21981
rect 24118 21972 24124 21984
rect 24176 21972 24182 22024
rect 26237 22015 26295 22021
rect 26237 21981 26249 22015
rect 26283 22012 26295 22015
rect 26602 22012 26608 22024
rect 26283 21984 26608 22012
rect 26283 21981 26295 21984
rect 26237 21975 26295 21981
rect 26602 21972 26608 21984
rect 26660 21972 26666 22024
rect 27985 22015 28043 22021
rect 27985 21981 27997 22015
rect 28031 22012 28043 22015
rect 28258 22012 28264 22024
rect 28031 21984 28264 22012
rect 28031 21981 28043 21984
rect 27985 21975 28043 21981
rect 28258 21972 28264 21984
rect 28316 21972 28322 22024
rect 28905 22015 28963 22021
rect 28905 21981 28917 22015
rect 28951 22012 28963 22015
rect 29270 22012 29276 22024
rect 28951 21984 29276 22012
rect 28951 21981 28963 21984
rect 28905 21975 28963 21981
rect 29270 21972 29276 21984
rect 29328 21972 29334 22024
rect 30285 22015 30343 22021
rect 30285 21981 30297 22015
rect 30331 22012 30343 22015
rect 30926 22012 30932 22024
rect 30331 21984 30932 22012
rect 30331 21981 30343 21984
rect 30285 21975 30343 21981
rect 30926 21972 30932 21984
rect 30984 21972 30990 22024
rect 31205 22015 31263 22021
rect 31205 21981 31217 22015
rect 31251 22012 31263 22015
rect 31312 22012 31340 22052
rect 33686 22040 33692 22052
rect 33744 22040 33750 22092
rect 31251 21984 31340 22012
rect 31251 21981 31263 21984
rect 31205 21975 31263 21981
rect 31386 21972 31392 22024
rect 31444 21972 31450 22024
rect 32033 22015 32091 22021
rect 32033 22012 32045 22015
rect 31496 21984 32045 22012
rect 31018 21904 31024 21956
rect 31076 21904 31082 21956
rect 31496 21944 31524 21984
rect 32033 21981 32045 21984
rect 32079 21981 32091 22015
rect 32033 21975 32091 21981
rect 32766 21972 32772 22024
rect 32824 21972 32830 22024
rect 33042 21972 33048 22024
rect 33100 22012 33106 22024
rect 33505 22015 33563 22021
rect 33505 22012 33517 22015
rect 33100 21984 33517 22012
rect 33100 21972 33106 21984
rect 33505 21981 33517 21984
rect 33551 22012 33563 22015
rect 34790 22012 34796 22024
rect 33551 21984 34796 22012
rect 33551 21981 33563 21984
rect 33505 21975 33563 21981
rect 34790 21972 34796 21984
rect 34848 21972 34854 22024
rect 35801 22021 35829 22108
rect 38948 22080 38976 22108
rect 38948 22052 39160 22080
rect 35693 22015 35751 22021
rect 35693 22012 35705 22015
rect 35636 21984 35705 22012
rect 31225 21916 31524 21944
rect 31680 21916 33732 21944
rect 23934 21876 23940 21888
rect 6886 21848 23940 21876
rect 23934 21836 23940 21848
rect 23992 21836 23998 21888
rect 25222 21836 25228 21888
rect 25280 21876 25286 21888
rect 26421 21879 26479 21885
rect 26421 21876 26433 21879
rect 25280 21848 26433 21876
rect 25280 21836 25286 21848
rect 26421 21845 26433 21848
rect 26467 21845 26479 21879
rect 26421 21839 26479 21845
rect 28166 21836 28172 21888
rect 28224 21836 28230 21888
rect 30469 21879 30527 21885
rect 30469 21845 30481 21879
rect 30515 21876 30527 21879
rect 31225 21876 31253 21916
rect 30515 21848 31253 21876
rect 31297 21879 31355 21885
rect 30515 21845 30527 21848
rect 30469 21839 30527 21845
rect 31297 21845 31309 21879
rect 31343 21876 31355 21879
rect 31386 21876 31392 21888
rect 31343 21848 31392 21876
rect 31343 21845 31355 21848
rect 31297 21839 31355 21845
rect 31386 21836 31392 21848
rect 31444 21876 31450 21888
rect 31680 21876 31708 21916
rect 31444 21848 31708 21876
rect 31444 21836 31450 21848
rect 32858 21836 32864 21888
rect 32916 21876 32922 21888
rect 33704 21885 33732 21916
rect 32953 21879 33011 21885
rect 32953 21876 32965 21879
rect 32916 21848 32965 21876
rect 32916 21836 32922 21848
rect 32953 21845 32965 21848
rect 32999 21845 33011 21879
rect 32953 21839 33011 21845
rect 33689 21879 33747 21885
rect 33689 21845 33701 21879
rect 33735 21845 33747 21879
rect 35636 21876 35664 21984
rect 35693 21981 35705 21984
rect 35739 21981 35751 22015
rect 35801 22015 35863 22021
rect 35801 21986 35817 22015
rect 35693 21975 35751 21981
rect 35805 21981 35817 21986
rect 35851 21981 35863 22015
rect 35805 21975 35863 21981
rect 35894 21972 35900 22024
rect 35952 22018 35958 22024
rect 35952 22012 35976 22018
rect 35964 21978 35976 22012
rect 35952 21972 35976 21978
rect 36081 22015 36139 22021
rect 36081 21981 36093 22015
rect 36127 22012 36139 22015
rect 36262 22012 36268 22024
rect 36127 21984 36268 22012
rect 36127 21981 36139 21984
rect 36081 21975 36139 21981
rect 36262 21972 36268 21984
rect 36320 21972 36326 22024
rect 36541 22015 36599 22021
rect 36541 21981 36553 22015
rect 36587 22012 36599 22015
rect 36906 22012 36912 22024
rect 36587 21984 36912 22012
rect 36587 21981 36599 21984
rect 36541 21975 36599 21981
rect 36906 21972 36912 21984
rect 36964 21972 36970 22024
rect 37277 22015 37335 22021
rect 37277 21981 37289 22015
rect 37323 21981 37335 22015
rect 37277 21975 37335 21981
rect 37921 22015 37979 22021
rect 37921 21981 37933 22015
rect 37967 22012 37979 22015
rect 37967 22006 38654 22012
rect 38746 22006 38752 22024
rect 37967 21984 38752 22006
rect 37967 21981 37979 21984
rect 37921 21975 37979 21981
rect 38626 21978 38752 21984
rect 37090 21944 37096 21956
rect 36280 21916 37096 21944
rect 36280 21876 36308 21916
rect 37090 21904 37096 21916
rect 37148 21904 37154 21956
rect 37292 21944 37320 21975
rect 38746 21972 38752 21978
rect 38804 21972 38810 22024
rect 39022 21972 39028 22024
rect 39080 21972 39086 22024
rect 39132 22015 39160 22052
rect 39230 22015 39288 22021
rect 39114 22009 39172 22015
rect 39114 21975 39126 22009
rect 39160 21975 39172 22009
rect 39230 21981 39242 22015
rect 39276 22012 39288 22015
rect 39316 22012 39344 22120
rect 47121 22117 47133 22151
rect 47167 22148 47179 22151
rect 47167 22120 47201 22148
rect 47167 22117 47179 22120
rect 47121 22111 47179 22117
rect 39666 22040 39672 22092
rect 39724 22080 39730 22092
rect 42061 22083 42119 22089
rect 42061 22080 42073 22083
rect 39724 22052 42073 22080
rect 39724 22040 39730 22052
rect 42061 22049 42073 22052
rect 42107 22080 42119 22083
rect 42794 22080 42800 22092
rect 42107 22052 42800 22080
rect 42107 22049 42119 22052
rect 42061 22043 42119 22049
rect 42794 22040 42800 22052
rect 42852 22040 42858 22092
rect 43441 22083 43499 22089
rect 43441 22049 43453 22083
rect 43487 22049 43499 22083
rect 47136 22080 47164 22111
rect 51718 22108 51724 22160
rect 51776 22108 51782 22160
rect 53024 22148 53052 22188
rect 53098 22176 53104 22228
rect 53156 22176 53162 22228
rect 54110 22176 54116 22228
rect 54168 22176 54174 22228
rect 57146 22216 57152 22228
rect 54220 22188 57152 22216
rect 54220 22148 54248 22188
rect 57146 22176 57152 22188
rect 57204 22176 57210 22228
rect 58250 22176 58256 22228
rect 58308 22176 58314 22228
rect 53024 22120 54248 22148
rect 47136 22052 47624 22080
rect 43441 22043 43499 22049
rect 39276 21984 39344 22012
rect 39393 22015 39451 22021
rect 39276 21981 39288 21984
rect 39230 21975 39288 21981
rect 39393 21981 39405 22015
rect 39439 22012 39451 22015
rect 39574 22012 39580 22024
rect 39439 21984 39580 22012
rect 39439 21981 39451 21984
rect 39393 21975 39451 21981
rect 39114 21969 39172 21975
rect 39574 21972 39580 21984
rect 39632 21972 39638 22024
rect 39850 21972 39856 22024
rect 39908 22012 39914 22024
rect 40037 22015 40095 22021
rect 40037 22012 40049 22015
rect 39908 21984 40049 22012
rect 39908 21972 39914 21984
rect 40037 21981 40049 21984
rect 40083 22012 40095 22015
rect 40494 22012 40500 22024
rect 40083 21984 40500 22012
rect 40083 21981 40095 21984
rect 40037 21975 40095 21981
rect 40494 21972 40500 21984
rect 40552 21972 40558 22024
rect 41322 21972 41328 22024
rect 41380 21972 41386 22024
rect 42334 21972 42340 22024
rect 42392 21972 42398 22024
rect 42610 21972 42616 22024
rect 42668 22012 42674 22024
rect 43456 22012 43484 22043
rect 42668 21984 43484 22012
rect 42668 21972 42674 21984
rect 44082 21972 44088 22024
rect 44140 22012 44146 22024
rect 44634 22012 44640 22024
rect 44140 21984 44640 22012
rect 44140 21972 44146 21984
rect 44634 21972 44640 21984
rect 44692 22012 44698 22024
rect 45189 22015 45247 22021
rect 45189 22012 45201 22015
rect 44692 21984 45201 22012
rect 44692 21972 44698 21984
rect 45189 21981 45201 21984
rect 45235 21981 45247 22015
rect 47596 22012 47624 22052
rect 47670 22040 47676 22092
rect 47728 22040 47734 22092
rect 51074 22080 51080 22092
rect 48424 22052 51080 22080
rect 48424 22012 48452 22052
rect 51074 22040 51080 22052
rect 51132 22040 51138 22092
rect 51736 22080 51764 22108
rect 51644 22052 51764 22080
rect 47596 21984 48452 22012
rect 45189 21975 45247 21981
rect 48590 21972 48596 22024
rect 48648 21972 48654 22024
rect 48682 21972 48688 22024
rect 48740 21972 48746 22024
rect 37292 21916 38056 21944
rect 35636 21848 36308 21876
rect 33689 21839 33747 21845
rect 36630 21836 36636 21888
rect 36688 21876 36694 21888
rect 36725 21879 36783 21885
rect 36725 21876 36737 21879
rect 36688 21848 36737 21876
rect 36688 21836 36694 21848
rect 36725 21845 36737 21848
rect 36771 21845 36783 21879
rect 36725 21839 36783 21845
rect 37369 21879 37427 21885
rect 37369 21845 37381 21879
rect 37415 21876 37427 21879
rect 37642 21876 37648 21888
rect 37415 21848 37648 21876
rect 37415 21845 37427 21848
rect 37369 21839 37427 21845
rect 37642 21836 37648 21848
rect 37700 21836 37706 21888
rect 38028 21876 38056 21916
rect 38102 21904 38108 21956
rect 38160 21904 38166 21956
rect 38289 21947 38347 21953
rect 38289 21913 38301 21947
rect 38335 21944 38347 21947
rect 38335 21916 38884 21944
rect 38335 21913 38347 21916
rect 38289 21907 38347 21913
rect 38562 21876 38568 21888
rect 38028 21848 38568 21876
rect 38562 21836 38568 21848
rect 38620 21836 38626 21888
rect 38856 21876 38884 21916
rect 40402 21904 40408 21956
rect 40460 21944 40466 21956
rect 40957 21947 41015 21953
rect 40957 21944 40969 21947
rect 40460 21916 40969 21944
rect 40460 21904 40466 21916
rect 40957 21913 40969 21916
rect 41003 21913 41015 21947
rect 40957 21907 41015 21913
rect 41141 21947 41199 21953
rect 41141 21913 41153 21947
rect 41187 21944 41199 21947
rect 41414 21944 41420 21956
rect 41187 21916 41420 21944
rect 41187 21913 41199 21916
rect 41141 21907 41199 21913
rect 41414 21904 41420 21916
rect 41472 21904 41478 21956
rect 43438 21904 43444 21956
rect 43496 21944 43502 21956
rect 44177 21947 44235 21953
rect 44177 21944 44189 21947
rect 43496 21916 44189 21944
rect 43496 21904 43502 21916
rect 44177 21913 44189 21916
rect 44223 21913 44235 21947
rect 44177 21907 44235 21913
rect 44358 21904 44364 21956
rect 44416 21904 44422 21956
rect 45278 21904 45284 21956
rect 45336 21944 45342 21956
rect 45434 21947 45492 21953
rect 45434 21944 45446 21947
rect 45336 21916 45446 21944
rect 45336 21904 45342 21916
rect 45434 21913 45446 21916
rect 45480 21913 45492 21947
rect 47489 21947 47547 21953
rect 47489 21944 47501 21947
rect 45434 21907 45492 21913
rect 46584 21916 47501 21944
rect 46584 21888 46612 21916
rect 47489 21913 47501 21916
rect 47535 21913 47547 21947
rect 47489 21907 47547 21913
rect 47581 21947 47639 21953
rect 47581 21913 47593 21947
rect 47627 21944 47639 21947
rect 47854 21944 47860 21956
rect 47627 21916 47860 21944
rect 47627 21913 47639 21916
rect 47581 21907 47639 21913
rect 47854 21904 47860 21916
rect 47912 21904 47918 21956
rect 39114 21876 39120 21888
rect 38856 21848 39120 21876
rect 39114 21836 39120 21848
rect 39172 21836 39178 21888
rect 40218 21836 40224 21888
rect 40276 21836 40282 21888
rect 41598 21836 41604 21888
rect 41656 21876 41662 21888
rect 43346 21876 43352 21888
rect 41656 21848 43352 21876
rect 41656 21836 41662 21848
rect 43346 21836 43352 21848
rect 43404 21836 43410 21888
rect 44542 21836 44548 21888
rect 44600 21836 44606 21888
rect 46566 21836 46572 21888
rect 46624 21836 46630 21888
rect 51644 21876 51672 22052
rect 53006 22040 53012 22092
rect 53064 22080 53070 22092
rect 53742 22080 53748 22092
rect 53064 22052 53748 22080
rect 53064 22040 53070 22052
rect 53742 22040 53748 22052
rect 53800 22040 53806 22092
rect 54018 22040 54024 22092
rect 54076 22080 54082 22092
rect 54076 22052 54248 22080
rect 54076 22040 54082 22052
rect 54220 22024 54248 22052
rect 57054 22040 57060 22092
rect 57112 22080 57118 22092
rect 57790 22080 57796 22092
rect 57112 22052 57796 22080
rect 57112 22040 57118 22052
rect 57790 22040 57796 22052
rect 57848 22080 57854 22092
rect 57848 22052 58020 22080
rect 57848 22040 57854 22052
rect 51721 22015 51779 22021
rect 51721 21981 51733 22015
rect 51767 22012 51779 22015
rect 52362 22012 52368 22024
rect 51767 21984 52368 22012
rect 51767 21981 51779 21984
rect 51721 21975 51779 21981
rect 52362 21972 52368 21984
rect 52420 21972 52426 22024
rect 53558 21972 53564 22024
rect 53616 21972 53622 22024
rect 53926 22012 53932 22024
rect 53668 21984 53932 22012
rect 51994 21953 52000 21956
rect 51988 21907 52000 21953
rect 51994 21904 52000 21907
rect 52052 21904 52058 21956
rect 53668 21876 53696 21984
rect 53926 21972 53932 21984
rect 53984 21972 53990 22024
rect 54202 21972 54208 22024
rect 54260 21972 54266 22024
rect 55766 21972 55772 22024
rect 55824 22012 55830 22024
rect 55861 22015 55919 22021
rect 55861 22012 55873 22015
rect 55824 21984 55873 22012
rect 55824 21972 55830 21984
rect 55861 21981 55873 21984
rect 55907 21981 55919 22015
rect 55861 21975 55919 21981
rect 57146 21972 57152 22024
rect 57204 22012 57210 22024
rect 57992 22021 58020 22052
rect 57701 22015 57759 22021
rect 57701 22012 57713 22015
rect 57204 21984 57713 22012
rect 57204 21972 57210 21984
rect 57701 21981 57713 21984
rect 57747 21981 57759 22015
rect 57701 21975 57759 21981
rect 57977 22015 58035 22021
rect 57977 21981 57989 22015
rect 58023 21981 58035 22015
rect 57977 21975 58035 21981
rect 58069 22015 58127 22021
rect 58069 21981 58081 22015
rect 58115 21981 58127 22015
rect 58069 21975 58127 21981
rect 53742 21904 53748 21956
rect 53800 21904 53806 21956
rect 53837 21947 53895 21953
rect 53837 21913 53849 21947
rect 53883 21944 53895 21947
rect 54018 21944 54024 21956
rect 53883 21916 54024 21944
rect 53883 21913 53895 21916
rect 53837 21907 53895 21913
rect 54018 21904 54024 21916
rect 54076 21904 54082 21956
rect 55674 21904 55680 21956
rect 55732 21944 55738 21956
rect 56106 21947 56164 21953
rect 56106 21944 56118 21947
rect 55732 21916 56118 21944
rect 55732 21904 55738 21916
rect 56106 21913 56118 21916
rect 56152 21913 56164 21947
rect 56106 21907 56164 21913
rect 56318 21904 56324 21956
rect 56376 21944 56382 21956
rect 56376 21916 57376 21944
rect 56376 21904 56382 21916
rect 51644 21848 53696 21876
rect 53760 21876 53788 21904
rect 55858 21876 55864 21888
rect 53760 21848 55864 21876
rect 55858 21836 55864 21848
rect 55916 21836 55922 21888
rect 56778 21836 56784 21888
rect 56836 21876 56842 21888
rect 57241 21879 57299 21885
rect 57241 21876 57253 21879
rect 56836 21848 57253 21876
rect 56836 21836 56842 21848
rect 57241 21845 57253 21848
rect 57287 21845 57299 21879
rect 57348 21876 57376 21916
rect 57422 21904 57428 21956
rect 57480 21944 57486 21956
rect 57885 21947 57943 21953
rect 57885 21944 57897 21947
rect 57480 21916 57897 21944
rect 57480 21904 57486 21916
rect 57885 21913 57897 21916
rect 57931 21913 57943 21947
rect 58084 21944 58112 21975
rect 57885 21907 57943 21913
rect 57992 21916 58112 21944
rect 57992 21876 58020 21916
rect 57348 21848 58020 21876
rect 57241 21839 57299 21845
rect 1104 21786 58880 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 50294 21786
rect 50346 21734 50358 21786
rect 50410 21734 50422 21786
rect 50474 21734 50486 21786
rect 50538 21734 50550 21786
rect 50602 21734 58880 21786
rect 1104 21712 58880 21734
rect 24026 21672 24032 21684
rect 23952 21644 24032 21672
rect 23198 21564 23204 21616
rect 23256 21604 23262 21616
rect 23293 21607 23351 21613
rect 23293 21604 23305 21607
rect 23256 21576 23305 21604
rect 23256 21564 23262 21576
rect 23293 21573 23305 21576
rect 23339 21573 23351 21607
rect 23293 21567 23351 21573
rect 23385 21607 23443 21613
rect 23385 21573 23397 21607
rect 23431 21604 23443 21607
rect 23474 21604 23480 21616
rect 23431 21576 23480 21604
rect 23431 21573 23443 21576
rect 23385 21567 23443 21573
rect 23474 21564 23480 21576
rect 23532 21564 23538 21616
rect 23952 21613 23980 21644
rect 24026 21632 24032 21644
rect 24084 21672 24090 21684
rect 24765 21675 24823 21681
rect 24765 21672 24777 21675
rect 24084 21644 24777 21672
rect 24084 21632 24090 21644
rect 24765 21641 24777 21644
rect 24811 21641 24823 21675
rect 24765 21635 24823 21641
rect 28258 21632 28264 21684
rect 28316 21632 28322 21684
rect 30282 21632 30288 21684
rect 30340 21632 30346 21684
rect 30926 21632 30932 21684
rect 30984 21632 30990 21684
rect 31018 21632 31024 21684
rect 31076 21672 31082 21684
rect 35253 21675 35311 21681
rect 35253 21672 35265 21675
rect 31076 21644 35265 21672
rect 31076 21632 31082 21644
rect 23937 21607 23995 21613
rect 23937 21573 23949 21607
rect 23983 21573 23995 21607
rect 24854 21604 24860 21616
rect 23937 21567 23995 21573
rect 24228 21576 24860 21604
rect 1581 21539 1639 21545
rect 1581 21505 1593 21539
rect 1627 21536 1639 21539
rect 11698 21536 11704 21548
rect 1627 21508 11704 21536
rect 1627 21505 1639 21508
rect 1581 21499 1639 21505
rect 11698 21496 11704 21508
rect 11756 21496 11762 21548
rect 22094 21496 22100 21548
rect 22152 21536 22158 21548
rect 22278 21536 22284 21548
rect 22152 21508 22284 21536
rect 22152 21496 22158 21508
rect 22278 21496 22284 21508
rect 22336 21496 22342 21548
rect 23753 21539 23811 21545
rect 23753 21505 23765 21539
rect 23799 21505 23811 21539
rect 23753 21499 23811 21505
rect 23845 21539 23903 21545
rect 23845 21505 23857 21539
rect 23891 21536 23903 21539
rect 24228 21536 24256 21576
rect 24854 21564 24860 21576
rect 24912 21564 24918 21616
rect 27706 21564 27712 21616
rect 27764 21604 27770 21616
rect 28074 21604 28080 21616
rect 27764 21576 28080 21604
rect 27764 21564 27770 21576
rect 28074 21564 28080 21576
rect 28132 21564 28138 21616
rect 30834 21604 30840 21616
rect 29932 21576 30840 21604
rect 23891 21508 24256 21536
rect 23891 21505 23903 21508
rect 23845 21499 23903 21505
rect 934 21428 940 21480
rect 992 21468 998 21480
rect 1765 21471 1823 21477
rect 1765 21468 1777 21471
rect 992 21440 1777 21468
rect 992 21428 998 21440
rect 1765 21437 1777 21440
rect 1811 21437 1823 21471
rect 1765 21431 1823 21437
rect 22649 21471 22707 21477
rect 22649 21437 22661 21471
rect 22695 21437 22707 21471
rect 23768 21468 23796 21499
rect 24578 21496 24584 21548
rect 24636 21536 24642 21548
rect 24673 21539 24731 21545
rect 24673 21536 24685 21539
rect 24636 21508 24685 21536
rect 24636 21496 24642 21508
rect 24673 21505 24685 21508
rect 24719 21505 24731 21539
rect 24673 21499 24731 21505
rect 25406 21496 25412 21548
rect 25464 21536 25470 21548
rect 26329 21539 26387 21545
rect 26329 21536 26341 21539
rect 25464 21508 26341 21536
rect 25464 21496 25470 21508
rect 26329 21505 26341 21508
rect 26375 21505 26387 21539
rect 26329 21499 26387 21505
rect 27801 21539 27859 21545
rect 27801 21505 27813 21539
rect 27847 21536 27859 21539
rect 28905 21539 28963 21545
rect 27847 21508 28856 21536
rect 27847 21505 27859 21508
rect 27801 21499 27859 21505
rect 24486 21468 24492 21480
rect 23768 21440 24492 21468
rect 22649 21431 22707 21437
rect 22462 21360 22468 21412
rect 22520 21400 22526 21412
rect 22664 21400 22692 21431
rect 24486 21428 24492 21440
rect 24544 21428 24550 21480
rect 28442 21468 28448 21480
rect 27908 21440 28448 21468
rect 27908 21400 27936 21440
rect 28442 21428 28448 21440
rect 28500 21428 28506 21480
rect 28828 21468 28856 21508
rect 28905 21505 28917 21539
rect 28951 21536 28963 21539
rect 29730 21536 29736 21548
rect 28951 21508 29736 21536
rect 28951 21505 28963 21508
rect 28905 21499 28963 21505
rect 29730 21496 29736 21508
rect 29788 21496 29794 21548
rect 29932 21545 29960 21576
rect 30834 21564 30840 21576
rect 30892 21604 30898 21616
rect 30892 21576 31340 21604
rect 30892 21564 30898 21576
rect 29917 21539 29975 21545
rect 29917 21505 29929 21539
rect 29963 21505 29975 21539
rect 31110 21536 31116 21548
rect 29917 21499 29975 21505
rect 30015 21508 31116 21536
rect 28997 21471 29055 21477
rect 28997 21468 29009 21471
rect 28828 21440 29009 21468
rect 28997 21437 29009 21440
rect 29043 21437 29055 21471
rect 28997 21431 29055 21437
rect 22520 21372 27936 21400
rect 28169 21403 28227 21409
rect 22520 21360 22526 21372
rect 28169 21369 28181 21403
rect 28215 21400 28227 21403
rect 28350 21400 28356 21412
rect 28215 21372 28356 21400
rect 28215 21369 28227 21372
rect 28169 21363 28227 21369
rect 28350 21360 28356 21372
rect 28408 21360 28414 21412
rect 29012 21400 29040 21431
rect 29270 21428 29276 21480
rect 29328 21428 29334 21480
rect 29822 21428 29828 21480
rect 29880 21428 29886 21480
rect 29086 21400 29092 21412
rect 29012 21372 29092 21400
rect 29086 21360 29092 21372
rect 29144 21400 29150 21412
rect 30015 21400 30043 21508
rect 31110 21496 31116 21508
rect 31168 21496 31174 21548
rect 31312 21545 31340 21576
rect 31297 21539 31355 21545
rect 31297 21505 31309 21539
rect 31343 21505 31355 21539
rect 31297 21499 31355 21505
rect 30650 21428 30656 21480
rect 30708 21468 30714 21480
rect 31205 21471 31263 21477
rect 31205 21468 31217 21471
rect 30708 21440 31217 21468
rect 30708 21428 30714 21440
rect 31205 21437 31217 21440
rect 31251 21437 31263 21471
rect 31205 21431 31263 21437
rect 31389 21471 31447 21477
rect 31389 21437 31401 21471
rect 31435 21468 31447 21471
rect 31496 21468 31524 21644
rect 35253 21641 35265 21644
rect 35299 21641 35311 21675
rect 35253 21635 35311 21641
rect 36722 21632 36728 21684
rect 36780 21632 36786 21684
rect 36998 21632 37004 21684
rect 37056 21672 37062 21684
rect 41598 21672 41604 21684
rect 37056 21644 41604 21672
rect 37056 21632 37062 21644
rect 41598 21632 41604 21644
rect 41656 21632 41662 21684
rect 41693 21675 41751 21681
rect 41693 21641 41705 21675
rect 41739 21672 41751 21675
rect 42058 21672 42064 21684
rect 41739 21644 42064 21672
rect 41739 21641 41751 21644
rect 41693 21635 41751 21641
rect 42058 21632 42064 21644
rect 42116 21632 42122 21684
rect 42610 21672 42616 21684
rect 42536 21644 42616 21672
rect 31570 21564 31576 21616
rect 31628 21604 31634 21616
rect 33042 21604 33048 21616
rect 31628 21576 33048 21604
rect 31628 21564 31634 21576
rect 33042 21564 33048 21576
rect 33100 21564 33106 21616
rect 36354 21604 36360 21616
rect 35084 21576 36360 21604
rect 32306 21496 32312 21548
rect 32364 21496 32370 21548
rect 33312 21539 33370 21545
rect 33312 21505 33324 21539
rect 33358 21536 33370 21539
rect 33686 21536 33692 21548
rect 33358 21508 33692 21536
rect 33358 21505 33370 21508
rect 33312 21499 33370 21505
rect 33686 21496 33692 21508
rect 33744 21496 33750 21548
rect 35084 21545 35112 21576
rect 36354 21564 36360 21576
rect 36412 21564 36418 21616
rect 38838 21604 38844 21616
rect 37292 21576 38844 21604
rect 35069 21539 35127 21545
rect 35069 21505 35081 21539
rect 35115 21505 35127 21539
rect 35069 21499 35127 21505
rect 35805 21539 35863 21545
rect 35805 21505 35817 21539
rect 35851 21505 35863 21539
rect 35805 21499 35863 21505
rect 36541 21539 36599 21545
rect 36541 21505 36553 21539
rect 36587 21536 36599 21539
rect 37182 21536 37188 21548
rect 36587 21508 37188 21536
rect 36587 21505 36599 21508
rect 36541 21499 36599 21505
rect 31435 21440 31524 21468
rect 31435 21437 31447 21440
rect 31389 21431 31447 21437
rect 29144 21372 30043 21400
rect 31220 21400 31248 21431
rect 33042 21428 33048 21480
rect 33100 21428 33106 21480
rect 34146 21428 34152 21480
rect 34204 21468 34210 21480
rect 35820 21468 35848 21499
rect 37182 21496 37188 21508
rect 37240 21496 37246 21548
rect 34204 21440 35848 21468
rect 34204 21428 34210 21440
rect 31570 21400 31576 21412
rect 31220 21372 31576 21400
rect 29144 21360 29150 21372
rect 31570 21360 31576 21372
rect 31628 21360 31634 21412
rect 37292 21400 37320 21576
rect 38838 21564 38844 21576
rect 38896 21564 38902 21616
rect 39666 21604 39672 21616
rect 39132 21576 39672 21604
rect 37366 21496 37372 21548
rect 37424 21536 37430 21548
rect 39132 21545 39160 21576
rect 39666 21564 39672 21576
rect 39724 21564 39730 21616
rect 40862 21564 40868 21616
rect 40920 21604 40926 21616
rect 41230 21604 41236 21616
rect 40920 21576 41236 21604
rect 40920 21564 40926 21576
rect 41230 21564 41236 21576
rect 41288 21604 41294 21616
rect 41509 21607 41567 21613
rect 41509 21604 41521 21607
rect 41288 21576 41521 21604
rect 41288 21564 41294 21576
rect 41509 21573 41521 21576
rect 41555 21604 41567 21607
rect 42536 21604 42564 21644
rect 42610 21632 42616 21644
rect 42668 21632 42674 21684
rect 42794 21632 42800 21684
rect 42852 21632 42858 21684
rect 43346 21632 43352 21684
rect 43404 21672 43410 21684
rect 45557 21675 45615 21681
rect 43404 21644 44772 21672
rect 43404 21632 43410 21644
rect 42812 21604 42840 21632
rect 44082 21604 44088 21616
rect 41555 21576 42564 21604
rect 42628 21576 44088 21604
rect 41555 21573 41567 21576
rect 41509 21567 41567 21573
rect 39390 21545 39396 21548
rect 37461 21539 37519 21545
rect 37461 21536 37473 21539
rect 37424 21508 37473 21536
rect 37424 21496 37430 21508
rect 37461 21505 37473 21508
rect 37507 21505 37519 21539
rect 38197 21539 38255 21545
rect 38197 21536 38209 21539
rect 37461 21499 37519 21505
rect 37660 21508 38209 21536
rect 37660 21409 37688 21508
rect 38197 21505 38209 21508
rect 38243 21505 38255 21539
rect 38197 21499 38255 21505
rect 39117 21539 39175 21545
rect 39117 21505 39129 21539
rect 39163 21505 39175 21539
rect 39117 21499 39175 21505
rect 39373 21539 39396 21545
rect 39373 21505 39385 21539
rect 39373 21499 39396 21505
rect 39390 21496 39396 21499
rect 39448 21496 39454 21548
rect 40402 21496 40408 21548
rect 40460 21536 40466 21548
rect 41325 21539 41383 21545
rect 41325 21536 41337 21539
rect 40460 21508 41337 21536
rect 40460 21496 40466 21508
rect 41325 21505 41337 21508
rect 41371 21536 41383 21539
rect 42518 21536 42524 21548
rect 41371 21508 42524 21536
rect 41371 21505 41383 21508
rect 41325 21499 41383 21505
rect 42518 21496 42524 21508
rect 42576 21496 42582 21548
rect 42628 21545 42656 21576
rect 44082 21564 44088 21576
rect 44140 21564 44146 21616
rect 44744 21613 44772 21644
rect 45557 21641 45569 21675
rect 45603 21672 45615 21675
rect 53558 21672 53564 21684
rect 45603 21644 53564 21672
rect 45603 21641 45615 21644
rect 45557 21635 45615 21641
rect 53558 21632 53564 21644
rect 53616 21632 53622 21684
rect 54018 21632 54024 21684
rect 54076 21672 54082 21684
rect 54297 21675 54355 21681
rect 54297 21672 54309 21675
rect 54076 21644 54309 21672
rect 54076 21632 54082 21644
rect 54297 21641 54309 21644
rect 54343 21641 54355 21675
rect 54297 21635 54355 21641
rect 44729 21607 44787 21613
rect 44729 21573 44741 21607
rect 44775 21604 44787 21607
rect 46566 21604 46572 21616
rect 44775 21576 46572 21604
rect 44775 21573 44787 21576
rect 44729 21567 44787 21573
rect 46566 21564 46572 21576
rect 46624 21564 46630 21616
rect 53184 21607 53242 21613
rect 53184 21573 53196 21607
rect 53230 21604 53242 21607
rect 53282 21604 53288 21616
rect 53230 21576 53288 21604
rect 53230 21573 53242 21576
rect 53184 21567 53242 21573
rect 53282 21564 53288 21576
rect 53340 21564 53346 21616
rect 54312 21604 54340 21635
rect 55674 21632 55680 21684
rect 55732 21632 55738 21684
rect 55858 21632 55864 21684
rect 55916 21672 55922 21684
rect 57422 21672 57428 21684
rect 55916 21644 57428 21672
rect 55916 21632 55922 21644
rect 57422 21632 57428 21644
rect 57480 21632 57486 21684
rect 56594 21604 56600 21616
rect 54312 21576 56600 21604
rect 56594 21564 56600 21576
rect 56652 21564 56658 21616
rect 42613 21539 42671 21545
rect 42613 21505 42625 21539
rect 42659 21505 42671 21539
rect 42613 21499 42671 21505
rect 42702 21496 42708 21548
rect 42760 21536 42766 21548
rect 42869 21539 42927 21545
rect 42869 21536 42881 21539
rect 42760 21508 42881 21536
rect 42760 21496 42766 21508
rect 42869 21505 42881 21508
rect 42915 21505 42927 21539
rect 42869 21499 42927 21505
rect 43438 21496 43444 21548
rect 43496 21536 43502 21548
rect 44545 21539 44603 21545
rect 44545 21536 44557 21539
rect 43496 21508 44557 21536
rect 43496 21496 43502 21508
rect 44545 21505 44557 21508
rect 44591 21505 44603 21539
rect 45925 21539 45983 21545
rect 45925 21536 45937 21539
rect 44545 21499 44603 21505
rect 45526 21508 45937 21536
rect 45526 21468 45554 21508
rect 45925 21505 45937 21508
rect 45971 21505 45983 21539
rect 45925 21499 45983 21505
rect 48774 21496 48780 21548
rect 48832 21496 48838 21548
rect 48961 21539 49019 21545
rect 48961 21505 48973 21539
rect 49007 21536 49019 21539
rect 49786 21536 49792 21548
rect 49007 21508 49792 21536
rect 49007 21505 49019 21508
rect 48961 21499 49019 21505
rect 49786 21496 49792 21508
rect 49844 21496 49850 21548
rect 55398 21496 55404 21548
rect 55456 21496 55462 21548
rect 55490 21496 55496 21548
rect 55548 21496 55554 21548
rect 56226 21496 56232 21548
rect 56284 21536 56290 21548
rect 56393 21539 56451 21545
rect 56393 21536 56405 21539
rect 56284 21508 56405 21536
rect 56284 21496 56290 21508
rect 56393 21505 56405 21508
rect 56439 21505 56451 21539
rect 56393 21499 56451 21505
rect 57422 21496 57428 21548
rect 57480 21536 57486 21548
rect 57698 21536 57704 21548
rect 57480 21508 57704 21536
rect 57480 21496 57486 21508
rect 57698 21496 57704 21508
rect 57756 21496 57762 21548
rect 58066 21496 58072 21548
rect 58124 21496 58130 21548
rect 44008 21440 45554 21468
rect 35912 21372 37320 21400
rect 37645 21403 37703 21409
rect 26234 21292 26240 21344
rect 26292 21332 26298 21344
rect 26513 21335 26571 21341
rect 26513 21332 26525 21335
rect 26292 21304 26525 21332
rect 26292 21292 26298 21304
rect 26513 21301 26525 21304
rect 26559 21301 26571 21335
rect 26513 21295 26571 21301
rect 27338 21292 27344 21344
rect 27396 21332 27402 21344
rect 30282 21332 30288 21344
rect 27396 21304 30288 21332
rect 27396 21292 27402 21304
rect 30282 21292 30288 21304
rect 30340 21292 30346 21344
rect 30834 21292 30840 21344
rect 30892 21332 30898 21344
rect 32493 21335 32551 21341
rect 32493 21332 32505 21335
rect 30892 21304 32505 21332
rect 30892 21292 30898 21304
rect 32493 21301 32505 21304
rect 32539 21301 32551 21335
rect 32493 21295 32551 21301
rect 34425 21335 34483 21341
rect 34425 21301 34437 21335
rect 34471 21332 34483 21335
rect 35912 21332 35940 21372
rect 37645 21369 37657 21403
rect 37691 21369 37703 21403
rect 37645 21363 37703 21369
rect 37734 21360 37740 21412
rect 37792 21400 37798 21412
rect 41414 21400 41420 21412
rect 37792 21372 38516 21400
rect 37792 21360 37798 21372
rect 34471 21304 35940 21332
rect 35989 21335 36047 21341
rect 34471 21301 34483 21304
rect 34425 21295 34483 21301
rect 35989 21301 36001 21335
rect 36035 21332 36047 21335
rect 36722 21332 36728 21344
rect 36035 21304 36728 21332
rect 36035 21301 36047 21304
rect 35989 21295 36047 21301
rect 36722 21292 36728 21304
rect 36780 21292 36786 21344
rect 37550 21292 37556 21344
rect 37608 21332 37614 21344
rect 38381 21335 38439 21341
rect 38381 21332 38393 21335
rect 37608 21304 38393 21332
rect 37608 21292 37614 21304
rect 38381 21301 38393 21304
rect 38427 21301 38439 21335
rect 38488 21332 38516 21372
rect 40052 21372 41420 21400
rect 40052 21332 40080 21372
rect 41414 21360 41420 21372
rect 41472 21360 41478 21412
rect 38488 21304 40080 21332
rect 38381 21295 38439 21301
rect 40494 21292 40500 21344
rect 40552 21292 40558 21344
rect 41432 21332 41460 21360
rect 44008 21341 44036 21440
rect 46014 21428 46020 21480
rect 46072 21428 46078 21480
rect 46201 21471 46259 21477
rect 46201 21437 46213 21471
rect 46247 21468 46259 21471
rect 46934 21468 46940 21480
rect 46247 21440 46940 21468
rect 46247 21437 46259 21440
rect 46201 21431 46259 21437
rect 46934 21428 46940 21440
rect 46992 21468 46998 21480
rect 47670 21468 47676 21480
rect 46992 21440 47676 21468
rect 46992 21428 46998 21440
rect 47670 21428 47676 21440
rect 47728 21428 47734 21480
rect 52362 21428 52368 21480
rect 52420 21468 52426 21480
rect 52917 21471 52975 21477
rect 52917 21468 52929 21471
rect 52420 21440 52929 21468
rect 52420 21428 52426 21440
rect 52917 21437 52929 21440
rect 52963 21437 52975 21471
rect 52917 21431 52975 21437
rect 56134 21428 56140 21480
rect 56192 21428 56198 21480
rect 44913 21403 44971 21409
rect 44913 21369 44925 21403
rect 44959 21400 44971 21403
rect 45646 21400 45652 21412
rect 44959 21372 45652 21400
rect 44959 21369 44971 21372
rect 44913 21363 44971 21369
rect 45646 21360 45652 21372
rect 45704 21360 45710 21412
rect 43993 21335 44051 21341
rect 43993 21332 44005 21335
rect 41432 21304 44005 21332
rect 43993 21301 44005 21304
rect 44039 21301 44051 21335
rect 43993 21295 44051 21301
rect 48682 21292 48688 21344
rect 48740 21332 48746 21344
rect 48777 21335 48835 21341
rect 48777 21332 48789 21335
rect 48740 21304 48789 21332
rect 48740 21292 48746 21304
rect 48777 21301 48789 21304
rect 48823 21301 48835 21335
rect 48777 21295 48835 21301
rect 57514 21292 57520 21344
rect 57572 21292 57578 21344
rect 57606 21292 57612 21344
rect 57664 21332 57670 21344
rect 58253 21335 58311 21341
rect 58253 21332 58265 21335
rect 57664 21304 58265 21332
rect 57664 21292 57670 21304
rect 58253 21301 58265 21304
rect 58299 21301 58311 21335
rect 58253 21295 58311 21301
rect 1104 21242 58880 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 58880 21242
rect 1104 21168 58880 21190
rect 23198 21088 23204 21140
rect 23256 21088 23262 21140
rect 23937 21131 23995 21137
rect 23937 21097 23949 21131
rect 23983 21128 23995 21131
rect 24854 21128 24860 21140
rect 23983 21100 24860 21128
rect 23983 21097 23995 21100
rect 23937 21091 23995 21097
rect 24854 21088 24860 21100
rect 24912 21088 24918 21140
rect 25406 21088 25412 21140
rect 25464 21088 25470 21140
rect 27338 21088 27344 21140
rect 27396 21088 27402 21140
rect 30650 21128 30656 21140
rect 28552 21100 30656 21128
rect 28552 21069 28580 21100
rect 30650 21088 30656 21100
rect 30708 21088 30714 21140
rect 31113 21131 31171 21137
rect 31113 21097 31125 21131
rect 31159 21128 31171 21131
rect 31159 21100 32904 21128
rect 31159 21097 31171 21100
rect 31113 21091 31171 21097
rect 28537 21063 28595 21069
rect 28537 21029 28549 21063
rect 28583 21029 28595 21063
rect 28537 21023 28595 21029
rect 29086 21020 29092 21072
rect 29144 21020 29150 21072
rect 31202 21020 31208 21072
rect 31260 21060 31266 21072
rect 31386 21060 31392 21072
rect 31260 21032 31392 21060
rect 31260 21020 31266 21032
rect 31386 21020 31392 21032
rect 31444 21020 31450 21072
rect 32876 21060 32904 21100
rect 32950 21088 32956 21140
rect 33008 21128 33014 21140
rect 33045 21131 33103 21137
rect 33045 21128 33057 21131
rect 33008 21100 33057 21128
rect 33008 21088 33014 21100
rect 33045 21097 33057 21100
rect 33091 21097 33103 21131
rect 33045 21091 33103 21097
rect 33686 21088 33692 21140
rect 33744 21088 33750 21140
rect 33796 21100 36032 21128
rect 33796 21060 33824 21100
rect 32876 21032 33824 21060
rect 36004 21060 36032 21100
rect 36078 21088 36084 21140
rect 36136 21128 36142 21140
rect 36265 21131 36323 21137
rect 36265 21128 36277 21131
rect 36136 21100 36277 21128
rect 36136 21088 36142 21100
rect 36265 21097 36277 21100
rect 36311 21097 36323 21131
rect 36265 21091 36323 21097
rect 36906 21088 36912 21140
rect 36964 21088 36970 21140
rect 37182 21088 37188 21140
rect 37240 21128 37246 21140
rect 37645 21131 37703 21137
rect 37645 21128 37657 21131
rect 37240 21100 37657 21128
rect 37240 21088 37246 21100
rect 37645 21097 37657 21100
rect 37691 21097 37703 21131
rect 37645 21091 37703 21097
rect 38378 21088 38384 21140
rect 38436 21128 38442 21140
rect 43530 21128 43536 21140
rect 38436 21100 43536 21128
rect 38436 21088 38442 21100
rect 43530 21088 43536 21100
rect 43588 21088 43594 21140
rect 43625 21131 43683 21137
rect 43625 21097 43637 21131
rect 43671 21128 43683 21131
rect 44174 21128 44180 21140
rect 43671 21100 44180 21128
rect 43671 21097 43683 21100
rect 43625 21091 43683 21097
rect 44174 21088 44180 21100
rect 44232 21088 44238 21140
rect 45189 21131 45247 21137
rect 45189 21097 45201 21131
rect 45235 21128 45247 21131
rect 45278 21128 45284 21140
rect 45235 21100 45284 21128
rect 45235 21097 45247 21100
rect 45189 21091 45247 21097
rect 45278 21088 45284 21100
rect 45336 21088 45342 21140
rect 49789 21131 49847 21137
rect 49789 21097 49801 21131
rect 49835 21128 49847 21131
rect 49878 21128 49884 21140
rect 49835 21100 49884 21128
rect 49835 21097 49847 21100
rect 49789 21091 49847 21097
rect 49878 21088 49884 21100
rect 49936 21088 49942 21140
rect 55490 21088 55496 21140
rect 55548 21128 55554 21140
rect 55769 21131 55827 21137
rect 55769 21128 55781 21131
rect 55548 21100 55781 21128
rect 55548 21088 55554 21100
rect 55769 21097 55781 21100
rect 55815 21097 55827 21131
rect 55769 21091 55827 21097
rect 57790 21088 57796 21140
rect 57848 21128 57854 21140
rect 58253 21131 58311 21137
rect 58253 21128 58265 21131
rect 57848 21100 58265 21128
rect 57848 21088 57854 21100
rect 58253 21097 58265 21100
rect 58299 21097 58311 21131
rect 58253 21091 58311 21097
rect 37734 21060 37740 21072
rect 36004 21032 37740 21060
rect 37734 21020 37740 21032
rect 37792 21020 37798 21072
rect 40310 21060 40316 21072
rect 38626 21032 40316 21060
rect 934 20952 940 21004
rect 992 20992 998 21004
rect 1765 20995 1823 21001
rect 1765 20992 1777 20995
rect 992 20964 1777 20992
rect 992 20952 998 20964
rect 1765 20961 1777 20964
rect 1811 20961 1823 20995
rect 28626 20992 28632 21004
rect 1765 20955 1823 20961
rect 27908 20964 28632 20992
rect 1581 20927 1639 20933
rect 1581 20893 1593 20927
rect 1627 20924 1639 20927
rect 1627 20896 6914 20924
rect 1627 20893 1639 20896
rect 1581 20887 1639 20893
rect 6886 20856 6914 20896
rect 22002 20884 22008 20936
rect 22060 20884 22066 20936
rect 22462 20884 22468 20936
rect 22520 20884 22526 20936
rect 23017 20927 23075 20933
rect 23017 20893 23029 20927
rect 23063 20893 23075 20927
rect 23017 20887 23075 20893
rect 22189 20859 22247 20865
rect 22189 20856 22201 20859
rect 6886 20828 22201 20856
rect 22189 20825 22201 20828
rect 22235 20825 22247 20859
rect 23032 20856 23060 20887
rect 23750 20884 23756 20936
rect 23808 20884 23814 20936
rect 25222 20884 25228 20936
rect 25280 20884 25286 20936
rect 27908 20933 27936 20964
rect 28626 20952 28632 20964
rect 28684 20992 28690 21004
rect 28684 20964 28948 20992
rect 28684 20952 28690 20964
rect 25961 20927 26019 20933
rect 25961 20893 25973 20927
rect 26007 20924 26019 20927
rect 27893 20927 27951 20933
rect 26007 20896 26372 20924
rect 26007 20893 26019 20896
rect 25961 20887 26019 20893
rect 26344 20868 26372 20896
rect 27893 20893 27905 20927
rect 27939 20893 27951 20927
rect 27893 20887 27951 20893
rect 28077 20927 28135 20933
rect 28077 20893 28089 20927
rect 28123 20924 28135 20927
rect 28534 20924 28540 20936
rect 28123 20896 28540 20924
rect 28123 20893 28135 20896
rect 28077 20887 28135 20893
rect 28534 20884 28540 20896
rect 28592 20924 28598 20936
rect 28920 20933 28948 20964
rect 33042 20952 33048 21004
rect 33100 20992 33106 21004
rect 34885 20995 34943 21001
rect 34885 20992 34897 20995
rect 33100 20964 34897 20992
rect 33100 20952 33106 20964
rect 34885 20961 34897 20964
rect 34931 20961 34943 20995
rect 38626 20992 38654 21032
rect 40310 21020 40316 21032
rect 40368 21020 40374 21072
rect 40494 21020 40500 21072
rect 40552 21060 40558 21072
rect 43254 21060 43260 21072
rect 40552 21032 43260 21060
rect 40552 21020 40558 21032
rect 43254 21020 43260 21032
rect 43312 21020 43318 21072
rect 45830 21060 45836 21072
rect 45480 21032 45836 21060
rect 34885 20955 34943 20961
rect 36832 20964 38654 20992
rect 39005 20995 39063 21001
rect 28813 20927 28871 20933
rect 28813 20924 28825 20927
rect 28592 20896 28825 20924
rect 28592 20884 28598 20896
rect 28813 20893 28825 20896
rect 28859 20893 28871 20927
rect 28813 20887 28871 20893
rect 28905 20927 28963 20933
rect 28905 20893 28917 20927
rect 28951 20893 28963 20927
rect 28905 20887 28963 20893
rect 29730 20884 29736 20936
rect 29788 20924 29794 20936
rect 31665 20927 31723 20933
rect 30668 20924 30880 20926
rect 31665 20924 31677 20927
rect 29788 20898 31677 20924
rect 29788 20896 30696 20898
rect 30852 20896 31677 20898
rect 29788 20884 29794 20896
rect 31665 20893 31677 20896
rect 31711 20924 31723 20927
rect 33060 20924 33088 20952
rect 31711 20896 33088 20924
rect 31711 20893 31723 20896
rect 31665 20887 31723 20893
rect 33502 20884 33508 20936
rect 33560 20884 33566 20936
rect 35152 20927 35210 20933
rect 35152 20893 35164 20927
rect 35198 20924 35210 20927
rect 36630 20924 36636 20936
rect 35198 20896 36636 20924
rect 35198 20893 35210 20896
rect 35152 20887 35210 20893
rect 36630 20884 36636 20896
rect 36688 20884 36694 20936
rect 36722 20884 36728 20936
rect 36780 20884 36786 20936
rect 24118 20856 24124 20868
rect 23032 20828 24124 20856
rect 22189 20819 22247 20825
rect 24118 20816 24124 20828
rect 24176 20816 24182 20868
rect 26234 20865 26240 20868
rect 26228 20856 26240 20865
rect 26195 20828 26240 20856
rect 26228 20819 26240 20828
rect 26234 20816 26240 20819
rect 26292 20816 26298 20868
rect 26326 20816 26332 20868
rect 26384 20816 26390 20868
rect 30006 20865 30012 20868
rect 28721 20859 28779 20865
rect 28721 20825 28733 20859
rect 28767 20856 28779 20859
rect 28767 20828 29960 20856
rect 28767 20825 28779 20828
rect 28721 20819 28779 20825
rect 27614 20748 27620 20800
rect 27672 20788 27678 20800
rect 27985 20791 28043 20797
rect 27985 20788 27997 20791
rect 27672 20760 27997 20788
rect 27672 20748 27678 20760
rect 27985 20757 27997 20760
rect 28031 20757 28043 20791
rect 29932 20788 29960 20828
rect 30000 20819 30012 20865
rect 30006 20816 30012 20819
rect 30064 20816 30070 20868
rect 31932 20859 31990 20865
rect 31036 20828 31754 20856
rect 31036 20788 31064 20828
rect 29932 20760 31064 20788
rect 31726 20788 31754 20828
rect 31932 20825 31944 20859
rect 31978 20856 31990 20859
rect 32858 20856 32864 20868
rect 31978 20828 32864 20856
rect 31978 20825 31990 20828
rect 31932 20819 31990 20825
rect 32858 20816 32864 20828
rect 32916 20816 32922 20868
rect 32950 20816 32956 20868
rect 33008 20856 33014 20868
rect 36832 20856 36860 20964
rect 39005 20961 39017 20995
rect 39051 20992 39063 20995
rect 44542 20992 44548 21004
rect 39051 20964 40816 20992
rect 39051 20961 39063 20964
rect 39005 20955 39063 20961
rect 37458 20884 37464 20936
rect 37516 20884 37522 20936
rect 38197 20927 38255 20933
rect 38197 20893 38209 20927
rect 38243 20924 38255 20927
rect 38378 20924 38384 20936
rect 38243 20896 38384 20924
rect 38243 20893 38255 20896
rect 38197 20887 38255 20893
rect 38378 20884 38384 20896
rect 38436 20884 38442 20936
rect 38562 20884 38568 20936
rect 38620 20924 38626 20936
rect 38838 20924 38844 20936
rect 38620 20896 38844 20924
rect 38620 20884 38626 20896
rect 38838 20884 38844 20896
rect 38896 20884 38902 20936
rect 39209 20927 39267 20933
rect 39209 20893 39221 20927
rect 39255 20893 39267 20927
rect 39209 20887 39267 20893
rect 40037 20927 40095 20933
rect 40037 20893 40049 20927
rect 40083 20924 40095 20927
rect 40218 20924 40224 20936
rect 40083 20896 40224 20924
rect 40083 20893 40095 20896
rect 40037 20887 40095 20893
rect 33008 20828 36860 20856
rect 33008 20816 33014 20828
rect 37826 20816 37832 20868
rect 37884 20856 37890 20868
rect 37884 20828 38516 20856
rect 37884 20816 37890 20828
rect 32306 20788 32312 20800
rect 31726 20760 32312 20788
rect 27985 20751 28043 20757
rect 32306 20748 32312 20760
rect 32364 20788 32370 20800
rect 38381 20791 38439 20797
rect 38381 20788 38393 20791
rect 32364 20760 38393 20788
rect 32364 20748 32370 20760
rect 38381 20757 38393 20760
rect 38427 20757 38439 20791
rect 38488 20788 38516 20828
rect 38654 20816 38660 20868
rect 38712 20856 38718 20868
rect 38933 20859 38991 20865
rect 38933 20856 38945 20859
rect 38712 20828 38945 20856
rect 38712 20816 38718 20828
rect 38933 20825 38945 20828
rect 38979 20825 38991 20859
rect 38933 20819 38991 20825
rect 39022 20816 39028 20868
rect 39080 20856 39086 20868
rect 39117 20859 39175 20865
rect 39117 20856 39129 20859
rect 39080 20828 39129 20856
rect 39080 20816 39086 20828
rect 39117 20825 39129 20828
rect 39163 20825 39175 20859
rect 39117 20819 39175 20825
rect 39224 20788 39252 20887
rect 40218 20884 40224 20896
rect 40276 20884 40282 20936
rect 40310 20884 40316 20936
rect 40368 20924 40374 20936
rect 40788 20933 40816 20964
rect 41386 20964 43484 20992
rect 40773 20927 40831 20933
rect 40368 20896 40724 20924
rect 40368 20884 40374 20896
rect 40696 20856 40724 20896
rect 40773 20893 40785 20927
rect 40819 20893 40831 20927
rect 40773 20887 40831 20893
rect 41230 20856 41236 20868
rect 40696 20828 41236 20856
rect 41230 20816 41236 20828
rect 41288 20856 41294 20868
rect 41386 20856 41414 20964
rect 41506 20884 41512 20936
rect 41564 20884 41570 20936
rect 42518 20884 42524 20936
rect 42576 20924 42582 20936
rect 42613 20927 42671 20933
rect 42613 20924 42625 20927
rect 42576 20896 42625 20924
rect 42576 20884 42582 20896
rect 42613 20893 42625 20896
rect 42659 20924 42671 20927
rect 43346 20924 43352 20936
rect 42659 20896 43352 20924
rect 42659 20893 42671 20896
rect 42613 20887 42671 20893
rect 43346 20884 43352 20896
rect 43404 20884 43410 20936
rect 41288 20828 41414 20856
rect 41785 20859 41843 20865
rect 41288 20816 41294 20828
rect 41785 20825 41797 20859
rect 41831 20856 41843 20859
rect 42150 20856 42156 20868
rect 41831 20828 42156 20856
rect 41831 20825 41843 20828
rect 41785 20819 41843 20825
rect 42150 20816 42156 20828
rect 42208 20816 42214 20868
rect 42794 20816 42800 20868
rect 42852 20816 42858 20868
rect 38488 20760 39252 20788
rect 38381 20751 38439 20757
rect 40218 20748 40224 20800
rect 40276 20748 40282 20800
rect 40310 20748 40316 20800
rect 40368 20788 40374 20800
rect 40957 20791 41015 20797
rect 40957 20788 40969 20791
rect 40368 20760 40969 20788
rect 40368 20748 40374 20760
rect 40957 20757 40969 20760
rect 41003 20757 41015 20791
rect 40957 20751 41015 20757
rect 42981 20791 43039 20797
rect 42981 20757 42993 20791
rect 43027 20788 43039 20791
rect 43346 20788 43352 20800
rect 43027 20760 43352 20788
rect 43027 20757 43039 20760
rect 42981 20751 43039 20757
rect 43346 20748 43352 20760
rect 43404 20748 43410 20800
rect 43456 20788 43484 20964
rect 44100 20964 44548 20992
rect 43622 20884 43628 20936
rect 43680 20924 43686 20936
rect 43898 20924 43904 20936
rect 43680 20896 43904 20924
rect 43680 20884 43686 20896
rect 43898 20884 43904 20896
rect 43956 20884 43962 20936
rect 43990 20884 43996 20936
rect 44048 20884 44054 20936
rect 44100 20933 44128 20964
rect 44542 20952 44548 20964
rect 44600 20952 44606 21004
rect 44085 20927 44143 20933
rect 44085 20893 44097 20927
rect 44131 20893 44143 20927
rect 44085 20887 44143 20893
rect 44266 20884 44272 20936
rect 44324 20884 44330 20936
rect 45480 20933 45508 21032
rect 45830 21020 45836 21032
rect 45888 21060 45894 21072
rect 46750 21060 46756 21072
rect 45888 21032 46756 21060
rect 45888 21020 45894 21032
rect 46750 21020 46756 21032
rect 46808 21020 46814 21072
rect 55766 20952 55772 21004
rect 55824 20992 55830 21004
rect 56134 20992 56140 21004
rect 55824 20964 56140 20992
rect 55824 20952 55830 20964
rect 56134 20952 56140 20964
rect 56192 20992 56198 21004
rect 56873 20995 56931 21001
rect 56873 20992 56885 20995
rect 56192 20964 56885 20992
rect 56192 20952 56198 20964
rect 56873 20961 56885 20964
rect 56919 20961 56931 20995
rect 56873 20955 56931 20961
rect 45465 20927 45523 20933
rect 45465 20893 45477 20927
rect 45511 20893 45523 20927
rect 45465 20887 45523 20893
rect 45554 20884 45560 20936
rect 45612 20884 45618 20936
rect 45646 20884 45652 20936
rect 45704 20884 45710 20936
rect 45833 20927 45891 20933
rect 45833 20893 45845 20927
rect 45879 20893 45891 20927
rect 45833 20887 45891 20893
rect 44284 20856 44312 20884
rect 45848 20856 45876 20887
rect 48406 20884 48412 20936
rect 48464 20884 48470 20936
rect 48682 20933 48688 20936
rect 48676 20924 48688 20933
rect 48643 20896 48688 20924
rect 48676 20887 48688 20896
rect 48682 20884 48688 20887
rect 48740 20884 48746 20936
rect 55858 20884 55864 20936
rect 55916 20924 55922 20936
rect 55953 20927 56011 20933
rect 55953 20924 55965 20927
rect 55916 20896 55965 20924
rect 55916 20884 55922 20896
rect 55953 20893 55965 20896
rect 55999 20893 56011 20927
rect 55953 20887 56011 20893
rect 56413 20927 56471 20933
rect 56413 20893 56425 20927
rect 56459 20924 56471 20927
rect 56778 20924 56784 20936
rect 56459 20896 56784 20924
rect 56459 20893 56471 20896
rect 56413 20887 56471 20893
rect 56778 20884 56784 20896
rect 56836 20884 56842 20936
rect 56962 20884 56968 20936
rect 57020 20924 57026 20936
rect 57129 20927 57187 20933
rect 57129 20924 57141 20927
rect 57020 20896 57141 20924
rect 57020 20884 57026 20896
rect 57129 20893 57141 20896
rect 57175 20893 57187 20927
rect 57129 20887 57187 20893
rect 44284 20828 45876 20856
rect 56042 20816 56048 20868
rect 56100 20816 56106 20868
rect 56318 20865 56324 20868
rect 56137 20859 56195 20865
rect 56137 20825 56149 20859
rect 56183 20825 56195 20859
rect 56137 20819 56195 20825
rect 56275 20859 56324 20865
rect 56275 20825 56287 20859
rect 56321 20825 56324 20859
rect 56275 20819 56324 20825
rect 48130 20788 48136 20800
rect 43456 20760 48136 20788
rect 48130 20748 48136 20760
rect 48188 20748 48194 20800
rect 56152 20788 56180 20819
rect 56318 20816 56324 20819
rect 56376 20816 56382 20868
rect 56410 20788 56416 20800
rect 56152 20760 56416 20788
rect 56410 20748 56416 20760
rect 56468 20748 56474 20800
rect 1104 20698 58880 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 50294 20698
rect 50346 20646 50358 20698
rect 50410 20646 50422 20698
rect 50474 20646 50486 20698
rect 50538 20646 50550 20698
rect 50602 20646 58880 20698
rect 1104 20624 58880 20646
rect 24302 20544 24308 20596
rect 24360 20544 24366 20596
rect 26602 20544 26608 20596
rect 26660 20544 26666 20596
rect 28810 20584 28816 20596
rect 28000 20556 28816 20584
rect 23658 20476 23664 20528
rect 23716 20476 23722 20528
rect 23934 20476 23940 20528
rect 23992 20516 23998 20528
rect 24320 20516 24348 20544
rect 28000 20516 28028 20556
rect 28810 20544 28816 20556
rect 28868 20544 28874 20596
rect 29273 20587 29331 20593
rect 29273 20553 29285 20587
rect 29319 20584 29331 20587
rect 34422 20584 34428 20596
rect 29319 20556 34428 20584
rect 29319 20553 29331 20556
rect 29273 20547 29331 20553
rect 34422 20544 34428 20556
rect 34480 20544 34486 20596
rect 37458 20544 37464 20596
rect 37516 20584 37522 20596
rect 37645 20587 37703 20593
rect 37645 20584 37657 20587
rect 37516 20556 37657 20584
rect 37516 20544 37522 20556
rect 37645 20553 37657 20556
rect 37691 20553 37703 20587
rect 37645 20547 37703 20553
rect 38838 20544 38844 20596
rect 38896 20584 38902 20596
rect 40402 20584 40408 20596
rect 38896 20556 40408 20584
rect 38896 20544 38902 20556
rect 40402 20544 40408 20556
rect 40460 20544 40466 20596
rect 40862 20544 40868 20596
rect 40920 20584 40926 20596
rect 46109 20587 46167 20593
rect 46109 20584 46121 20587
rect 40920 20556 46121 20584
rect 40920 20544 40926 20556
rect 46109 20553 46121 20556
rect 46155 20553 46167 20587
rect 46109 20547 46167 20553
rect 47762 20544 47768 20596
rect 47820 20584 47826 20596
rect 47949 20587 48007 20593
rect 47949 20584 47961 20587
rect 47820 20556 47961 20584
rect 47820 20544 47826 20556
rect 47949 20553 47961 20556
rect 47995 20553 48007 20587
rect 47949 20547 48007 20553
rect 48774 20544 48780 20596
rect 48832 20584 48838 20596
rect 48961 20587 49019 20593
rect 48961 20584 48973 20587
rect 48832 20556 48973 20584
rect 48832 20544 48838 20556
rect 48961 20553 48973 20556
rect 49007 20553 49019 20587
rect 48961 20547 49019 20553
rect 49142 20544 49148 20596
rect 49200 20544 49206 20596
rect 50522 20544 50528 20596
rect 50580 20584 50586 20596
rect 51445 20587 51503 20593
rect 51445 20584 51457 20587
rect 50580 20556 51457 20584
rect 50580 20544 50586 20556
rect 51445 20553 51457 20556
rect 51491 20553 51503 20587
rect 51445 20547 51503 20553
rect 28166 20525 28172 20528
rect 28160 20516 28172 20525
rect 23992 20488 24808 20516
rect 23992 20476 23998 20488
rect 1581 20451 1639 20457
rect 1581 20417 1593 20451
rect 1627 20448 1639 20451
rect 2958 20448 2964 20460
rect 1627 20420 2964 20448
rect 1627 20417 1639 20420
rect 1581 20411 1639 20417
rect 2958 20408 2964 20420
rect 3016 20408 3022 20460
rect 24305 20451 24363 20457
rect 24305 20417 24317 20451
rect 24351 20417 24363 20451
rect 24305 20411 24363 20417
rect 934 20340 940 20392
rect 992 20380 998 20392
rect 1765 20383 1823 20389
rect 1765 20380 1777 20383
rect 992 20352 1777 20380
rect 992 20340 998 20352
rect 1765 20349 1777 20352
rect 1811 20349 1823 20383
rect 24320 20380 24348 20411
rect 24394 20408 24400 20460
rect 24452 20408 24458 20460
rect 24670 20408 24676 20460
rect 24728 20408 24734 20460
rect 24780 20457 24808 20488
rect 26252 20488 28028 20516
rect 28127 20488 28172 20516
rect 26252 20457 26280 20488
rect 28160 20479 28172 20488
rect 28166 20476 28172 20479
rect 28224 20476 28230 20528
rect 38657 20519 38715 20525
rect 32600 20488 37596 20516
rect 24765 20451 24823 20457
rect 24765 20417 24777 20451
rect 24811 20417 24823 20451
rect 24765 20411 24823 20417
rect 26237 20451 26295 20457
rect 26237 20417 26249 20451
rect 26283 20417 26295 20451
rect 26237 20411 26295 20417
rect 27157 20451 27215 20457
rect 27157 20417 27169 20451
rect 27203 20448 27215 20451
rect 28442 20448 28448 20460
rect 27203 20420 28448 20448
rect 27203 20417 27215 20420
rect 27157 20411 27215 20417
rect 28442 20408 28448 20420
rect 28500 20408 28506 20460
rect 28718 20408 28724 20460
rect 28776 20448 28782 20460
rect 29730 20448 29736 20460
rect 28776 20420 29736 20448
rect 28776 20408 28782 20420
rect 29730 20408 29736 20420
rect 29788 20448 29794 20460
rect 30009 20451 30067 20457
rect 30009 20448 30021 20451
rect 29788 20420 30021 20448
rect 29788 20408 29794 20420
rect 30009 20417 30021 20420
rect 30055 20417 30067 20451
rect 30009 20411 30067 20417
rect 30650 20408 30656 20460
rect 30708 20448 30714 20460
rect 32600 20457 32628 20488
rect 32585 20451 32643 20457
rect 32585 20448 32597 20451
rect 30708 20420 32597 20448
rect 30708 20408 30714 20420
rect 32585 20417 32597 20420
rect 32631 20417 32643 20451
rect 32585 20411 32643 20417
rect 33042 20408 33048 20460
rect 33100 20448 33106 20460
rect 33321 20451 33379 20457
rect 33321 20448 33333 20451
rect 33100 20420 33333 20448
rect 33100 20408 33106 20420
rect 33321 20417 33333 20420
rect 33367 20417 33379 20451
rect 33321 20411 33379 20417
rect 33588 20451 33646 20457
rect 33588 20417 33600 20451
rect 33634 20448 33646 20451
rect 34790 20448 34796 20460
rect 33634 20420 34796 20448
rect 33634 20417 33646 20420
rect 33588 20411 33646 20417
rect 34790 20408 34796 20420
rect 34848 20408 34854 20460
rect 35250 20408 35256 20460
rect 35308 20408 35314 20460
rect 35526 20408 35532 20460
rect 35584 20448 35590 20460
rect 35584 20420 36676 20448
rect 35584 20408 35590 20420
rect 26329 20383 26387 20389
rect 24320 20352 24716 20380
rect 1765 20343 1823 20349
rect 24688 20324 24716 20352
rect 26329 20349 26341 20383
rect 26375 20380 26387 20383
rect 27614 20380 27620 20392
rect 26375 20352 27620 20380
rect 26375 20349 26387 20352
rect 26329 20343 26387 20349
rect 27614 20340 27620 20352
rect 27672 20340 27678 20392
rect 27890 20340 27896 20392
rect 27948 20340 27954 20392
rect 30285 20383 30343 20389
rect 30285 20349 30297 20383
rect 30331 20380 30343 20383
rect 31202 20380 31208 20392
rect 30331 20352 31208 20380
rect 30331 20349 30343 20352
rect 30285 20343 30343 20349
rect 31202 20340 31208 20352
rect 31260 20340 31266 20392
rect 31665 20383 31723 20389
rect 31665 20349 31677 20383
rect 31711 20380 31723 20383
rect 32950 20380 32956 20392
rect 31711 20352 32956 20380
rect 31711 20349 31723 20352
rect 31665 20343 31723 20349
rect 32950 20340 32956 20352
rect 33008 20340 33014 20392
rect 35986 20340 35992 20392
rect 36044 20380 36050 20392
rect 36541 20383 36599 20389
rect 36541 20380 36553 20383
rect 36044 20352 36553 20380
rect 36044 20340 36050 20352
rect 36541 20349 36553 20352
rect 36587 20349 36599 20383
rect 36648 20380 36676 20420
rect 36722 20408 36728 20460
rect 36780 20448 36786 20460
rect 37182 20448 37188 20460
rect 36780 20420 37188 20448
rect 36780 20408 36786 20420
rect 37182 20408 37188 20420
rect 37240 20408 37246 20460
rect 37458 20408 37464 20460
rect 37516 20408 37522 20460
rect 37568 20448 37596 20488
rect 38657 20485 38669 20519
rect 38703 20516 38715 20519
rect 40006 20519 40064 20525
rect 40006 20516 40018 20519
rect 38703 20488 40018 20516
rect 38703 20485 38715 20488
rect 38657 20479 38715 20485
rect 40006 20485 40018 20488
rect 40052 20485 40064 20519
rect 40006 20479 40064 20485
rect 41966 20476 41972 20528
rect 42024 20476 42030 20528
rect 44634 20516 44640 20528
rect 43272 20488 44640 20516
rect 38838 20448 38844 20460
rect 37568 20420 38844 20448
rect 38838 20408 38844 20420
rect 38896 20408 38902 20460
rect 38930 20408 38936 20460
rect 38988 20408 38994 20460
rect 39025 20451 39083 20457
rect 39025 20417 39037 20451
rect 39071 20417 39083 20451
rect 39025 20411 39083 20417
rect 38562 20380 38568 20392
rect 36648 20352 38568 20380
rect 36541 20343 36599 20349
rect 38562 20340 38568 20352
rect 38620 20340 38626 20392
rect 38746 20340 38752 20392
rect 38804 20380 38810 20392
rect 39040 20380 39068 20411
rect 39114 20408 39120 20460
rect 39172 20408 39178 20460
rect 39301 20451 39359 20457
rect 39301 20417 39313 20451
rect 39347 20448 39359 20451
rect 39574 20448 39580 20460
rect 39347 20420 39580 20448
rect 39347 20417 39359 20420
rect 39301 20411 39359 20417
rect 39574 20408 39580 20420
rect 39632 20408 39638 20460
rect 39666 20408 39672 20460
rect 39724 20448 39730 20460
rect 39761 20451 39819 20457
rect 39761 20448 39773 20451
rect 39724 20420 39773 20448
rect 39724 20408 39730 20420
rect 39761 20417 39773 20420
rect 39807 20417 39819 20451
rect 39761 20411 39819 20417
rect 40494 20408 40500 20460
rect 40552 20448 40558 20460
rect 41046 20448 41052 20460
rect 40552 20420 41052 20448
rect 40552 20408 40558 20420
rect 41046 20408 41052 20420
rect 41104 20408 41110 20460
rect 41690 20408 41696 20460
rect 41748 20408 41754 20460
rect 41984 20448 42012 20476
rect 42610 20448 42616 20460
rect 41984 20420 42616 20448
rect 42610 20408 42616 20420
rect 42668 20408 42674 20460
rect 43272 20457 43300 20488
rect 44634 20476 44640 20488
rect 44692 20476 44698 20528
rect 48406 20476 48412 20528
rect 48464 20516 48470 20528
rect 51074 20516 51080 20528
rect 48464 20488 51080 20516
rect 48464 20476 48470 20488
rect 43530 20457 43536 20460
rect 42797 20451 42855 20457
rect 42797 20417 42809 20451
rect 42843 20417 42855 20451
rect 42797 20411 42855 20417
rect 43257 20451 43315 20457
rect 43257 20417 43269 20451
rect 43303 20417 43315 20451
rect 43257 20411 43315 20417
rect 43524 20411 43536 20457
rect 38804 20352 39068 20380
rect 38804 20340 38810 20352
rect 41966 20340 41972 20392
rect 42024 20380 42030 20392
rect 42812 20380 42840 20411
rect 43530 20408 43536 20411
rect 43588 20408 43594 20460
rect 45189 20451 45247 20457
rect 45189 20448 45201 20451
rect 44284 20420 45201 20448
rect 42024 20352 42840 20380
rect 42024 20340 42030 20352
rect 24670 20272 24676 20324
rect 24728 20272 24734 20324
rect 32769 20315 32827 20321
rect 32769 20312 32781 20315
rect 30944 20284 32781 20312
rect 17402 20204 17408 20256
rect 17460 20244 17466 20256
rect 23658 20244 23664 20256
rect 17460 20216 23664 20244
rect 17460 20204 17466 20216
rect 23658 20204 23664 20216
rect 23716 20204 23722 20256
rect 27341 20247 27399 20253
rect 27341 20213 27353 20247
rect 27387 20244 27399 20247
rect 28258 20244 28264 20256
rect 27387 20216 28264 20244
rect 27387 20213 27399 20216
rect 27341 20207 27399 20213
rect 28258 20204 28264 20216
rect 28316 20204 28322 20256
rect 28902 20204 28908 20256
rect 28960 20244 28966 20256
rect 30944 20244 30972 20284
rect 32769 20281 32781 20284
rect 32815 20281 32827 20315
rect 36262 20312 36268 20324
rect 32769 20275 32827 20281
rect 34256 20284 36268 20312
rect 28960 20216 30972 20244
rect 28960 20204 28966 20216
rect 34054 20204 34060 20256
rect 34112 20244 34118 20256
rect 34256 20244 34284 20284
rect 36262 20272 36268 20284
rect 36320 20272 36326 20324
rect 36630 20272 36636 20324
rect 36688 20312 36694 20324
rect 37826 20312 37832 20324
rect 36688 20284 37832 20312
rect 36688 20272 36694 20284
rect 37826 20272 37832 20284
rect 37884 20272 37890 20324
rect 41506 20272 41512 20324
rect 41564 20312 41570 20324
rect 42705 20315 42763 20321
rect 42705 20312 42717 20315
rect 41564 20284 42717 20312
rect 41564 20272 41570 20284
rect 42705 20281 42717 20284
rect 42751 20281 42763 20315
rect 42705 20275 42763 20281
rect 34112 20216 34284 20244
rect 34112 20204 34118 20216
rect 34698 20204 34704 20256
rect 34756 20204 34762 20256
rect 35434 20204 35440 20256
rect 35492 20204 35498 20256
rect 36909 20247 36967 20253
rect 36909 20213 36921 20247
rect 36955 20244 36967 20247
rect 36998 20244 37004 20256
rect 36955 20216 37004 20244
rect 36955 20213 36967 20216
rect 36909 20207 36967 20213
rect 36998 20204 37004 20216
rect 37056 20204 37062 20256
rect 41138 20204 41144 20256
rect 41196 20204 41202 20256
rect 41874 20204 41880 20256
rect 41932 20204 41938 20256
rect 42058 20204 42064 20256
rect 42116 20244 42122 20256
rect 44284 20244 44312 20420
rect 45189 20417 45201 20420
rect 45235 20417 45247 20451
rect 45189 20411 45247 20417
rect 45922 20408 45928 20460
rect 45980 20408 45986 20460
rect 47946 20448 47952 20460
rect 47907 20420 47952 20448
rect 47946 20408 47952 20420
rect 48004 20408 48010 20460
rect 48317 20451 48375 20457
rect 48317 20417 48329 20451
rect 48363 20448 48375 20451
rect 48682 20448 48688 20460
rect 48363 20420 48688 20448
rect 48363 20417 48375 20420
rect 48317 20411 48375 20417
rect 48682 20408 48688 20420
rect 48740 20408 48746 20460
rect 49142 20451 49200 20457
rect 49142 20417 49154 20451
rect 49188 20448 49200 20451
rect 49878 20448 49884 20460
rect 49188 20420 49884 20448
rect 49188 20417 49200 20420
rect 49142 20411 49200 20417
rect 49878 20408 49884 20420
rect 49936 20408 49942 20460
rect 50080 20457 50108 20488
rect 51074 20476 51080 20488
rect 51132 20476 51138 20528
rect 51460 20516 51488 20547
rect 53098 20544 53104 20596
rect 53156 20544 53162 20596
rect 57422 20584 57428 20596
rect 53484 20556 57428 20584
rect 53484 20550 53512 20556
rect 53208 20522 53512 20550
rect 57422 20544 57428 20556
rect 57480 20544 57486 20596
rect 53208 20516 53236 20522
rect 51460 20488 53236 20516
rect 55214 20476 55220 20528
rect 55272 20516 55278 20528
rect 56137 20519 56195 20525
rect 56137 20516 56149 20519
rect 55272 20488 56149 20516
rect 55272 20476 55278 20488
rect 56137 20485 56149 20488
rect 56183 20485 56195 20519
rect 56137 20479 56195 20485
rect 50065 20451 50123 20457
rect 50065 20417 50077 20451
rect 50111 20417 50123 20451
rect 50065 20411 50123 20417
rect 50154 20408 50160 20460
rect 50212 20448 50218 20460
rect 50321 20451 50379 20457
rect 50321 20448 50333 20451
rect 50212 20420 50333 20448
rect 50212 20408 50218 20420
rect 50321 20417 50333 20420
rect 50367 20417 50379 20451
rect 50321 20411 50379 20417
rect 52181 20451 52239 20457
rect 52181 20417 52193 20451
rect 52227 20417 52239 20451
rect 52181 20411 52239 20417
rect 44542 20340 44548 20392
rect 44600 20380 44606 20392
rect 45370 20380 45376 20392
rect 44600 20352 45376 20380
rect 44600 20340 44606 20352
rect 45370 20340 45376 20352
rect 45428 20340 45434 20392
rect 48409 20383 48467 20389
rect 48409 20380 48421 20383
rect 45526 20352 48421 20380
rect 44358 20272 44364 20324
rect 44416 20312 44422 20324
rect 45526 20312 45554 20352
rect 48409 20349 48421 20352
rect 48455 20349 48467 20383
rect 48409 20343 48467 20349
rect 49605 20383 49663 20389
rect 49605 20349 49617 20383
rect 49651 20349 49663 20383
rect 52196 20380 52224 20411
rect 52270 20408 52276 20460
rect 52328 20448 52334 20460
rect 52365 20451 52423 20457
rect 52365 20448 52377 20451
rect 52328 20420 52377 20448
rect 52328 20408 52334 20420
rect 52365 20417 52377 20420
rect 52411 20417 52423 20451
rect 52365 20411 52423 20417
rect 53098 20451 53156 20457
rect 53098 20417 53110 20451
rect 53144 20448 53156 20451
rect 53834 20448 53840 20460
rect 53144 20420 53840 20448
rect 53144 20417 53156 20420
rect 53098 20411 53156 20417
rect 53834 20408 53840 20420
rect 53892 20408 53898 20460
rect 55674 20408 55680 20460
rect 55732 20448 55738 20460
rect 55858 20448 55864 20460
rect 55732 20420 55864 20448
rect 55732 20408 55738 20420
rect 55858 20408 55864 20420
rect 55916 20448 55922 20460
rect 56045 20451 56103 20457
rect 56045 20448 56057 20451
rect 55916 20420 56057 20448
rect 55916 20408 55922 20420
rect 56045 20417 56057 20420
rect 56091 20417 56103 20451
rect 56045 20411 56103 20417
rect 56229 20451 56287 20457
rect 56229 20417 56241 20451
rect 56275 20417 56287 20451
rect 56229 20411 56287 20417
rect 53466 20380 53472 20392
rect 52196 20352 53472 20380
rect 49605 20343 49663 20349
rect 44416 20284 45554 20312
rect 47765 20315 47823 20321
rect 44416 20272 44422 20284
rect 47765 20281 47777 20315
rect 47811 20312 47823 20315
rect 49513 20315 49571 20321
rect 49513 20312 49525 20315
rect 47811 20284 49525 20312
rect 47811 20281 47823 20284
rect 47765 20275 47823 20281
rect 49513 20281 49525 20284
rect 49559 20281 49571 20315
rect 49513 20275 49571 20281
rect 42116 20216 44312 20244
rect 42116 20204 42122 20216
rect 44542 20204 44548 20256
rect 44600 20244 44606 20256
rect 44637 20247 44695 20253
rect 44637 20244 44649 20247
rect 44600 20216 44649 20244
rect 44600 20204 44606 20216
rect 44637 20213 44649 20216
rect 44683 20213 44695 20247
rect 44637 20207 44695 20213
rect 44726 20204 44732 20256
rect 44784 20244 44790 20256
rect 45373 20247 45431 20253
rect 45373 20244 45385 20247
rect 44784 20216 45385 20244
rect 44784 20204 44790 20216
rect 45373 20213 45385 20216
rect 45419 20213 45431 20247
rect 49620 20244 49648 20343
rect 53466 20340 53472 20352
rect 53524 20340 53530 20392
rect 53558 20340 53564 20392
rect 53616 20340 53622 20392
rect 52181 20315 52239 20321
rect 52181 20281 52193 20315
rect 52227 20312 52239 20315
rect 53006 20312 53012 20324
rect 52227 20284 53012 20312
rect 52227 20281 52239 20284
rect 52181 20275 52239 20281
rect 53006 20272 53012 20284
rect 53064 20272 53070 20324
rect 53098 20272 53104 20324
rect 53156 20312 53162 20324
rect 56244 20312 56272 20411
rect 56318 20408 56324 20460
rect 56376 20457 56382 20460
rect 56376 20451 56405 20457
rect 56393 20417 56405 20451
rect 56376 20411 56405 20417
rect 56505 20451 56563 20457
rect 56505 20417 56517 20451
rect 56551 20448 56563 20451
rect 57514 20448 57520 20460
rect 56551 20420 57520 20448
rect 56551 20417 56563 20420
rect 56505 20411 56563 20417
rect 56376 20408 56382 20411
rect 57514 20408 57520 20420
rect 57572 20408 57578 20460
rect 58158 20408 58164 20460
rect 58216 20408 58222 20460
rect 56410 20312 56416 20324
rect 53156 20284 53604 20312
rect 53156 20272 53162 20284
rect 51258 20244 51264 20256
rect 49620 20216 51264 20244
rect 45373 20207 45431 20213
rect 51258 20204 51264 20216
rect 51316 20204 51322 20256
rect 51994 20204 52000 20256
rect 52052 20244 52058 20256
rect 52917 20247 52975 20253
rect 52917 20244 52929 20247
rect 52052 20216 52929 20244
rect 52052 20204 52058 20216
rect 52917 20213 52929 20216
rect 52963 20213 52975 20247
rect 52917 20207 52975 20213
rect 53466 20204 53472 20256
rect 53524 20204 53530 20256
rect 53576 20244 53604 20284
rect 53944 20284 56180 20312
rect 56244 20284 56416 20312
rect 53944 20244 53972 20284
rect 53576 20216 53972 20244
rect 55861 20247 55919 20253
rect 55861 20213 55873 20247
rect 55907 20244 55919 20247
rect 56042 20244 56048 20256
rect 55907 20216 56048 20244
rect 55907 20213 55919 20216
rect 55861 20207 55919 20213
rect 56042 20204 56048 20216
rect 56100 20204 56106 20256
rect 56152 20244 56180 20284
rect 56410 20272 56416 20284
rect 56468 20272 56474 20324
rect 56318 20244 56324 20256
rect 56152 20216 56324 20244
rect 56318 20204 56324 20216
rect 56376 20204 56382 20256
rect 57974 20204 57980 20256
rect 58032 20244 58038 20256
rect 58253 20247 58311 20253
rect 58253 20244 58265 20247
rect 58032 20216 58265 20244
rect 58032 20204 58038 20216
rect 58253 20213 58265 20216
rect 58299 20213 58311 20247
rect 58253 20207 58311 20213
rect 1104 20154 58880 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 58880 20154
rect 1104 20080 58880 20102
rect 28442 20000 28448 20052
rect 28500 20000 28506 20052
rect 28626 20040 28632 20052
rect 28552 20012 28632 20040
rect 22005 19975 22063 19981
rect 22005 19972 22017 19975
rect 6886 19944 22017 19972
rect 934 19864 940 19916
rect 992 19904 998 19916
rect 1765 19907 1823 19913
rect 1765 19904 1777 19907
rect 992 19876 1777 19904
rect 992 19864 998 19876
rect 1765 19873 1777 19876
rect 1811 19873 1823 19907
rect 1765 19867 1823 19873
rect 1581 19839 1639 19845
rect 1581 19805 1593 19839
rect 1627 19836 1639 19839
rect 6886 19836 6914 19944
rect 22005 19941 22017 19944
rect 22051 19941 22063 19975
rect 22005 19935 22063 19941
rect 22186 19904 22192 19916
rect 22066 19876 22192 19904
rect 1627 19808 6914 19836
rect 21821 19839 21879 19845
rect 1627 19805 1639 19808
rect 1581 19799 1639 19805
rect 21821 19805 21833 19839
rect 21867 19836 21879 19839
rect 22066 19836 22094 19876
rect 22186 19864 22192 19876
rect 22244 19904 22250 19916
rect 23106 19904 23112 19916
rect 22244 19876 23112 19904
rect 22244 19864 22250 19876
rect 23106 19864 23112 19876
rect 23164 19864 23170 19916
rect 28552 19904 28580 20012
rect 28626 20000 28632 20012
rect 28684 20000 28690 20052
rect 28810 20000 28816 20052
rect 28868 20040 28874 20052
rect 30834 20040 30840 20052
rect 28868 20012 30840 20040
rect 28868 20000 28874 20012
rect 30834 20000 30840 20012
rect 30892 20000 30898 20052
rect 31202 20000 31208 20052
rect 31260 20000 31266 20052
rect 35434 20040 35440 20052
rect 32048 20012 35440 20040
rect 30469 19975 30527 19981
rect 30469 19941 30481 19975
rect 30515 19941 30527 19975
rect 30469 19935 30527 19941
rect 28621 19907 28679 19913
rect 28621 19904 28633 19907
rect 28552 19876 28633 19904
rect 28621 19873 28633 19876
rect 28667 19873 28679 19907
rect 28621 19867 28679 19873
rect 28810 19864 28816 19916
rect 28868 19864 28874 19916
rect 28902 19864 28908 19916
rect 28960 19864 28966 19916
rect 21867 19808 22094 19836
rect 22281 19839 22339 19845
rect 21867 19805 21879 19808
rect 21821 19799 21879 19805
rect 22281 19805 22293 19839
rect 22327 19836 22339 19839
rect 22370 19836 22376 19848
rect 22327 19808 22376 19836
rect 22327 19805 22339 19808
rect 22281 19799 22339 19805
rect 22370 19796 22376 19808
rect 22428 19796 22434 19848
rect 24486 19796 24492 19848
rect 24544 19836 24550 19848
rect 24673 19839 24731 19845
rect 24673 19836 24685 19839
rect 24544 19808 24685 19836
rect 24544 19796 24550 19808
rect 24673 19805 24685 19808
rect 24719 19836 24731 19839
rect 24762 19836 24768 19848
rect 24719 19808 24768 19836
rect 24719 19805 24731 19808
rect 24673 19799 24731 19805
rect 24762 19796 24768 19808
rect 24820 19796 24826 19848
rect 24857 19839 24915 19845
rect 24857 19805 24869 19839
rect 24903 19805 24915 19839
rect 24857 19799 24915 19805
rect 2593 19771 2651 19777
rect 2593 19737 2605 19771
rect 2639 19768 2651 19771
rect 17218 19768 17224 19780
rect 2639 19740 17224 19768
rect 2639 19737 2651 19740
rect 2593 19731 2651 19737
rect 17218 19728 17224 19740
rect 17276 19728 17282 19780
rect 24118 19728 24124 19780
rect 24176 19768 24182 19780
rect 24872 19768 24900 19799
rect 25314 19796 25320 19848
rect 25372 19836 25378 19848
rect 25409 19839 25467 19845
rect 25409 19836 25421 19839
rect 25372 19808 25421 19836
rect 25372 19796 25378 19808
rect 25409 19805 25421 19808
rect 25455 19805 25467 19839
rect 25409 19799 25467 19805
rect 26326 19796 26332 19848
rect 26384 19836 26390 19848
rect 27890 19836 27896 19848
rect 26384 19808 27896 19836
rect 26384 19796 26390 19808
rect 27890 19796 27896 19808
rect 27948 19796 27954 19848
rect 28710 19839 28768 19845
rect 28710 19814 28722 19839
rect 28644 19805 28722 19814
rect 28756 19805 28768 19839
rect 28644 19799 28768 19805
rect 25498 19768 25504 19780
rect 24176 19740 25504 19768
rect 24176 19728 24182 19740
rect 25498 19728 25504 19740
rect 25556 19728 25562 19780
rect 26596 19771 26654 19777
rect 26596 19737 26608 19771
rect 26642 19768 26654 19771
rect 27062 19768 27068 19780
rect 26642 19740 27068 19768
rect 26642 19737 26654 19740
rect 26596 19731 26654 19737
rect 27062 19728 27068 19740
rect 27120 19728 27126 19780
rect 934 19660 940 19712
rect 992 19700 998 19712
rect 2685 19703 2743 19709
rect 2685 19700 2697 19703
rect 992 19672 2697 19700
rect 992 19660 998 19672
rect 2685 19669 2697 19672
rect 2731 19669 2743 19703
rect 2685 19663 2743 19669
rect 24670 19660 24676 19712
rect 24728 19660 24734 19712
rect 27709 19703 27767 19709
rect 27709 19669 27721 19703
rect 27755 19700 27767 19703
rect 27798 19700 27804 19712
rect 27755 19672 27804 19700
rect 27755 19669 27767 19672
rect 27709 19663 27767 19669
rect 27798 19660 27804 19672
rect 27856 19660 27862 19712
rect 27908 19700 27936 19796
rect 28644 19786 28764 19799
rect 30282 19796 30288 19848
rect 30340 19796 30346 19848
rect 30484 19836 30512 19935
rect 30650 19932 30656 19984
rect 30708 19972 30714 19984
rect 31941 19975 31999 19981
rect 31941 19972 31953 19975
rect 30708 19944 31953 19972
rect 30708 19932 30714 19944
rect 31941 19941 31953 19944
rect 31987 19941 31999 19975
rect 31941 19935 31999 19941
rect 31021 19839 31079 19845
rect 31021 19836 31033 19839
rect 30484 19808 31033 19836
rect 31021 19805 31033 19808
rect 31067 19805 31079 19839
rect 31021 19799 31079 19805
rect 31757 19839 31815 19845
rect 31757 19805 31769 19839
rect 31803 19836 31815 19839
rect 32048 19836 32076 20012
rect 35434 20000 35440 20012
rect 35492 20000 35498 20052
rect 36909 20043 36967 20049
rect 36909 20009 36921 20043
rect 36955 20040 36967 20043
rect 36955 20012 37044 20040
rect 36955 20009 36967 20012
rect 36909 20003 36967 20009
rect 34333 19975 34391 19981
rect 34333 19941 34345 19975
rect 34379 19972 34391 19975
rect 36814 19972 36820 19984
rect 34379 19944 36820 19972
rect 34379 19941 34391 19944
rect 34333 19935 34391 19941
rect 36814 19932 36820 19944
rect 36872 19932 36878 19984
rect 37016 19972 37044 20012
rect 37366 20000 37372 20052
rect 37424 20040 37430 20052
rect 37550 20040 37556 20052
rect 37424 20012 37556 20040
rect 37424 20000 37430 20012
rect 37550 20000 37556 20012
rect 37608 20000 37614 20052
rect 37734 20000 37740 20052
rect 37792 20040 37798 20052
rect 38470 20040 38476 20052
rect 37792 20012 38476 20040
rect 37792 20000 37798 20012
rect 38470 20000 38476 20012
rect 38528 20000 38534 20052
rect 39114 20000 39120 20052
rect 39172 20040 39178 20052
rect 40405 20043 40463 20049
rect 40405 20040 40417 20043
rect 39172 20012 40417 20040
rect 39172 20000 39178 20012
rect 40405 20009 40417 20012
rect 40451 20009 40463 20043
rect 40405 20003 40463 20009
rect 42889 20043 42947 20049
rect 42889 20009 42901 20043
rect 42935 20040 42947 20043
rect 43530 20040 43536 20052
rect 42935 20012 43536 20040
rect 42935 20009 42947 20012
rect 42889 20003 42947 20009
rect 43530 20000 43536 20012
rect 43588 20000 43594 20052
rect 44174 20000 44180 20052
rect 44232 20040 44238 20052
rect 44542 20040 44548 20052
rect 44232 20012 44548 20040
rect 44232 20000 44238 20012
rect 44542 20000 44548 20012
rect 44600 20000 44606 20052
rect 48314 20000 48320 20052
rect 48372 20040 48378 20052
rect 49142 20040 49148 20052
rect 48372 20012 49148 20040
rect 48372 20000 48378 20012
rect 49142 20000 49148 20012
rect 49200 20040 49206 20052
rect 50430 20040 50436 20052
rect 49200 20012 50436 20040
rect 49200 20000 49206 20012
rect 50430 20000 50436 20012
rect 50488 20040 50494 20052
rect 51166 20040 51172 20052
rect 50488 20012 51172 20040
rect 50488 20000 50494 20012
rect 51166 20000 51172 20012
rect 51224 20000 51230 20052
rect 53466 20040 53472 20052
rect 52012 20012 53472 20040
rect 41874 19972 41880 19984
rect 37016 19944 41880 19972
rect 41874 19932 41880 19944
rect 41932 19932 41938 19984
rect 42150 19932 42156 19984
rect 42208 19972 42214 19984
rect 44358 19972 44364 19984
rect 42208 19944 44364 19972
rect 42208 19932 42214 19944
rect 44358 19932 44364 19944
rect 44416 19932 44422 19984
rect 52012 19972 52040 20012
rect 53466 20000 53472 20012
rect 53524 20000 53530 20052
rect 53650 20000 53656 20052
rect 53708 20040 53714 20052
rect 53837 20043 53895 20049
rect 53837 20040 53849 20043
rect 53708 20012 53849 20040
rect 53708 20000 53714 20012
rect 53837 20009 53849 20012
rect 53883 20009 53895 20043
rect 53837 20003 53895 20009
rect 56226 20000 56232 20052
rect 56284 20000 56290 20052
rect 47965 19944 52040 19972
rect 53377 19975 53435 19981
rect 35253 19907 35311 19913
rect 35253 19873 35265 19907
rect 35299 19904 35311 19907
rect 37366 19904 37372 19916
rect 35299 19876 37372 19904
rect 35299 19873 35311 19876
rect 35253 19867 35311 19873
rect 37366 19864 37372 19876
rect 37424 19864 37430 19916
rect 37553 19907 37611 19913
rect 37553 19873 37565 19907
rect 37599 19873 37611 19907
rect 40034 19904 40040 19916
rect 37553 19867 37611 19873
rect 38396 19876 40040 19904
rect 31803 19808 32076 19836
rect 32953 19839 33011 19845
rect 31803 19805 31815 19808
rect 31757 19799 31815 19805
rect 32953 19805 32965 19839
rect 32999 19836 33011 19839
rect 33042 19836 33048 19848
rect 32999 19808 33048 19836
rect 32999 19805 33011 19808
rect 32953 19799 33011 19805
rect 28534 19728 28540 19780
rect 28592 19768 28598 19780
rect 28644 19768 28672 19786
rect 28592 19740 28672 19768
rect 28592 19728 28598 19740
rect 28810 19728 28816 19780
rect 28868 19768 28874 19780
rect 30466 19768 30472 19780
rect 28868 19740 30472 19768
rect 28868 19728 28874 19740
rect 30466 19728 30472 19740
rect 30524 19728 30530 19780
rect 28718 19700 28724 19712
rect 27908 19672 28724 19700
rect 28718 19660 28724 19672
rect 28776 19660 28782 19712
rect 28994 19660 29000 19712
rect 29052 19700 29058 19712
rect 31772 19700 31800 19799
rect 33042 19796 33048 19808
rect 33100 19796 33106 19848
rect 33220 19839 33278 19845
rect 33220 19805 33232 19839
rect 33266 19836 33278 19839
rect 33266 19808 35940 19836
rect 33266 19805 33278 19808
rect 33220 19799 33278 19805
rect 34330 19728 34336 19780
rect 34388 19768 34394 19780
rect 35805 19771 35863 19777
rect 35805 19768 35817 19771
rect 34388 19740 35817 19768
rect 34388 19728 34394 19740
rect 35805 19737 35817 19740
rect 35851 19737 35863 19771
rect 35912 19768 35940 19808
rect 36170 19796 36176 19848
rect 36228 19836 36234 19848
rect 36538 19839 36596 19845
rect 36538 19836 36550 19839
rect 36228 19808 36550 19836
rect 36228 19796 36234 19808
rect 36538 19805 36550 19808
rect 36584 19836 36596 19839
rect 36630 19836 36636 19848
rect 36584 19808 36636 19836
rect 36584 19805 36596 19808
rect 36538 19799 36596 19805
rect 36630 19796 36636 19808
rect 36688 19796 36694 19848
rect 36998 19845 37004 19848
rect 36995 19799 37004 19845
rect 37056 19836 37062 19848
rect 37056 19808 37095 19836
rect 36998 19796 37004 19799
rect 37056 19796 37062 19808
rect 37182 19796 37188 19848
rect 37240 19836 37246 19848
rect 37568 19836 37596 19867
rect 37240 19808 37596 19836
rect 37645 19839 37703 19845
rect 37240 19796 37246 19808
rect 37645 19805 37657 19839
rect 37691 19836 37703 19839
rect 38396 19836 38424 19876
rect 40034 19864 40040 19876
rect 40092 19864 40098 19916
rect 41138 19904 41144 19916
rect 40236 19876 41144 19904
rect 40236 19848 40264 19876
rect 41138 19864 41144 19876
rect 41196 19904 41202 19916
rect 42058 19904 42064 19916
rect 41196 19876 42064 19904
rect 41196 19864 41202 19876
rect 42058 19864 42064 19876
rect 42116 19864 42122 19916
rect 42610 19864 42616 19916
rect 42668 19904 42674 19916
rect 43990 19904 43996 19916
rect 42668 19876 43996 19904
rect 42668 19864 42674 19876
rect 37691 19808 38424 19836
rect 37691 19805 37703 19808
rect 37645 19799 37703 19805
rect 38470 19796 38476 19848
rect 38528 19796 38534 19848
rect 38654 19796 38660 19848
rect 38712 19836 38718 19848
rect 39209 19839 39267 19845
rect 38712 19808 38792 19836
rect 38712 19796 38718 19808
rect 38764 19768 38792 19808
rect 39209 19805 39221 19839
rect 39255 19836 39267 19839
rect 40126 19836 40132 19848
rect 39255 19808 40132 19836
rect 39255 19805 39267 19808
rect 39209 19799 39267 19805
rect 40126 19796 40132 19808
rect 40184 19796 40190 19848
rect 40218 19796 40224 19848
rect 40276 19796 40282 19848
rect 40862 19796 40868 19848
rect 40920 19796 40926 19848
rect 41414 19796 41420 19848
rect 41472 19836 41478 19848
rect 41601 19839 41659 19845
rect 41601 19836 41613 19839
rect 41472 19808 41613 19836
rect 41472 19796 41478 19808
rect 41601 19805 41613 19808
rect 41647 19805 41659 19839
rect 41601 19799 41659 19805
rect 42978 19796 42984 19848
rect 43036 19836 43042 19848
rect 43162 19836 43168 19848
rect 43036 19808 43168 19836
rect 43036 19796 43042 19808
rect 43162 19796 43168 19808
rect 43220 19796 43226 19848
rect 43272 19845 43300 19876
rect 43990 19864 43996 19876
rect 44048 19904 44054 19916
rect 45373 19907 45431 19913
rect 45373 19904 45385 19907
rect 44048 19876 45385 19904
rect 44048 19864 44054 19876
rect 43257 19839 43315 19845
rect 43257 19805 43269 19839
rect 43303 19805 43315 19839
rect 43257 19799 43315 19805
rect 43346 19796 43352 19848
rect 43404 19796 43410 19848
rect 43533 19839 43591 19845
rect 43533 19805 43545 19839
rect 43579 19836 43591 19839
rect 44174 19836 44180 19848
rect 43579 19808 44180 19836
rect 43579 19805 43591 19808
rect 43533 19799 43591 19805
rect 44174 19796 44180 19808
rect 44232 19796 44238 19848
rect 44266 19796 44272 19848
rect 44324 19796 44330 19848
rect 44376 19845 44404 19876
rect 45373 19873 45385 19876
rect 45419 19873 45431 19907
rect 45373 19867 45431 19873
rect 44361 19839 44419 19845
rect 44361 19805 44373 19839
rect 44407 19805 44419 19839
rect 44361 19799 44419 19805
rect 44450 19796 44456 19848
rect 44508 19796 44514 19848
rect 44542 19796 44548 19848
rect 44600 19836 44606 19848
rect 44637 19839 44695 19845
rect 44637 19836 44649 19839
rect 44600 19808 44649 19836
rect 44600 19796 44606 19808
rect 44637 19805 44649 19808
rect 44683 19805 44695 19839
rect 44637 19799 44695 19805
rect 45189 19839 45247 19845
rect 45189 19805 45201 19839
rect 45235 19836 45247 19839
rect 45554 19836 45560 19848
rect 45235 19808 45560 19836
rect 45235 19805 45247 19808
rect 45189 19799 45247 19805
rect 45554 19796 45560 19808
rect 45612 19796 45618 19848
rect 47762 19796 47768 19848
rect 47820 19796 47826 19848
rect 47854 19796 47860 19848
rect 47912 19796 47918 19848
rect 40037 19771 40095 19777
rect 35912 19740 38700 19768
rect 38764 19740 39528 19768
rect 35805 19731 35863 19737
rect 29052 19672 31800 19700
rect 29052 19660 29058 19672
rect 35434 19660 35440 19712
rect 35492 19660 35498 19712
rect 35526 19660 35532 19712
rect 35584 19660 35590 19712
rect 35621 19703 35679 19709
rect 35621 19669 35633 19703
rect 35667 19700 35679 19703
rect 35894 19700 35900 19712
rect 35667 19672 35900 19700
rect 35667 19669 35679 19672
rect 35621 19663 35679 19669
rect 35894 19660 35900 19672
rect 35952 19660 35958 19712
rect 36357 19703 36415 19709
rect 36357 19669 36369 19703
rect 36403 19700 36415 19703
rect 36446 19700 36452 19712
rect 36403 19672 36452 19700
rect 36403 19669 36415 19672
rect 36357 19663 36415 19669
rect 36446 19660 36452 19672
rect 36504 19660 36510 19712
rect 36538 19660 36544 19712
rect 36596 19660 36602 19712
rect 37366 19660 37372 19712
rect 37424 19700 37430 19712
rect 38672 19709 38700 19740
rect 38013 19703 38071 19709
rect 38013 19700 38025 19703
rect 37424 19672 38025 19700
rect 37424 19660 37430 19672
rect 38013 19669 38025 19672
rect 38059 19669 38071 19703
rect 38013 19663 38071 19669
rect 38657 19703 38715 19709
rect 38657 19669 38669 19703
rect 38703 19669 38715 19703
rect 38657 19663 38715 19669
rect 38838 19660 38844 19712
rect 38896 19700 38902 19712
rect 39393 19703 39451 19709
rect 39393 19700 39405 19703
rect 38896 19672 39405 19700
rect 38896 19660 38902 19672
rect 39393 19669 39405 19672
rect 39439 19669 39451 19703
rect 39500 19700 39528 19740
rect 40037 19737 40049 19771
rect 40083 19768 40095 19771
rect 40494 19768 40500 19780
rect 40083 19740 40500 19768
rect 40083 19737 40095 19740
rect 40037 19731 40095 19737
rect 40494 19728 40500 19740
rect 40552 19728 40558 19780
rect 40954 19728 40960 19780
rect 41012 19768 41018 19780
rect 41012 19740 45048 19768
rect 41012 19728 41018 19740
rect 41049 19703 41107 19709
rect 41049 19700 41061 19703
rect 39500 19672 41061 19700
rect 39393 19663 39451 19669
rect 41049 19669 41061 19672
rect 41095 19669 41107 19703
rect 41049 19663 41107 19669
rect 41322 19660 41328 19712
rect 41380 19700 41386 19712
rect 41690 19700 41696 19712
rect 41380 19672 41696 19700
rect 41380 19660 41386 19672
rect 41690 19660 41696 19672
rect 41748 19700 41754 19712
rect 41785 19703 41843 19709
rect 41785 19700 41797 19703
rect 41748 19672 41797 19700
rect 41748 19660 41754 19672
rect 41785 19669 41797 19672
rect 41831 19669 41843 19703
rect 41785 19663 41843 19669
rect 42150 19660 42156 19712
rect 42208 19700 42214 19712
rect 43714 19700 43720 19712
rect 42208 19672 43720 19700
rect 42208 19660 42214 19672
rect 43714 19660 43720 19672
rect 43772 19660 43778 19712
rect 43993 19703 44051 19709
rect 43993 19669 44005 19703
rect 44039 19700 44051 19703
rect 44910 19700 44916 19712
rect 44039 19672 44916 19700
rect 44039 19669 44051 19672
rect 43993 19663 44051 19669
rect 44910 19660 44916 19672
rect 44968 19660 44974 19712
rect 45020 19700 45048 19740
rect 47965 19700 47993 19944
rect 53377 19941 53389 19975
rect 53423 19972 53435 19975
rect 53926 19972 53932 19984
rect 53423 19944 53932 19972
rect 53423 19941 53435 19944
rect 53377 19935 53435 19941
rect 53926 19932 53932 19944
rect 53984 19932 53990 19984
rect 48041 19907 48099 19913
rect 48041 19873 48053 19907
rect 48087 19904 48099 19907
rect 50893 19907 50951 19913
rect 50893 19904 50905 19907
rect 48087 19876 50905 19904
rect 48087 19873 48099 19876
rect 48041 19867 48099 19873
rect 50893 19873 50905 19876
rect 50939 19873 50951 19907
rect 50893 19867 50951 19873
rect 53558 19864 53564 19916
rect 53616 19904 53622 19916
rect 54481 19907 54539 19913
rect 54481 19904 54493 19907
rect 53616 19876 54493 19904
rect 53616 19864 53622 19876
rect 54481 19873 54493 19876
rect 54527 19873 54539 19907
rect 54481 19867 54539 19873
rect 55398 19864 55404 19916
rect 55456 19904 55462 19916
rect 55861 19907 55919 19913
rect 55861 19904 55873 19907
rect 55456 19876 55873 19904
rect 55456 19864 55462 19876
rect 55861 19873 55873 19876
rect 55907 19873 55919 19907
rect 55861 19867 55919 19873
rect 58161 19907 58219 19913
rect 58161 19873 58173 19907
rect 58207 19904 58219 19907
rect 58250 19904 58256 19916
rect 58207 19876 58256 19904
rect 58207 19873 58219 19876
rect 58161 19867 58219 19873
rect 58250 19864 58256 19876
rect 58308 19864 58314 19916
rect 48130 19796 48136 19848
rect 48188 19796 48194 19848
rect 48501 19839 48559 19845
rect 48501 19805 48513 19839
rect 48547 19805 48559 19839
rect 48501 19799 48559 19805
rect 48516 19768 48544 19799
rect 48590 19796 48596 19848
rect 48648 19836 48654 19848
rect 49053 19839 49111 19845
rect 49053 19836 49065 19839
rect 48648 19808 49065 19836
rect 48648 19796 48654 19808
rect 49053 19805 49065 19808
rect 49099 19805 49111 19839
rect 49053 19799 49111 19805
rect 48958 19768 48964 19780
rect 48516 19740 48964 19768
rect 48958 19728 48964 19740
rect 49016 19728 49022 19780
rect 49068 19768 49096 19799
rect 49142 19796 49148 19848
rect 49200 19796 49206 19848
rect 50522 19836 50528 19848
rect 50483 19808 50528 19836
rect 50522 19796 50528 19808
rect 50580 19796 50586 19848
rect 50985 19839 51043 19845
rect 50985 19805 50997 19839
rect 51031 19836 51043 19839
rect 51258 19836 51264 19848
rect 51031 19808 51264 19836
rect 51031 19805 51043 19808
rect 50985 19799 51043 19805
rect 51258 19796 51264 19808
rect 51316 19836 51322 19848
rect 51902 19836 51908 19848
rect 51316 19808 51908 19836
rect 51316 19796 51322 19808
rect 51902 19796 51908 19808
rect 51960 19796 51966 19848
rect 51997 19839 52055 19845
rect 51997 19805 52009 19839
rect 52043 19836 52055 19839
rect 54018 19839 54076 19845
rect 52043 19808 52408 19836
rect 52043 19805 52055 19808
rect 51997 19799 52055 19805
rect 49234 19768 49240 19780
rect 49068 19740 49240 19768
rect 49234 19728 49240 19740
rect 49292 19728 49298 19780
rect 49510 19728 49516 19780
rect 49568 19768 49574 19780
rect 49568 19740 50660 19768
rect 49568 19728 49574 19740
rect 45020 19672 47993 19700
rect 49326 19660 49332 19712
rect 49384 19660 49390 19712
rect 50154 19660 50160 19712
rect 50212 19700 50218 19712
rect 50341 19703 50399 19709
rect 50341 19700 50353 19703
rect 50212 19672 50353 19700
rect 50212 19660 50218 19672
rect 50341 19669 50353 19672
rect 50387 19669 50399 19703
rect 50341 19663 50399 19669
rect 50430 19660 50436 19712
rect 50488 19700 50494 19712
rect 50525 19703 50583 19709
rect 50525 19700 50537 19703
rect 50488 19672 50537 19700
rect 50488 19660 50494 19672
rect 50525 19669 50537 19672
rect 50571 19669 50583 19703
rect 50632 19700 50660 19740
rect 51074 19728 51080 19780
rect 51132 19768 51138 19780
rect 52012 19768 52040 19799
rect 52380 19780 52408 19808
rect 54018 19805 54030 19839
rect 54064 19836 54076 19839
rect 54110 19836 54116 19848
rect 54064 19808 54116 19836
rect 54064 19805 54076 19808
rect 54018 19799 54076 19805
rect 54110 19796 54116 19808
rect 54168 19796 54174 19848
rect 54386 19796 54392 19848
rect 54444 19796 54450 19848
rect 56042 19796 56048 19848
rect 56100 19796 56106 19848
rect 57885 19839 57943 19845
rect 57885 19805 57897 19839
rect 57931 19805 57943 19839
rect 57885 19799 57943 19805
rect 51132 19740 52040 19768
rect 51132 19728 51138 19740
rect 52086 19728 52092 19780
rect 52144 19768 52150 19780
rect 52242 19771 52300 19777
rect 52242 19768 52254 19771
rect 52144 19740 52254 19768
rect 52144 19728 52150 19740
rect 52242 19737 52254 19740
rect 52288 19737 52300 19771
rect 52242 19731 52300 19737
rect 52362 19728 52368 19780
rect 52420 19728 52426 19780
rect 57900 19768 57928 19799
rect 53300 19740 57928 19768
rect 53300 19700 53328 19740
rect 50632 19672 53328 19700
rect 50525 19663 50583 19669
rect 54018 19660 54024 19712
rect 54076 19660 54082 19712
rect 1104 19610 58880 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 50294 19610
rect 50346 19558 50358 19610
rect 50410 19558 50422 19610
rect 50474 19558 50486 19610
rect 50538 19558 50550 19610
rect 50602 19558 58880 19610
rect 1104 19536 58880 19558
rect 20625 19499 20683 19505
rect 20625 19465 20637 19499
rect 20671 19465 20683 19499
rect 20625 19459 20683 19465
rect 21361 19499 21419 19505
rect 21361 19465 21373 19499
rect 21407 19465 21419 19499
rect 21361 19459 21419 19465
rect 1026 19388 1032 19440
rect 1084 19428 1090 19440
rect 1857 19431 1915 19437
rect 1857 19428 1869 19431
rect 1084 19400 1869 19428
rect 1084 19388 1090 19400
rect 1857 19397 1869 19400
rect 1903 19397 1915 19431
rect 1857 19391 1915 19397
rect 1581 19363 1639 19369
rect 1581 19329 1593 19363
rect 1627 19360 1639 19363
rect 18782 19360 18788 19372
rect 1627 19332 18788 19360
rect 1627 19329 1639 19332
rect 1581 19323 1639 19329
rect 18782 19320 18788 19332
rect 18840 19320 18846 19372
rect 20441 19363 20499 19369
rect 20441 19329 20453 19363
rect 20487 19360 20499 19363
rect 20530 19360 20536 19372
rect 20487 19332 20536 19360
rect 20487 19329 20499 19332
rect 20441 19323 20499 19329
rect 20530 19320 20536 19332
rect 20588 19320 20594 19372
rect 20640 19360 20668 19459
rect 21177 19363 21235 19369
rect 21177 19360 21189 19363
rect 20640 19332 21189 19360
rect 21177 19329 21189 19332
rect 21223 19329 21235 19363
rect 21376 19360 21404 19459
rect 22370 19456 22376 19508
rect 22428 19496 22434 19508
rect 26513 19499 26571 19505
rect 22428 19468 24532 19496
rect 22428 19456 22434 19468
rect 24394 19428 24400 19440
rect 22848 19400 24400 19428
rect 22848 19369 22876 19400
rect 24394 19388 24400 19400
rect 24452 19388 24458 19440
rect 24504 19428 24532 19468
rect 26513 19465 26525 19499
rect 26559 19496 26571 19499
rect 27614 19496 27620 19508
rect 26559 19468 27620 19496
rect 26559 19465 26571 19468
rect 26513 19459 26571 19465
rect 27614 19456 27620 19468
rect 27672 19456 27678 19508
rect 28350 19456 28356 19508
rect 28408 19496 28414 19508
rect 28445 19499 28503 19505
rect 28445 19496 28457 19499
rect 28408 19468 28457 19496
rect 28408 19456 28414 19468
rect 28445 19465 28457 19468
rect 28491 19465 28503 19499
rect 28445 19459 28503 19465
rect 28626 19456 28632 19508
rect 28684 19496 28690 19508
rect 34330 19496 34336 19508
rect 28684 19468 34336 19496
rect 28684 19456 28690 19468
rect 34330 19456 34336 19468
rect 34388 19456 34394 19508
rect 34609 19499 34667 19505
rect 34609 19465 34621 19499
rect 34655 19465 34667 19499
rect 34609 19459 34667 19465
rect 29362 19428 29368 19440
rect 24504 19400 29368 19428
rect 29362 19388 29368 19400
rect 29420 19388 29426 19440
rect 34624 19428 34652 19459
rect 34790 19456 34796 19508
rect 34848 19496 34854 19508
rect 35253 19499 35311 19505
rect 35253 19496 35265 19499
rect 34848 19468 35265 19496
rect 34848 19456 34854 19468
rect 35253 19465 35265 19468
rect 35299 19465 35311 19499
rect 35253 19459 35311 19465
rect 36078 19456 36084 19508
rect 36136 19456 36142 19508
rect 36173 19499 36231 19505
rect 36173 19465 36185 19499
rect 36219 19496 36231 19499
rect 37182 19496 37188 19508
rect 36219 19468 37188 19496
rect 36219 19465 36231 19468
rect 36173 19459 36231 19465
rect 37182 19456 37188 19468
rect 37240 19456 37246 19508
rect 37458 19456 37464 19508
rect 37516 19496 37522 19508
rect 37559 19499 37617 19505
rect 37559 19496 37571 19499
rect 37516 19468 37571 19496
rect 37516 19456 37522 19468
rect 37559 19465 37571 19468
rect 37605 19465 37617 19499
rect 37559 19459 37617 19465
rect 37645 19499 37703 19505
rect 37645 19465 37657 19499
rect 37691 19496 37703 19499
rect 37826 19496 37832 19508
rect 37691 19468 37832 19496
rect 37691 19465 37703 19468
rect 37645 19459 37703 19465
rect 37826 19456 37832 19468
rect 37884 19456 37890 19508
rect 39577 19499 39635 19505
rect 39577 19496 39589 19499
rect 38212 19468 39589 19496
rect 34624 19400 35848 19428
rect 22005 19363 22063 19369
rect 22005 19360 22017 19363
rect 21376 19332 22017 19360
rect 21177 19323 21235 19329
rect 22005 19329 22017 19332
rect 22051 19329 22063 19363
rect 22005 19323 22063 19329
rect 22833 19363 22891 19369
rect 22833 19329 22845 19363
rect 22879 19329 22891 19363
rect 22833 19323 22891 19329
rect 23106 19320 23112 19372
rect 23164 19320 23170 19372
rect 24029 19363 24087 19369
rect 24029 19329 24041 19363
rect 24075 19329 24087 19363
rect 24029 19323 24087 19329
rect 11698 19252 11704 19304
rect 11756 19292 11762 19304
rect 23293 19295 23351 19301
rect 23293 19292 23305 19295
rect 11756 19264 23305 19292
rect 11756 19252 11762 19264
rect 23293 19261 23305 19264
rect 23339 19261 23351 19295
rect 24044 19292 24072 19323
rect 24118 19320 24124 19372
rect 24176 19360 24182 19372
rect 24578 19360 24584 19372
rect 24176 19332 24221 19360
rect 24320 19332 24584 19360
rect 24176 19320 24182 19332
rect 24320 19292 24348 19332
rect 24578 19320 24584 19332
rect 24636 19360 24642 19372
rect 25314 19360 25320 19372
rect 24636 19332 25320 19360
rect 24636 19320 24642 19332
rect 25314 19320 25320 19332
rect 25372 19320 25378 19372
rect 26329 19363 26387 19369
rect 26329 19329 26341 19363
rect 26375 19360 26387 19363
rect 27341 19363 27399 19369
rect 26375 19332 27292 19360
rect 26375 19329 26387 19332
rect 26329 19323 26387 19329
rect 24044 19264 24348 19292
rect 23293 19255 23351 19261
rect 22922 19184 22928 19236
rect 22980 19184 22986 19236
rect 22094 19116 22100 19168
rect 22152 19156 22158 19168
rect 22189 19159 22247 19165
rect 22189 19156 22201 19159
rect 22152 19128 22201 19156
rect 22152 19116 22158 19128
rect 22189 19125 22201 19128
rect 22235 19125 22247 19159
rect 27264 19156 27292 19332
rect 27341 19329 27353 19363
rect 27387 19360 27399 19363
rect 27387 19332 28212 19360
rect 27387 19329 27399 19332
rect 27341 19323 27399 19329
rect 27433 19295 27491 19301
rect 27433 19261 27445 19295
rect 27479 19261 27491 19295
rect 28184 19292 28212 19332
rect 28258 19320 28264 19372
rect 28316 19320 28322 19372
rect 30650 19360 30656 19372
rect 28368 19332 30656 19360
rect 28368 19292 28396 19332
rect 30650 19320 30656 19332
rect 30708 19320 30714 19372
rect 33042 19320 33048 19372
rect 33100 19360 33106 19372
rect 33229 19363 33287 19369
rect 33229 19360 33241 19363
rect 33100 19332 33241 19360
rect 33100 19320 33106 19332
rect 33229 19329 33241 19332
rect 33275 19329 33287 19363
rect 33229 19323 33287 19329
rect 33496 19363 33554 19369
rect 33496 19329 33508 19363
rect 33542 19360 33554 19363
rect 34606 19360 34612 19372
rect 33542 19332 34612 19360
rect 33542 19329 33554 19332
rect 33496 19323 33554 19329
rect 34606 19320 34612 19332
rect 34664 19320 34670 19372
rect 35069 19363 35127 19369
rect 35069 19329 35081 19363
rect 35115 19360 35127 19363
rect 35342 19360 35348 19372
rect 35115 19332 35348 19360
rect 35115 19329 35127 19332
rect 35069 19323 35127 19329
rect 35342 19320 35348 19332
rect 35400 19320 35406 19372
rect 35820 19360 35848 19400
rect 35894 19388 35900 19440
rect 35952 19428 35958 19440
rect 36357 19431 36415 19437
rect 36357 19428 36369 19431
rect 35952 19400 36369 19428
rect 35952 19388 35958 19400
rect 36357 19397 36369 19400
rect 36403 19428 36415 19431
rect 36538 19428 36544 19440
rect 36403 19400 36544 19428
rect 36403 19397 36415 19400
rect 36357 19391 36415 19397
rect 36538 19388 36544 19400
rect 36596 19428 36602 19440
rect 38212 19428 38240 19468
rect 39577 19465 39589 19468
rect 39623 19465 39635 19499
rect 39577 19459 39635 19465
rect 38470 19437 38476 19440
rect 36596 19400 37780 19428
rect 36596 19388 36602 19400
rect 35820 19332 35940 19360
rect 28184 19264 28396 19292
rect 35912 19292 35940 19332
rect 35986 19320 35992 19372
rect 36044 19320 36050 19372
rect 37461 19363 37519 19369
rect 36096 19332 37412 19360
rect 36096 19292 36124 19332
rect 35912 19264 36124 19292
rect 37384 19292 37412 19332
rect 37461 19329 37473 19363
rect 37507 19360 37519 19363
rect 37550 19360 37556 19372
rect 37507 19332 37556 19360
rect 37507 19329 37519 19332
rect 37461 19323 37519 19329
rect 37550 19320 37556 19332
rect 37608 19320 37614 19372
rect 37752 19369 37780 19400
rect 37844 19400 38240 19428
rect 37737 19363 37795 19369
rect 37737 19329 37749 19363
rect 37783 19329 37795 19363
rect 37737 19323 37795 19329
rect 37844 19292 37872 19400
rect 38464 19391 38476 19437
rect 38470 19388 38476 19391
rect 38528 19388 38534 19440
rect 39592 19428 39620 19459
rect 40034 19456 40040 19508
rect 40092 19496 40098 19508
rect 40221 19499 40279 19505
rect 40221 19496 40233 19499
rect 40092 19468 40233 19496
rect 40092 19456 40098 19468
rect 40221 19465 40233 19468
rect 40267 19465 40279 19499
rect 40221 19459 40279 19465
rect 40954 19456 40960 19508
rect 41012 19456 41018 19508
rect 41138 19456 41144 19508
rect 41196 19456 41202 19508
rect 44177 19499 44235 19505
rect 44177 19465 44189 19499
rect 44223 19496 44235 19499
rect 44450 19496 44456 19508
rect 44223 19468 44456 19496
rect 44223 19465 44235 19468
rect 44177 19459 44235 19465
rect 44450 19456 44456 19468
rect 44508 19456 44514 19508
rect 46014 19496 46020 19508
rect 44560 19468 46020 19496
rect 39592 19400 42656 19428
rect 38194 19320 38200 19372
rect 38252 19320 38258 19372
rect 38304 19332 39252 19360
rect 38304 19292 38332 19332
rect 37384 19264 37872 19292
rect 37936 19264 38332 19292
rect 27433 19255 27491 19261
rect 27448 19224 27476 19255
rect 28626 19224 28632 19236
rect 27448 19196 28632 19224
rect 28626 19184 28632 19196
rect 28684 19184 28690 19236
rect 35805 19227 35863 19233
rect 35805 19193 35817 19227
rect 35851 19193 35863 19227
rect 35805 19187 35863 19193
rect 27709 19159 27767 19165
rect 27709 19156 27721 19159
rect 27264 19128 27721 19156
rect 22189 19119 22247 19125
rect 27709 19125 27721 19128
rect 27755 19125 27767 19159
rect 35820 19156 35848 19187
rect 36354 19184 36360 19236
rect 36412 19224 36418 19236
rect 36906 19224 36912 19236
rect 36412 19196 36912 19224
rect 36412 19184 36418 19196
rect 36906 19184 36912 19196
rect 36964 19224 36970 19236
rect 37936 19224 37964 19264
rect 36964 19196 37964 19224
rect 39224 19224 39252 19332
rect 40034 19320 40040 19372
rect 40092 19320 40098 19372
rect 40218 19320 40224 19372
rect 40276 19360 40282 19372
rect 41082 19363 41140 19369
rect 41082 19360 41094 19363
rect 40276 19332 41094 19360
rect 40276 19320 40282 19332
rect 41082 19329 41094 19332
rect 41128 19360 41140 19363
rect 41230 19360 41236 19372
rect 41128 19332 41236 19360
rect 41128 19329 41140 19332
rect 41082 19323 41140 19329
rect 41230 19320 41236 19332
rect 41288 19320 41294 19372
rect 42628 19369 42656 19400
rect 42702 19388 42708 19440
rect 42760 19428 42766 19440
rect 43438 19428 43444 19440
rect 42760 19400 43444 19428
rect 42760 19388 42766 19400
rect 43438 19388 43444 19400
rect 43496 19428 43502 19440
rect 43809 19431 43867 19437
rect 43809 19428 43821 19431
rect 43496 19400 43821 19428
rect 43496 19388 43502 19400
rect 43809 19397 43821 19400
rect 43855 19397 43867 19431
rect 43809 19391 43867 19397
rect 42613 19363 42671 19369
rect 41524 19332 42104 19360
rect 39666 19252 39672 19304
rect 39724 19292 39730 19304
rect 41524 19292 41552 19332
rect 39724 19264 41552 19292
rect 41601 19295 41659 19301
rect 39724 19252 39730 19264
rect 41601 19261 41613 19295
rect 41647 19292 41659 19295
rect 41966 19292 41972 19304
rect 41647 19264 41972 19292
rect 41647 19261 41659 19264
rect 41601 19255 41659 19261
rect 41966 19252 41972 19264
rect 42024 19252 42030 19304
rect 42076 19292 42104 19332
rect 42613 19329 42625 19363
rect 42659 19329 42671 19363
rect 43824 19360 43852 19391
rect 43990 19388 43996 19440
rect 44048 19428 44054 19440
rect 44560 19428 44588 19468
rect 46014 19456 46020 19468
rect 46072 19456 46078 19508
rect 46569 19499 46627 19505
rect 46569 19465 46581 19499
rect 46615 19496 46627 19499
rect 49142 19496 49148 19508
rect 46615 19468 49148 19496
rect 46615 19465 46627 19468
rect 46569 19459 46627 19465
rect 49142 19456 49148 19468
rect 49200 19456 49206 19508
rect 49510 19456 49516 19508
rect 49568 19496 49574 19508
rect 49697 19499 49755 19505
rect 49697 19496 49709 19499
rect 49568 19468 49709 19496
rect 49568 19456 49574 19468
rect 49697 19465 49709 19468
rect 49743 19465 49755 19499
rect 49697 19459 49755 19465
rect 50062 19456 50068 19508
rect 50120 19496 50126 19508
rect 50249 19499 50307 19505
rect 50249 19496 50261 19499
rect 50120 19468 50261 19496
rect 50120 19456 50126 19468
rect 50249 19465 50261 19468
rect 50295 19465 50307 19499
rect 50249 19459 50307 19465
rect 50356 19468 51074 19496
rect 44910 19437 44916 19440
rect 44904 19428 44916 19437
rect 44048 19400 44588 19428
rect 44871 19400 44916 19428
rect 44048 19388 44054 19400
rect 44904 19391 44916 19400
rect 44910 19388 44916 19391
rect 44968 19388 44974 19440
rect 46842 19388 46848 19440
rect 46900 19388 46906 19440
rect 46937 19431 46995 19437
rect 46937 19397 46949 19431
rect 46983 19428 46995 19431
rect 48038 19428 48044 19440
rect 46983 19400 48044 19428
rect 46983 19397 46995 19400
rect 46937 19391 46995 19397
rect 48038 19388 48044 19400
rect 48096 19388 48102 19440
rect 48584 19431 48642 19437
rect 48240 19400 48544 19428
rect 44450 19360 44456 19372
rect 43824 19332 44456 19360
rect 42613 19323 42671 19329
rect 44450 19320 44456 19332
rect 44508 19320 44514 19372
rect 44634 19320 44640 19372
rect 44692 19320 44698 19372
rect 46753 19363 46811 19369
rect 46753 19329 46765 19363
rect 46799 19360 46811 19363
rect 47075 19363 47133 19369
rect 46799 19332 46888 19360
rect 46799 19329 46811 19332
rect 46753 19323 46811 19329
rect 44358 19292 44364 19304
rect 42076 19264 44364 19292
rect 44358 19252 44364 19264
rect 44416 19252 44422 19304
rect 46860 19292 46888 19332
rect 47075 19329 47087 19363
rect 47121 19360 47133 19363
rect 48130 19360 48136 19372
rect 47121 19332 48136 19360
rect 47121 19329 47133 19332
rect 47075 19323 47133 19329
rect 48130 19320 48136 19332
rect 48188 19320 48194 19372
rect 47213 19295 47271 19301
rect 46860 19264 47164 19292
rect 47136 19236 47164 19264
rect 47213 19261 47225 19295
rect 47259 19292 47271 19295
rect 48240 19292 48268 19400
rect 48317 19363 48375 19369
rect 48317 19329 48329 19363
rect 48363 19360 48375 19363
rect 48406 19360 48412 19372
rect 48363 19332 48412 19360
rect 48363 19329 48375 19332
rect 48317 19323 48375 19329
rect 48406 19320 48412 19332
rect 48464 19320 48470 19372
rect 48516 19360 48544 19400
rect 48584 19397 48596 19431
rect 48630 19428 48642 19431
rect 49326 19428 49332 19440
rect 48630 19400 49332 19428
rect 48630 19397 48642 19400
rect 48584 19391 48642 19397
rect 49326 19388 49332 19400
rect 49384 19388 49390 19440
rect 49528 19360 49556 19456
rect 49786 19388 49792 19440
rect 49844 19428 49850 19440
rect 50356 19428 50384 19468
rect 49844 19400 50384 19428
rect 49844 19388 49850 19400
rect 48516 19332 49556 19360
rect 50154 19320 50160 19372
rect 50212 19320 50218 19372
rect 50356 19369 50384 19400
rect 50341 19363 50399 19369
rect 50341 19329 50353 19363
rect 50387 19329 50399 19363
rect 50341 19323 50399 19329
rect 47259 19264 48268 19292
rect 51046 19292 51074 19468
rect 52086 19456 52092 19508
rect 52144 19456 52150 19508
rect 53558 19496 53564 19508
rect 52196 19468 53564 19496
rect 51902 19388 51908 19440
rect 51960 19428 51966 19440
rect 52196 19428 52224 19468
rect 53558 19456 53564 19468
rect 53616 19456 53622 19508
rect 54110 19456 54116 19508
rect 54168 19496 54174 19508
rect 54297 19499 54355 19505
rect 54297 19496 54309 19499
rect 54168 19468 54309 19496
rect 54168 19456 54174 19468
rect 54297 19465 54309 19468
rect 54343 19496 54355 19499
rect 56502 19496 56508 19508
rect 54343 19468 56508 19496
rect 54343 19465 54355 19468
rect 54297 19459 54355 19465
rect 56502 19456 56508 19468
rect 56560 19456 56566 19508
rect 56594 19456 56600 19508
rect 56652 19496 56658 19508
rect 57149 19499 57207 19505
rect 57149 19496 57161 19499
rect 56652 19468 57161 19496
rect 56652 19456 56658 19468
rect 57149 19465 57161 19468
rect 57195 19496 57207 19499
rect 57882 19496 57888 19508
rect 57195 19468 57888 19496
rect 57195 19465 57207 19468
rect 57149 19459 57207 19465
rect 57882 19456 57888 19468
rect 57940 19456 57946 19508
rect 51960 19400 52224 19428
rect 51960 19388 51966 19400
rect 52362 19388 52368 19440
rect 52420 19428 52426 19440
rect 52420 19400 55812 19428
rect 52420 19388 52426 19400
rect 51994 19320 52000 19372
rect 52052 19320 52058 19372
rect 52086 19320 52092 19372
rect 52144 19360 52150 19372
rect 52932 19369 52960 19400
rect 55784 19372 55812 19400
rect 52181 19363 52239 19369
rect 52181 19360 52193 19363
rect 52144 19332 52193 19360
rect 52144 19320 52150 19332
rect 52181 19329 52193 19332
rect 52227 19329 52239 19363
rect 52181 19323 52239 19329
rect 52917 19363 52975 19369
rect 52917 19329 52929 19363
rect 52963 19329 52975 19363
rect 52917 19323 52975 19329
rect 53006 19320 53012 19372
rect 53064 19360 53070 19372
rect 53173 19363 53231 19369
rect 53173 19360 53185 19363
rect 53064 19332 53185 19360
rect 53064 19320 53070 19332
rect 53173 19329 53185 19332
rect 53219 19329 53231 19363
rect 53173 19323 53231 19329
rect 55766 19320 55772 19372
rect 55824 19320 55830 19372
rect 55858 19320 55864 19372
rect 55916 19360 55922 19372
rect 56025 19363 56083 19369
rect 56025 19360 56037 19363
rect 55916 19332 56037 19360
rect 55916 19320 55922 19332
rect 56025 19329 56037 19332
rect 56071 19329 56083 19363
rect 56025 19323 56083 19329
rect 58161 19363 58219 19369
rect 58161 19329 58173 19363
rect 58207 19360 58219 19363
rect 58986 19360 58992 19372
rect 58207 19332 58992 19360
rect 58207 19329 58219 19332
rect 58161 19323 58219 19329
rect 58986 19320 58992 19332
rect 59044 19320 59050 19372
rect 52270 19292 52276 19304
rect 51046 19264 52276 19292
rect 47259 19261 47271 19264
rect 47213 19255 47271 19261
rect 52270 19252 52276 19264
rect 52328 19252 52334 19304
rect 39224 19196 41552 19224
rect 36964 19184 36970 19196
rect 41322 19156 41328 19168
rect 35820 19128 41328 19156
rect 27709 19119 27767 19125
rect 41322 19116 41328 19128
rect 41380 19116 41386 19168
rect 41524 19165 41552 19196
rect 45940 19196 46704 19224
rect 41509 19159 41567 19165
rect 41509 19125 41521 19159
rect 41555 19125 41567 19159
rect 41509 19119 41567 19125
rect 41598 19116 41604 19168
rect 41656 19156 41662 19168
rect 42797 19159 42855 19165
rect 42797 19156 42809 19159
rect 41656 19128 42809 19156
rect 41656 19116 41662 19128
rect 42797 19125 42809 19128
rect 42843 19125 42855 19159
rect 42797 19119 42855 19125
rect 44266 19116 44272 19168
rect 44324 19156 44330 19168
rect 45940 19156 45968 19196
rect 44324 19128 45968 19156
rect 44324 19116 44330 19128
rect 46014 19116 46020 19168
rect 46072 19116 46078 19168
rect 46676 19156 46704 19196
rect 47118 19184 47124 19236
rect 47176 19184 47182 19236
rect 58345 19227 58403 19233
rect 58345 19224 58357 19227
rect 49620 19196 49832 19224
rect 49620 19156 49648 19196
rect 46676 19128 49648 19156
rect 49804 19156 49832 19196
rect 54220 19196 54432 19224
rect 54220 19156 54248 19196
rect 49804 19128 54248 19156
rect 54404 19156 54432 19196
rect 56704 19196 58357 19224
rect 56704 19156 56732 19196
rect 58345 19193 58357 19196
rect 58391 19193 58403 19227
rect 58345 19187 58403 19193
rect 54404 19128 56732 19156
rect 1104 19066 58880 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 58880 19066
rect 1104 18992 58880 19014
rect 20714 18912 20720 18964
rect 20772 18952 20778 18964
rect 21085 18955 21143 18961
rect 21085 18952 21097 18955
rect 20772 18924 21097 18952
rect 20772 18912 20778 18924
rect 21085 18921 21097 18924
rect 21131 18921 21143 18955
rect 21085 18915 21143 18921
rect 23201 18955 23259 18961
rect 23201 18921 23213 18955
rect 23247 18952 23259 18955
rect 26418 18952 26424 18964
rect 23247 18924 26424 18952
rect 23247 18921 23259 18924
rect 23201 18915 23259 18921
rect 26418 18912 26424 18924
rect 26476 18912 26482 18964
rect 27062 18912 27068 18964
rect 27120 18912 27126 18964
rect 29733 18955 29791 18961
rect 29733 18921 29745 18955
rect 29779 18952 29791 18955
rect 34422 18952 34428 18964
rect 29779 18924 34428 18952
rect 29779 18921 29791 18924
rect 29733 18915 29791 18921
rect 34422 18912 34428 18924
rect 34480 18912 34486 18964
rect 35161 18955 35219 18961
rect 35161 18921 35173 18955
rect 35207 18952 35219 18955
rect 35342 18952 35348 18964
rect 35207 18924 35348 18952
rect 35207 18921 35219 18924
rect 35161 18915 35219 18921
rect 35342 18912 35348 18924
rect 35400 18912 35406 18964
rect 36538 18912 36544 18964
rect 36596 18912 36602 18964
rect 38381 18955 38439 18961
rect 36639 18924 37504 18952
rect 24762 18844 24768 18896
rect 24820 18884 24826 18896
rect 33410 18884 33416 18896
rect 24820 18856 25268 18884
rect 24820 18844 24826 18856
rect 20901 18819 20959 18825
rect 20901 18785 20913 18819
rect 20947 18816 20959 18819
rect 21913 18819 21971 18825
rect 20947 18788 21772 18816
rect 20947 18785 20959 18788
rect 20901 18779 20959 18785
rect 21744 18760 21772 18788
rect 21913 18785 21925 18819
rect 21959 18816 21971 18819
rect 22094 18816 22100 18828
rect 21959 18788 22100 18816
rect 21959 18785 21971 18788
rect 21913 18779 21971 18785
rect 22094 18776 22100 18788
rect 22152 18776 22158 18828
rect 24394 18776 24400 18828
rect 24452 18816 24458 18828
rect 25240 18816 25268 18856
rect 29932 18856 33416 18884
rect 25869 18819 25927 18825
rect 25869 18816 25881 18819
rect 24452 18788 25084 18816
rect 24452 18776 24458 18788
rect 1581 18751 1639 18757
rect 1581 18717 1593 18751
rect 1627 18748 1639 18751
rect 12250 18748 12256 18760
rect 1627 18720 12256 18748
rect 1627 18717 1639 18720
rect 1581 18711 1639 18717
rect 12250 18708 12256 18720
rect 12308 18708 12314 18760
rect 20806 18708 20812 18760
rect 20864 18708 20870 18760
rect 21542 18708 21548 18760
rect 21600 18748 21606 18760
rect 21637 18751 21695 18757
rect 21637 18748 21649 18751
rect 21600 18720 21649 18748
rect 21600 18708 21606 18720
rect 21637 18717 21649 18720
rect 21683 18717 21695 18751
rect 21637 18711 21695 18717
rect 21726 18708 21732 18760
rect 21784 18708 21790 18760
rect 24578 18708 24584 18760
rect 24636 18748 24642 18760
rect 25056 18757 25084 18788
rect 25240 18788 25881 18816
rect 25240 18757 25268 18788
rect 25869 18785 25881 18788
rect 25915 18785 25927 18819
rect 25869 18779 25927 18785
rect 24765 18751 24823 18757
rect 24765 18748 24777 18751
rect 24636 18720 24777 18748
rect 24636 18708 24642 18720
rect 24765 18717 24777 18720
rect 24811 18717 24823 18751
rect 24765 18711 24823 18717
rect 25041 18751 25099 18757
rect 25041 18717 25053 18751
rect 25087 18717 25099 18751
rect 25041 18711 25099 18717
rect 25225 18751 25283 18757
rect 25225 18717 25237 18751
rect 25271 18717 25283 18751
rect 25225 18711 25283 18717
rect 25685 18751 25743 18757
rect 25685 18717 25697 18751
rect 25731 18717 25743 18751
rect 25685 18711 25743 18717
rect 26881 18751 26939 18757
rect 26881 18717 26893 18751
rect 26927 18717 26939 18751
rect 26881 18711 26939 18717
rect 934 18640 940 18692
rect 992 18680 998 18692
rect 1857 18683 1915 18689
rect 1857 18680 1869 18683
rect 992 18652 1869 18680
rect 992 18640 998 18652
rect 1857 18649 1869 18652
rect 1903 18649 1915 18683
rect 1857 18643 1915 18649
rect 24854 18640 24860 18692
rect 24912 18680 24918 18692
rect 25700 18680 25728 18711
rect 24912 18652 25728 18680
rect 26896 18680 26924 18711
rect 27614 18708 27620 18760
rect 27672 18708 27678 18760
rect 29932 18757 29960 18856
rect 33410 18844 33416 18856
rect 33468 18844 33474 18896
rect 33505 18887 33563 18893
rect 33505 18853 33517 18887
rect 33551 18884 33563 18887
rect 34790 18884 34796 18896
rect 33551 18856 34796 18884
rect 33551 18853 33563 18856
rect 33505 18847 33563 18853
rect 34790 18844 34796 18856
rect 34848 18844 34854 18896
rect 35986 18844 35992 18896
rect 36044 18884 36050 18896
rect 36639 18884 36667 18924
rect 36044 18856 36667 18884
rect 37369 18887 37427 18893
rect 36044 18844 36050 18856
rect 37369 18853 37381 18887
rect 37415 18853 37427 18887
rect 37476 18884 37504 18924
rect 38381 18921 38393 18955
rect 38427 18952 38439 18955
rect 38470 18952 38476 18964
rect 38427 18924 38476 18952
rect 38427 18921 38439 18924
rect 38381 18915 38439 18921
rect 38470 18912 38476 18924
rect 38528 18912 38534 18964
rect 40221 18955 40279 18961
rect 40221 18921 40233 18955
rect 40267 18952 40279 18955
rect 40402 18952 40408 18964
rect 40267 18924 40408 18952
rect 40267 18921 40279 18924
rect 40221 18915 40279 18921
rect 40402 18912 40408 18924
rect 40460 18912 40466 18964
rect 44545 18955 44603 18961
rect 44545 18921 44557 18955
rect 44591 18952 44603 18955
rect 45922 18952 45928 18964
rect 44591 18924 45928 18952
rect 44591 18921 44603 18924
rect 44545 18915 44603 18921
rect 45922 18912 45928 18924
rect 45980 18912 45986 18964
rect 47118 18912 47124 18964
rect 47176 18952 47182 18964
rect 47305 18955 47363 18961
rect 47305 18952 47317 18955
rect 47176 18924 47317 18952
rect 47176 18912 47182 18924
rect 47305 18921 47317 18924
rect 47351 18921 47363 18955
rect 47305 18915 47363 18921
rect 55674 18912 55680 18964
rect 55732 18952 55738 18964
rect 55732 18924 56180 18952
rect 55732 18912 55738 18924
rect 56152 18896 56180 18924
rect 37476 18856 40080 18884
rect 37369 18847 37427 18853
rect 33870 18816 33876 18828
rect 32324 18788 33876 18816
rect 32324 18757 32352 18788
rect 33870 18776 33876 18788
rect 33928 18776 33934 18828
rect 37384 18816 37412 18847
rect 34992 18788 37412 18816
rect 38856 18788 39988 18816
rect 29917 18751 29975 18757
rect 29917 18717 29929 18751
rect 29963 18717 29975 18751
rect 29917 18711 29975 18717
rect 30193 18751 30251 18757
rect 30193 18717 30205 18751
rect 30239 18717 30251 18751
rect 30193 18711 30251 18717
rect 32309 18751 32367 18757
rect 32309 18717 32321 18751
rect 32355 18717 32367 18751
rect 32309 18711 32367 18717
rect 26896 18652 27844 18680
rect 24912 18640 24918 18652
rect 24581 18615 24639 18621
rect 24581 18581 24593 18615
rect 24627 18612 24639 18615
rect 26326 18612 26332 18624
rect 24627 18584 26332 18612
rect 24627 18581 24639 18584
rect 24581 18575 24639 18581
rect 26326 18572 26332 18584
rect 26384 18572 26390 18624
rect 27816 18621 27844 18652
rect 29546 18640 29552 18692
rect 29604 18680 29610 18692
rect 30208 18680 30236 18711
rect 32490 18708 32496 18760
rect 32548 18708 32554 18760
rect 33321 18751 33379 18757
rect 33321 18717 33333 18751
rect 33367 18717 33379 18751
rect 33321 18711 33379 18717
rect 34057 18751 34115 18757
rect 34057 18717 34069 18751
rect 34103 18748 34115 18751
rect 34882 18748 34888 18760
rect 34103 18720 34888 18748
rect 34103 18717 34115 18720
rect 34057 18711 34115 18717
rect 29604 18652 30236 18680
rect 33336 18680 33364 18711
rect 34882 18708 34888 18720
rect 34940 18708 34946 18760
rect 34992 18757 35020 18788
rect 34977 18751 35035 18757
rect 34977 18717 34989 18751
rect 35023 18717 35035 18751
rect 34977 18711 35035 18717
rect 35710 18708 35716 18760
rect 35768 18708 35774 18760
rect 35897 18751 35955 18757
rect 35897 18717 35909 18751
rect 35943 18748 35955 18751
rect 36170 18748 36176 18760
rect 35943 18720 36176 18748
rect 35943 18717 35955 18720
rect 35897 18711 35955 18717
rect 36170 18708 36176 18720
rect 36228 18708 36234 18760
rect 36446 18708 36452 18760
rect 36504 18748 36510 18760
rect 37185 18751 37243 18757
rect 37185 18748 37197 18751
rect 36504 18720 37197 18748
rect 36504 18708 36510 18720
rect 37185 18717 37197 18720
rect 37231 18717 37243 18751
rect 37185 18711 37243 18717
rect 38657 18751 38715 18757
rect 38657 18717 38669 18751
rect 38703 18717 38715 18751
rect 38657 18711 38715 18717
rect 35805 18683 35863 18689
rect 35805 18680 35817 18683
rect 33336 18652 35817 18680
rect 29604 18640 29610 18652
rect 35805 18649 35817 18652
rect 35851 18649 35863 18683
rect 35805 18643 35863 18649
rect 27801 18615 27859 18621
rect 27801 18581 27813 18615
rect 27847 18581 27859 18615
rect 27801 18575 27859 18581
rect 27890 18572 27896 18624
rect 27948 18612 27954 18624
rect 30101 18615 30159 18621
rect 30101 18612 30113 18615
rect 27948 18584 30113 18612
rect 27948 18572 27954 18584
rect 30101 18581 30113 18584
rect 30147 18581 30159 18615
rect 30101 18575 30159 18581
rect 32214 18572 32220 18624
rect 32272 18612 32278 18624
rect 32401 18615 32459 18621
rect 32401 18612 32413 18615
rect 32272 18584 32413 18612
rect 32272 18572 32278 18584
rect 32401 18581 32413 18584
rect 32447 18581 32459 18615
rect 32401 18575 32459 18581
rect 34241 18615 34299 18621
rect 34241 18581 34253 18615
rect 34287 18612 34299 18615
rect 34698 18612 34704 18624
rect 34287 18584 34704 18612
rect 34287 18581 34299 18584
rect 34241 18575 34299 18581
rect 34698 18572 34704 18584
rect 34756 18572 34762 18624
rect 36188 18612 36216 18708
rect 36357 18683 36415 18689
rect 36357 18649 36369 18683
rect 36403 18680 36415 18683
rect 38672 18680 38700 18711
rect 38746 18708 38752 18760
rect 38804 18708 38810 18760
rect 38856 18757 38884 18788
rect 38841 18751 38899 18757
rect 38841 18717 38853 18751
rect 38887 18717 38899 18751
rect 38841 18711 38899 18717
rect 39025 18751 39083 18757
rect 39025 18717 39037 18751
rect 39071 18748 39083 18751
rect 39666 18748 39672 18760
rect 39071 18720 39672 18748
rect 39071 18717 39083 18720
rect 39025 18711 39083 18717
rect 39666 18708 39672 18720
rect 39724 18708 39730 18760
rect 39574 18680 39580 18692
rect 36403 18652 38608 18680
rect 38672 18652 39580 18680
rect 36403 18649 36415 18652
rect 36357 18643 36415 18649
rect 36557 18615 36615 18621
rect 36557 18612 36569 18615
rect 36188 18584 36569 18612
rect 36557 18581 36569 18584
rect 36603 18581 36615 18615
rect 36557 18575 36615 18581
rect 36722 18572 36728 18624
rect 36780 18572 36786 18624
rect 38580 18612 38608 18652
rect 38856 18624 38884 18652
rect 39574 18640 39580 18652
rect 39632 18640 39638 18692
rect 39960 18680 39988 18788
rect 40052 18757 40080 18856
rect 40862 18844 40868 18896
rect 40920 18884 40926 18896
rect 40920 18856 42748 18884
rect 40920 18844 40926 18856
rect 41506 18816 41512 18828
rect 40236 18788 41512 18816
rect 40037 18751 40095 18757
rect 40037 18717 40049 18751
rect 40083 18748 40095 18751
rect 40126 18748 40132 18760
rect 40083 18720 40132 18748
rect 40083 18717 40095 18720
rect 40037 18711 40095 18717
rect 40126 18708 40132 18720
rect 40184 18708 40190 18760
rect 40236 18680 40264 18788
rect 41506 18776 41512 18788
rect 41564 18776 41570 18828
rect 41690 18776 41696 18828
rect 41748 18776 41754 18828
rect 42720 18760 42748 18856
rect 45002 18844 45008 18896
rect 45060 18884 45066 18896
rect 52454 18884 52460 18896
rect 45060 18856 52460 18884
rect 45060 18844 45066 18856
rect 52454 18844 52460 18856
rect 52512 18844 52518 18896
rect 56134 18844 56140 18896
rect 56192 18844 56198 18896
rect 43809 18819 43867 18825
rect 43809 18785 43821 18819
rect 43855 18816 43867 18819
rect 46750 18816 46756 18828
rect 43855 18788 46756 18816
rect 43855 18785 43867 18788
rect 43809 18779 43867 18785
rect 46750 18776 46756 18788
rect 46808 18776 46814 18828
rect 48498 18776 48504 18828
rect 48556 18776 48562 18828
rect 49050 18776 49056 18828
rect 49108 18776 49114 18828
rect 55674 18776 55680 18828
rect 55732 18776 55738 18828
rect 56152 18816 56180 18844
rect 55968 18788 56180 18816
rect 40402 18708 40408 18760
rect 40460 18748 40466 18760
rect 41138 18748 41144 18760
rect 40460 18720 41144 18748
rect 40460 18708 40466 18720
rect 41138 18708 41144 18720
rect 41196 18748 41202 18760
rect 41417 18751 41475 18757
rect 41417 18748 41429 18751
rect 41196 18720 41429 18748
rect 41196 18708 41202 18720
rect 41417 18717 41429 18720
rect 41463 18717 41475 18751
rect 41417 18711 41475 18717
rect 41969 18751 42027 18757
rect 41969 18717 41981 18751
rect 42015 18717 42027 18751
rect 41969 18711 42027 18717
rect 39960 18652 40264 18680
rect 41984 18680 42012 18711
rect 42058 18708 42064 18760
rect 42116 18708 42122 18760
rect 42702 18708 42708 18760
rect 42760 18708 42766 18760
rect 43438 18708 43444 18760
rect 43496 18748 43502 18760
rect 43625 18751 43683 18757
rect 43625 18748 43637 18751
rect 43496 18720 43637 18748
rect 43496 18708 43502 18720
rect 43625 18717 43637 18720
rect 43671 18717 43683 18751
rect 43625 18711 43683 18717
rect 44361 18751 44419 18757
rect 44361 18717 44373 18751
rect 44407 18748 44419 18751
rect 46014 18748 46020 18760
rect 44407 18720 46020 18748
rect 44407 18717 44419 18720
rect 44361 18711 44419 18717
rect 46014 18708 46020 18720
rect 46072 18708 46078 18760
rect 48593 18751 48651 18757
rect 46860 18720 48084 18748
rect 46860 18680 46888 18720
rect 41984 18652 42104 18680
rect 42076 18624 42104 18652
rect 43180 18652 46888 18680
rect 38654 18612 38660 18624
rect 38580 18584 38660 18612
rect 38654 18572 38660 18584
rect 38712 18572 38718 18624
rect 38838 18572 38844 18624
rect 38896 18572 38902 18624
rect 39114 18572 39120 18624
rect 39172 18612 39178 18624
rect 41966 18612 41972 18624
rect 39172 18584 41972 18612
rect 39172 18572 39178 18584
rect 41966 18572 41972 18584
rect 42024 18572 42030 18624
rect 42058 18572 42064 18624
rect 42116 18572 42122 18624
rect 43180 18621 43208 18652
rect 46934 18640 46940 18692
rect 46992 18640 46998 18692
rect 47121 18683 47179 18689
rect 47121 18649 47133 18683
rect 47167 18649 47179 18683
rect 47121 18643 47179 18649
rect 43165 18615 43223 18621
rect 43165 18581 43177 18615
rect 43211 18581 43223 18615
rect 43165 18575 43223 18581
rect 43254 18572 43260 18624
rect 43312 18612 43318 18624
rect 43533 18615 43591 18621
rect 43533 18612 43545 18615
rect 43312 18584 43545 18612
rect 43312 18572 43318 18584
rect 43533 18581 43545 18584
rect 43579 18581 43591 18615
rect 43533 18575 43591 18581
rect 46014 18572 46020 18624
rect 46072 18612 46078 18624
rect 47136 18612 47164 18643
rect 47946 18640 47952 18692
rect 48004 18640 48010 18692
rect 48056 18680 48084 18720
rect 48593 18717 48605 18751
rect 48639 18748 48651 18751
rect 48774 18748 48780 18760
rect 48639 18720 48780 18748
rect 48639 18717 48651 18720
rect 48593 18711 48651 18717
rect 48774 18708 48780 18720
rect 48832 18708 48838 18760
rect 48961 18751 49019 18757
rect 48961 18717 48973 18751
rect 49007 18748 49019 18751
rect 54202 18748 54208 18760
rect 49007 18720 54208 18748
rect 49007 18717 49019 18720
rect 48961 18711 49019 18717
rect 54202 18708 54208 18720
rect 54260 18708 54266 18760
rect 55861 18751 55919 18757
rect 55861 18717 55873 18751
rect 55907 18748 55919 18751
rect 55968 18748 55996 18788
rect 58158 18776 58164 18828
rect 58216 18776 58222 18828
rect 55907 18720 55996 18748
rect 55907 18717 55919 18720
rect 55861 18711 55919 18717
rect 56042 18708 56048 18760
rect 56100 18757 56106 18760
rect 56100 18748 56108 18757
rect 56318 18748 56324 18760
rect 56100 18720 56324 18748
rect 56100 18711 56108 18720
rect 56100 18708 56106 18711
rect 56318 18708 56324 18720
rect 56376 18708 56382 18760
rect 56778 18708 56784 18760
rect 56836 18748 56842 18760
rect 56965 18751 57023 18757
rect 56965 18748 56977 18751
rect 56836 18720 56977 18748
rect 56836 18708 56842 18720
rect 56965 18717 56977 18720
rect 57011 18717 57023 18751
rect 57885 18751 57943 18757
rect 57885 18748 57897 18751
rect 56965 18711 57023 18717
rect 57052 18720 57897 18748
rect 55677 18683 55735 18689
rect 55677 18680 55689 18683
rect 48056 18652 55689 18680
rect 55677 18649 55689 18652
rect 55723 18649 55735 18683
rect 55677 18643 55735 18649
rect 55953 18683 56011 18689
rect 55953 18649 55965 18683
rect 55999 18680 56011 18683
rect 56594 18680 56600 18692
rect 55999 18652 56600 18680
rect 55999 18649 56011 18652
rect 55953 18643 56011 18649
rect 56594 18640 56600 18652
rect 56652 18640 56658 18692
rect 46072 18584 47164 18612
rect 46072 18572 46078 18584
rect 49510 18572 49516 18624
rect 49568 18612 49574 18624
rect 57052 18612 57080 18720
rect 57885 18717 57897 18720
rect 57931 18717 57943 18751
rect 57885 18711 57943 18717
rect 57241 18683 57299 18689
rect 57241 18649 57253 18683
rect 57287 18649 57299 18683
rect 57241 18643 57299 18649
rect 49568 18584 57080 18612
rect 57256 18612 57284 18643
rect 58986 18612 58992 18624
rect 57256 18584 58992 18612
rect 49568 18572 49574 18584
rect 58986 18572 58992 18584
rect 59044 18572 59050 18624
rect 1104 18522 58880 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 50294 18522
rect 50346 18470 50358 18522
rect 50410 18470 50422 18522
rect 50474 18470 50486 18522
rect 50538 18470 50550 18522
rect 50602 18470 58880 18522
rect 1104 18448 58880 18470
rect 20898 18368 20904 18420
rect 20956 18408 20962 18420
rect 29546 18408 29552 18420
rect 20956 18380 29552 18408
rect 20956 18368 20962 18380
rect 29546 18368 29552 18380
rect 29604 18368 29610 18420
rect 29638 18368 29644 18420
rect 29696 18368 29702 18420
rect 29748 18380 34560 18408
rect 20530 18300 20536 18352
rect 20588 18340 20594 18352
rect 29748 18340 29776 18380
rect 20588 18312 29776 18340
rect 34532 18340 34560 18380
rect 34606 18368 34612 18420
rect 34664 18408 34670 18420
rect 34885 18411 34943 18417
rect 34885 18408 34897 18411
rect 34664 18380 34897 18408
rect 34664 18368 34670 18380
rect 34885 18377 34897 18380
rect 34931 18377 34943 18411
rect 34885 18371 34943 18377
rect 34974 18368 34980 18420
rect 35032 18408 35038 18420
rect 36817 18411 36875 18417
rect 36817 18408 36829 18411
rect 35032 18380 36829 18408
rect 35032 18368 35038 18380
rect 36817 18377 36829 18380
rect 36863 18377 36875 18411
rect 39117 18411 39175 18417
rect 36817 18371 36875 18377
rect 37568 18380 39068 18408
rect 36081 18343 36139 18349
rect 34532 18312 36032 18340
rect 20588 18300 20594 18312
rect 1581 18275 1639 18281
rect 1581 18241 1593 18275
rect 1627 18272 1639 18275
rect 1627 18244 2452 18272
rect 1627 18241 1639 18244
rect 1581 18235 1639 18241
rect 934 18164 940 18216
rect 992 18204 998 18216
rect 1765 18207 1823 18213
rect 1765 18204 1777 18207
rect 992 18176 1777 18204
rect 992 18164 998 18176
rect 1765 18173 1777 18176
rect 1811 18173 1823 18207
rect 1765 18167 1823 18173
rect 2424 18145 2452 18244
rect 22278 18232 22284 18284
rect 22336 18272 22342 18284
rect 24213 18275 24271 18281
rect 24213 18272 24225 18275
rect 22336 18244 24225 18272
rect 22336 18232 22342 18244
rect 24213 18241 24225 18244
rect 24259 18241 24271 18275
rect 24213 18235 24271 18241
rect 24302 18232 24308 18284
rect 24360 18272 24366 18284
rect 25501 18275 25559 18281
rect 25501 18272 25513 18275
rect 24360 18244 25513 18272
rect 24360 18232 24366 18244
rect 25501 18241 25513 18244
rect 25547 18241 25559 18275
rect 25501 18235 25559 18241
rect 26326 18232 26332 18284
rect 26384 18272 26390 18284
rect 27890 18272 27896 18284
rect 26384 18244 27896 18272
rect 26384 18232 26390 18244
rect 27890 18232 27896 18244
rect 27948 18232 27954 18284
rect 28721 18275 28779 18281
rect 28721 18241 28733 18275
rect 28767 18272 28779 18275
rect 28994 18272 29000 18284
rect 28767 18244 29000 18272
rect 28767 18241 28779 18244
rect 28721 18235 28779 18241
rect 28994 18232 29000 18244
rect 29052 18232 29058 18284
rect 29086 18232 29092 18284
rect 29144 18272 29150 18284
rect 29457 18275 29515 18281
rect 29457 18272 29469 18275
rect 29144 18244 29469 18272
rect 29144 18232 29150 18244
rect 29457 18241 29469 18244
rect 29503 18241 29515 18275
rect 29457 18235 29515 18241
rect 29638 18232 29644 18284
rect 29696 18272 29702 18284
rect 30193 18275 30251 18281
rect 30193 18272 30205 18275
rect 29696 18244 30205 18272
rect 29696 18232 29702 18244
rect 30193 18241 30205 18244
rect 30239 18241 30251 18275
rect 30193 18235 30251 18241
rect 30374 18232 30380 18284
rect 30432 18232 30438 18284
rect 32398 18232 32404 18284
rect 32456 18232 32462 18284
rect 33137 18275 33195 18281
rect 33137 18241 33149 18275
rect 33183 18241 33195 18275
rect 33137 18235 33195 18241
rect 33873 18275 33931 18281
rect 33873 18241 33885 18275
rect 33919 18272 33931 18275
rect 34606 18272 34612 18284
rect 33919 18244 34612 18272
rect 33919 18241 33931 18244
rect 33873 18235 33931 18241
rect 24394 18164 24400 18216
rect 24452 18164 24458 18216
rect 24762 18164 24768 18216
rect 24820 18204 24826 18216
rect 25317 18207 25375 18213
rect 25317 18204 25329 18207
rect 24820 18176 25329 18204
rect 24820 18164 24826 18176
rect 25317 18173 25329 18176
rect 25363 18173 25375 18207
rect 25317 18167 25375 18173
rect 25685 18207 25743 18213
rect 25685 18173 25697 18207
rect 25731 18204 25743 18207
rect 26694 18204 26700 18216
rect 25731 18176 26700 18204
rect 25731 18173 25743 18176
rect 25685 18167 25743 18173
rect 26694 18164 26700 18176
rect 26752 18164 26758 18216
rect 33152 18204 33180 18235
rect 34606 18232 34612 18244
rect 34664 18232 34670 18284
rect 34698 18232 34704 18284
rect 34756 18232 34762 18284
rect 35526 18232 35532 18284
rect 35584 18272 35590 18284
rect 35897 18275 35955 18281
rect 35897 18272 35909 18275
rect 35584 18244 35909 18272
rect 35584 18232 35590 18244
rect 35897 18241 35909 18244
rect 35943 18241 35955 18275
rect 36004 18272 36032 18312
rect 36081 18309 36093 18343
rect 36127 18340 36139 18343
rect 36170 18340 36176 18352
rect 36127 18312 36176 18340
rect 36127 18309 36139 18312
rect 36081 18303 36139 18309
rect 36170 18300 36176 18312
rect 36228 18300 36234 18352
rect 37568 18340 37596 18380
rect 36556 18312 37596 18340
rect 36556 18272 36584 18312
rect 37642 18300 37648 18352
rect 37700 18340 37706 18352
rect 39040 18340 39068 18380
rect 39117 18377 39129 18411
rect 39163 18408 39175 18411
rect 39942 18408 39948 18420
rect 39163 18380 39948 18408
rect 39163 18377 39175 18380
rect 39117 18371 39175 18377
rect 39942 18368 39948 18380
rect 40000 18368 40006 18420
rect 40218 18408 40224 18420
rect 40052 18380 40224 18408
rect 40052 18340 40080 18380
rect 40218 18368 40224 18380
rect 40276 18368 40282 18420
rect 40313 18411 40371 18417
rect 40313 18377 40325 18411
rect 40359 18408 40371 18411
rect 41414 18408 41420 18420
rect 40359 18380 41420 18408
rect 40359 18377 40371 18380
rect 40313 18371 40371 18377
rect 41414 18368 41420 18380
rect 41472 18368 41478 18420
rect 41616 18380 42656 18408
rect 41616 18340 41644 18380
rect 37700 18312 38654 18340
rect 39040 18312 40080 18340
rect 40227 18312 41644 18340
rect 42628 18340 42656 18380
rect 42702 18368 42708 18420
rect 42760 18408 42766 18420
rect 42760 18380 44864 18408
rect 42760 18368 42766 18380
rect 44726 18340 44732 18352
rect 42628 18312 44732 18340
rect 37700 18300 37706 18312
rect 36004 18244 36584 18272
rect 36633 18275 36691 18281
rect 35897 18235 35955 18241
rect 36633 18241 36645 18275
rect 36679 18272 36691 18275
rect 37366 18272 37372 18284
rect 36679 18244 37372 18272
rect 36679 18241 36691 18244
rect 36633 18235 36691 18241
rect 37366 18232 37372 18244
rect 37424 18232 37430 18284
rect 37461 18275 37519 18281
rect 37461 18241 37473 18275
rect 37507 18241 37519 18275
rect 37461 18235 37519 18241
rect 35713 18207 35771 18213
rect 33152 18176 34100 18204
rect 34072 18145 34100 18176
rect 35713 18173 35725 18207
rect 35759 18204 35771 18207
rect 36814 18204 36820 18216
rect 35759 18176 36820 18204
rect 35759 18173 35771 18176
rect 35713 18167 35771 18173
rect 36814 18164 36820 18176
rect 36872 18164 36878 18216
rect 37476 18204 37504 18235
rect 37918 18232 37924 18284
rect 37976 18272 37982 18284
rect 38197 18275 38255 18281
rect 38197 18272 38209 18275
rect 37976 18244 38209 18272
rect 37976 18232 37982 18244
rect 38197 18241 38209 18244
rect 38243 18241 38255 18275
rect 38626 18272 38654 18312
rect 38933 18275 38991 18281
rect 38933 18272 38945 18275
rect 38626 18244 38945 18272
rect 38197 18235 38255 18241
rect 38933 18241 38945 18244
rect 38979 18272 38991 18275
rect 39114 18272 39120 18284
rect 38979 18244 39120 18272
rect 38979 18241 38991 18244
rect 38933 18235 38991 18241
rect 39114 18232 39120 18244
rect 39172 18232 39178 18284
rect 40135 18275 40193 18281
rect 40135 18241 40147 18275
rect 40181 18261 40193 18275
rect 40227 18261 40255 18312
rect 44726 18300 44732 18312
rect 44784 18300 44790 18352
rect 44836 18340 44864 18380
rect 45002 18368 45008 18420
rect 45060 18368 45066 18420
rect 45370 18368 45376 18420
rect 45428 18368 45434 18420
rect 46934 18368 46940 18420
rect 46992 18408 46998 18420
rect 47670 18408 47676 18420
rect 46992 18380 47676 18408
rect 46992 18368 46998 18380
rect 47670 18368 47676 18380
rect 47728 18368 47734 18420
rect 48958 18408 48964 18420
rect 48056 18380 48964 18408
rect 48056 18340 48084 18380
rect 48958 18368 48964 18380
rect 49016 18368 49022 18420
rect 50893 18411 50951 18417
rect 50893 18377 50905 18411
rect 50939 18408 50951 18411
rect 51074 18408 51080 18420
rect 50939 18380 51080 18408
rect 50939 18377 50951 18380
rect 50893 18371 50951 18377
rect 51074 18368 51080 18380
rect 51132 18368 51138 18420
rect 55858 18368 55864 18420
rect 55916 18368 55922 18420
rect 56042 18368 56048 18420
rect 56100 18408 56106 18420
rect 56100 18380 57100 18408
rect 56100 18368 56106 18380
rect 50982 18340 50988 18352
rect 44836 18312 48084 18340
rect 48792 18312 50988 18340
rect 40181 18241 40255 18261
rect 40135 18235 40255 18241
rect 40865 18275 40923 18281
rect 40865 18241 40877 18275
rect 40911 18272 40923 18275
rect 41598 18272 41604 18284
rect 40911 18244 41604 18272
rect 40911 18241 40923 18244
rect 40865 18235 40923 18241
rect 40144 18233 40255 18235
rect 41598 18232 41604 18244
rect 41656 18232 41662 18284
rect 41693 18275 41751 18281
rect 41693 18241 41705 18275
rect 41739 18241 41751 18275
rect 41693 18235 41751 18241
rect 40310 18204 40316 18216
rect 37476 18176 40316 18204
rect 40310 18164 40316 18176
rect 40368 18164 40374 18216
rect 41708 18204 41736 18235
rect 41874 18232 41880 18284
rect 41932 18232 41938 18284
rect 43990 18232 43996 18284
rect 44048 18232 44054 18284
rect 44361 18275 44419 18281
rect 44361 18241 44373 18275
rect 44407 18272 44419 18275
rect 44910 18272 44916 18284
rect 44407 18244 44916 18272
rect 44407 18241 44419 18244
rect 44361 18235 44419 18241
rect 44910 18232 44916 18244
rect 44968 18232 44974 18284
rect 48409 18275 48467 18281
rect 48409 18241 48421 18275
rect 48455 18272 48467 18275
rect 48682 18272 48688 18284
rect 48455 18244 48688 18272
rect 48455 18241 48467 18244
rect 48409 18235 48467 18241
rect 48682 18232 48688 18244
rect 48740 18232 48746 18284
rect 48792 18281 48820 18312
rect 50982 18300 50988 18312
rect 51040 18300 51046 18352
rect 52270 18300 52276 18352
rect 52328 18340 52334 18352
rect 56410 18340 56416 18352
rect 52328 18312 56416 18340
rect 52328 18300 52334 18312
rect 48777 18275 48835 18281
rect 48777 18241 48789 18275
rect 48823 18241 48835 18275
rect 48777 18235 48835 18241
rect 48866 18232 48872 18284
rect 48924 18272 48930 18284
rect 48961 18275 49019 18281
rect 48961 18272 48973 18275
rect 48924 18244 48973 18272
rect 48924 18232 48930 18244
rect 48961 18241 48973 18244
rect 49007 18272 49019 18275
rect 49050 18272 49056 18284
rect 49007 18244 49056 18272
rect 49007 18241 49019 18244
rect 48961 18235 49019 18241
rect 49050 18232 49056 18244
rect 49108 18232 49114 18284
rect 49418 18232 49424 18284
rect 49476 18232 49482 18284
rect 55674 18232 55680 18284
rect 55732 18262 55738 18284
rect 55968 18281 55996 18312
rect 56410 18300 56416 18312
rect 56468 18300 56474 18352
rect 56686 18300 56692 18352
rect 56744 18300 56750 18352
rect 56962 18300 56968 18352
rect 57020 18300 57026 18352
rect 57072 18303 57100 18380
rect 57062 18297 57120 18303
rect 55769 18275 55827 18281
rect 55769 18262 55781 18275
rect 55732 18241 55781 18262
rect 55815 18241 55827 18275
rect 55732 18235 55827 18241
rect 55953 18275 56011 18281
rect 55953 18241 55965 18275
rect 55999 18241 56011 18275
rect 56873 18275 56931 18281
rect 56873 18272 56885 18275
rect 55953 18235 56011 18241
rect 56040 18244 56885 18272
rect 55732 18234 55812 18235
rect 55732 18232 55738 18234
rect 41966 18204 41972 18216
rect 41708 18176 41972 18204
rect 41966 18164 41972 18176
rect 42024 18204 42030 18216
rect 42610 18204 42616 18216
rect 42024 18176 42616 18204
rect 42024 18164 42030 18176
rect 42610 18164 42616 18176
rect 42668 18164 42674 18216
rect 43070 18164 43076 18216
rect 43128 18204 43134 18216
rect 43898 18204 43904 18216
rect 43128 18176 43904 18204
rect 43128 18164 43134 18176
rect 43898 18164 43904 18176
rect 43956 18164 43962 18216
rect 44453 18207 44511 18213
rect 44453 18173 44465 18207
rect 44499 18204 44511 18207
rect 45094 18204 45100 18216
rect 44499 18176 45100 18204
rect 44499 18173 44511 18176
rect 44453 18167 44511 18173
rect 45094 18164 45100 18176
rect 45152 18164 45158 18216
rect 45462 18164 45468 18216
rect 45520 18164 45526 18216
rect 45649 18207 45707 18213
rect 45649 18173 45661 18207
rect 45695 18204 45707 18207
rect 46934 18204 46940 18216
rect 45695 18176 46940 18204
rect 45695 18173 45707 18176
rect 45649 18167 45707 18173
rect 46934 18164 46940 18176
rect 46992 18164 46998 18216
rect 48498 18164 48504 18216
rect 48556 18164 48562 18216
rect 56040 18204 56068 18244
rect 56873 18241 56885 18244
rect 56919 18241 56931 18275
rect 57062 18263 57074 18297
rect 57108 18263 57120 18297
rect 57062 18257 57120 18263
rect 58069 18275 58127 18281
rect 56873 18235 56931 18241
rect 58069 18241 58081 18275
rect 58115 18241 58127 18275
rect 58069 18235 58127 18241
rect 58084 18204 58112 18235
rect 55324 18176 56068 18204
rect 56096 18176 58112 18204
rect 2409 18139 2467 18145
rect 2409 18105 2421 18139
rect 2455 18136 2467 18139
rect 34057 18139 34115 18145
rect 2455 18108 34008 18136
rect 2455 18105 2467 18108
rect 2409 18099 2467 18105
rect 18598 18028 18604 18080
rect 18656 18068 18662 18080
rect 24118 18068 24124 18080
rect 18656 18040 24124 18068
rect 18656 18028 18662 18040
rect 24118 18028 24124 18040
rect 24176 18068 24182 18080
rect 24762 18068 24768 18080
rect 24176 18040 24768 18068
rect 24176 18028 24182 18040
rect 24762 18028 24768 18040
rect 24820 18068 24826 18080
rect 24949 18071 25007 18077
rect 24949 18068 24961 18071
rect 24820 18040 24961 18068
rect 24820 18028 24826 18040
rect 24949 18037 24961 18040
rect 24995 18037 25007 18071
rect 24949 18031 25007 18037
rect 26329 18071 26387 18077
rect 26329 18037 26341 18071
rect 26375 18068 26387 18071
rect 26878 18068 26884 18080
rect 26375 18040 26884 18068
rect 26375 18037 26387 18040
rect 26329 18031 26387 18037
rect 26878 18028 26884 18040
rect 26936 18028 26942 18080
rect 28905 18071 28963 18077
rect 28905 18037 28917 18071
rect 28951 18068 28963 18071
rect 30098 18068 30104 18080
rect 28951 18040 30104 18068
rect 28951 18037 28963 18040
rect 28905 18031 28963 18037
rect 30098 18028 30104 18040
rect 30156 18028 30162 18080
rect 30193 18071 30251 18077
rect 30193 18037 30205 18071
rect 30239 18068 30251 18071
rect 30650 18068 30656 18080
rect 30239 18040 30656 18068
rect 30239 18037 30251 18040
rect 30193 18031 30251 18037
rect 30650 18028 30656 18040
rect 30708 18028 30714 18080
rect 32582 18028 32588 18080
rect 32640 18028 32646 18080
rect 32674 18028 32680 18080
rect 32732 18068 32738 18080
rect 33321 18071 33379 18077
rect 33321 18068 33333 18071
rect 32732 18040 33333 18068
rect 32732 18028 32738 18040
rect 33321 18037 33333 18040
rect 33367 18037 33379 18071
rect 33980 18068 34008 18108
rect 34057 18105 34069 18139
rect 34103 18105 34115 18139
rect 34057 18099 34115 18105
rect 37458 18096 37464 18148
rect 37516 18136 37522 18148
rect 38381 18139 38439 18145
rect 38381 18136 38393 18139
rect 37516 18108 38393 18136
rect 37516 18096 37522 18108
rect 38381 18105 38393 18108
rect 38427 18105 38439 18139
rect 38381 18099 38439 18105
rect 40126 18096 40132 18148
rect 40184 18136 40190 18148
rect 41049 18139 41107 18145
rect 41049 18136 41061 18139
rect 40184 18108 41061 18136
rect 40184 18096 40190 18108
rect 41049 18105 41061 18108
rect 41095 18105 41107 18139
rect 41049 18099 41107 18105
rect 41690 18096 41696 18148
rect 41748 18136 41754 18148
rect 54386 18136 54392 18148
rect 41748 18108 54392 18136
rect 41748 18096 41754 18108
rect 54386 18096 54392 18108
rect 54444 18096 54450 18148
rect 36630 18068 36636 18080
rect 33980 18040 36636 18068
rect 33321 18031 33379 18037
rect 36630 18028 36636 18040
rect 36688 18028 36694 18080
rect 37550 18028 37556 18080
rect 37608 18068 37614 18080
rect 37645 18071 37703 18077
rect 37645 18068 37657 18071
rect 37608 18040 37657 18068
rect 37608 18028 37614 18040
rect 37645 18037 37657 18040
rect 37691 18037 37703 18071
rect 37645 18031 37703 18037
rect 37826 18028 37832 18080
rect 37884 18068 37890 18080
rect 40862 18068 40868 18080
rect 37884 18040 40868 18068
rect 37884 18028 37890 18040
rect 40862 18028 40868 18040
rect 40920 18028 40926 18080
rect 42061 18071 42119 18077
rect 42061 18037 42073 18071
rect 42107 18068 42119 18071
rect 43070 18068 43076 18080
rect 42107 18040 43076 18068
rect 42107 18037 42119 18040
rect 42061 18031 42119 18037
rect 43070 18028 43076 18040
rect 43128 18028 43134 18080
rect 43438 18028 43444 18080
rect 43496 18028 43502 18080
rect 46474 18028 46480 18080
rect 46532 18068 46538 18080
rect 47854 18068 47860 18080
rect 46532 18040 47860 18068
rect 46532 18028 46538 18040
rect 47854 18028 47860 18040
rect 47912 18028 47918 18080
rect 48314 18028 48320 18080
rect 48372 18068 48378 18080
rect 54938 18068 54944 18080
rect 48372 18040 54944 18068
rect 48372 18028 48378 18040
rect 54938 18028 54944 18040
rect 54996 18068 55002 18080
rect 55324 18068 55352 18176
rect 55398 18096 55404 18148
rect 55456 18136 55462 18148
rect 56096 18136 56124 18176
rect 55456 18108 56124 18136
rect 55456 18096 55462 18108
rect 56410 18096 56416 18148
rect 56468 18136 56474 18148
rect 58253 18139 58311 18145
rect 58253 18136 58265 18139
rect 56468 18108 58265 18136
rect 56468 18096 56474 18108
rect 58253 18105 58265 18108
rect 58299 18105 58311 18139
rect 58253 18099 58311 18105
rect 54996 18040 55352 18068
rect 54996 18028 55002 18040
rect 56686 18028 56692 18080
rect 56744 18028 56750 18080
rect 1104 17978 58880 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 58880 17978
rect 1104 17904 58880 17926
rect 2409 17867 2467 17873
rect 2409 17833 2421 17867
rect 2455 17864 2467 17867
rect 35618 17864 35624 17876
rect 2455 17836 35624 17864
rect 2455 17833 2467 17836
rect 2409 17827 2467 17833
rect 1581 17663 1639 17669
rect 1581 17629 1593 17663
rect 1627 17660 1639 17663
rect 2424 17660 2452 17827
rect 35618 17824 35624 17836
rect 35676 17824 35682 17876
rect 36814 17824 36820 17876
rect 36872 17864 36878 17876
rect 38657 17867 38715 17873
rect 38657 17864 38669 17867
rect 36872 17836 38669 17864
rect 36872 17824 36878 17836
rect 38657 17833 38669 17836
rect 38703 17833 38715 17867
rect 38657 17827 38715 17833
rect 39022 17824 39028 17876
rect 39080 17864 39086 17876
rect 39393 17867 39451 17873
rect 39393 17864 39405 17867
rect 39080 17836 39405 17864
rect 39080 17824 39086 17836
rect 39393 17833 39405 17836
rect 39439 17833 39451 17867
rect 39393 17827 39451 17833
rect 41874 17824 41880 17876
rect 41932 17864 41938 17876
rect 43625 17867 43683 17873
rect 43625 17864 43637 17867
rect 41932 17836 43637 17864
rect 41932 17824 41938 17836
rect 43625 17833 43637 17836
rect 43671 17833 43683 17867
rect 43625 17827 43683 17833
rect 43714 17824 43720 17876
rect 43772 17864 43778 17876
rect 44174 17864 44180 17876
rect 43772 17836 44180 17864
rect 43772 17824 43778 17836
rect 44174 17824 44180 17836
rect 44232 17824 44238 17876
rect 44358 17824 44364 17876
rect 44416 17864 44422 17876
rect 45554 17864 45560 17876
rect 44416 17836 45560 17864
rect 44416 17824 44422 17836
rect 45554 17824 45560 17836
rect 45612 17864 45618 17876
rect 46293 17867 46351 17873
rect 46293 17864 46305 17867
rect 45612 17836 46305 17864
rect 45612 17824 45618 17836
rect 46293 17833 46305 17836
rect 46339 17833 46351 17867
rect 46293 17827 46351 17833
rect 47762 17824 47768 17876
rect 47820 17864 47826 17876
rect 49053 17867 49111 17873
rect 49053 17864 49065 17867
rect 47820 17836 49065 17864
rect 47820 17824 47826 17836
rect 49053 17833 49065 17836
rect 49099 17833 49111 17867
rect 49053 17827 49111 17833
rect 56870 17824 56876 17876
rect 56928 17864 56934 17876
rect 58253 17867 58311 17873
rect 58253 17864 58265 17867
rect 56928 17836 58265 17864
rect 56928 17824 56934 17836
rect 58253 17833 58265 17836
rect 58299 17833 58311 17867
rect 58253 17827 58311 17833
rect 24670 17756 24676 17808
rect 24728 17756 24734 17808
rect 27522 17796 27528 17808
rect 25792 17768 27528 17796
rect 22738 17688 22744 17740
rect 22796 17728 22802 17740
rect 25792 17728 25820 17768
rect 27522 17756 27528 17768
rect 27580 17756 27586 17808
rect 28994 17756 29000 17808
rect 29052 17796 29058 17808
rect 29917 17799 29975 17805
rect 29917 17796 29929 17799
rect 29052 17768 29929 17796
rect 29052 17756 29058 17768
rect 29917 17765 29929 17768
rect 29963 17765 29975 17799
rect 29917 17759 29975 17765
rect 34241 17799 34299 17805
rect 34241 17765 34253 17799
rect 34287 17796 34299 17799
rect 36170 17796 36176 17808
rect 34287 17768 36176 17796
rect 34287 17765 34299 17768
rect 34241 17759 34299 17765
rect 36170 17756 36176 17768
rect 36228 17796 36234 17808
rect 36228 17768 36860 17796
rect 36228 17756 36234 17768
rect 28258 17728 28264 17740
rect 22796 17700 25820 17728
rect 22796 17688 22802 17700
rect 1627 17632 2452 17660
rect 17865 17663 17923 17669
rect 1627 17629 1639 17632
rect 1581 17623 1639 17629
rect 17865 17629 17877 17663
rect 17911 17660 17923 17663
rect 17954 17660 17960 17672
rect 17911 17632 17960 17660
rect 17911 17629 17923 17632
rect 17865 17623 17923 17629
rect 17954 17620 17960 17632
rect 18012 17620 18018 17672
rect 18049 17663 18107 17669
rect 18049 17629 18061 17663
rect 18095 17660 18107 17663
rect 18414 17660 18420 17672
rect 18095 17632 18420 17660
rect 18095 17629 18107 17632
rect 18049 17623 18107 17629
rect 18414 17620 18420 17632
rect 18472 17620 18478 17672
rect 20533 17663 20591 17669
rect 20533 17629 20545 17663
rect 20579 17660 20591 17663
rect 21174 17660 21180 17672
rect 20579 17632 21180 17660
rect 20579 17629 20591 17632
rect 20533 17623 20591 17629
rect 21174 17620 21180 17632
rect 21232 17620 21238 17672
rect 21269 17663 21327 17669
rect 21269 17629 21281 17663
rect 21315 17629 21327 17663
rect 21269 17623 21327 17629
rect 21453 17663 21511 17669
rect 21453 17629 21465 17663
rect 21499 17660 21511 17663
rect 22646 17660 22652 17672
rect 21499 17632 22652 17660
rect 21499 17629 21511 17632
rect 21453 17623 21511 17629
rect 934 17552 940 17604
rect 992 17592 998 17604
rect 1857 17595 1915 17601
rect 1857 17592 1869 17595
rect 992 17564 1869 17592
rect 992 17552 998 17564
rect 1857 17561 1869 17564
rect 1903 17561 1915 17595
rect 21284 17592 21312 17623
rect 22646 17620 22652 17632
rect 22704 17620 22710 17672
rect 24578 17620 24584 17672
rect 24636 17620 24642 17672
rect 24762 17620 24768 17672
rect 24820 17660 24826 17672
rect 25792 17669 25820 17700
rect 25976 17700 28264 17728
rect 25976 17669 26004 17700
rect 28258 17688 28264 17700
rect 28316 17688 28322 17740
rect 28350 17688 28356 17740
rect 28408 17728 28414 17740
rect 28445 17731 28503 17737
rect 28445 17728 28457 17731
rect 28408 17700 28457 17728
rect 28408 17688 28414 17700
rect 28445 17697 28457 17700
rect 28491 17697 28503 17731
rect 28445 17691 28503 17697
rect 28905 17731 28963 17737
rect 28905 17697 28917 17731
rect 28951 17697 28963 17731
rect 32674 17728 32680 17740
rect 28905 17691 28963 17697
rect 31496 17700 32680 17728
rect 24857 17663 24915 17669
rect 24857 17660 24869 17663
rect 24820 17632 24869 17660
rect 24820 17620 24826 17632
rect 24857 17629 24869 17632
rect 24903 17629 24915 17663
rect 24857 17623 24915 17629
rect 25777 17663 25835 17669
rect 25777 17629 25789 17663
rect 25823 17629 25835 17663
rect 25777 17623 25835 17629
rect 25961 17663 26019 17669
rect 25961 17629 25973 17663
rect 26007 17629 26019 17663
rect 25961 17623 26019 17629
rect 26142 17620 26148 17672
rect 26200 17620 26206 17672
rect 26234 17620 26240 17672
rect 26292 17660 26298 17672
rect 26789 17663 26847 17669
rect 26789 17660 26801 17663
rect 26292 17632 26801 17660
rect 26292 17620 26298 17632
rect 26789 17629 26801 17632
rect 26835 17629 26847 17663
rect 26789 17623 26847 17629
rect 28534 17620 28540 17672
rect 28592 17620 28598 17672
rect 28920 17660 28948 17691
rect 29733 17663 29791 17669
rect 29733 17660 29745 17663
rect 28920 17632 29745 17660
rect 29733 17629 29745 17632
rect 29779 17629 29791 17663
rect 29733 17623 29791 17629
rect 30098 17620 30104 17672
rect 30156 17660 30162 17672
rect 31496 17669 31524 17700
rect 32674 17688 32680 17700
rect 32732 17688 32738 17740
rect 35989 17731 36047 17737
rect 35989 17697 36001 17731
rect 36035 17728 36047 17731
rect 36078 17728 36084 17740
rect 36035 17700 36084 17728
rect 36035 17697 36047 17700
rect 35989 17691 36047 17697
rect 36078 17688 36084 17700
rect 36136 17688 36142 17740
rect 36262 17688 36268 17740
rect 36320 17688 36326 17740
rect 36832 17728 36860 17768
rect 36906 17756 36912 17808
rect 36964 17756 36970 17808
rect 37108 17768 38516 17796
rect 37108 17728 37136 17768
rect 36832 17700 37136 17728
rect 37182 17688 37188 17740
rect 37240 17728 37246 17740
rect 38488 17728 38516 17768
rect 38562 17756 38568 17808
rect 38620 17796 38626 17808
rect 41966 17796 41972 17808
rect 38620 17768 41972 17796
rect 38620 17756 38626 17768
rect 41966 17756 41972 17768
rect 42024 17756 42030 17808
rect 43898 17756 43904 17808
rect 43956 17796 43962 17808
rect 43956 17768 47992 17796
rect 43956 17756 43962 17768
rect 37240 17700 38424 17728
rect 38488 17700 40356 17728
rect 37240 17688 37246 17700
rect 30469 17663 30527 17669
rect 30469 17660 30481 17663
rect 30156 17632 30481 17660
rect 30156 17620 30162 17632
rect 30469 17629 30481 17632
rect 30515 17629 30527 17663
rect 30469 17623 30527 17629
rect 31481 17663 31539 17669
rect 31481 17629 31493 17663
rect 31527 17629 31539 17663
rect 31481 17623 31539 17629
rect 31665 17663 31723 17669
rect 31665 17629 31677 17663
rect 31711 17660 31723 17663
rect 31754 17660 31760 17672
rect 31711 17632 31760 17660
rect 31711 17629 31723 17632
rect 31665 17623 31723 17629
rect 31754 17620 31760 17632
rect 31812 17620 31818 17672
rect 32122 17620 32128 17672
rect 32180 17620 32186 17672
rect 32861 17663 32919 17669
rect 32861 17629 32873 17663
rect 32907 17660 32919 17663
rect 32950 17660 32956 17672
rect 32907 17632 32956 17660
rect 32907 17629 32919 17632
rect 32861 17623 32919 17629
rect 32950 17620 32956 17632
rect 33008 17620 33014 17672
rect 34790 17620 34796 17672
rect 34848 17660 34854 17672
rect 34885 17663 34943 17669
rect 34885 17660 34897 17663
rect 34848 17632 34897 17660
rect 34848 17620 34854 17632
rect 34885 17629 34897 17632
rect 34931 17629 34943 17663
rect 34885 17623 34943 17629
rect 35897 17663 35955 17669
rect 35897 17629 35909 17663
rect 35943 17660 35955 17663
rect 36538 17660 36544 17672
rect 35943 17632 36544 17660
rect 35943 17629 35955 17632
rect 35897 17623 35955 17629
rect 36538 17620 36544 17632
rect 36596 17620 36602 17672
rect 36725 17663 36783 17669
rect 36725 17629 36737 17663
rect 36771 17629 36783 17663
rect 36725 17623 36783 17629
rect 21634 17592 21640 17604
rect 21284 17564 21640 17592
rect 1857 17555 1915 17561
rect 21634 17552 21640 17564
rect 21692 17552 21698 17604
rect 23750 17552 23756 17604
rect 23808 17592 23814 17604
rect 24210 17592 24216 17604
rect 23808 17564 24216 17592
rect 23808 17552 23814 17564
rect 24210 17552 24216 17564
rect 24268 17592 24274 17604
rect 26053 17595 26111 17601
rect 24268 17564 26004 17592
rect 24268 17552 24274 17564
rect 18049 17527 18107 17533
rect 18049 17493 18061 17527
rect 18095 17524 18107 17527
rect 18322 17524 18328 17536
rect 18095 17496 18328 17524
rect 18095 17493 18107 17496
rect 18049 17487 18107 17493
rect 18322 17484 18328 17496
rect 18380 17484 18386 17536
rect 20346 17484 20352 17536
rect 20404 17524 20410 17536
rect 20717 17527 20775 17533
rect 20717 17524 20729 17527
rect 20404 17496 20729 17524
rect 20404 17484 20410 17496
rect 20717 17493 20729 17496
rect 20763 17493 20775 17527
rect 20717 17487 20775 17493
rect 21358 17484 21364 17536
rect 21416 17484 21422 17536
rect 24026 17484 24032 17536
rect 24084 17524 24090 17536
rect 24762 17524 24768 17536
rect 24084 17496 24768 17524
rect 24084 17484 24090 17496
rect 24762 17484 24768 17496
rect 24820 17484 24826 17536
rect 25041 17527 25099 17533
rect 25041 17493 25053 17527
rect 25087 17524 25099 17527
rect 25866 17524 25872 17536
rect 25087 17496 25872 17524
rect 25087 17493 25099 17496
rect 25041 17487 25099 17493
rect 25866 17484 25872 17496
rect 25924 17484 25930 17536
rect 25976 17524 26004 17564
rect 26053 17561 26065 17595
rect 26099 17592 26111 17595
rect 26602 17592 26608 17604
rect 26099 17564 26608 17592
rect 26099 17561 26111 17564
rect 26053 17555 26111 17561
rect 26602 17552 26608 17564
rect 26660 17592 26666 17604
rect 26881 17595 26939 17601
rect 26881 17592 26893 17595
rect 26660 17564 26893 17592
rect 26660 17552 26666 17564
rect 26881 17561 26893 17564
rect 26927 17561 26939 17595
rect 26881 17555 26939 17561
rect 33128 17595 33186 17601
rect 33128 17561 33140 17595
rect 33174 17592 33186 17595
rect 33174 17564 35112 17592
rect 33174 17561 33186 17564
rect 33128 17555 33186 17561
rect 26234 17524 26240 17536
rect 25976 17496 26240 17524
rect 26234 17484 26240 17496
rect 26292 17484 26298 17536
rect 26329 17527 26387 17533
rect 26329 17493 26341 17527
rect 26375 17524 26387 17527
rect 26510 17524 26516 17536
rect 26375 17496 26516 17524
rect 26375 17493 26387 17496
rect 26329 17487 26387 17493
rect 26510 17484 26516 17496
rect 26568 17484 26574 17536
rect 30006 17484 30012 17536
rect 30064 17524 30070 17536
rect 30653 17527 30711 17533
rect 30653 17524 30665 17527
rect 30064 17496 30665 17524
rect 30064 17484 30070 17496
rect 30653 17493 30665 17496
rect 30699 17493 30711 17527
rect 30653 17487 30711 17493
rect 31570 17484 31576 17536
rect 31628 17484 31634 17536
rect 32306 17484 32312 17536
rect 32364 17484 32370 17536
rect 35084 17533 35112 17564
rect 35069 17527 35127 17533
rect 35069 17493 35081 17527
rect 35115 17493 35127 17527
rect 36740 17524 36768 17623
rect 37366 17620 37372 17672
rect 37424 17660 37430 17672
rect 37461 17663 37519 17669
rect 37461 17660 37473 17663
rect 37424 17632 37473 17660
rect 37424 17620 37430 17632
rect 37461 17629 37473 17632
rect 37507 17629 37519 17663
rect 37461 17623 37519 17629
rect 38396 17592 38424 17700
rect 38470 17620 38476 17672
rect 38528 17620 38534 17672
rect 39209 17663 39267 17669
rect 39209 17629 39221 17663
rect 39255 17629 39267 17663
rect 39209 17623 39267 17629
rect 40129 17663 40187 17669
rect 40129 17629 40141 17663
rect 40175 17629 40187 17663
rect 40129 17623 40187 17629
rect 39224 17592 39252 17623
rect 39666 17592 39672 17604
rect 38396 17564 39672 17592
rect 39666 17552 39672 17564
rect 39724 17552 39730 17604
rect 40144 17592 40172 17623
rect 40218 17620 40224 17672
rect 40276 17620 40282 17672
rect 40328 17660 40356 17700
rect 40402 17688 40408 17740
rect 40460 17688 40466 17740
rect 40494 17688 40500 17740
rect 40552 17728 40558 17740
rect 41322 17728 41328 17740
rect 40552 17700 41328 17728
rect 40552 17688 40558 17700
rect 41322 17688 41328 17700
rect 41380 17728 41386 17740
rect 41380 17700 42380 17728
rect 41380 17688 41386 17700
rect 41049 17663 41107 17669
rect 41049 17660 41061 17663
rect 40328 17632 41061 17660
rect 41049 17629 41061 17632
rect 41095 17660 41107 17663
rect 41874 17660 41880 17672
rect 41095 17632 41880 17660
rect 41095 17629 41107 17632
rect 41049 17623 41107 17629
rect 41874 17620 41880 17632
rect 41932 17620 41938 17672
rect 42242 17620 42248 17672
rect 42300 17620 42306 17672
rect 42352 17660 42380 17700
rect 44174 17688 44180 17740
rect 44232 17728 44238 17740
rect 45462 17728 45468 17740
rect 44232 17700 45468 17728
rect 44232 17688 44238 17700
rect 45462 17688 45468 17700
rect 45520 17728 45526 17740
rect 47964 17737 47992 17768
rect 55766 17756 55772 17808
rect 55824 17796 55830 17808
rect 55824 17768 56732 17796
rect 55824 17756 55830 17768
rect 47397 17731 47455 17737
rect 47397 17728 47409 17731
rect 45520 17700 47409 17728
rect 45520 17688 45526 17700
rect 47397 17697 47409 17700
rect 47443 17697 47455 17731
rect 47397 17691 47455 17697
rect 47949 17731 48007 17737
rect 47949 17697 47961 17731
rect 47995 17697 48007 17731
rect 47949 17691 48007 17697
rect 48958 17688 48964 17740
rect 49016 17728 49022 17740
rect 49016 17700 49280 17728
rect 49016 17688 49022 17700
rect 49252 17672 49280 17700
rect 51074 17688 51080 17740
rect 51132 17728 51138 17740
rect 56704 17728 56732 17768
rect 56873 17731 56931 17737
rect 56873 17728 56885 17731
rect 51132 17700 56548 17728
rect 56704 17700 56885 17728
rect 51132 17688 51138 17700
rect 44082 17660 44088 17672
rect 42352 17632 44088 17660
rect 44082 17620 44088 17632
rect 44140 17660 44146 17672
rect 44269 17663 44327 17669
rect 44269 17660 44281 17663
rect 44140 17632 44281 17660
rect 44140 17620 44146 17632
rect 44269 17629 44281 17632
rect 44315 17629 44327 17663
rect 44269 17623 44327 17629
rect 44450 17620 44456 17672
rect 44508 17660 44514 17672
rect 44637 17663 44695 17669
rect 44637 17660 44649 17663
rect 44508 17632 44649 17660
rect 44508 17620 44514 17632
rect 44637 17629 44649 17632
rect 44683 17629 44695 17663
rect 44637 17623 44695 17629
rect 45646 17620 45652 17672
rect 45704 17660 45710 17672
rect 46109 17663 46167 17669
rect 46109 17660 46121 17663
rect 45704 17632 46121 17660
rect 45704 17620 45710 17632
rect 46109 17629 46121 17632
rect 46155 17629 46167 17663
rect 46109 17623 46167 17629
rect 47578 17620 47584 17672
rect 47636 17660 47642 17672
rect 48041 17663 48099 17669
rect 48041 17660 48053 17663
rect 47636 17632 48053 17660
rect 47636 17620 47642 17632
rect 48041 17629 48053 17632
rect 48087 17629 48099 17663
rect 48041 17623 48099 17629
rect 48406 17620 48412 17672
rect 48464 17620 48470 17672
rect 48593 17663 48651 17669
rect 48593 17629 48605 17663
rect 48639 17660 48651 17663
rect 48866 17660 48872 17672
rect 48639 17632 48872 17660
rect 48639 17629 48651 17632
rect 48593 17623 48651 17629
rect 48866 17620 48872 17632
rect 48924 17620 48930 17672
rect 49050 17620 49056 17672
rect 49108 17620 49114 17672
rect 49234 17620 49240 17672
rect 49292 17620 49298 17672
rect 51718 17620 51724 17672
rect 51776 17660 51782 17672
rect 51905 17663 51963 17669
rect 51905 17660 51917 17663
rect 51776 17632 51917 17660
rect 51776 17620 51782 17632
rect 51905 17629 51917 17632
rect 51951 17629 51963 17663
rect 51905 17623 51963 17629
rect 51994 17620 52000 17672
rect 52052 17660 52058 17672
rect 52089 17663 52147 17669
rect 52089 17660 52101 17663
rect 52052 17632 52101 17660
rect 52052 17620 52058 17632
rect 52089 17629 52101 17632
rect 52135 17629 52147 17663
rect 52089 17623 52147 17629
rect 56229 17663 56287 17669
rect 56229 17629 56241 17663
rect 56275 17629 56287 17663
rect 56229 17623 56287 17629
rect 42512 17595 42570 17601
rect 40144 17564 41414 17592
rect 37645 17527 37703 17533
rect 37645 17524 37657 17527
rect 36740 17496 37657 17524
rect 35069 17487 35127 17493
rect 37645 17493 37657 17496
rect 37691 17493 37703 17527
rect 37645 17487 37703 17493
rect 38102 17484 38108 17536
rect 38160 17524 38166 17536
rect 40862 17524 40868 17536
rect 38160 17496 40868 17524
rect 38160 17484 38166 17496
rect 40862 17484 40868 17496
rect 40920 17484 40926 17536
rect 41230 17484 41236 17536
rect 41288 17484 41294 17536
rect 41386 17524 41414 17564
rect 42512 17561 42524 17595
rect 42558 17592 42570 17595
rect 42610 17592 42616 17604
rect 42558 17564 42616 17592
rect 42558 17561 42570 17564
rect 42512 17555 42570 17561
rect 42610 17552 42616 17564
rect 42668 17552 42674 17604
rect 45278 17552 45284 17604
rect 45336 17552 45342 17604
rect 42702 17524 42708 17536
rect 41386 17496 42708 17524
rect 42702 17484 42708 17496
rect 42760 17484 42766 17536
rect 51997 17527 52055 17533
rect 51997 17493 52009 17527
rect 52043 17524 52055 17527
rect 52086 17524 52092 17536
rect 52043 17496 52092 17524
rect 52043 17493 52055 17496
rect 51997 17487 52055 17493
rect 52086 17484 52092 17496
rect 52144 17484 52150 17536
rect 56244 17524 56272 17623
rect 56410 17620 56416 17672
rect 56468 17620 56474 17672
rect 56520 17660 56548 17700
rect 56873 17697 56885 17700
rect 56919 17697 56931 17731
rect 56873 17691 56931 17697
rect 59446 17660 59452 17672
rect 56520 17632 59452 17660
rect 59446 17620 59452 17632
rect 59504 17620 59510 17672
rect 56321 17595 56379 17601
rect 56321 17561 56333 17595
rect 56367 17592 56379 17595
rect 57118 17595 57176 17601
rect 57118 17592 57130 17595
rect 56367 17564 57130 17592
rect 56367 17561 56379 17564
rect 56321 17555 56379 17561
rect 57118 17561 57130 17564
rect 57164 17561 57176 17595
rect 57118 17555 57176 17561
rect 56686 17524 56692 17536
rect 56244 17496 56692 17524
rect 56686 17484 56692 17496
rect 56744 17484 56750 17536
rect 1104 17434 58880 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 50294 17434
rect 50346 17382 50358 17434
rect 50410 17382 50422 17434
rect 50474 17382 50486 17434
rect 50538 17382 50550 17434
rect 50602 17382 58880 17434
rect 1104 17360 58880 17382
rect 20349 17323 20407 17329
rect 20349 17289 20361 17323
rect 20395 17289 20407 17323
rect 20349 17283 20407 17289
rect 20993 17323 21051 17329
rect 20993 17289 21005 17323
rect 21039 17289 21051 17323
rect 20993 17283 21051 17289
rect 3510 17212 3516 17264
rect 3568 17252 3574 17264
rect 11698 17252 11704 17264
rect 3568 17224 11704 17252
rect 3568 17212 3574 17224
rect 11698 17212 11704 17224
rect 11756 17212 11762 17264
rect 1581 17187 1639 17193
rect 1581 17153 1593 17187
rect 1627 17184 1639 17187
rect 12342 17184 12348 17196
rect 1627 17156 12348 17184
rect 1627 17153 1639 17156
rect 1581 17147 1639 17153
rect 12342 17144 12348 17156
rect 12400 17144 12406 17196
rect 17586 17144 17592 17196
rect 17644 17144 17650 17196
rect 18322 17144 18328 17196
rect 18380 17144 18386 17196
rect 19981 17187 20039 17193
rect 19981 17153 19993 17187
rect 20027 17153 20039 17187
rect 20364 17184 20392 17283
rect 20809 17187 20867 17193
rect 20809 17184 20821 17187
rect 20364 17156 20821 17184
rect 19981 17147 20039 17153
rect 20809 17153 20821 17156
rect 20855 17153 20867 17187
rect 21008 17184 21036 17283
rect 21174 17280 21180 17332
rect 21232 17320 21238 17332
rect 22189 17323 22247 17329
rect 22189 17320 22201 17323
rect 21232 17292 22201 17320
rect 21232 17280 21238 17292
rect 22189 17289 22201 17292
rect 22235 17289 22247 17323
rect 22189 17283 22247 17289
rect 24118 17280 24124 17332
rect 24176 17280 24182 17332
rect 24762 17280 24768 17332
rect 24820 17320 24826 17332
rect 28626 17320 28632 17332
rect 24820 17292 28632 17320
rect 24820 17280 24826 17292
rect 28626 17280 28632 17292
rect 28684 17280 28690 17332
rect 31665 17323 31723 17329
rect 31665 17289 31677 17323
rect 31711 17320 31723 17323
rect 32122 17320 32128 17332
rect 31711 17292 32128 17320
rect 31711 17289 31723 17292
rect 31665 17283 31723 17289
rect 32122 17280 32128 17292
rect 32180 17280 32186 17332
rect 32398 17280 32404 17332
rect 32456 17320 32462 17332
rect 32493 17323 32551 17329
rect 32493 17320 32505 17323
rect 32456 17292 32505 17320
rect 32456 17280 32462 17292
rect 32493 17289 32505 17292
rect 32539 17289 32551 17323
rect 36078 17320 36084 17332
rect 32493 17283 32551 17289
rect 33612 17292 36084 17320
rect 23753 17255 23811 17261
rect 23753 17221 23765 17255
rect 23799 17252 23811 17255
rect 28988 17255 29046 17261
rect 23799 17224 24624 17252
rect 23799 17221 23811 17224
rect 23753 17215 23811 17221
rect 24136 17196 24164 17224
rect 24596 17196 24624 17224
rect 26344 17224 27752 17252
rect 22005 17187 22063 17193
rect 22005 17184 22017 17187
rect 21008 17156 22017 17184
rect 20809 17147 20867 17153
rect 22005 17153 22017 17156
rect 22051 17153 22063 17187
rect 22005 17147 22063 17153
rect 22925 17187 22983 17193
rect 22925 17153 22937 17187
rect 22971 17184 22983 17187
rect 23566 17184 23572 17196
rect 22971 17156 23572 17184
rect 22971 17153 22983 17156
rect 22925 17147 22983 17153
rect 934 17076 940 17128
rect 992 17116 998 17128
rect 1765 17119 1823 17125
rect 1765 17116 1777 17119
rect 992 17088 1777 17116
rect 992 17076 998 17088
rect 1765 17085 1777 17088
rect 1811 17085 1823 17119
rect 1765 17079 1823 17085
rect 19996 17048 20024 17147
rect 23566 17144 23572 17156
rect 23624 17144 23630 17196
rect 23937 17153 23995 17159
rect 23937 17128 23949 17153
rect 23983 17128 23995 17153
rect 24118 17144 24124 17196
rect 24176 17144 24182 17196
rect 24213 17187 24271 17193
rect 24213 17153 24225 17187
rect 24259 17184 24271 17187
rect 24302 17184 24308 17196
rect 24259 17156 24308 17184
rect 24259 17153 24271 17156
rect 24213 17147 24271 17153
rect 24302 17144 24308 17156
rect 24360 17144 24366 17196
rect 24578 17144 24584 17196
rect 24636 17184 24642 17196
rect 25133 17187 25191 17193
rect 25133 17184 25145 17187
rect 24636 17156 25145 17184
rect 24636 17144 24642 17156
rect 25133 17153 25145 17156
rect 25179 17153 25191 17187
rect 25133 17147 25191 17153
rect 25501 17187 25559 17193
rect 25501 17153 25513 17187
rect 25547 17153 25559 17187
rect 25501 17147 25559 17153
rect 20073 17119 20131 17125
rect 20073 17085 20085 17119
rect 20119 17116 20131 17119
rect 21358 17116 21364 17128
rect 20119 17088 21364 17116
rect 20119 17085 20131 17088
rect 20073 17079 20131 17085
rect 21358 17076 21364 17088
rect 21416 17076 21422 17128
rect 23014 17076 23020 17128
rect 23072 17116 23078 17128
rect 23072 17088 23888 17116
rect 23072 17076 23078 17088
rect 23658 17048 23664 17060
rect 19996 17020 23664 17048
rect 23658 17008 23664 17020
rect 23716 17008 23722 17060
rect 23860 17048 23888 17088
rect 23934 17076 23940 17128
rect 23992 17076 23998 17128
rect 25516 17116 25544 17147
rect 25682 17144 25688 17196
rect 25740 17184 25746 17196
rect 26344 17193 26372 17224
rect 26329 17187 26387 17193
rect 26329 17184 26341 17187
rect 25740 17156 26341 17184
rect 25740 17144 25746 17156
rect 26329 17153 26341 17156
rect 26375 17153 26387 17187
rect 26329 17147 26387 17153
rect 26602 17144 26608 17196
rect 26660 17144 26666 17196
rect 27341 17187 27399 17193
rect 27341 17153 27353 17187
rect 27387 17153 27399 17187
rect 27341 17147 27399 17153
rect 27433 17187 27491 17193
rect 27433 17153 27445 17187
rect 27479 17184 27491 17187
rect 27522 17184 27528 17196
rect 27479 17156 27528 17184
rect 27479 17153 27491 17156
rect 27433 17147 27491 17153
rect 24872 17088 25544 17116
rect 25593 17119 25651 17125
rect 24872 17048 24900 17088
rect 25593 17085 25605 17119
rect 25639 17116 25651 17119
rect 25774 17116 25780 17128
rect 25639 17088 25780 17116
rect 25639 17085 25651 17088
rect 25593 17079 25651 17085
rect 25774 17076 25780 17088
rect 25832 17116 25838 17128
rect 26142 17116 26148 17128
rect 25832 17088 26148 17116
rect 25832 17076 25838 17088
rect 26142 17076 26148 17088
rect 26200 17076 26206 17128
rect 26513 17119 26571 17125
rect 26513 17085 26525 17119
rect 26559 17116 26571 17119
rect 26786 17116 26792 17128
rect 26559 17088 26792 17116
rect 26559 17085 26571 17088
rect 26513 17079 26571 17085
rect 26786 17076 26792 17088
rect 26844 17076 26850 17128
rect 27356 17116 27384 17147
rect 27522 17144 27528 17156
rect 27580 17144 27586 17196
rect 27614 17144 27620 17196
rect 27672 17144 27678 17196
rect 27724 17193 27752 17224
rect 28988 17221 29000 17255
rect 29034 17252 29046 17255
rect 30006 17252 30012 17264
rect 29034 17224 30012 17252
rect 29034 17221 29046 17224
rect 28988 17215 29046 17221
rect 30006 17212 30012 17224
rect 30064 17212 30070 17264
rect 32214 17252 32220 17264
rect 31496 17224 32220 17252
rect 27709 17187 27767 17193
rect 27709 17153 27721 17187
rect 27755 17153 27767 17187
rect 27709 17147 27767 17153
rect 28368 17156 29776 17184
rect 28258 17116 28264 17128
rect 27356 17088 28264 17116
rect 28258 17076 28264 17088
rect 28316 17076 28322 17128
rect 23860 17020 24900 17048
rect 24949 17051 25007 17057
rect 24949 17017 24961 17051
rect 24995 17048 25007 17051
rect 28368 17048 28396 17156
rect 28718 17076 28724 17128
rect 28776 17076 28782 17128
rect 29748 17116 29776 17156
rect 30650 17144 30656 17196
rect 30708 17144 30714 17196
rect 31496 17193 31524 17224
rect 32214 17212 32220 17224
rect 32272 17212 32278 17264
rect 31481 17187 31539 17193
rect 31481 17153 31493 17187
rect 31527 17153 31539 17187
rect 31481 17147 31539 17153
rect 31570 17144 31576 17196
rect 31628 17184 31634 17196
rect 32309 17187 32367 17193
rect 32309 17184 32321 17187
rect 31628 17156 32321 17184
rect 31628 17144 31634 17156
rect 32309 17153 32321 17156
rect 32355 17153 32367 17187
rect 32309 17147 32367 17153
rect 32950 17144 32956 17196
rect 33008 17184 33014 17196
rect 33505 17187 33563 17193
rect 33505 17184 33517 17187
rect 33008 17156 33517 17184
rect 33008 17144 33014 17156
rect 33505 17153 33517 17156
rect 33551 17153 33563 17187
rect 33505 17147 33563 17153
rect 33612 17116 33640 17292
rect 36078 17280 36084 17292
rect 36136 17280 36142 17332
rect 36538 17280 36544 17332
rect 36596 17320 36602 17332
rect 39022 17320 39028 17332
rect 36596 17292 39028 17320
rect 36596 17280 36602 17292
rect 39022 17280 39028 17292
rect 39080 17280 39086 17332
rect 39577 17323 39635 17329
rect 39577 17289 39589 17323
rect 39623 17289 39635 17323
rect 39577 17283 39635 17289
rect 33772 17255 33830 17261
rect 33772 17221 33784 17255
rect 33818 17252 33830 17255
rect 36906 17252 36912 17264
rect 33818 17224 36912 17252
rect 33818 17221 33830 17224
rect 33772 17215 33830 17221
rect 36906 17212 36912 17224
rect 36964 17212 36970 17264
rect 39592 17252 39620 17283
rect 39666 17280 39672 17332
rect 39724 17320 39730 17332
rect 41601 17323 41659 17329
rect 41601 17320 41613 17323
rect 39724 17292 41613 17320
rect 39724 17280 39730 17292
rect 41601 17289 41613 17292
rect 41647 17289 41659 17323
rect 41601 17283 41659 17289
rect 42610 17280 42616 17332
rect 42668 17280 42674 17332
rect 42702 17280 42708 17332
rect 42760 17320 42766 17332
rect 46106 17320 46112 17332
rect 42760 17292 46112 17320
rect 42760 17280 42766 17292
rect 46106 17280 46112 17292
rect 46164 17280 46170 17332
rect 48498 17280 48504 17332
rect 48556 17320 48562 17332
rect 48556 17292 48912 17320
rect 48556 17280 48562 17292
rect 37476 17224 39620 17252
rect 34790 17144 34796 17196
rect 34848 17184 34854 17196
rect 35437 17187 35495 17193
rect 35437 17184 35449 17187
rect 34848 17156 35449 17184
rect 34848 17144 34854 17156
rect 35437 17153 35449 17156
rect 35483 17153 35495 17187
rect 35989 17187 36047 17193
rect 35989 17184 36001 17187
rect 35437 17147 35495 17153
rect 35544 17156 36001 17184
rect 35544 17116 35572 17156
rect 35989 17153 36001 17156
rect 36035 17153 36047 17187
rect 35989 17147 36047 17153
rect 36170 17144 36176 17196
rect 36228 17184 36234 17196
rect 37476 17193 37504 17224
rect 40310 17212 40316 17264
rect 40368 17252 40374 17264
rect 40770 17252 40776 17264
rect 40368 17224 40776 17252
rect 40368 17212 40374 17224
rect 40770 17212 40776 17224
rect 40828 17212 40834 17264
rect 40862 17212 40868 17264
rect 40920 17252 40926 17264
rect 45646 17252 45652 17264
rect 40920 17224 45652 17252
rect 40920 17212 40926 17224
rect 45646 17212 45652 17224
rect 45704 17212 45710 17264
rect 45738 17212 45744 17264
rect 45796 17252 45802 17264
rect 45922 17252 45928 17264
rect 45796 17224 45928 17252
rect 45796 17212 45802 17224
rect 45922 17212 45928 17224
rect 45980 17252 45986 17264
rect 46385 17255 46443 17261
rect 46385 17252 46397 17255
rect 45980 17224 46397 17252
rect 45980 17212 45986 17224
rect 46385 17221 46397 17224
rect 46431 17221 46443 17255
rect 46385 17215 46443 17221
rect 36265 17187 36323 17193
rect 36265 17184 36277 17187
rect 36228 17156 36277 17184
rect 36228 17144 36234 17156
rect 36265 17153 36277 17156
rect 36311 17153 36323 17187
rect 36265 17147 36323 17153
rect 36633 17187 36691 17193
rect 36633 17153 36645 17187
rect 36679 17153 36691 17187
rect 36633 17147 36691 17153
rect 37461 17187 37519 17193
rect 37461 17153 37473 17187
rect 37507 17153 37519 17187
rect 37461 17147 37519 17153
rect 29748 17088 33640 17116
rect 34532 17088 35572 17116
rect 24995 17020 28396 17048
rect 29656 17020 31754 17048
rect 24995 17017 25007 17020
rect 24949 17011 25007 17017
rect 14918 16940 14924 16992
rect 14976 16980 14982 16992
rect 17402 16980 17408 16992
rect 14976 16952 17408 16980
rect 14976 16940 14982 16952
rect 17402 16940 17408 16952
rect 17460 16940 17466 16992
rect 17494 16940 17500 16992
rect 17552 16980 17558 16992
rect 17773 16983 17831 16989
rect 17773 16980 17785 16983
rect 17552 16952 17785 16980
rect 17552 16940 17558 16952
rect 17773 16949 17785 16952
rect 17819 16949 17831 16983
rect 17773 16943 17831 16949
rect 17862 16940 17868 16992
rect 17920 16980 17926 16992
rect 18509 16983 18567 16989
rect 18509 16980 18521 16983
rect 17920 16952 18521 16980
rect 17920 16940 17926 16952
rect 18509 16949 18521 16952
rect 18555 16949 18567 16983
rect 18509 16943 18567 16949
rect 22462 16940 22468 16992
rect 22520 16980 22526 16992
rect 23109 16983 23167 16989
rect 23109 16980 23121 16983
rect 22520 16952 23121 16980
rect 22520 16940 22526 16952
rect 23109 16949 23121 16952
rect 23155 16949 23167 16983
rect 23109 16943 23167 16949
rect 23474 16940 23480 16992
rect 23532 16980 23538 16992
rect 24964 16980 24992 17011
rect 23532 16952 24992 16980
rect 26145 16983 26203 16989
rect 23532 16940 23538 16952
rect 26145 16949 26157 16983
rect 26191 16980 26203 16983
rect 26326 16980 26332 16992
rect 26191 16952 26332 16980
rect 26191 16949 26203 16952
rect 26145 16943 26203 16949
rect 26326 16940 26332 16952
rect 26384 16940 26390 16992
rect 27154 16940 27160 16992
rect 27212 16940 27218 16992
rect 27246 16940 27252 16992
rect 27304 16980 27310 16992
rect 29656 16980 29684 17020
rect 27304 16952 29684 16980
rect 27304 16940 27310 16952
rect 29730 16940 29736 16992
rect 29788 16980 29794 16992
rect 30101 16983 30159 16989
rect 30101 16980 30113 16983
rect 29788 16952 30113 16980
rect 29788 16940 29794 16952
rect 30101 16949 30113 16952
rect 30147 16949 30159 16983
rect 30101 16943 30159 16949
rect 30834 16940 30840 16992
rect 30892 16940 30898 16992
rect 31726 16980 31754 17020
rect 33318 16980 33324 16992
rect 31726 16952 33324 16980
rect 33318 16940 33324 16952
rect 33376 16980 33382 16992
rect 34532 16980 34560 17088
rect 35894 17076 35900 17128
rect 35952 17076 35958 17128
rect 36639 17116 36667 17147
rect 38562 17144 38568 17196
rect 38620 17144 38626 17196
rect 38746 17144 38752 17196
rect 38804 17184 38810 17196
rect 39393 17187 39451 17193
rect 39393 17184 39405 17187
rect 38804 17156 39405 17184
rect 38804 17144 38810 17156
rect 39393 17153 39405 17156
rect 39439 17153 39451 17187
rect 39393 17147 39451 17153
rect 40129 17187 40187 17193
rect 40129 17153 40141 17187
rect 40175 17184 40187 17187
rect 41230 17184 41236 17196
rect 40175 17156 41236 17184
rect 40175 17153 40187 17156
rect 40129 17147 40187 17153
rect 41230 17144 41236 17156
rect 41288 17144 41294 17196
rect 41417 17187 41475 17193
rect 41417 17153 41429 17187
rect 41463 17184 41475 17187
rect 42794 17184 42800 17196
rect 41463 17156 42800 17184
rect 41463 17153 41475 17156
rect 41417 17147 41475 17153
rect 42794 17144 42800 17156
rect 42852 17144 42858 17196
rect 42889 17187 42947 17193
rect 42889 17153 42901 17187
rect 42935 17153 42947 17187
rect 42889 17147 42947 17153
rect 42981 17187 43039 17193
rect 42981 17153 42993 17187
rect 43027 17153 43039 17187
rect 42981 17147 43039 17153
rect 37826 17116 37832 17128
rect 36639 17088 37832 17116
rect 34885 17051 34943 17057
rect 34885 17017 34897 17051
rect 34931 17048 34943 17051
rect 36538 17048 36544 17060
rect 34931 17020 36544 17048
rect 34931 17017 34943 17020
rect 34885 17011 34943 17017
rect 36538 17008 36544 17020
rect 36596 17008 36602 17060
rect 33376 16952 34560 16980
rect 33376 16940 33382 16952
rect 35894 16940 35900 16992
rect 35952 16980 35958 16992
rect 36639 16980 36667 17088
rect 37826 17076 37832 17088
rect 37884 17076 37890 17128
rect 41874 17076 41880 17128
rect 41932 17116 41938 17128
rect 42904 17116 42932 17147
rect 41932 17088 42932 17116
rect 41932 17076 41938 17088
rect 38470 17008 38476 17060
rect 38528 17048 38534 17060
rect 40313 17051 40371 17057
rect 40313 17048 40325 17051
rect 38528 17020 40325 17048
rect 38528 17008 38534 17020
rect 40313 17017 40325 17020
rect 40359 17017 40371 17051
rect 40313 17011 40371 17017
rect 35952 16952 36667 16980
rect 35952 16940 35958 16952
rect 37642 16940 37648 16992
rect 37700 16940 37706 16992
rect 38654 16940 38660 16992
rect 38712 16980 38718 16992
rect 38933 16983 38991 16989
rect 38933 16980 38945 16983
rect 38712 16952 38945 16980
rect 38712 16940 38718 16952
rect 38933 16949 38945 16952
rect 38979 16949 38991 16983
rect 42904 16980 42932 17088
rect 42996 17048 43024 17147
rect 43070 17144 43076 17196
rect 43128 17144 43134 17196
rect 43254 17144 43260 17196
rect 43312 17184 43318 17196
rect 43714 17184 43720 17196
rect 43312 17156 43720 17184
rect 43312 17144 43318 17156
rect 43714 17144 43720 17156
rect 43772 17144 43778 17196
rect 43809 17187 43867 17193
rect 43809 17153 43821 17187
rect 43855 17153 43867 17187
rect 43809 17147 43867 17153
rect 43070 17048 43076 17060
rect 42996 17020 43076 17048
rect 43070 17008 43076 17020
rect 43128 17008 43134 17060
rect 43824 17048 43852 17147
rect 44082 17144 44088 17196
rect 44140 17144 44146 17196
rect 44729 17187 44787 17193
rect 44729 17153 44741 17187
rect 44775 17184 44787 17187
rect 46109 17187 46167 17193
rect 44775 17156 45692 17184
rect 44775 17153 44787 17156
rect 44729 17147 44787 17153
rect 45664 17128 45692 17156
rect 46109 17153 46121 17187
rect 46155 17184 46167 17187
rect 48314 17184 48320 17196
rect 46155 17156 48320 17184
rect 46155 17153 46167 17156
rect 46109 17147 46167 17153
rect 48314 17144 48320 17156
rect 48372 17144 48378 17196
rect 48498 17144 48504 17196
rect 48556 17184 48562 17196
rect 48884 17193 48912 17292
rect 51718 17280 51724 17332
rect 51776 17280 51782 17332
rect 51905 17323 51963 17329
rect 51905 17320 51917 17323
rect 51828 17292 51917 17320
rect 51074 17252 51080 17264
rect 49160 17224 51080 17252
rect 49160 17193 49188 17224
rect 51074 17212 51080 17224
rect 51132 17212 51138 17264
rect 51166 17212 51172 17264
rect 51224 17252 51230 17264
rect 51828 17252 51856 17292
rect 51905 17289 51917 17292
rect 51951 17289 51963 17323
rect 53006 17320 53012 17332
rect 51905 17283 51963 17289
rect 52012 17292 53012 17320
rect 52012 17252 52040 17292
rect 53006 17280 53012 17292
rect 53064 17280 53070 17332
rect 58253 17323 58311 17329
rect 58253 17320 58265 17323
rect 53116 17292 58265 17320
rect 51224 17224 51856 17252
rect 51917 17224 52040 17252
rect 51224 17212 51230 17224
rect 51917 17193 51945 17224
rect 48777 17187 48835 17193
rect 48777 17184 48789 17187
rect 48556 17156 48789 17184
rect 48556 17144 48562 17156
rect 48777 17153 48789 17156
rect 48823 17153 48835 17187
rect 48777 17147 48835 17153
rect 48869 17187 48927 17193
rect 48869 17153 48881 17187
rect 48915 17153 48927 17187
rect 48869 17147 48927 17153
rect 49145 17187 49203 17193
rect 49145 17153 49157 17187
rect 49191 17153 49203 17187
rect 49145 17147 49203 17153
rect 51902 17187 51960 17193
rect 51902 17153 51914 17187
rect 51948 17153 51960 17187
rect 53116 17184 53144 17292
rect 58253 17289 58265 17292
rect 58299 17289 58311 17323
rect 58253 17283 58311 17289
rect 56229 17255 56287 17261
rect 56229 17221 56241 17255
rect 56275 17252 56287 17255
rect 56275 17224 57100 17252
rect 56275 17221 56287 17224
rect 56229 17215 56287 17221
rect 51902 17147 51960 17153
rect 52196 17156 53144 17184
rect 44174 17076 44180 17128
rect 44232 17116 44238 17128
rect 45278 17116 45284 17128
rect 44232 17088 45284 17116
rect 44232 17076 44238 17088
rect 45278 17076 45284 17088
rect 45336 17116 45342 17128
rect 45465 17119 45523 17125
rect 45465 17116 45477 17119
rect 45336 17088 45477 17116
rect 45336 17076 45342 17088
rect 45465 17085 45477 17088
rect 45511 17085 45523 17119
rect 45465 17079 45523 17085
rect 45646 17076 45652 17128
rect 45704 17076 45710 17128
rect 48222 17076 48228 17128
rect 48280 17116 48286 17128
rect 48406 17116 48412 17128
rect 48280 17088 48412 17116
rect 48280 17076 48286 17088
rect 48406 17076 48412 17088
rect 48464 17076 48470 17128
rect 48608 17088 48820 17116
rect 45554 17048 45560 17060
rect 43824 17020 45560 17048
rect 45554 17008 45560 17020
rect 45612 17008 45618 17060
rect 48608 17048 48636 17088
rect 48148 17020 48636 17048
rect 48792 17048 48820 17088
rect 48958 17076 48964 17128
rect 49016 17116 49022 17128
rect 49237 17119 49295 17125
rect 49237 17116 49249 17119
rect 49016 17088 49249 17116
rect 49016 17076 49022 17088
rect 49237 17085 49249 17088
rect 49283 17085 49295 17119
rect 49237 17079 49295 17085
rect 52196 17048 52224 17156
rect 53466 17144 53472 17196
rect 53524 17184 53530 17196
rect 55953 17187 56011 17193
rect 55953 17184 55965 17187
rect 53524 17156 55965 17184
rect 53524 17144 53530 17156
rect 55953 17153 55965 17156
rect 55999 17153 56011 17187
rect 55953 17147 56011 17153
rect 56134 17144 56140 17196
rect 56192 17144 56198 17196
rect 57072 17193 57100 17224
rect 58158 17212 58164 17264
rect 58216 17212 58222 17264
rect 56321 17187 56379 17193
rect 56321 17153 56333 17187
rect 56367 17153 56379 17187
rect 56321 17147 56379 17153
rect 57057 17187 57115 17193
rect 57057 17153 57069 17187
rect 57103 17184 57115 17187
rect 58250 17184 58256 17196
rect 57103 17156 58256 17184
rect 57103 17153 57115 17156
rect 57057 17147 57115 17153
rect 52365 17119 52423 17125
rect 52365 17085 52377 17119
rect 52411 17085 52423 17119
rect 52365 17079 52423 17085
rect 48792 17020 52224 17048
rect 48148 16980 48176 17020
rect 52270 17008 52276 17060
rect 52328 17008 52334 17060
rect 42904 16952 48176 16980
rect 48225 16983 48283 16989
rect 38933 16943 38991 16949
rect 48225 16949 48237 16983
rect 48271 16980 48283 16983
rect 48406 16980 48412 16992
rect 48271 16952 48412 16980
rect 48271 16949 48283 16952
rect 48225 16943 48283 16949
rect 48406 16940 48412 16952
rect 48464 16940 48470 16992
rect 51534 16940 51540 16992
rect 51592 16980 51598 16992
rect 51902 16980 51908 16992
rect 51592 16952 51908 16980
rect 51592 16940 51598 16952
rect 51902 16940 51908 16952
rect 51960 16980 51966 16992
rect 52380 16980 52408 17079
rect 54662 17076 54668 17128
rect 54720 17116 54726 17128
rect 56042 17116 56048 17128
rect 54720 17088 56048 17116
rect 54720 17076 54726 17088
rect 56042 17076 56048 17088
rect 56100 17116 56106 17128
rect 56336 17116 56364 17147
rect 58250 17144 58256 17156
rect 58308 17144 58314 17196
rect 56100 17088 56364 17116
rect 57333 17119 57391 17125
rect 56100 17076 56106 17088
rect 57333 17085 57345 17119
rect 57379 17116 57391 17119
rect 58986 17116 58992 17128
rect 57379 17088 58992 17116
rect 57379 17085 57391 17088
rect 57333 17079 57391 17085
rect 58986 17076 58992 17088
rect 59044 17076 59050 17128
rect 51960 16952 52408 16980
rect 51960 16940 51966 16952
rect 56226 16940 56232 16992
rect 56284 16980 56290 16992
rect 56505 16983 56563 16989
rect 56505 16980 56517 16983
rect 56284 16952 56517 16980
rect 56284 16940 56290 16952
rect 56505 16949 56517 16952
rect 56551 16949 56563 16983
rect 56505 16943 56563 16949
rect 1104 16890 58880 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 58880 16890
rect 1104 16816 58880 16838
rect 16669 16779 16727 16785
rect 16669 16745 16681 16779
rect 16715 16776 16727 16779
rect 17586 16776 17592 16788
rect 16715 16748 17592 16776
rect 16715 16745 16727 16748
rect 16669 16739 16727 16745
rect 17586 16736 17592 16748
rect 17644 16736 17650 16788
rect 25038 16776 25044 16788
rect 22204 16748 25044 16776
rect 17218 16600 17224 16652
rect 17276 16640 17282 16652
rect 19426 16640 19432 16652
rect 17276 16612 19432 16640
rect 17276 16600 17282 16612
rect 19426 16600 19432 16612
rect 19484 16640 19490 16652
rect 20073 16643 20131 16649
rect 20073 16640 20085 16643
rect 19484 16612 20085 16640
rect 19484 16600 19490 16612
rect 20073 16609 20085 16612
rect 20119 16640 20131 16643
rect 21542 16640 21548 16652
rect 20119 16612 21548 16640
rect 20119 16609 20131 16612
rect 20073 16603 20131 16609
rect 21542 16600 21548 16612
rect 21600 16640 21606 16652
rect 22204 16649 22232 16748
rect 25038 16736 25044 16748
rect 25096 16736 25102 16788
rect 27246 16776 27252 16788
rect 26528 16748 27252 16776
rect 26528 16708 26556 16748
rect 27246 16736 27252 16748
rect 27304 16736 27310 16788
rect 27632 16748 32812 16776
rect 27632 16717 27660 16748
rect 23216 16680 26556 16708
rect 26605 16711 26663 16717
rect 22189 16643 22247 16649
rect 22189 16640 22201 16643
rect 21600 16612 22201 16640
rect 21600 16600 21606 16612
rect 22189 16609 22201 16612
rect 22235 16609 22247 16643
rect 22189 16603 22247 16609
rect 1578 16532 1584 16584
rect 1636 16532 1642 16584
rect 16206 16532 16212 16584
rect 16264 16572 16270 16584
rect 16485 16575 16543 16581
rect 16485 16572 16497 16575
rect 16264 16544 16497 16572
rect 16264 16532 16270 16544
rect 16485 16541 16497 16544
rect 16531 16541 16543 16575
rect 16485 16535 16543 16541
rect 17494 16532 17500 16584
rect 17552 16532 17558 16584
rect 20346 16532 20352 16584
rect 20404 16532 20410 16584
rect 22462 16581 22468 16584
rect 22456 16572 22468 16581
rect 22423 16544 22468 16572
rect 22456 16535 22468 16544
rect 22462 16532 22468 16535
rect 22520 16532 22526 16584
rect 22830 16532 22836 16584
rect 22888 16572 22894 16584
rect 23216 16572 23244 16680
rect 26605 16677 26617 16711
rect 26651 16708 26663 16711
rect 27617 16711 27675 16717
rect 27617 16708 27629 16711
rect 26651 16680 27629 16708
rect 26651 16677 26663 16680
rect 26605 16671 26663 16677
rect 27617 16677 27629 16680
rect 27663 16677 27675 16711
rect 32784 16708 32812 16748
rect 35710 16736 35716 16788
rect 35768 16776 35774 16788
rect 36909 16779 36967 16785
rect 36909 16776 36921 16779
rect 35768 16748 36921 16776
rect 35768 16736 35774 16748
rect 36909 16745 36921 16748
rect 36955 16745 36967 16779
rect 36909 16739 36967 16745
rect 37461 16779 37519 16785
rect 37461 16745 37473 16779
rect 37507 16776 37519 16779
rect 37734 16776 37740 16788
rect 37507 16748 37740 16776
rect 37507 16745 37519 16748
rect 37461 16739 37519 16745
rect 37734 16736 37740 16748
rect 37792 16736 37798 16788
rect 38746 16736 38752 16788
rect 38804 16776 38810 16788
rect 39485 16779 39543 16785
rect 39485 16776 39497 16779
rect 38804 16748 39497 16776
rect 38804 16736 38810 16748
rect 39485 16745 39497 16748
rect 39531 16745 39543 16779
rect 39485 16739 39543 16745
rect 39574 16736 39580 16788
rect 39632 16776 39638 16788
rect 44174 16776 44180 16788
rect 39632 16748 44180 16776
rect 39632 16736 39638 16748
rect 44174 16736 44180 16748
rect 44232 16736 44238 16788
rect 44542 16736 44548 16788
rect 44600 16776 44606 16788
rect 48501 16779 48559 16785
rect 48501 16776 48513 16779
rect 44600 16748 48513 16776
rect 44600 16736 44606 16748
rect 48501 16745 48513 16748
rect 48547 16776 48559 16779
rect 49050 16776 49056 16788
rect 48547 16748 49056 16776
rect 48547 16745 48559 16748
rect 48501 16739 48559 16745
rect 49050 16736 49056 16748
rect 49108 16736 49114 16788
rect 51077 16779 51135 16785
rect 51077 16745 51089 16779
rect 51123 16776 51135 16779
rect 51166 16776 51172 16788
rect 51123 16748 51172 16776
rect 51123 16745 51135 16748
rect 51077 16739 51135 16745
rect 51166 16736 51172 16748
rect 51224 16736 51230 16788
rect 53466 16776 53472 16788
rect 51736 16748 53472 16776
rect 36078 16708 36084 16720
rect 32784 16680 36084 16708
rect 27617 16671 27675 16677
rect 36078 16668 36084 16680
rect 36136 16668 36142 16720
rect 36173 16711 36231 16717
rect 36173 16677 36185 16711
rect 36219 16708 36231 16711
rect 36219 16680 36492 16708
rect 36219 16677 36231 16680
rect 36173 16671 36231 16677
rect 25498 16600 25504 16652
rect 25556 16600 25562 16652
rect 26510 16649 26516 16652
rect 26476 16643 26516 16649
rect 26476 16609 26488 16643
rect 26476 16603 26516 16609
rect 26510 16600 26516 16603
rect 26568 16600 26574 16652
rect 26694 16600 26700 16652
rect 26752 16640 26758 16652
rect 26752 16612 27108 16640
rect 26752 16600 26758 16612
rect 22888 16544 23244 16572
rect 22888 16532 22894 16544
rect 24854 16532 24860 16584
rect 24912 16572 24918 16584
rect 25041 16575 25099 16581
rect 25041 16572 25053 16575
rect 24912 16544 25053 16572
rect 24912 16532 24918 16544
rect 25041 16541 25053 16544
rect 25087 16541 25099 16575
rect 25041 16535 25099 16541
rect 25314 16532 25320 16584
rect 25372 16532 25378 16584
rect 25682 16532 25688 16584
rect 25740 16532 25746 16584
rect 26326 16532 26332 16584
rect 26384 16532 26390 16584
rect 27080 16572 27108 16612
rect 27154 16600 27160 16652
rect 27212 16640 27218 16652
rect 27212 16612 27568 16640
rect 27212 16600 27218 16612
rect 27540 16581 27568 16612
rect 28718 16600 28724 16652
rect 28776 16640 28782 16652
rect 29733 16643 29791 16649
rect 29733 16640 29745 16643
rect 28776 16612 29745 16640
rect 28776 16600 28782 16612
rect 29733 16609 29745 16612
rect 29779 16609 29791 16643
rect 29733 16603 29791 16609
rect 33410 16600 33416 16652
rect 33468 16640 33474 16652
rect 33468 16612 35020 16640
rect 33468 16600 33474 16612
rect 27525 16575 27583 16581
rect 27080 16544 27476 16572
rect 934 16464 940 16516
rect 992 16504 998 16516
rect 1857 16507 1915 16513
rect 1857 16504 1869 16507
rect 992 16476 1869 16504
rect 992 16464 998 16476
rect 1857 16473 1869 16476
rect 1903 16473 1915 16507
rect 1857 16467 1915 16473
rect 21729 16507 21787 16513
rect 21729 16473 21741 16507
rect 21775 16504 21787 16507
rect 25590 16504 25596 16516
rect 21775 16476 25596 16504
rect 21775 16473 21787 16476
rect 21729 16467 21787 16473
rect 25590 16464 25596 16476
rect 25648 16464 25654 16516
rect 27065 16507 27123 16513
rect 27065 16473 27077 16507
rect 27111 16504 27123 16507
rect 27246 16504 27252 16516
rect 27111 16476 27252 16504
rect 27111 16473 27123 16476
rect 27065 16467 27123 16473
rect 27246 16464 27252 16476
rect 27304 16464 27310 16516
rect 27448 16504 27476 16544
rect 27525 16541 27537 16575
rect 27571 16541 27583 16575
rect 27525 16535 27583 16541
rect 27801 16575 27859 16581
rect 27801 16541 27813 16575
rect 27847 16541 27859 16575
rect 27801 16535 27859 16541
rect 27816 16504 27844 16535
rect 28350 16532 28356 16584
rect 28408 16572 28414 16584
rect 28905 16575 28963 16581
rect 28905 16572 28917 16575
rect 28408 16544 28917 16572
rect 28408 16532 28414 16544
rect 28905 16541 28917 16544
rect 28951 16541 28963 16575
rect 31849 16575 31907 16581
rect 28905 16535 28963 16541
rect 29932 16544 31754 16572
rect 29932 16504 29960 16544
rect 27448 16476 27844 16504
rect 28000 16476 29960 16504
rect 30000 16507 30058 16513
rect 18690 16396 18696 16448
rect 18748 16436 18754 16448
rect 18785 16439 18843 16445
rect 18785 16436 18797 16439
rect 18748 16408 18797 16436
rect 18748 16396 18754 16408
rect 18785 16405 18797 16408
rect 18831 16405 18843 16439
rect 18785 16399 18843 16405
rect 23569 16439 23627 16445
rect 23569 16405 23581 16439
rect 23615 16436 23627 16439
rect 24762 16436 24768 16448
rect 23615 16408 24768 16436
rect 23615 16405 23627 16408
rect 23569 16399 23627 16405
rect 24762 16396 24768 16408
rect 24820 16396 24826 16448
rect 25866 16396 25872 16448
rect 25924 16436 25930 16448
rect 28000 16445 28028 16476
rect 30000 16473 30012 16507
rect 30046 16504 30058 16507
rect 30098 16504 30104 16516
rect 30046 16476 30104 16504
rect 30046 16473 30058 16476
rect 30000 16467 30058 16473
rect 30098 16464 30104 16476
rect 30156 16464 30162 16516
rect 27985 16439 28043 16445
rect 27985 16436 27997 16439
rect 25924 16408 27997 16436
rect 25924 16396 25930 16408
rect 27985 16405 27997 16408
rect 28031 16405 28043 16439
rect 27985 16399 28043 16405
rect 28166 16396 28172 16448
rect 28224 16436 28230 16448
rect 28534 16436 28540 16448
rect 28224 16408 28540 16436
rect 28224 16396 28230 16408
rect 28534 16396 28540 16408
rect 28592 16396 28598 16448
rect 29086 16396 29092 16448
rect 29144 16396 29150 16448
rect 31110 16396 31116 16448
rect 31168 16396 31174 16448
rect 31726 16436 31754 16544
rect 31849 16541 31861 16575
rect 31895 16572 31907 16575
rect 32674 16572 32680 16584
rect 31895 16544 32680 16572
rect 31895 16541 31907 16544
rect 31849 16535 31907 16541
rect 32674 16532 32680 16544
rect 32732 16572 32738 16584
rect 32950 16572 32956 16584
rect 32732 16544 32956 16572
rect 32732 16532 32738 16544
rect 32950 16532 32956 16544
rect 33008 16532 33014 16584
rect 33686 16532 33692 16584
rect 33744 16532 33750 16584
rect 34790 16532 34796 16584
rect 34848 16572 34854 16584
rect 34885 16575 34943 16581
rect 34885 16572 34897 16575
rect 34848 16544 34897 16572
rect 34848 16532 34854 16544
rect 34885 16541 34897 16544
rect 34931 16541 34943 16575
rect 34992 16572 35020 16612
rect 35258 16575 35316 16581
rect 35258 16572 35270 16575
rect 34992 16544 35270 16572
rect 34885 16535 34943 16541
rect 35258 16541 35270 16544
rect 35304 16572 35316 16575
rect 35894 16572 35900 16584
rect 35304 16544 35900 16572
rect 35304 16541 35316 16544
rect 35258 16535 35316 16541
rect 35894 16532 35900 16544
rect 35952 16532 35958 16584
rect 35989 16575 36047 16581
rect 35989 16541 36001 16575
rect 36035 16572 36047 16575
rect 36262 16572 36268 16584
rect 36035 16544 36268 16572
rect 36035 16541 36047 16544
rect 35989 16535 36047 16541
rect 36262 16532 36268 16544
rect 36320 16532 36326 16584
rect 36464 16572 36492 16680
rect 36722 16668 36728 16720
rect 36780 16708 36786 16720
rect 43533 16711 43591 16717
rect 36780 16680 37688 16708
rect 36780 16668 36786 16680
rect 37550 16640 37556 16652
rect 37476 16612 37556 16640
rect 36725 16575 36783 16581
rect 36464 16544 36676 16572
rect 32116 16507 32174 16513
rect 32116 16473 32128 16507
rect 32162 16504 32174 16507
rect 32306 16504 32312 16516
rect 32162 16476 32312 16504
rect 32162 16473 32174 16476
rect 32116 16467 32174 16473
rect 32306 16464 32312 16476
rect 32364 16464 32370 16516
rect 34514 16504 34520 16516
rect 33244 16476 34520 16504
rect 32766 16436 32772 16448
rect 31726 16408 32772 16436
rect 32766 16396 32772 16408
rect 32824 16396 32830 16448
rect 33244 16445 33272 16476
rect 34514 16464 34520 16476
rect 34572 16464 34578 16516
rect 35069 16507 35127 16513
rect 35069 16473 35081 16507
rect 35115 16473 35127 16507
rect 35069 16467 35127 16473
rect 33229 16439 33287 16445
rect 33229 16405 33241 16439
rect 33275 16405 33287 16439
rect 33229 16399 33287 16405
rect 33870 16396 33876 16448
rect 33928 16396 33934 16448
rect 34238 16396 34244 16448
rect 34296 16436 34302 16448
rect 35084 16436 35112 16467
rect 35158 16464 35164 16516
rect 35216 16464 35222 16516
rect 36648 16504 36676 16544
rect 36725 16541 36737 16575
rect 36771 16572 36783 16575
rect 36906 16572 36912 16584
rect 36771 16544 36912 16572
rect 36771 16541 36783 16544
rect 36725 16535 36783 16541
rect 36906 16532 36912 16544
rect 36964 16532 36970 16584
rect 37476 16581 37504 16612
rect 37550 16600 37556 16612
rect 37608 16600 37614 16652
rect 37660 16581 37688 16680
rect 43533 16677 43545 16711
rect 43579 16708 43591 16711
rect 44450 16708 44456 16720
rect 43579 16680 44456 16708
rect 43579 16677 43591 16680
rect 43533 16671 43591 16677
rect 44450 16668 44456 16680
rect 44508 16668 44514 16720
rect 44634 16668 44640 16720
rect 44692 16668 44698 16720
rect 51534 16708 51540 16720
rect 48792 16680 51540 16708
rect 38102 16600 38108 16652
rect 38160 16600 38166 16652
rect 40681 16643 40739 16649
rect 40681 16609 40693 16643
rect 40727 16640 40739 16643
rect 41138 16640 41144 16652
rect 40727 16612 41144 16640
rect 40727 16609 40739 16612
rect 40681 16603 40739 16609
rect 41138 16600 41144 16612
rect 41196 16600 41202 16652
rect 44652 16640 44680 16668
rect 45186 16640 45192 16652
rect 44192 16612 45192 16640
rect 37461 16575 37519 16581
rect 37461 16541 37473 16575
rect 37507 16541 37519 16575
rect 37461 16535 37519 16541
rect 37645 16575 37703 16581
rect 37645 16541 37657 16575
rect 37691 16541 37703 16575
rect 37645 16535 37703 16541
rect 40405 16575 40463 16581
rect 40405 16541 40417 16575
rect 40451 16572 40463 16575
rect 41046 16572 41052 16584
rect 40451 16544 41052 16572
rect 40451 16541 40463 16544
rect 40405 16535 40463 16541
rect 41046 16532 41052 16544
rect 41104 16532 41110 16584
rect 42242 16532 42248 16584
rect 42300 16572 42306 16584
rect 44192 16572 44220 16612
rect 45186 16600 45192 16612
rect 45244 16600 45250 16652
rect 48792 16649 48820 16680
rect 51534 16668 51540 16680
rect 51592 16668 51598 16720
rect 48777 16643 48835 16649
rect 48777 16609 48789 16643
rect 48823 16609 48835 16643
rect 48777 16603 48835 16609
rect 42300 16544 44220 16572
rect 42300 16532 42306 16544
rect 44266 16532 44272 16584
rect 44324 16532 44330 16584
rect 44358 16532 44364 16584
rect 44416 16532 44422 16584
rect 44450 16532 44456 16584
rect 44508 16532 44514 16584
rect 44637 16575 44695 16581
rect 44637 16541 44649 16575
rect 44683 16572 44695 16575
rect 44726 16572 44732 16584
rect 44683 16544 44732 16572
rect 44683 16541 44695 16544
rect 44637 16535 44695 16541
rect 44726 16532 44732 16544
rect 44784 16532 44790 16584
rect 48869 16575 48927 16581
rect 45526 16544 48544 16572
rect 37366 16504 37372 16516
rect 36648 16476 37372 16504
rect 37366 16464 37372 16476
rect 37424 16464 37430 16516
rect 37476 16476 37688 16504
rect 34296 16408 35112 16436
rect 35454 16439 35512 16445
rect 34296 16396 34302 16408
rect 35454 16405 35466 16439
rect 35500 16436 35512 16439
rect 37476 16436 37504 16476
rect 35500 16408 37504 16436
rect 37660 16436 37688 16476
rect 37734 16464 37740 16516
rect 37792 16504 37798 16516
rect 38350 16507 38408 16513
rect 38350 16504 38362 16507
rect 37792 16476 38362 16504
rect 37792 16464 37798 16476
rect 38350 16473 38362 16476
rect 38396 16473 38408 16507
rect 38350 16467 38408 16473
rect 38562 16464 38568 16516
rect 38620 16504 38626 16516
rect 38746 16504 38752 16516
rect 38620 16476 38752 16504
rect 38620 16464 38626 16476
rect 38746 16464 38752 16476
rect 38804 16464 38810 16516
rect 39408 16476 41414 16504
rect 39408 16436 39436 16476
rect 37660 16408 39436 16436
rect 35500 16405 35512 16408
rect 35454 16399 35512 16405
rect 40034 16396 40040 16448
rect 40092 16396 40098 16448
rect 40126 16396 40132 16448
rect 40184 16436 40190 16448
rect 40497 16439 40555 16445
rect 40497 16436 40509 16439
rect 40184 16408 40509 16436
rect 40184 16396 40190 16408
rect 40497 16405 40509 16408
rect 40543 16405 40555 16439
rect 41386 16436 41414 16476
rect 41966 16464 41972 16516
rect 42024 16504 42030 16516
rect 43165 16507 43223 16513
rect 43165 16504 43177 16507
rect 42024 16476 43177 16504
rect 42024 16464 42030 16476
rect 43165 16473 43177 16476
rect 43211 16473 43223 16507
rect 43165 16467 43223 16473
rect 43346 16464 43352 16516
rect 43404 16464 43410 16516
rect 43993 16507 44051 16513
rect 43993 16473 44005 16507
rect 44039 16504 44051 16507
rect 45434 16507 45492 16513
rect 45434 16504 45446 16507
rect 44039 16476 45446 16504
rect 44039 16473 44051 16476
rect 43993 16467 44051 16473
rect 45434 16473 45446 16476
rect 45480 16473 45492 16507
rect 45434 16467 45492 16473
rect 45526 16436 45554 16544
rect 47118 16464 47124 16516
rect 47176 16464 47182 16516
rect 47305 16507 47363 16513
rect 47305 16473 47317 16507
rect 47351 16473 47363 16507
rect 47305 16467 47363 16473
rect 41386 16408 45554 16436
rect 40497 16399 40555 16405
rect 46566 16396 46572 16448
rect 46624 16436 46630 16448
rect 47320 16436 47348 16467
rect 48406 16464 48412 16516
rect 48464 16464 48470 16516
rect 48516 16504 48544 16544
rect 48869 16541 48881 16575
rect 48915 16572 48927 16575
rect 49234 16572 49240 16584
rect 48915 16544 49240 16572
rect 48915 16541 48927 16544
rect 48869 16535 48927 16541
rect 49234 16532 49240 16544
rect 49292 16532 49298 16584
rect 51736 16572 51764 16748
rect 53466 16736 53472 16748
rect 53524 16736 53530 16788
rect 56778 16736 56784 16788
rect 56836 16736 56842 16788
rect 58250 16736 58256 16788
rect 58308 16736 58314 16788
rect 53006 16668 53012 16720
rect 53064 16708 53070 16720
rect 53193 16711 53251 16717
rect 53193 16708 53205 16711
rect 53064 16680 53205 16708
rect 53064 16668 53070 16680
rect 53193 16677 53205 16680
rect 53239 16708 53251 16711
rect 56796 16708 56824 16736
rect 53239 16680 56824 16708
rect 53239 16677 53251 16680
rect 53193 16671 53251 16677
rect 55950 16640 55956 16652
rect 54864 16612 55956 16640
rect 49344 16544 51764 16572
rect 49344 16504 49372 16544
rect 51810 16532 51816 16584
rect 51868 16532 51874 16584
rect 52086 16581 52092 16584
rect 52080 16572 52092 16581
rect 52047 16544 52092 16572
rect 52080 16535 52092 16544
rect 52086 16532 52092 16535
rect 52144 16532 52150 16584
rect 54662 16532 54668 16584
rect 54720 16532 54726 16584
rect 54864 16581 54892 16612
rect 55950 16600 55956 16612
rect 56008 16600 56014 16652
rect 56042 16600 56048 16652
rect 56100 16600 56106 16652
rect 56413 16643 56471 16649
rect 56413 16609 56425 16643
rect 56459 16640 56471 16643
rect 56459 16612 56732 16640
rect 56459 16609 56471 16612
rect 56413 16603 56471 16609
rect 54849 16575 54907 16581
rect 54849 16541 54861 16575
rect 54895 16541 54907 16575
rect 54849 16535 54907 16541
rect 56226 16532 56232 16584
rect 56284 16532 56290 16584
rect 56704 16572 56732 16612
rect 56870 16600 56876 16652
rect 56928 16600 56934 16652
rect 57129 16575 57187 16581
rect 57129 16572 57141 16575
rect 56704 16544 57141 16572
rect 57129 16541 57141 16544
rect 57175 16541 57187 16575
rect 57129 16535 57187 16541
rect 48516 16476 49372 16504
rect 50801 16507 50859 16513
rect 50801 16473 50813 16507
rect 50847 16504 50859 16507
rect 50982 16504 50988 16516
rect 50847 16476 50988 16504
rect 50847 16473 50859 16476
rect 50801 16467 50859 16473
rect 50982 16464 50988 16476
rect 51040 16464 51046 16516
rect 46624 16408 47348 16436
rect 47489 16439 47547 16445
rect 46624 16396 46630 16408
rect 47489 16405 47501 16439
rect 47535 16436 47547 16439
rect 47670 16436 47676 16448
rect 47535 16408 47676 16436
rect 47535 16405 47547 16408
rect 47489 16399 47547 16405
rect 47670 16396 47676 16408
rect 47728 16396 47734 16448
rect 49053 16439 49111 16445
rect 49053 16405 49065 16439
rect 49099 16436 49111 16439
rect 51074 16436 51080 16448
rect 49099 16408 51080 16436
rect 49099 16405 49111 16408
rect 49053 16399 49111 16405
rect 51074 16396 51080 16408
rect 51132 16396 51138 16448
rect 53650 16396 53656 16448
rect 53708 16436 53714 16448
rect 54757 16439 54815 16445
rect 54757 16436 54769 16439
rect 53708 16408 54769 16436
rect 53708 16396 53714 16408
rect 54757 16405 54769 16408
rect 54803 16405 54815 16439
rect 54757 16399 54815 16405
rect 1104 16346 58880 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 50294 16346
rect 50346 16294 50358 16346
rect 50410 16294 50422 16346
rect 50474 16294 50486 16346
rect 50538 16294 50550 16346
rect 50602 16294 58880 16346
rect 1104 16272 58880 16294
rect 16206 16192 16212 16244
rect 16264 16192 16270 16244
rect 16546 16204 21404 16232
rect 11330 16124 11336 16176
rect 11388 16164 11394 16176
rect 16546 16164 16574 16204
rect 11388 16136 16574 16164
rect 21376 16164 21404 16204
rect 23566 16192 23572 16244
rect 23624 16192 23630 16244
rect 28083 16235 28141 16241
rect 28083 16201 28095 16235
rect 28129 16232 28141 16235
rect 28350 16232 28356 16244
rect 28129 16204 28356 16232
rect 28129 16201 28141 16204
rect 28083 16195 28141 16201
rect 28350 16192 28356 16204
rect 28408 16192 28414 16244
rect 31757 16235 31815 16241
rect 28460 16204 31530 16232
rect 25866 16164 25872 16176
rect 21376 16136 25872 16164
rect 11388 16124 11394 16136
rect 25866 16124 25872 16136
rect 25924 16124 25930 16176
rect 25961 16167 26019 16173
rect 25961 16133 25973 16167
rect 26007 16164 26019 16167
rect 27798 16164 27804 16176
rect 26007 16136 27804 16164
rect 26007 16133 26019 16136
rect 25961 16127 26019 16133
rect 27798 16124 27804 16136
rect 27856 16124 27862 16176
rect 28460 16164 28488 16204
rect 27908 16136 28488 16164
rect 28988 16167 29046 16173
rect 1581 16099 1639 16105
rect 1581 16065 1593 16099
rect 1627 16096 1639 16099
rect 14550 16096 14556 16108
rect 1627 16068 14556 16096
rect 1627 16065 1639 16068
rect 1581 16059 1639 16065
rect 14550 16056 14556 16068
rect 14608 16056 14614 16108
rect 16025 16099 16083 16105
rect 16025 16065 16037 16099
rect 16071 16096 16083 16099
rect 17770 16096 17776 16108
rect 16071 16068 17776 16096
rect 16071 16065 16083 16068
rect 16025 16059 16083 16065
rect 17770 16056 17776 16068
rect 17828 16056 17834 16108
rect 19426 16056 19432 16108
rect 19484 16096 19490 16108
rect 19613 16099 19671 16105
rect 19613 16096 19625 16099
rect 19484 16068 19625 16096
rect 19484 16056 19490 16068
rect 19613 16065 19625 16068
rect 19659 16065 19671 16099
rect 19613 16059 19671 16065
rect 20714 16056 20720 16108
rect 20772 16096 20778 16108
rect 22465 16099 22523 16105
rect 22465 16096 22477 16099
rect 20772 16068 22477 16096
rect 20772 16056 20778 16068
rect 22465 16065 22477 16068
rect 22511 16065 22523 16099
rect 22465 16059 22523 16065
rect 22557 16099 22615 16105
rect 22557 16065 22569 16099
rect 22603 16096 22615 16099
rect 24029 16099 24087 16105
rect 22603 16068 23796 16096
rect 22603 16065 22615 16068
rect 22557 16059 22615 16065
rect 934 15988 940 16040
rect 992 16028 998 16040
rect 1765 16031 1823 16037
rect 1765 16028 1777 16031
rect 992 16000 1777 16028
rect 992 15988 998 16000
rect 1765 15997 1777 16000
rect 1811 15997 1823 16031
rect 1765 15991 1823 15997
rect 17037 16031 17095 16037
rect 17037 15997 17049 16031
rect 17083 16028 17095 16031
rect 17218 16028 17224 16040
rect 17083 16000 17224 16028
rect 17083 15997 17095 16000
rect 17037 15991 17095 15997
rect 17218 15988 17224 16000
rect 17276 15988 17282 16040
rect 17313 16031 17371 16037
rect 17313 15997 17325 16031
rect 17359 16028 17371 16031
rect 17678 16028 17684 16040
rect 17359 16000 17684 16028
rect 17359 15997 17371 16000
rect 17313 15991 17371 15997
rect 17678 15988 17684 16000
rect 17736 15988 17742 16040
rect 18414 15988 18420 16040
rect 18472 15988 18478 16040
rect 19889 16031 19947 16037
rect 19889 15997 19901 16031
rect 19935 16028 19947 16031
rect 20346 16028 20352 16040
rect 19935 16000 20352 16028
rect 19935 15997 19947 16000
rect 19889 15991 19947 15997
rect 20346 15988 20352 16000
rect 20404 15988 20410 16040
rect 20622 15988 20628 16040
rect 20680 16028 20686 16040
rect 22278 16028 22284 16040
rect 20680 16000 22284 16028
rect 20680 15988 20686 16000
rect 22278 15988 22284 16000
rect 22336 15988 22342 16040
rect 22373 16031 22431 16037
rect 22373 15997 22385 16031
rect 22419 15997 22431 16031
rect 22373 15991 22431 15997
rect 18432 15960 18460 15988
rect 21358 15960 21364 15972
rect 18432 15932 19656 15960
rect 18230 15852 18236 15904
rect 18288 15892 18294 15904
rect 18417 15895 18475 15901
rect 18417 15892 18429 15895
rect 18288 15864 18429 15892
rect 18288 15852 18294 15864
rect 18417 15861 18429 15864
rect 18463 15861 18475 15895
rect 19628 15892 19656 15932
rect 21100 15932 21364 15960
rect 21100 15892 21128 15932
rect 21358 15920 21364 15932
rect 21416 15960 21422 15972
rect 22388 15960 22416 15991
rect 23106 15988 23112 16040
rect 23164 16028 23170 16040
rect 23164 16000 23704 16028
rect 23164 15988 23170 16000
rect 21416 15932 22416 15960
rect 21416 15920 21422 15932
rect 23382 15920 23388 15972
rect 23440 15920 23446 15972
rect 19628 15864 21128 15892
rect 18417 15855 18475 15861
rect 21174 15852 21180 15904
rect 21232 15852 21238 15904
rect 22097 15895 22155 15901
rect 22097 15861 22109 15895
rect 22143 15892 22155 15895
rect 23474 15892 23480 15904
rect 22143 15864 23480 15892
rect 22143 15861 22155 15864
rect 22097 15855 22155 15861
rect 23474 15852 23480 15864
rect 23532 15852 23538 15904
rect 23676 15892 23704 16000
rect 23768 15960 23796 16068
rect 24029 16065 24041 16099
rect 24075 16096 24087 16099
rect 24118 16096 24124 16108
rect 24075 16068 24124 16096
rect 24075 16065 24087 16068
rect 24029 16059 24087 16065
rect 24118 16056 24124 16068
rect 24176 16056 24182 16108
rect 24213 16099 24271 16105
rect 24213 16065 24225 16099
rect 24259 16096 24271 16099
rect 24394 16096 24400 16108
rect 24259 16068 24400 16096
rect 24259 16065 24271 16068
rect 24213 16059 24271 16065
rect 23842 15988 23848 16040
rect 23900 16028 23906 16040
rect 24228 16028 24256 16059
rect 24394 16056 24400 16068
rect 24452 16056 24458 16108
rect 24581 16099 24639 16105
rect 24581 16065 24593 16099
rect 24627 16096 24639 16099
rect 27908 16096 27936 16136
rect 28988 16133 29000 16167
rect 29034 16164 29046 16167
rect 30834 16164 30840 16176
rect 29034 16136 30840 16164
rect 29034 16133 29046 16136
rect 28988 16127 29046 16133
rect 30834 16124 30840 16136
rect 30892 16124 30898 16176
rect 31386 16164 31392 16176
rect 31128 16136 31392 16164
rect 24627 16068 27936 16096
rect 27985 16099 28043 16105
rect 24627 16065 24639 16068
rect 24581 16059 24639 16065
rect 27985 16065 27997 16099
rect 28031 16065 28043 16099
rect 27985 16059 28043 16065
rect 23900 16000 24256 16028
rect 23900 15988 23906 16000
rect 24302 15988 24308 16040
rect 24360 16028 24366 16040
rect 24596 16028 24624 16059
rect 25498 16037 25504 16040
rect 24360 16000 24624 16028
rect 25483 16031 25504 16037
rect 24360 15988 24366 16000
rect 25483 15997 25495 16031
rect 25483 15991 25504 15997
rect 25498 15988 25504 15991
rect 25556 15988 25562 16040
rect 25958 15988 25964 16040
rect 26016 15988 26022 16040
rect 26053 16031 26111 16037
rect 26053 15997 26065 16031
rect 26099 16028 26111 16031
rect 27890 16028 27896 16040
rect 26099 16000 27896 16028
rect 26099 15997 26111 16000
rect 26053 15991 26111 15997
rect 27890 15988 27896 16000
rect 27948 15988 27954 16040
rect 28000 16028 28028 16059
rect 28166 16056 28172 16108
rect 28224 16056 28230 16108
rect 28258 16056 28264 16108
rect 28316 16096 28322 16108
rect 30561 16099 30619 16105
rect 30561 16096 30573 16099
rect 28316 16068 30573 16096
rect 28316 16056 28322 16068
rect 30561 16065 30573 16068
rect 30607 16065 30619 16099
rect 30561 16059 30619 16065
rect 30765 16089 30823 16095
rect 28350 16028 28356 16040
rect 28000 16000 28356 16028
rect 28350 15988 28356 16000
rect 28408 15988 28414 16040
rect 28718 15988 28724 16040
rect 28776 15988 28782 16040
rect 24946 15960 24952 15972
rect 23768 15932 24952 15960
rect 24946 15920 24952 15932
rect 25004 15920 25010 15972
rect 25038 15920 25044 15972
rect 25096 15960 25102 15972
rect 28736 15960 28764 15988
rect 25096 15932 28764 15960
rect 30576 15960 30604 16059
rect 30765 16055 30777 16089
rect 30811 16086 30823 16089
rect 30811 16058 30880 16086
rect 30811 16055 30823 16058
rect 30765 16049 30823 16055
rect 30852 16028 30880 16058
rect 31018 16028 31024 16040
rect 30852 16000 31024 16028
rect 31018 15988 31024 16000
rect 31076 15988 31082 16040
rect 31128 15960 31156 16136
rect 31386 16124 31392 16136
rect 31444 16124 31450 16176
rect 31502 16096 31530 16204
rect 31757 16201 31769 16235
rect 31803 16232 31815 16235
rect 32490 16232 32496 16244
rect 31803 16204 32496 16232
rect 31803 16201 31815 16204
rect 31757 16195 31815 16201
rect 32490 16192 32496 16204
rect 32548 16232 32554 16244
rect 32548 16204 34560 16232
rect 32548 16192 32554 16204
rect 31605 16167 31663 16173
rect 31605 16133 31617 16167
rect 31651 16164 31663 16167
rect 32122 16164 32128 16176
rect 31651 16136 32128 16164
rect 31651 16133 31663 16136
rect 31605 16127 31663 16133
rect 32122 16124 32128 16136
rect 32180 16124 32186 16176
rect 32582 16124 32588 16176
rect 32640 16164 32646 16176
rect 32922 16167 32980 16173
rect 32922 16164 32934 16167
rect 32640 16136 32934 16164
rect 32640 16124 32646 16136
rect 32922 16133 32934 16136
rect 32968 16133 32980 16167
rect 32922 16127 32980 16133
rect 31502 16068 31800 16096
rect 31772 16028 31800 16068
rect 32674 16056 32680 16108
rect 32732 16056 32738 16108
rect 33502 16096 33508 16108
rect 32784 16068 33508 16096
rect 32784 16028 32812 16068
rect 33502 16056 33508 16068
rect 33560 16056 33566 16108
rect 34532 16105 34560 16204
rect 34606 16192 34612 16244
rect 34664 16192 34670 16244
rect 36906 16192 36912 16244
rect 36964 16232 36970 16244
rect 37458 16232 37464 16244
rect 36964 16204 37464 16232
rect 36964 16192 36970 16204
rect 37458 16192 37464 16204
rect 37516 16192 37522 16244
rect 37553 16235 37611 16241
rect 37553 16201 37565 16235
rect 37599 16232 37611 16235
rect 37734 16232 37740 16244
rect 37599 16204 37740 16232
rect 37599 16201 37611 16204
rect 37553 16195 37611 16201
rect 37734 16192 37740 16204
rect 37792 16192 37798 16244
rect 41601 16235 41659 16241
rect 37936 16204 41552 16232
rect 37642 16164 37648 16176
rect 35469 16136 37648 16164
rect 34517 16099 34575 16105
rect 34517 16065 34529 16099
rect 34563 16065 34575 16099
rect 34517 16059 34575 16065
rect 34698 16056 34704 16108
rect 34756 16056 34762 16108
rect 35469 16105 35497 16136
rect 37642 16124 37648 16136
rect 37700 16124 37706 16176
rect 35437 16099 35497 16105
rect 35437 16065 35449 16099
rect 35483 16066 35497 16099
rect 35483 16065 35495 16066
rect 35437 16059 35495 16065
rect 35526 16056 35532 16108
rect 35584 16096 35590 16108
rect 36725 16099 36783 16105
rect 36725 16096 36737 16099
rect 35584 16068 36737 16096
rect 35584 16056 35590 16068
rect 36725 16065 36737 16068
rect 36771 16065 36783 16099
rect 36725 16059 36783 16065
rect 36814 16056 36820 16108
rect 36872 16096 36878 16108
rect 36909 16099 36967 16105
rect 36909 16096 36921 16099
rect 36872 16068 36921 16096
rect 36872 16056 36878 16068
rect 36909 16065 36921 16068
rect 36955 16065 36967 16099
rect 36909 16059 36967 16065
rect 37826 16056 37832 16108
rect 37884 16056 37890 16108
rect 37936 16105 37964 16204
rect 38654 16164 38660 16176
rect 38028 16136 38660 16164
rect 38028 16105 38056 16136
rect 38654 16124 38660 16136
rect 38712 16124 38718 16176
rect 38924 16167 38982 16173
rect 38924 16133 38936 16167
rect 38970 16164 38982 16167
rect 40034 16164 40040 16176
rect 38970 16136 40040 16164
rect 38970 16133 38982 16136
rect 38924 16127 38982 16133
rect 40034 16124 40040 16136
rect 40092 16124 40098 16176
rect 41524 16164 41552 16204
rect 41601 16201 41613 16235
rect 41647 16232 41659 16235
rect 41782 16232 41788 16244
rect 41647 16204 41788 16232
rect 41647 16201 41659 16204
rect 41601 16195 41659 16201
rect 41782 16192 41788 16204
rect 41840 16192 41846 16244
rect 42794 16192 42800 16244
rect 42852 16232 42858 16244
rect 43625 16235 43683 16241
rect 43625 16232 43637 16235
rect 42852 16204 43637 16232
rect 42852 16192 42858 16204
rect 43625 16201 43637 16204
rect 43671 16201 43683 16235
rect 43625 16195 43683 16201
rect 45465 16235 45523 16241
rect 45465 16201 45477 16235
rect 45511 16232 45523 16235
rect 45511 16204 45545 16232
rect 45511 16201 45523 16204
rect 45465 16195 45523 16201
rect 43070 16164 43076 16176
rect 41524 16136 43076 16164
rect 43070 16124 43076 16136
rect 43128 16164 43134 16176
rect 44358 16164 44364 16176
rect 43128 16136 44364 16164
rect 43128 16124 43134 16136
rect 44358 16124 44364 16136
rect 44416 16124 44422 16176
rect 45186 16124 45192 16176
rect 45244 16164 45250 16176
rect 45480 16164 45508 16195
rect 47118 16192 47124 16244
rect 47176 16232 47182 16244
rect 47762 16232 47768 16244
rect 47176 16204 47768 16232
rect 47176 16192 47182 16204
rect 47762 16192 47768 16204
rect 47820 16232 47826 16244
rect 47820 16204 48084 16232
rect 47820 16192 47826 16204
rect 48056 16164 48084 16204
rect 48130 16192 48136 16244
rect 48188 16232 48194 16244
rect 49145 16235 49203 16241
rect 49145 16232 49157 16235
rect 48188 16204 49157 16232
rect 48188 16192 48194 16204
rect 49145 16201 49157 16204
rect 49191 16232 49203 16235
rect 49510 16232 49516 16244
rect 49191 16204 49516 16232
rect 49191 16201 49203 16204
rect 49145 16195 49203 16201
rect 49510 16192 49516 16204
rect 49568 16192 49574 16244
rect 53650 16192 53656 16244
rect 53708 16192 53714 16244
rect 55585 16235 55643 16241
rect 55585 16201 55597 16235
rect 55631 16232 55643 16235
rect 55950 16232 55956 16244
rect 55631 16204 55956 16232
rect 55631 16201 55643 16204
rect 55585 16195 55643 16201
rect 55950 16192 55956 16204
rect 56008 16192 56014 16244
rect 48314 16164 48320 16176
rect 45244 16136 47808 16164
rect 48056 16136 48320 16164
rect 45244 16124 45250 16136
rect 37921 16099 37979 16105
rect 37921 16065 37933 16099
rect 37967 16065 37979 16099
rect 37921 16059 37979 16065
rect 38013 16099 38071 16105
rect 38013 16065 38025 16099
rect 38059 16065 38071 16099
rect 38013 16059 38071 16065
rect 38197 16099 38255 16105
rect 38197 16065 38209 16099
rect 38243 16096 38255 16099
rect 39758 16096 39764 16108
rect 38243 16068 39764 16096
rect 38243 16065 38255 16068
rect 38197 16059 38255 16065
rect 39758 16056 39764 16068
rect 39816 16056 39822 16108
rect 43346 16096 43352 16108
rect 39868 16068 43352 16096
rect 38562 16028 38568 16040
rect 31772 16000 32812 16028
rect 35176 16000 38568 16028
rect 35176 15972 35204 16000
rect 38562 15988 38568 16000
rect 38620 15988 38626 16040
rect 38654 15988 38660 16040
rect 38712 15988 38718 16040
rect 30576 15932 31156 15960
rect 34057 15963 34115 15969
rect 25096 15920 25102 15932
rect 34057 15929 34069 15963
rect 34103 15960 34115 15963
rect 35158 15960 35164 15972
rect 34103 15932 35164 15960
rect 34103 15929 34115 15932
rect 34057 15923 34115 15929
rect 35158 15920 35164 15932
rect 35216 15920 35222 15972
rect 36725 15963 36783 15969
rect 36725 15929 36737 15963
rect 36771 15960 36783 15963
rect 37918 15960 37924 15972
rect 36771 15932 37924 15960
rect 36771 15929 36783 15932
rect 36725 15923 36783 15929
rect 37918 15920 37924 15932
rect 37976 15920 37982 15972
rect 28258 15892 28264 15904
rect 23676 15864 28264 15892
rect 28258 15852 28264 15864
rect 28316 15852 28322 15904
rect 30101 15895 30159 15901
rect 30101 15861 30113 15895
rect 30147 15892 30159 15895
rect 30282 15892 30288 15904
rect 30147 15864 30288 15892
rect 30147 15861 30159 15864
rect 30101 15855 30159 15861
rect 30282 15852 30288 15864
rect 30340 15852 30346 15904
rect 30374 15852 30380 15904
rect 30432 15892 30438 15904
rect 30650 15892 30656 15904
rect 30432 15864 30656 15892
rect 30432 15852 30438 15864
rect 30650 15852 30656 15864
rect 30708 15892 30714 15904
rect 30929 15895 30987 15901
rect 30929 15892 30941 15895
rect 30708 15864 30941 15892
rect 30708 15852 30714 15864
rect 30929 15861 30941 15864
rect 30975 15861 30987 15895
rect 30929 15855 30987 15861
rect 31018 15852 31024 15904
rect 31076 15892 31082 15904
rect 31573 15895 31631 15901
rect 31573 15892 31585 15895
rect 31076 15864 31585 15892
rect 31076 15852 31082 15864
rect 31573 15861 31585 15864
rect 31619 15861 31631 15895
rect 31573 15855 31631 15861
rect 34698 15852 34704 15904
rect 34756 15892 34762 15904
rect 35621 15895 35679 15901
rect 35621 15892 35633 15895
rect 34756 15864 35633 15892
rect 34756 15852 34762 15864
rect 35621 15861 35633 15864
rect 35667 15861 35679 15895
rect 35621 15855 35679 15861
rect 36078 15852 36084 15904
rect 36136 15892 36142 15904
rect 37734 15892 37740 15904
rect 36136 15864 37740 15892
rect 36136 15852 36142 15864
rect 37734 15852 37740 15864
rect 37792 15852 37798 15904
rect 38194 15852 38200 15904
rect 38252 15892 38258 15904
rect 39868 15892 39896 16068
rect 43346 16056 43352 16068
rect 43404 16096 43410 16108
rect 43441 16099 43499 16105
rect 43441 16096 43453 16099
rect 43404 16068 43453 16096
rect 43404 16056 43410 16068
rect 43441 16065 43453 16068
rect 43487 16065 43499 16099
rect 43441 16059 43499 16065
rect 39942 15988 39948 16040
rect 40000 16028 40006 16040
rect 41690 16028 41696 16040
rect 40000 16000 41696 16028
rect 40000 15988 40006 16000
rect 41690 15988 41696 16000
rect 41748 15988 41754 16040
rect 41877 16031 41935 16037
rect 41877 15997 41889 16031
rect 41923 15997 41935 16031
rect 43456 16028 43484 16059
rect 44174 16056 44180 16108
rect 44232 16056 44238 16108
rect 46750 16056 46756 16108
rect 46808 16056 46814 16108
rect 47780 16105 47808 16136
rect 48314 16124 48320 16136
rect 48372 16124 48378 16176
rect 52454 16124 52460 16176
rect 52512 16164 52518 16176
rect 53469 16167 53527 16173
rect 53469 16164 53481 16167
rect 52512 16136 53481 16164
rect 52512 16124 52518 16136
rect 53469 16133 53481 16136
rect 53515 16133 53527 16167
rect 53469 16127 53527 16133
rect 53558 16124 53564 16176
rect 53616 16164 53622 16176
rect 54450 16167 54508 16173
rect 54450 16164 54462 16167
rect 53616 16136 54462 16164
rect 53616 16124 53622 16136
rect 54450 16133 54462 16136
rect 54496 16133 54508 16167
rect 54450 16127 54508 16133
rect 58158 16124 58164 16176
rect 58216 16124 58222 16176
rect 59078 16124 59084 16176
rect 59136 16164 59142 16176
rect 59722 16164 59728 16176
rect 59136 16136 59728 16164
rect 59136 16124 59142 16136
rect 59722 16124 59728 16136
rect 59780 16124 59786 16176
rect 48038 16105 48044 16108
rect 47765 16099 47823 16105
rect 47765 16065 47777 16099
rect 47811 16065 47823 16099
rect 47765 16059 47823 16065
rect 48032 16059 48044 16105
rect 48038 16056 48044 16059
rect 48096 16056 48102 16108
rect 50065 16099 50123 16105
rect 50065 16065 50077 16099
rect 50111 16096 50123 16099
rect 50154 16096 50160 16108
rect 50111 16068 50160 16096
rect 50111 16065 50123 16068
rect 50065 16059 50123 16065
rect 50154 16056 50160 16068
rect 50212 16056 50218 16108
rect 50332 16099 50390 16105
rect 50332 16065 50344 16099
rect 50378 16096 50390 16099
rect 50614 16096 50620 16108
rect 50378 16068 50620 16096
rect 50378 16065 50390 16068
rect 50332 16059 50390 16065
rect 50614 16056 50620 16068
rect 50672 16056 50678 16108
rect 51074 16056 51080 16108
rect 51132 16096 51138 16108
rect 53745 16099 53803 16105
rect 53745 16096 53757 16099
rect 51132 16068 53757 16096
rect 51132 16056 51138 16068
rect 53745 16065 53757 16068
rect 53791 16065 53803 16099
rect 56870 16096 56876 16108
rect 53745 16059 53803 16065
rect 54220 16068 56876 16096
rect 46566 16028 46572 16040
rect 43456 16000 46572 16028
rect 41877 15991 41935 15997
rect 41892 15960 41920 15991
rect 46566 15988 46572 16000
rect 46624 15988 46630 16040
rect 46842 15988 46848 16040
rect 46900 15988 46906 16040
rect 46937 16031 46995 16037
rect 46937 15997 46949 16031
rect 46983 15997 46995 16031
rect 46937 15991 46995 15997
rect 44082 15960 44088 15972
rect 41892 15932 44088 15960
rect 44082 15920 44088 15932
rect 44140 15960 44146 15972
rect 46952 15960 46980 15991
rect 51810 15988 51816 16040
rect 51868 16028 51874 16040
rect 54220 16037 54248 16068
rect 56870 16056 56876 16068
rect 56928 16056 56934 16108
rect 54205 16031 54263 16037
rect 54205 16028 54217 16031
rect 51868 16000 54217 16028
rect 51868 15988 51874 16000
rect 54205 15997 54217 16000
rect 54251 15997 54263 16031
rect 54205 15991 54263 15997
rect 58345 15963 58403 15969
rect 58345 15960 58357 15963
rect 44140 15932 46980 15960
rect 51046 15932 53604 15960
rect 44140 15920 44146 15932
rect 38252 15864 39896 15892
rect 38252 15852 38258 15864
rect 40034 15852 40040 15904
rect 40092 15852 40098 15904
rect 41230 15852 41236 15904
rect 41288 15852 41294 15904
rect 43070 15852 43076 15904
rect 43128 15892 43134 15904
rect 43254 15892 43260 15904
rect 43128 15864 43260 15892
rect 43128 15852 43134 15864
rect 43254 15852 43260 15864
rect 43312 15892 43318 15904
rect 44726 15892 44732 15904
rect 43312 15864 44732 15892
rect 43312 15852 43318 15864
rect 44726 15852 44732 15864
rect 44784 15852 44790 15904
rect 46382 15852 46388 15904
rect 46440 15852 46446 15904
rect 46566 15852 46572 15904
rect 46624 15892 46630 15904
rect 51046 15892 51074 15932
rect 46624 15864 51074 15892
rect 51445 15895 51503 15901
rect 46624 15852 46630 15864
rect 51445 15861 51457 15895
rect 51491 15892 51503 15895
rect 51534 15892 51540 15904
rect 51491 15864 51540 15892
rect 51491 15861 51503 15864
rect 51445 15855 51503 15861
rect 51534 15852 51540 15864
rect 51592 15852 51598 15904
rect 53466 15852 53472 15904
rect 53524 15852 53530 15904
rect 53576 15892 53604 15932
rect 55140 15932 58357 15960
rect 55140 15892 55168 15932
rect 58345 15929 58357 15932
rect 58391 15929 58403 15963
rect 58345 15923 58403 15929
rect 53576 15864 55168 15892
rect 1104 15802 58880 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 58880 15802
rect 1104 15728 58880 15750
rect 14550 15648 14556 15700
rect 14608 15648 14614 15700
rect 23198 15688 23204 15700
rect 14844 15660 23204 15688
rect 11422 15512 11428 15564
rect 11480 15512 11486 15564
rect 11790 15512 11796 15564
rect 11848 15512 11854 15564
rect 14844 15561 14872 15660
rect 23198 15648 23204 15660
rect 23256 15648 23262 15700
rect 23382 15648 23388 15700
rect 23440 15688 23446 15700
rect 23661 15691 23719 15697
rect 23661 15688 23673 15691
rect 23440 15660 23673 15688
rect 23440 15648 23446 15660
rect 23661 15657 23673 15660
rect 23707 15657 23719 15691
rect 23661 15651 23719 15657
rect 25038 15648 25044 15700
rect 25096 15648 25102 15700
rect 25590 15648 25596 15700
rect 25648 15688 25654 15700
rect 28994 15688 29000 15700
rect 25648 15660 29000 15688
rect 25648 15648 25654 15660
rect 28994 15648 29000 15660
rect 29052 15648 29058 15700
rect 29178 15648 29184 15700
rect 29236 15688 29242 15700
rect 30006 15688 30012 15700
rect 29236 15660 30012 15688
rect 29236 15648 29242 15660
rect 30006 15648 30012 15660
rect 30064 15648 30070 15700
rect 31018 15648 31024 15700
rect 31076 15688 31082 15700
rect 31113 15691 31171 15697
rect 31113 15688 31125 15691
rect 31076 15660 31125 15688
rect 31076 15648 31082 15660
rect 31113 15657 31125 15660
rect 31159 15657 31171 15691
rect 31113 15651 31171 15657
rect 32214 15648 32220 15700
rect 32272 15648 32278 15700
rect 32953 15691 33011 15697
rect 32953 15657 32965 15691
rect 32999 15688 33011 15691
rect 33686 15688 33692 15700
rect 32999 15660 33692 15688
rect 32999 15657 33011 15660
rect 32953 15651 33011 15657
rect 33686 15648 33692 15660
rect 33744 15648 33750 15700
rect 39942 15688 39948 15700
rect 34624 15660 39948 15688
rect 15470 15620 15476 15632
rect 14936 15592 15476 15620
rect 14936 15561 14964 15592
rect 15470 15580 15476 15592
rect 15528 15620 15534 15632
rect 15528 15592 15976 15620
rect 15528 15580 15534 15592
rect 14829 15555 14887 15561
rect 14829 15521 14841 15555
rect 14875 15521 14887 15555
rect 14829 15515 14887 15521
rect 14921 15555 14979 15561
rect 14921 15521 14933 15555
rect 14967 15521 14979 15555
rect 14921 15515 14979 15521
rect 15838 15512 15844 15564
rect 15896 15512 15902 15564
rect 15948 15561 15976 15592
rect 17770 15580 17776 15632
rect 17828 15580 17834 15632
rect 20257 15623 20315 15629
rect 20257 15589 20269 15623
rect 20303 15589 20315 15623
rect 20257 15583 20315 15589
rect 15933 15555 15991 15561
rect 15933 15521 15945 15555
rect 15979 15521 15991 15555
rect 15933 15515 15991 15521
rect 17497 15555 17555 15561
rect 17497 15521 17509 15555
rect 17543 15552 17555 15555
rect 17862 15552 17868 15564
rect 17543 15524 17868 15552
rect 17543 15521 17555 15524
rect 17497 15515 17555 15521
rect 17862 15512 17868 15524
rect 17920 15512 17926 15564
rect 20272 15552 20300 15583
rect 28718 15580 28724 15632
rect 28776 15620 28782 15632
rect 34624 15620 34652 15660
rect 39942 15648 39948 15660
rect 40000 15648 40006 15700
rect 42242 15688 42248 15700
rect 40696 15660 42248 15688
rect 28776 15592 34652 15620
rect 28776 15580 28782 15592
rect 38654 15580 38660 15632
rect 38712 15620 38718 15632
rect 40696 15620 40724 15660
rect 42242 15648 42248 15660
rect 42300 15648 42306 15700
rect 51813 15691 51871 15697
rect 47964 15660 51764 15688
rect 38712 15592 40724 15620
rect 38712 15580 38718 15592
rect 21266 15552 21272 15564
rect 20272 15524 21272 15552
rect 21266 15512 21272 15524
rect 21324 15512 21330 15564
rect 21637 15555 21695 15561
rect 21637 15521 21649 15555
rect 21683 15552 21695 15555
rect 22281 15555 22339 15561
rect 21683 15524 22232 15552
rect 21683 15521 21695 15524
rect 21637 15515 21695 15521
rect 1581 15487 1639 15493
rect 1581 15453 1593 15487
rect 1627 15484 1639 15487
rect 2682 15484 2688 15496
rect 1627 15456 2688 15484
rect 1627 15453 1639 15456
rect 1581 15447 1639 15453
rect 2682 15444 2688 15456
rect 2740 15444 2746 15496
rect 11330 15444 11336 15496
rect 11388 15444 11394 15496
rect 11698 15444 11704 15496
rect 11756 15444 11762 15496
rect 14737 15487 14795 15493
rect 14737 15453 14749 15487
rect 14783 15453 14795 15487
rect 14737 15447 14795 15453
rect 15013 15487 15071 15493
rect 15013 15453 15025 15487
rect 15059 15484 15071 15487
rect 15654 15484 15660 15496
rect 15059 15456 15660 15484
rect 15059 15453 15071 15456
rect 15013 15447 15071 15453
rect 934 15376 940 15428
rect 992 15416 998 15428
rect 1857 15419 1915 15425
rect 1857 15416 1869 15419
rect 992 15388 1869 15416
rect 992 15376 998 15388
rect 1857 15385 1869 15388
rect 1903 15385 1915 15419
rect 1857 15379 1915 15385
rect 10502 15376 10508 15428
rect 10560 15416 10566 15428
rect 10689 15419 10747 15425
rect 10689 15416 10701 15419
rect 10560 15388 10701 15416
rect 10560 15376 10566 15388
rect 10689 15385 10701 15388
rect 10735 15385 10747 15419
rect 14752 15416 14780 15447
rect 15654 15444 15660 15456
rect 15712 15444 15718 15496
rect 15746 15444 15752 15496
rect 15804 15444 15810 15496
rect 16025 15487 16083 15493
rect 16025 15453 16037 15487
rect 16071 15484 16083 15487
rect 16206 15484 16212 15496
rect 16071 15456 16212 15484
rect 16071 15453 16083 15456
rect 16025 15447 16083 15453
rect 16206 15444 16212 15456
rect 16264 15444 16270 15496
rect 17405 15487 17463 15493
rect 17405 15453 17417 15487
rect 17451 15484 17463 15487
rect 20714 15484 20720 15496
rect 17451 15456 20720 15484
rect 17451 15453 17463 15456
rect 17405 15447 17463 15453
rect 20714 15444 20720 15456
rect 20772 15444 20778 15496
rect 21361 15487 21419 15493
rect 21361 15453 21373 15487
rect 21407 15453 21419 15487
rect 21361 15447 21419 15453
rect 15764 15416 15792 15444
rect 14752 15388 15792 15416
rect 10689 15379 10747 15385
rect 17954 15376 17960 15428
rect 18012 15416 18018 15428
rect 18233 15419 18291 15425
rect 18233 15416 18245 15419
rect 18012 15388 18245 15416
rect 18012 15376 18018 15388
rect 18233 15385 18245 15388
rect 18279 15385 18291 15419
rect 18233 15379 18291 15385
rect 12250 15308 12256 15360
rect 12308 15348 12314 15360
rect 15565 15351 15623 15357
rect 15565 15348 15577 15351
rect 12308 15320 15577 15348
rect 12308 15308 12314 15320
rect 15565 15317 15577 15320
rect 15611 15317 15623 15351
rect 18248 15348 18276 15379
rect 18414 15376 18420 15428
rect 18472 15376 18478 15428
rect 19981 15419 20039 15425
rect 19981 15416 19993 15419
rect 18524 15388 19993 15416
rect 18524 15348 18552 15388
rect 19981 15385 19993 15388
rect 20027 15416 20039 15419
rect 20622 15416 20628 15428
rect 20027 15388 20628 15416
rect 20027 15385 20039 15388
rect 19981 15379 20039 15385
rect 20622 15376 20628 15388
rect 20680 15376 20686 15428
rect 21376 15416 21404 15447
rect 21450 15444 21456 15496
rect 21508 15444 21514 15496
rect 21545 15487 21603 15493
rect 21545 15453 21557 15487
rect 21591 15484 21603 15487
rect 22204 15484 22232 15524
rect 22281 15521 22293 15555
rect 22327 15552 22339 15555
rect 25038 15552 25044 15564
rect 22327 15524 25044 15552
rect 22327 15521 22339 15524
rect 22281 15515 22339 15521
rect 25038 15512 25044 15524
rect 25096 15512 25102 15564
rect 29270 15552 29276 15564
rect 28552 15524 29276 15552
rect 21591 15456 22094 15484
rect 22204 15456 23428 15484
rect 21591 15453 21603 15456
rect 21545 15447 21603 15453
rect 21634 15416 21640 15428
rect 21376 15388 21640 15416
rect 21634 15376 21640 15388
rect 21692 15376 21698 15428
rect 22066 15416 22094 15456
rect 22186 15416 22192 15428
rect 22066 15388 22192 15416
rect 22186 15376 22192 15388
rect 22244 15376 22250 15428
rect 22370 15376 22376 15428
rect 22428 15416 22434 15428
rect 22649 15419 22707 15425
rect 22649 15416 22661 15419
rect 22428 15388 22661 15416
rect 22428 15376 22434 15388
rect 22649 15385 22661 15388
rect 22695 15416 22707 15419
rect 22738 15416 22744 15428
rect 22695 15388 22744 15416
rect 22695 15385 22707 15388
rect 22649 15379 22707 15385
rect 22738 15376 22744 15388
rect 22796 15376 22802 15428
rect 23017 15419 23075 15425
rect 23017 15385 23029 15419
rect 23063 15416 23075 15419
rect 23106 15416 23112 15428
rect 23063 15388 23112 15416
rect 23063 15385 23075 15388
rect 23017 15379 23075 15385
rect 23106 15376 23112 15388
rect 23164 15376 23170 15428
rect 18248 15320 18552 15348
rect 15565 15311 15623 15317
rect 18598 15308 18604 15360
rect 18656 15308 18662 15360
rect 20254 15308 20260 15360
rect 20312 15348 20318 15360
rect 20441 15351 20499 15357
rect 20441 15348 20453 15351
rect 20312 15320 20453 15348
rect 20312 15308 20318 15320
rect 20441 15317 20453 15320
rect 20487 15317 20499 15351
rect 20441 15311 20499 15317
rect 20990 15308 20996 15360
rect 21048 15348 21054 15360
rect 21177 15351 21235 15357
rect 21177 15348 21189 15351
rect 21048 15320 21189 15348
rect 21048 15308 21054 15320
rect 21177 15317 21189 15320
rect 21223 15317 21235 15351
rect 21177 15311 21235 15317
rect 22462 15308 22468 15360
rect 22520 15308 22526 15360
rect 22554 15308 22560 15360
rect 22612 15308 22618 15360
rect 23400 15348 23428 15456
rect 23474 15444 23480 15496
rect 23532 15444 23538 15496
rect 28169 15487 28227 15493
rect 28169 15453 28181 15487
rect 28215 15453 28227 15487
rect 28169 15447 28227 15453
rect 23750 15376 23756 15428
rect 23808 15416 23814 15428
rect 25317 15419 25375 15425
rect 25317 15416 25329 15419
rect 23808 15388 25329 15416
rect 23808 15376 23814 15388
rect 25317 15385 25329 15388
rect 25363 15385 25375 15419
rect 25317 15379 25375 15385
rect 25498 15376 25504 15428
rect 25556 15376 25562 15428
rect 25593 15419 25651 15425
rect 25593 15385 25605 15419
rect 25639 15416 25651 15419
rect 26694 15416 26700 15428
rect 25639 15388 26700 15416
rect 25639 15385 25651 15388
rect 25593 15379 25651 15385
rect 26694 15376 26700 15388
rect 26752 15376 26758 15428
rect 28184 15416 28212 15447
rect 28552 15416 28580 15524
rect 29270 15512 29276 15524
rect 29328 15512 29334 15564
rect 30009 15555 30067 15561
rect 30009 15521 30021 15555
rect 30055 15552 30067 15555
rect 30650 15552 30656 15564
rect 30055 15524 30656 15552
rect 30055 15521 30067 15524
rect 30009 15515 30067 15521
rect 30650 15512 30656 15524
rect 30708 15512 30714 15564
rect 31665 15555 31723 15561
rect 31665 15521 31677 15555
rect 31711 15552 31723 15555
rect 34698 15552 34704 15564
rect 31711 15524 34704 15552
rect 31711 15521 31723 15524
rect 31665 15515 31723 15521
rect 34698 15512 34704 15524
rect 34756 15512 34762 15564
rect 40696 15561 40724 15592
rect 41690 15580 41696 15632
rect 41748 15620 41754 15632
rect 42061 15623 42119 15629
rect 42061 15620 42073 15623
rect 41748 15592 42073 15620
rect 41748 15580 41754 15592
rect 42061 15589 42073 15592
rect 42107 15589 42119 15623
rect 42061 15583 42119 15589
rect 38841 15555 38899 15561
rect 38841 15521 38853 15555
rect 38887 15521 38899 15555
rect 38841 15515 38899 15521
rect 40681 15555 40739 15561
rect 40681 15521 40693 15555
rect 40727 15521 40739 15555
rect 42260 15552 42288 15648
rect 46842 15580 46848 15632
rect 46900 15620 46906 15632
rect 46937 15623 46995 15629
rect 46937 15620 46949 15623
rect 46900 15592 46949 15620
rect 46900 15580 46906 15592
rect 46937 15589 46949 15592
rect 46983 15589 46995 15623
rect 46937 15583 46995 15589
rect 47486 15580 47492 15632
rect 47544 15620 47550 15632
rect 47762 15620 47768 15632
rect 47544 15592 47768 15620
rect 47544 15580 47550 15592
rect 47762 15580 47768 15592
rect 47820 15580 47826 15632
rect 42981 15555 43039 15561
rect 42981 15552 42993 15555
rect 42260 15524 42993 15552
rect 40681 15515 40739 15521
rect 42981 15521 42993 15524
rect 43027 15521 43039 15555
rect 42981 15515 43039 15521
rect 28902 15444 28908 15496
rect 28960 15444 28966 15496
rect 29917 15487 29975 15493
rect 29917 15453 29929 15487
rect 29963 15484 29975 15487
rect 30190 15484 30196 15496
rect 29963 15456 30196 15484
rect 29963 15453 29975 15456
rect 29917 15447 29975 15453
rect 30190 15444 30196 15456
rect 30248 15444 30254 15496
rect 30745 15487 30803 15493
rect 30745 15453 30757 15487
rect 30791 15453 30803 15487
rect 30745 15447 30803 15453
rect 30760 15416 30788 15447
rect 30926 15444 30932 15496
rect 30984 15444 30990 15496
rect 31018 15444 31024 15496
rect 31076 15484 31082 15496
rect 31941 15487 31999 15493
rect 31941 15484 31953 15487
rect 31076 15456 31953 15484
rect 31076 15444 31082 15456
rect 31941 15453 31953 15456
rect 31987 15453 31999 15487
rect 31941 15447 31999 15453
rect 32769 15487 32827 15493
rect 32769 15453 32781 15487
rect 32815 15453 32827 15487
rect 32769 15447 32827 15453
rect 32784 15416 32812 15447
rect 32950 15444 32956 15496
rect 33008 15484 33014 15496
rect 33597 15487 33655 15493
rect 33597 15484 33609 15487
rect 33008 15456 33609 15484
rect 33008 15444 33014 15456
rect 33597 15453 33609 15456
rect 33643 15453 33655 15487
rect 33597 15447 33655 15453
rect 33781 15487 33839 15493
rect 33781 15453 33793 15487
rect 33827 15453 33839 15487
rect 33781 15447 33839 15453
rect 33965 15487 34023 15493
rect 33965 15453 33977 15487
rect 34011 15484 34023 15487
rect 34790 15484 34796 15496
rect 34011 15456 34796 15484
rect 34011 15453 34023 15456
rect 33965 15447 34023 15453
rect 28184 15388 28580 15416
rect 28966 15388 30788 15416
rect 31036 15388 32812 15416
rect 26142 15348 26148 15360
rect 23400 15320 26148 15348
rect 26142 15308 26148 15320
rect 26200 15308 26206 15360
rect 27890 15308 27896 15360
rect 27948 15348 27954 15360
rect 28258 15348 28264 15360
rect 27948 15320 28264 15348
rect 27948 15308 27954 15320
rect 28258 15308 28264 15320
rect 28316 15308 28322 15360
rect 28350 15308 28356 15360
rect 28408 15348 28414 15360
rect 28966 15348 28994 15388
rect 31036 15360 31064 15388
rect 33502 15376 33508 15428
rect 33560 15416 33566 15428
rect 33796 15416 33824 15447
rect 34790 15444 34796 15456
rect 34848 15444 34854 15496
rect 38470 15444 38476 15496
rect 38528 15484 38534 15496
rect 38856 15484 38884 15515
rect 45186 15512 45192 15564
rect 45244 15552 45250 15564
rect 45557 15555 45615 15561
rect 45557 15552 45569 15555
rect 45244 15524 45569 15552
rect 45244 15512 45250 15524
rect 45557 15521 45569 15524
rect 45603 15521 45615 15555
rect 45557 15515 45615 15521
rect 40770 15484 40776 15496
rect 38528 15456 40776 15484
rect 38528 15444 38534 15456
rect 40770 15444 40776 15456
rect 40828 15444 40834 15496
rect 40948 15487 41006 15493
rect 40948 15453 40960 15487
rect 40994 15484 41006 15487
rect 41230 15484 41236 15496
rect 40994 15456 41236 15484
rect 40994 15453 41006 15456
rect 40948 15447 41006 15453
rect 41230 15444 41236 15456
rect 41288 15444 41294 15496
rect 45824 15487 45882 15493
rect 45824 15453 45836 15487
rect 45870 15484 45882 15487
rect 46382 15484 46388 15496
rect 45870 15456 46388 15484
rect 45870 15453 45882 15456
rect 45824 15447 45882 15453
rect 46382 15444 46388 15456
rect 46440 15444 46446 15496
rect 47486 15444 47492 15496
rect 47544 15444 47550 15496
rect 47670 15444 47676 15496
rect 47728 15444 47734 15496
rect 47857 15487 47915 15493
rect 47857 15453 47869 15487
rect 47903 15484 47915 15487
rect 47964 15484 47992 15660
rect 51736 15620 51764 15660
rect 51813 15657 51825 15691
rect 51859 15688 51871 15691
rect 51902 15688 51908 15700
rect 51859 15660 51908 15688
rect 51859 15657 51871 15660
rect 51813 15651 51871 15657
rect 51902 15648 51908 15660
rect 51960 15648 51966 15700
rect 55858 15620 55864 15632
rect 50724 15592 51074 15620
rect 51736 15592 55864 15620
rect 47903 15456 47992 15484
rect 47903 15453 47915 15456
rect 47857 15447 47915 15453
rect 48130 15444 48136 15496
rect 48188 15444 48194 15496
rect 50614 15487 50672 15493
rect 50614 15453 50626 15487
rect 50660 15484 50672 15487
rect 50724 15484 50752 15592
rect 51046 15552 51074 15592
rect 55858 15580 55864 15592
rect 55916 15620 55922 15632
rect 56134 15620 56140 15632
rect 55916 15592 56140 15620
rect 55916 15580 55922 15592
rect 56134 15580 56140 15592
rect 56192 15580 56198 15632
rect 51534 15552 51540 15564
rect 51046 15524 51540 15552
rect 51534 15512 51540 15524
rect 51592 15552 51598 15564
rect 51592 15524 57928 15552
rect 51592 15512 51598 15524
rect 50660 15456 50752 15484
rect 50985 15487 51043 15493
rect 50660 15453 50672 15456
rect 50614 15447 50672 15453
rect 50985 15453 50997 15487
rect 51031 15453 51043 15487
rect 50985 15447 51043 15453
rect 33560 15388 33824 15416
rect 33560 15376 33566 15388
rect 37826 15376 37832 15428
rect 37884 15416 37890 15428
rect 38565 15419 38623 15425
rect 38565 15416 38577 15419
rect 37884 15388 38577 15416
rect 37884 15376 37890 15388
rect 38565 15385 38577 15388
rect 38611 15416 38623 15419
rect 38611 15388 39252 15416
rect 38611 15385 38623 15388
rect 38565 15379 38623 15385
rect 28408 15320 28994 15348
rect 29089 15351 29147 15357
rect 28408 15308 28414 15320
rect 29089 15317 29101 15351
rect 29135 15348 29147 15351
rect 29822 15348 29828 15360
rect 29135 15320 29828 15348
rect 29135 15317 29147 15320
rect 29089 15311 29147 15317
rect 29822 15308 29828 15320
rect 29880 15308 29886 15360
rect 29914 15308 29920 15360
rect 29972 15348 29978 15360
rect 30285 15351 30343 15357
rect 30285 15348 30297 15351
rect 29972 15320 30297 15348
rect 29972 15308 29978 15320
rect 30285 15317 30297 15320
rect 30331 15317 30343 15351
rect 30285 15311 30343 15317
rect 31018 15308 31024 15360
rect 31076 15308 31082 15360
rect 31386 15308 31392 15360
rect 31444 15348 31450 15360
rect 31849 15351 31907 15357
rect 31849 15348 31861 15351
rect 31444 15320 31861 15348
rect 31444 15308 31450 15320
rect 31849 15317 31861 15320
rect 31895 15317 31907 15351
rect 31849 15311 31907 15317
rect 32033 15351 32091 15357
rect 32033 15317 32045 15351
rect 32079 15348 32091 15351
rect 32122 15348 32128 15360
rect 32079 15320 32128 15348
rect 32079 15317 32091 15320
rect 32033 15311 32091 15317
rect 32122 15308 32128 15320
rect 32180 15308 32186 15360
rect 38194 15308 38200 15360
rect 38252 15308 38258 15360
rect 38378 15308 38384 15360
rect 38436 15348 38442 15360
rect 38657 15351 38715 15357
rect 38657 15348 38669 15351
rect 38436 15320 38669 15348
rect 38436 15308 38442 15320
rect 38657 15317 38669 15320
rect 38703 15317 38715 15351
rect 39224 15348 39252 15388
rect 39758 15376 39764 15428
rect 39816 15416 39822 15428
rect 43070 15416 43076 15428
rect 39816 15388 43076 15416
rect 39816 15376 39822 15388
rect 43070 15376 43076 15388
rect 43128 15376 43134 15428
rect 43248 15419 43306 15425
rect 43248 15385 43260 15419
rect 43294 15416 43306 15419
rect 43530 15416 43536 15428
rect 43294 15388 43536 15416
rect 43294 15385 43306 15388
rect 43248 15379 43306 15385
rect 43530 15376 43536 15388
rect 43588 15376 43594 15428
rect 46566 15416 46572 15428
rect 43640 15388 46572 15416
rect 43640 15348 43668 15388
rect 46566 15376 46572 15388
rect 46624 15376 46630 15428
rect 47765 15419 47823 15425
rect 47765 15416 47777 15419
rect 46676 15388 47777 15416
rect 39224 15320 43668 15348
rect 38657 15311 38715 15317
rect 44358 15308 44364 15360
rect 44416 15308 44422 15360
rect 44450 15308 44456 15360
rect 44508 15348 44514 15360
rect 46676 15348 46704 15388
rect 47765 15385 47777 15388
rect 47811 15385 47823 15419
rect 47765 15379 47823 15385
rect 47946 15376 47952 15428
rect 48004 15425 48010 15428
rect 48004 15419 48033 15425
rect 48021 15385 48033 15419
rect 51000 15416 51028 15447
rect 51074 15444 51080 15496
rect 51132 15484 51138 15496
rect 51721 15487 51779 15493
rect 51132 15456 51672 15484
rect 51132 15444 51138 15456
rect 48004 15379 48033 15385
rect 48240 15388 51028 15416
rect 48004 15376 48010 15379
rect 44508 15320 46704 15348
rect 44508 15308 44514 15320
rect 46842 15308 46848 15360
rect 46900 15348 46906 15360
rect 48240 15348 48268 15388
rect 51166 15376 51172 15428
rect 51224 15416 51230 15428
rect 51537 15419 51595 15425
rect 51537 15416 51549 15419
rect 51224 15388 51549 15416
rect 51224 15376 51230 15388
rect 51537 15385 51549 15388
rect 51583 15385 51595 15419
rect 51644 15416 51672 15456
rect 51721 15453 51733 15487
rect 51767 15484 51779 15487
rect 52086 15484 52092 15496
rect 51767 15456 52092 15484
rect 51767 15453 51779 15456
rect 51721 15447 51779 15453
rect 52086 15444 52092 15456
rect 52144 15484 52150 15496
rect 54478 15484 54484 15496
rect 52144 15456 54484 15484
rect 52144 15444 52150 15456
rect 54478 15444 54484 15456
rect 54536 15444 54542 15496
rect 57900 15493 57928 15524
rect 57885 15487 57943 15493
rect 57885 15453 57897 15487
rect 57931 15453 57943 15487
rect 57885 15447 57943 15453
rect 51902 15416 51908 15428
rect 51644 15388 51908 15416
rect 51537 15379 51595 15385
rect 51902 15376 51908 15388
rect 51960 15376 51966 15428
rect 58158 15376 58164 15428
rect 58216 15376 58222 15428
rect 46900 15320 48268 15348
rect 46900 15308 46906 15320
rect 48866 15308 48872 15360
rect 48924 15348 48930 15360
rect 49234 15348 49240 15360
rect 48924 15320 49240 15348
rect 48924 15308 48930 15320
rect 49234 15308 49240 15320
rect 49292 15308 49298 15360
rect 50062 15308 50068 15360
rect 50120 15348 50126 15360
rect 50433 15351 50491 15357
rect 50433 15348 50445 15351
rect 50120 15320 50445 15348
rect 50120 15308 50126 15320
rect 50433 15317 50445 15320
rect 50479 15317 50491 15351
rect 50433 15311 50491 15317
rect 50617 15351 50675 15357
rect 50617 15317 50629 15351
rect 50663 15348 50675 15351
rect 51184 15348 51212 15376
rect 50663 15320 51212 15348
rect 50663 15317 50675 15320
rect 50617 15311 50675 15317
rect 1104 15258 58880 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 50294 15258
rect 50346 15206 50358 15258
rect 50410 15206 50422 15258
rect 50474 15206 50486 15258
rect 50538 15206 50550 15258
rect 50602 15206 58880 15258
rect 1104 15184 58880 15206
rect 12342 15104 12348 15156
rect 12400 15144 12406 15156
rect 15105 15147 15163 15153
rect 15105 15144 15117 15147
rect 12400 15116 15117 15144
rect 12400 15104 12406 15116
rect 15105 15113 15117 15116
rect 15151 15113 15163 15147
rect 15105 15107 15163 15113
rect 15746 15104 15752 15156
rect 15804 15144 15810 15156
rect 17402 15144 17408 15156
rect 15804 15116 17408 15144
rect 15804 15104 15810 15116
rect 17402 15104 17408 15116
rect 17460 15104 17466 15156
rect 17604 15116 18000 15144
rect 5442 15036 5448 15088
rect 5500 15076 5506 15088
rect 17604 15076 17632 15116
rect 17862 15076 17868 15088
rect 5500 15048 17632 15076
rect 17696 15048 17868 15076
rect 5500 15036 5506 15048
rect 1581 15011 1639 15017
rect 1581 14977 1593 15011
rect 1627 15008 1639 15011
rect 12434 15008 12440 15020
rect 1627 14980 12440 15008
rect 1627 14977 1639 14980
rect 1581 14971 1639 14977
rect 12434 14968 12440 14980
rect 12492 14968 12498 15020
rect 15289 15011 15347 15017
rect 15289 14977 15301 15011
rect 15335 15008 15347 15011
rect 15746 15008 15752 15020
rect 15335 14980 15752 15008
rect 15335 14977 15347 14980
rect 15289 14971 15347 14977
rect 15746 14968 15752 14980
rect 15804 14968 15810 15020
rect 17696 15017 17724 15048
rect 17862 15036 17868 15048
rect 17920 15036 17926 15088
rect 17972 15076 18000 15116
rect 20346 15104 20352 15156
rect 20404 15144 20410 15156
rect 20441 15147 20499 15153
rect 20441 15144 20453 15147
rect 20404 15116 20453 15144
rect 20404 15104 20410 15116
rect 20441 15113 20453 15116
rect 20487 15113 20499 15147
rect 20441 15107 20499 15113
rect 20806 15104 20812 15156
rect 20864 15144 20870 15156
rect 21450 15144 21456 15156
rect 20864 15116 21456 15144
rect 20864 15104 20870 15116
rect 21450 15104 21456 15116
rect 21508 15144 21514 15156
rect 23385 15147 23443 15153
rect 23385 15144 23397 15147
rect 21508 15116 23397 15144
rect 21508 15104 21514 15116
rect 23385 15113 23397 15116
rect 23431 15113 23443 15147
rect 23385 15107 23443 15113
rect 23934 15104 23940 15156
rect 23992 15144 23998 15156
rect 24118 15144 24124 15156
rect 23992 15116 24124 15144
rect 23992 15104 23998 15116
rect 24118 15104 24124 15116
rect 24176 15104 24182 15156
rect 27890 15144 27896 15156
rect 24504 15116 27896 15144
rect 22281 15079 22339 15085
rect 17972 15048 22094 15076
rect 17681 15011 17739 15017
rect 17681 14977 17693 15011
rect 17727 14977 17739 15011
rect 17681 14971 17739 14977
rect 17773 15011 17831 15017
rect 17773 14977 17785 15011
rect 17819 14977 17831 15011
rect 17773 14971 17831 14977
rect 18417 15011 18475 15017
rect 18417 14977 18429 15011
rect 18463 15008 18475 15011
rect 18598 15008 18604 15020
rect 18463 14980 18604 15008
rect 18463 14977 18475 14980
rect 18417 14971 18475 14977
rect 934 14900 940 14952
rect 992 14940 998 14952
rect 1765 14943 1823 14949
rect 1765 14940 1777 14943
rect 992 14912 1777 14940
rect 992 14900 998 14912
rect 1765 14909 1777 14912
rect 1811 14909 1823 14943
rect 1765 14903 1823 14909
rect 15381 14943 15439 14949
rect 15381 14909 15393 14943
rect 15427 14909 15439 14943
rect 15381 14903 15439 14909
rect 15396 14872 15424 14903
rect 15470 14900 15476 14952
rect 15528 14900 15534 14952
rect 15562 14900 15568 14952
rect 15620 14900 15626 14952
rect 17788 14940 17816 14971
rect 18598 14968 18604 14980
rect 18656 14968 18662 15020
rect 20254 14968 20260 15020
rect 20312 14968 20318 15020
rect 20990 14968 20996 15020
rect 21048 14968 21054 15020
rect 22066 15008 22094 15048
rect 22281 15045 22293 15079
rect 22327 15076 22339 15079
rect 22646 15076 22652 15088
rect 22327 15048 22652 15076
rect 22327 15045 22339 15048
rect 22281 15039 22339 15045
rect 22646 15036 22652 15048
rect 22704 15036 22710 15088
rect 22738 15036 22744 15088
rect 22796 15036 22802 15088
rect 24504 15076 24532 15116
rect 27890 15104 27896 15116
rect 27948 15104 27954 15156
rect 28534 15104 28540 15156
rect 28592 15144 28598 15156
rect 28629 15147 28687 15153
rect 28629 15144 28641 15147
rect 28592 15116 28641 15144
rect 28592 15104 28598 15116
rect 28629 15113 28641 15116
rect 28675 15113 28687 15147
rect 28629 15107 28687 15113
rect 30098 15104 30104 15156
rect 30156 15104 30162 15156
rect 32398 15144 32404 15156
rect 30208 15116 32404 15144
rect 22848 15048 24532 15076
rect 22848 15008 22876 15048
rect 24578 15036 24584 15088
rect 24636 15076 24642 15088
rect 30208 15076 30236 15116
rect 32398 15104 32404 15116
rect 32456 15104 32462 15156
rect 32493 15147 32551 15153
rect 32493 15113 32505 15147
rect 32539 15113 32551 15147
rect 32493 15107 32551 15113
rect 33888 15116 42932 15144
rect 32508 15076 32536 15107
rect 33888 15085 33916 15116
rect 24636 15048 30236 15076
rect 31128 15048 32536 15076
rect 33873 15079 33931 15085
rect 24636 15036 24642 15048
rect 22066 14980 22876 15008
rect 23198 14968 23204 15020
rect 23256 14968 23262 15020
rect 23934 14968 23940 15020
rect 23992 15008 23998 15020
rect 24857 15011 24915 15017
rect 24857 15008 24869 15011
rect 23992 14980 24869 15008
rect 23992 14968 23998 14980
rect 24857 14977 24869 14980
rect 24903 15008 24915 15011
rect 25406 15008 25412 15020
rect 24903 14980 25412 15008
rect 24903 14977 24915 14980
rect 24857 14971 24915 14977
rect 25406 14968 25412 14980
rect 25464 14968 25470 15020
rect 25866 14968 25872 15020
rect 25924 14968 25930 15020
rect 26145 15011 26203 15017
rect 26145 14977 26157 15011
rect 26191 14977 26203 15011
rect 26145 14971 26203 14977
rect 17788 14912 18644 14940
rect 18616 14881 18644 14912
rect 21726 14900 21732 14952
rect 21784 14940 21790 14952
rect 22002 14940 22008 14952
rect 21784 14912 22008 14940
rect 21784 14900 21790 14912
rect 22002 14900 22008 14912
rect 22060 14900 22066 14952
rect 22370 14900 22376 14952
rect 22428 14900 22434 14952
rect 22465 14943 22523 14949
rect 22465 14909 22477 14943
rect 22511 14940 22523 14943
rect 25130 14940 25136 14952
rect 22511 14912 25136 14940
rect 22511 14909 22523 14912
rect 22465 14903 22523 14909
rect 25130 14900 25136 14912
rect 25188 14900 25194 14952
rect 25225 14943 25283 14949
rect 25225 14909 25237 14943
rect 25271 14909 25283 14943
rect 25225 14903 25283 14909
rect 18601 14875 18659 14881
rect 15396 14844 18552 14872
rect 17494 14764 17500 14816
rect 17552 14804 17558 14816
rect 17957 14807 18015 14813
rect 17957 14804 17969 14807
rect 17552 14776 17969 14804
rect 17552 14764 17558 14776
rect 17957 14773 17969 14776
rect 18003 14773 18015 14807
rect 18524 14804 18552 14844
rect 18601 14841 18613 14875
rect 18647 14841 18659 14875
rect 24670 14872 24676 14884
rect 18601 14835 18659 14841
rect 18708 14844 24676 14872
rect 18708 14804 18736 14844
rect 24670 14832 24676 14844
rect 24728 14832 24734 14884
rect 25240 14872 25268 14903
rect 25314 14900 25320 14952
rect 25372 14900 25378 14952
rect 25682 14900 25688 14952
rect 25740 14940 25746 14952
rect 26160 14940 26188 14971
rect 28442 14968 28448 15020
rect 28500 14968 28506 15020
rect 29365 15011 29423 15017
rect 29365 14977 29377 15011
rect 29411 14977 29423 15011
rect 29365 14971 29423 14977
rect 25740 14912 26188 14940
rect 25740 14900 25746 14912
rect 26510 14900 26516 14952
rect 26568 14900 26574 14952
rect 28902 14900 28908 14952
rect 28960 14940 28966 14952
rect 28960 14900 28994 14940
rect 25866 14872 25872 14884
rect 25240 14844 25872 14872
rect 25866 14832 25872 14844
rect 25924 14832 25930 14884
rect 25961 14875 26019 14881
rect 25961 14841 25973 14875
rect 26007 14872 26019 14875
rect 27062 14872 27068 14884
rect 26007 14844 27068 14872
rect 26007 14841 26019 14844
rect 25961 14835 26019 14841
rect 18524 14776 18736 14804
rect 17957 14767 18015 14773
rect 21082 14764 21088 14816
rect 21140 14804 21146 14816
rect 21177 14807 21235 14813
rect 21177 14804 21189 14807
rect 21140 14776 21189 14804
rect 21140 14764 21146 14776
rect 21177 14773 21189 14776
rect 21223 14773 21235 14807
rect 21177 14767 21235 14773
rect 22646 14764 22652 14816
rect 22704 14804 22710 14816
rect 23198 14804 23204 14816
rect 22704 14776 23204 14804
rect 22704 14764 22710 14776
rect 23198 14764 23204 14776
rect 23256 14764 23262 14816
rect 24118 14764 24124 14816
rect 24176 14804 24182 14816
rect 24486 14804 24492 14816
rect 24176 14776 24492 14804
rect 24176 14764 24182 14776
rect 24486 14764 24492 14776
rect 24544 14804 24550 14816
rect 25976 14804 26004 14835
rect 27062 14832 27068 14844
rect 27120 14832 27126 14884
rect 24544 14776 26004 14804
rect 28966 14804 28994 14900
rect 29380 14872 29408 14971
rect 29914 14968 29920 15020
rect 29972 14968 29978 15020
rect 31128 15017 31156 15048
rect 33873 15045 33885 15079
rect 33919 15045 33931 15079
rect 33873 15039 33931 15045
rect 33965 15079 34023 15085
rect 33965 15045 33977 15079
rect 34011 15076 34023 15079
rect 36354 15076 36360 15088
rect 34011 15048 36360 15076
rect 34011 15045 34023 15048
rect 33965 15039 34023 15045
rect 31113 15011 31171 15017
rect 31113 14977 31125 15011
rect 31159 14977 31171 15011
rect 31113 14971 31171 14977
rect 31754 14968 31760 15020
rect 31812 15008 31818 15020
rect 32309 15011 32367 15017
rect 32309 15008 32321 15011
rect 31812 14980 32321 15008
rect 31812 14968 31818 14980
rect 32309 14977 32321 14980
rect 32355 14977 32367 15011
rect 32309 14971 32367 14977
rect 32398 14968 32404 15020
rect 32456 15008 32462 15020
rect 32456 14980 32996 15008
rect 32456 14968 32462 14980
rect 32968 14940 32996 14980
rect 33594 14968 33600 15020
rect 33652 14968 33658 15020
rect 33686 14968 33692 15020
rect 33744 15008 33750 15020
rect 33980 15008 34008 15039
rect 36354 15036 36360 15048
rect 36412 15036 36418 15088
rect 38102 15076 38108 15088
rect 37660 15048 38108 15076
rect 37660 15020 37688 15048
rect 38102 15036 38108 15048
rect 38160 15036 38166 15088
rect 42794 15076 42800 15088
rect 39960 15048 42800 15076
rect 33744 14980 34008 15008
rect 33744 14968 33750 14980
rect 34422 14968 34428 15020
rect 34480 14968 34486 15020
rect 37642 14968 37648 15020
rect 37700 14968 37706 15020
rect 37912 15011 37970 15017
rect 37912 14977 37924 15011
rect 37958 15008 37970 15011
rect 38194 15008 38200 15020
rect 37958 14980 38200 15008
rect 37958 14977 37970 14980
rect 37912 14971 37970 14977
rect 38194 14968 38200 14980
rect 38252 14968 38258 15020
rect 39960 15017 39988 15048
rect 42794 15036 42800 15048
rect 42852 15036 42858 15088
rect 42904 15076 42932 15116
rect 43530 15104 43536 15156
rect 43588 15104 43594 15156
rect 43901 15147 43959 15153
rect 43901 15113 43913 15147
rect 43947 15144 43959 15147
rect 44818 15144 44824 15156
rect 43947 15116 44824 15144
rect 43947 15113 43959 15116
rect 43901 15107 43959 15113
rect 44818 15104 44824 15116
rect 44876 15104 44882 15156
rect 44910 15104 44916 15156
rect 44968 15144 44974 15156
rect 44968 15116 45554 15144
rect 44968 15104 44974 15116
rect 44450 15076 44456 15088
rect 42904 15048 44456 15076
rect 44450 15036 44456 15048
rect 44508 15036 44514 15088
rect 44726 15036 44732 15088
rect 44784 15076 44790 15088
rect 45189 15079 45247 15085
rect 45189 15076 45201 15079
rect 44784 15048 45201 15076
rect 44784 15036 44790 15048
rect 39945 15011 40003 15017
rect 39945 14977 39957 15011
rect 39991 14977 40003 15011
rect 39945 14971 40003 14977
rect 40212 15011 40270 15017
rect 40212 14977 40224 15011
rect 40258 15008 40270 15011
rect 40494 15008 40500 15020
rect 40258 14980 40500 15008
rect 40258 14977 40270 14980
rect 40212 14971 40270 14977
rect 40494 14968 40500 14980
rect 40552 14968 40558 15020
rect 44358 15008 44364 15020
rect 44008 14980 44364 15008
rect 33781 14943 33839 14949
rect 33781 14940 33793 14943
rect 32968 14912 33793 14940
rect 33781 14909 33793 14912
rect 33827 14909 33839 14943
rect 33781 14903 33839 14909
rect 31297 14875 31355 14881
rect 31297 14872 31309 14875
rect 29380 14844 31309 14872
rect 31297 14841 31309 14844
rect 31343 14841 31355 14875
rect 31297 14835 31355 14841
rect 29365 14807 29423 14813
rect 29365 14804 29377 14807
rect 28966 14776 29377 14804
rect 24544 14764 24550 14776
rect 29365 14773 29377 14776
rect 29411 14804 29423 14807
rect 29546 14804 29552 14816
rect 29411 14776 29552 14804
rect 29411 14773 29423 14776
rect 29365 14767 29423 14773
rect 29546 14764 29552 14776
rect 29604 14764 29610 14816
rect 29638 14764 29644 14816
rect 29696 14804 29702 14816
rect 30834 14804 30840 14816
rect 29696 14776 30840 14804
rect 29696 14764 29702 14776
rect 30834 14764 30840 14776
rect 30892 14764 30898 14816
rect 31312 14804 31340 14835
rect 31386 14832 31392 14884
rect 31444 14872 31450 14884
rect 33796 14872 33824 14903
rect 43530 14900 43536 14952
rect 43588 14940 43594 14952
rect 44008 14949 44036 14980
rect 44358 14968 44364 14980
rect 44416 14968 44422 15020
rect 43993 14943 44051 14949
rect 43993 14940 44005 14943
rect 43588 14912 44005 14940
rect 43588 14900 43594 14912
rect 43993 14909 44005 14912
rect 44039 14909 44051 14943
rect 43993 14903 44051 14909
rect 44082 14900 44088 14952
rect 44140 14900 44146 14952
rect 44836 14940 44864 15048
rect 45189 15045 45201 15048
rect 45235 15045 45247 15079
rect 45526 15076 45554 15116
rect 48038 15104 48044 15156
rect 48096 15144 48102 15156
rect 48133 15147 48191 15153
rect 48133 15144 48145 15147
rect 48096 15116 48145 15144
rect 48096 15104 48102 15116
rect 48133 15113 48145 15116
rect 48179 15113 48191 15147
rect 48133 15107 48191 15113
rect 50249 15147 50307 15153
rect 50249 15113 50261 15147
rect 50295 15144 50307 15147
rect 50614 15144 50620 15156
rect 50295 15116 50620 15144
rect 50295 15113 50307 15116
rect 50249 15107 50307 15113
rect 50614 15104 50620 15116
rect 50672 15104 50678 15156
rect 49878 15076 49884 15088
rect 45526 15048 49884 15076
rect 45189 15039 45247 15045
rect 49878 15036 49884 15048
rect 49936 15036 49942 15088
rect 50982 15036 50988 15088
rect 51040 15076 51046 15088
rect 51077 15079 51135 15085
rect 51077 15076 51089 15079
rect 51040 15048 51089 15076
rect 51040 15036 51046 15048
rect 51077 15045 51089 15048
rect 51123 15076 51135 15079
rect 54662 15076 54668 15088
rect 51123 15048 54668 15076
rect 51123 15045 51135 15048
rect 51077 15039 51135 15045
rect 54662 15036 54668 15048
rect 54720 15076 54726 15088
rect 54720 15048 54800 15076
rect 54720 15036 54726 15048
rect 44913 15011 44971 15017
rect 44913 14977 44925 15011
rect 44959 15008 44971 15011
rect 45922 15008 45928 15020
rect 44959 14980 45928 15008
rect 44959 14977 44971 14980
rect 44913 14971 44971 14977
rect 45922 14968 45928 14980
rect 45980 14968 45986 15020
rect 47486 14968 47492 15020
rect 47544 15008 47550 15020
rect 47949 15011 48007 15017
rect 47949 15008 47961 15011
rect 47544 14980 47961 15008
rect 47544 14968 47550 14980
rect 47949 14977 47961 14980
rect 47995 14977 48007 15011
rect 47949 14971 48007 14977
rect 50062 14968 50068 15020
rect 50120 15008 50126 15020
rect 50157 15011 50215 15017
rect 50157 15008 50169 15011
rect 50120 14980 50169 15008
rect 50120 14968 50126 14980
rect 50157 14977 50169 14980
rect 50203 14977 50215 15011
rect 50157 14971 50215 14977
rect 50341 15011 50399 15017
rect 50341 14977 50353 15011
rect 50387 14977 50399 15011
rect 50341 14971 50399 14977
rect 50801 15011 50859 15017
rect 50801 14977 50813 15011
rect 50847 15008 50859 15011
rect 50890 15008 50896 15020
rect 50847 14980 50896 15008
rect 50847 14977 50859 14980
rect 50801 14971 50859 14977
rect 47765 14943 47823 14949
rect 47765 14940 47777 14943
rect 44836 14912 47777 14940
rect 47765 14909 47777 14912
rect 47811 14909 47823 14943
rect 47765 14903 47823 14909
rect 33962 14872 33968 14884
rect 31444 14844 32628 14872
rect 33796 14844 33968 14872
rect 31444 14832 31450 14844
rect 31662 14804 31668 14816
rect 31312 14776 31668 14804
rect 31662 14764 31668 14776
rect 31720 14764 31726 14816
rect 32600 14804 32628 14844
rect 33962 14832 33968 14844
rect 34020 14832 34026 14884
rect 49786 14832 49792 14884
rect 49844 14872 49850 14884
rect 50356 14872 50384 14971
rect 50890 14968 50896 14980
rect 50948 14968 50954 15020
rect 54478 14968 54484 15020
rect 54536 14968 54542 15020
rect 54772 15017 54800 15048
rect 54938 15036 54944 15088
rect 54996 15036 55002 15088
rect 54757 15011 54815 15017
rect 54757 14977 54769 15011
rect 54803 14977 54815 15011
rect 54757 14971 54815 14977
rect 58066 14968 58072 15020
rect 58124 14968 58130 15020
rect 51994 14872 52000 14884
rect 49844 14844 52000 14872
rect 49844 14832 49850 14844
rect 51994 14832 52000 14844
rect 52052 14872 52058 14884
rect 56042 14872 56048 14884
rect 52052 14844 56048 14872
rect 52052 14832 52058 14844
rect 56042 14832 56048 14844
rect 56100 14832 56106 14884
rect 34609 14807 34667 14813
rect 34609 14804 34621 14807
rect 32600 14776 34621 14804
rect 34609 14773 34621 14776
rect 34655 14773 34667 14807
rect 34609 14767 34667 14773
rect 34698 14764 34704 14816
rect 34756 14804 34762 14816
rect 38378 14804 38384 14816
rect 34756 14776 38384 14804
rect 34756 14764 34762 14776
rect 38378 14764 38384 14776
rect 38436 14804 38442 14816
rect 39025 14807 39083 14813
rect 39025 14804 39037 14807
rect 38436 14776 39037 14804
rect 38436 14764 38442 14776
rect 39025 14773 39037 14776
rect 39071 14773 39083 14807
rect 39025 14767 39083 14773
rect 39942 14764 39948 14816
rect 40000 14804 40006 14816
rect 40954 14804 40960 14816
rect 40000 14776 40960 14804
rect 40000 14764 40006 14776
rect 40954 14764 40960 14776
rect 41012 14804 41018 14816
rect 41325 14807 41383 14813
rect 41325 14804 41337 14807
rect 41012 14776 41337 14804
rect 41012 14764 41018 14776
rect 41325 14773 41337 14776
rect 41371 14773 41383 14807
rect 41325 14767 41383 14773
rect 58250 14764 58256 14816
rect 58308 14764 58314 14816
rect 1104 14714 58880 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 58880 14714
rect 1104 14640 58880 14662
rect 15654 14560 15660 14612
rect 15712 14600 15718 14612
rect 16301 14603 16359 14609
rect 16301 14600 16313 14603
rect 15712 14572 16313 14600
rect 15712 14560 15718 14572
rect 16301 14569 16313 14572
rect 16347 14569 16359 14603
rect 24578 14600 24584 14612
rect 16301 14563 16359 14569
rect 16408 14572 24584 14600
rect 13354 14492 13360 14544
rect 13412 14532 13418 14544
rect 16117 14535 16175 14541
rect 16117 14532 16129 14535
rect 13412 14504 16129 14532
rect 13412 14492 13418 14504
rect 16117 14501 16129 14504
rect 16163 14501 16175 14535
rect 16117 14495 16175 14501
rect 15102 14424 15108 14476
rect 15160 14464 15166 14476
rect 16408 14464 16436 14572
rect 24578 14560 24584 14572
rect 24636 14560 24642 14612
rect 24946 14560 24952 14612
rect 25004 14600 25010 14612
rect 25225 14603 25283 14609
rect 25225 14600 25237 14603
rect 25004 14572 25237 14600
rect 25004 14560 25010 14572
rect 25225 14569 25237 14572
rect 25271 14569 25283 14603
rect 25225 14563 25283 14569
rect 28442 14560 28448 14612
rect 28500 14600 28506 14612
rect 29089 14603 29147 14609
rect 29089 14600 29101 14603
rect 28500 14572 29101 14600
rect 28500 14560 28506 14572
rect 29089 14569 29101 14572
rect 29135 14600 29147 14603
rect 30926 14600 30932 14612
rect 29135 14572 30932 14600
rect 29135 14569 29147 14572
rect 29089 14563 29147 14569
rect 30926 14560 30932 14572
rect 30984 14560 30990 14612
rect 31110 14560 31116 14612
rect 31168 14560 31174 14612
rect 31754 14560 31760 14612
rect 31812 14560 31818 14612
rect 32122 14560 32128 14612
rect 32180 14600 32186 14612
rect 32309 14603 32367 14609
rect 32309 14600 32321 14603
rect 32180 14572 32321 14600
rect 32180 14560 32186 14572
rect 32309 14569 32321 14572
rect 32355 14569 32367 14603
rect 32309 14563 32367 14569
rect 32674 14560 32680 14612
rect 32732 14600 32738 14612
rect 33505 14603 33563 14609
rect 33505 14600 33517 14603
rect 32732 14572 33517 14600
rect 32732 14560 32738 14572
rect 33505 14569 33517 14572
rect 33551 14600 33563 14603
rect 33686 14600 33692 14612
rect 33551 14572 33692 14600
rect 33551 14569 33563 14572
rect 33505 14563 33563 14569
rect 33686 14560 33692 14572
rect 33744 14560 33750 14612
rect 33778 14560 33784 14612
rect 33836 14600 33842 14612
rect 35713 14603 35771 14609
rect 35713 14600 35725 14603
rect 33836 14572 35725 14600
rect 33836 14560 33842 14572
rect 35713 14569 35725 14572
rect 35759 14569 35771 14603
rect 35713 14563 35771 14569
rect 40494 14560 40500 14612
rect 40552 14560 40558 14612
rect 44910 14600 44916 14612
rect 40604 14572 44916 14600
rect 17678 14492 17684 14544
rect 17736 14492 17742 14544
rect 18782 14492 18788 14544
rect 18840 14532 18846 14544
rect 20073 14535 20131 14541
rect 20073 14532 20085 14535
rect 18840 14504 20085 14532
rect 18840 14492 18846 14504
rect 20073 14501 20085 14504
rect 20119 14501 20131 14535
rect 20073 14495 20131 14501
rect 21266 14492 21272 14544
rect 21324 14492 21330 14544
rect 21634 14492 21640 14544
rect 21692 14532 21698 14544
rect 29638 14532 29644 14544
rect 21692 14504 29644 14532
rect 21692 14492 21698 14504
rect 29638 14492 29644 14504
rect 29696 14492 29702 14544
rect 30834 14492 30840 14544
rect 30892 14532 30898 14544
rect 33045 14535 33103 14541
rect 30892 14504 32444 14532
rect 30892 14492 30898 14504
rect 17310 14464 17316 14476
rect 15160 14436 16436 14464
rect 16546 14436 17316 14464
rect 15160 14424 15166 14436
rect 1581 14399 1639 14405
rect 1581 14365 1593 14399
rect 1627 14396 1639 14399
rect 5442 14396 5448 14408
rect 1627 14368 5448 14396
rect 1627 14365 1639 14368
rect 1581 14359 1639 14365
rect 5442 14356 5448 14368
rect 5500 14356 5506 14408
rect 15010 14356 15016 14408
rect 15068 14356 15074 14408
rect 16546 14396 16574 14436
rect 17310 14424 17316 14436
rect 17368 14424 17374 14476
rect 17402 14424 17408 14476
rect 17460 14464 17466 14476
rect 22278 14464 22284 14476
rect 17460 14436 22284 14464
rect 17460 14424 17466 14436
rect 22278 14424 22284 14436
rect 22336 14424 22342 14476
rect 22370 14424 22376 14476
rect 22428 14464 22434 14476
rect 25406 14464 25412 14476
rect 22428 14436 25412 14464
rect 22428 14424 22434 14436
rect 15212 14368 16574 14396
rect 934 14288 940 14340
rect 992 14328 998 14340
rect 1857 14331 1915 14337
rect 1857 14328 1869 14331
rect 992 14300 1869 14328
rect 992 14288 998 14300
rect 1857 14297 1869 14300
rect 1903 14297 1915 14331
rect 1857 14291 1915 14297
rect 12526 14288 12532 14340
rect 12584 14328 12590 14340
rect 14829 14331 14887 14337
rect 14829 14328 14841 14331
rect 12584 14300 14841 14328
rect 12584 14288 12590 14300
rect 14829 14297 14841 14300
rect 14875 14328 14887 14331
rect 15212 14328 15240 14368
rect 17494 14356 17500 14408
rect 17552 14356 17558 14408
rect 20257 14399 20315 14405
rect 20257 14365 20269 14399
rect 20303 14396 20315 14399
rect 20303 14368 21036 14396
rect 20303 14365 20315 14368
rect 20257 14359 20315 14365
rect 14875 14300 15240 14328
rect 14875 14297 14887 14300
rect 14829 14291 14887 14297
rect 15838 14288 15844 14340
rect 15896 14288 15902 14340
rect 20438 14288 20444 14340
rect 20496 14337 20502 14340
rect 20496 14331 20539 14337
rect 20527 14297 20539 14331
rect 20496 14291 20539 14297
rect 20496 14288 20502 14291
rect 20622 14288 20628 14340
rect 20680 14288 20686 14340
rect 21008 14328 21036 14368
rect 21082 14356 21088 14408
rect 21140 14356 21146 14408
rect 23676 14405 23704 14436
rect 25406 14424 25412 14436
rect 25464 14424 25470 14476
rect 26878 14424 26884 14476
rect 26936 14424 26942 14476
rect 28276 14436 29868 14464
rect 23661 14399 23719 14405
rect 23661 14365 23673 14399
rect 23707 14365 23719 14399
rect 23661 14359 23719 14365
rect 25038 14356 25044 14408
rect 25096 14356 25102 14408
rect 26510 14396 26516 14408
rect 25148 14368 26516 14396
rect 25148 14328 25176 14368
rect 26510 14356 26516 14368
rect 26568 14356 26574 14408
rect 26602 14356 26608 14408
rect 26660 14396 26666 14408
rect 28276 14405 28304 14436
rect 26697 14399 26755 14405
rect 26697 14396 26709 14399
rect 26660 14368 26709 14396
rect 26660 14356 26666 14368
rect 26697 14365 26709 14368
rect 26743 14365 26755 14399
rect 26697 14359 26755 14365
rect 28261 14399 28319 14405
rect 28261 14365 28273 14399
rect 28307 14365 28319 14399
rect 28261 14359 28319 14365
rect 28445 14399 28503 14405
rect 28445 14365 28457 14399
rect 28491 14396 28503 14399
rect 28810 14396 28816 14408
rect 28491 14368 28816 14396
rect 28491 14365 28503 14368
rect 28445 14359 28503 14365
rect 28810 14356 28816 14368
rect 28868 14356 28874 14408
rect 28905 14399 28963 14405
rect 28905 14365 28917 14399
rect 28951 14396 28963 14399
rect 29454 14396 29460 14408
rect 28951 14368 29460 14396
rect 28951 14365 28963 14368
rect 28905 14359 28963 14365
rect 29454 14356 29460 14368
rect 29512 14356 29518 14408
rect 29733 14399 29791 14405
rect 29733 14365 29745 14399
rect 29779 14365 29791 14399
rect 29840 14396 29868 14436
rect 29840 14368 30144 14396
rect 29733 14359 29791 14365
rect 21008 14300 25176 14328
rect 25222 14288 25228 14340
rect 25280 14328 25286 14340
rect 27706 14328 27712 14340
rect 25280 14300 27712 14328
rect 25280 14288 25286 14300
rect 27706 14288 27712 14300
rect 27764 14288 27770 14340
rect 28353 14331 28411 14337
rect 28353 14297 28365 14331
rect 28399 14328 28411 14331
rect 29546 14328 29552 14340
rect 28399 14300 29552 14328
rect 28399 14297 28411 14300
rect 28353 14291 28411 14297
rect 29546 14288 29552 14300
rect 29604 14288 29610 14340
rect 29748 14328 29776 14359
rect 30116 14340 30144 14368
rect 31110 14356 31116 14408
rect 31168 14396 31174 14408
rect 31573 14399 31631 14405
rect 31573 14396 31585 14399
rect 31168 14368 31585 14396
rect 31168 14356 31174 14368
rect 31573 14365 31585 14368
rect 31619 14365 31631 14399
rect 32309 14399 32367 14405
rect 32309 14396 32321 14399
rect 31573 14359 31631 14365
rect 31726 14368 32321 14396
rect 29822 14328 29828 14340
rect 29748 14300 29828 14328
rect 29822 14288 29828 14300
rect 29880 14288 29886 14340
rect 29978 14331 30036 14337
rect 29978 14297 29990 14331
rect 30024 14328 30036 14331
rect 30024 14297 30052 14328
rect 29978 14291 30052 14297
rect 14458 14220 14464 14272
rect 14516 14260 14522 14272
rect 15102 14260 15108 14272
rect 14516 14232 15108 14260
rect 14516 14220 14522 14232
rect 15102 14220 15108 14232
rect 15160 14220 15166 14272
rect 20349 14263 20407 14269
rect 20349 14229 20361 14263
rect 20395 14260 20407 14263
rect 23382 14260 23388 14272
rect 20395 14232 23388 14260
rect 20395 14229 20407 14232
rect 20349 14223 20407 14229
rect 23382 14220 23388 14232
rect 23440 14220 23446 14272
rect 23658 14220 23664 14272
rect 23716 14260 23722 14272
rect 23845 14263 23903 14269
rect 23845 14260 23857 14263
rect 23716 14232 23857 14260
rect 23716 14220 23722 14232
rect 23845 14229 23857 14232
rect 23891 14229 23903 14263
rect 23845 14223 23903 14229
rect 26234 14220 26240 14272
rect 26292 14220 26298 14272
rect 26605 14263 26663 14269
rect 26605 14229 26617 14263
rect 26651 14260 26663 14263
rect 29086 14260 29092 14272
rect 26651 14232 29092 14260
rect 26651 14229 26663 14232
rect 26605 14223 26663 14229
rect 29086 14220 29092 14232
rect 29144 14220 29150 14272
rect 29178 14220 29184 14272
rect 29236 14260 29242 14272
rect 30024 14260 30052 14291
rect 30098 14288 30104 14340
rect 30156 14288 30162 14340
rect 30190 14288 30196 14340
rect 30248 14328 30254 14340
rect 31726 14328 31754 14368
rect 32309 14365 32321 14368
rect 32355 14365 32367 14399
rect 32309 14359 32367 14365
rect 30248 14300 31754 14328
rect 30248 14288 30254 14300
rect 29236 14232 30052 14260
rect 29236 14220 29242 14232
rect 31110 14220 31116 14272
rect 31168 14260 31174 14272
rect 31294 14260 31300 14272
rect 31168 14232 31300 14260
rect 31168 14220 31174 14232
rect 31294 14220 31300 14232
rect 31352 14220 31358 14272
rect 32416 14260 32444 14504
rect 33045 14501 33057 14535
rect 33091 14532 33103 14535
rect 34241 14535 34299 14541
rect 33091 14504 34192 14532
rect 33091 14501 33103 14504
rect 33045 14495 33103 14501
rect 34164 14464 34192 14504
rect 34241 14501 34253 14535
rect 34287 14532 34299 14535
rect 34422 14532 34428 14544
rect 34287 14504 34428 14532
rect 34287 14501 34299 14504
rect 34241 14495 34299 14501
rect 34422 14492 34428 14504
rect 34480 14532 34486 14544
rect 34480 14504 35664 14532
rect 34480 14492 34486 14504
rect 32508 14436 33640 14464
rect 34164 14436 35572 14464
rect 32508 14405 32536 14436
rect 32493 14399 32551 14405
rect 32493 14365 32505 14399
rect 32539 14365 32551 14399
rect 32493 14359 32551 14365
rect 33226 14356 33232 14408
rect 33284 14356 33290 14408
rect 33612 14405 33640 14436
rect 33321 14399 33379 14405
rect 33321 14365 33333 14399
rect 33367 14365 33379 14399
rect 33321 14359 33379 14365
rect 33597 14399 33655 14405
rect 33597 14365 33609 14399
rect 33643 14396 33655 14399
rect 33778 14396 33784 14408
rect 33643 14368 33784 14396
rect 33643 14365 33655 14368
rect 33597 14359 33655 14365
rect 32582 14288 32588 14340
rect 32640 14328 32646 14340
rect 33336 14328 33364 14359
rect 33778 14356 33784 14368
rect 33836 14356 33842 14408
rect 34057 14399 34115 14405
rect 34057 14365 34069 14399
rect 34103 14365 34115 14399
rect 34057 14359 34115 14365
rect 32640 14300 33364 14328
rect 34072 14328 34100 14359
rect 34514 14356 34520 14408
rect 34572 14396 34578 14408
rect 34885 14399 34943 14405
rect 34885 14396 34897 14399
rect 34572 14368 34897 14396
rect 34572 14356 34578 14368
rect 34885 14365 34897 14368
rect 34931 14396 34943 14399
rect 35342 14396 35348 14408
rect 34931 14368 35348 14396
rect 34931 14365 34943 14368
rect 34885 14359 34943 14365
rect 35342 14356 35348 14368
rect 35400 14356 35406 14408
rect 34072 14300 35112 14328
rect 32640 14288 32646 14300
rect 34054 14260 34060 14272
rect 32416 14232 34060 14260
rect 34054 14220 34060 14232
rect 34112 14220 34118 14272
rect 35084 14269 35112 14300
rect 35069 14263 35127 14269
rect 35069 14229 35081 14263
rect 35115 14229 35127 14263
rect 35544 14260 35572 14436
rect 35636 14405 35664 14504
rect 35802 14492 35808 14544
rect 35860 14532 35866 14544
rect 40604 14532 40632 14572
rect 44910 14560 44916 14572
rect 44968 14560 44974 14612
rect 59538 14600 59544 14612
rect 45526 14572 59544 14600
rect 45526 14532 45554 14572
rect 59538 14560 59544 14572
rect 59596 14560 59602 14612
rect 35860 14504 40632 14532
rect 40880 14504 45554 14532
rect 35860 14492 35866 14504
rect 35621 14399 35679 14405
rect 35621 14365 35633 14399
rect 35667 14365 35679 14399
rect 35621 14359 35679 14365
rect 40880 14337 40908 14504
rect 40954 14424 40960 14476
rect 41012 14424 41018 14476
rect 41138 14424 41144 14476
rect 41196 14424 41202 14476
rect 45278 14424 45284 14476
rect 45336 14464 45342 14476
rect 48406 14464 48412 14476
rect 45336 14436 48412 14464
rect 45336 14424 45342 14436
rect 48406 14424 48412 14436
rect 48464 14424 48470 14476
rect 49605 14399 49663 14405
rect 49605 14365 49617 14399
rect 49651 14365 49663 14399
rect 49605 14359 49663 14365
rect 40221 14331 40279 14337
rect 40221 14297 40233 14331
rect 40267 14328 40279 14331
rect 40865 14331 40923 14337
rect 40865 14328 40877 14331
rect 40267 14300 40877 14328
rect 40267 14297 40279 14300
rect 40221 14291 40279 14297
rect 40865 14297 40877 14300
rect 40911 14297 40923 14331
rect 46842 14328 46848 14340
rect 40865 14291 40923 14297
rect 41386 14300 46848 14328
rect 41386 14260 41414 14300
rect 46842 14288 46848 14300
rect 46900 14288 46906 14340
rect 35544 14232 41414 14260
rect 49620 14260 49648 14359
rect 49786 14356 49792 14408
rect 49844 14356 49850 14408
rect 50154 14356 50160 14408
rect 50212 14396 50218 14408
rect 50341 14399 50399 14405
rect 50341 14396 50353 14399
rect 50212 14368 50353 14396
rect 50212 14356 50218 14368
rect 50341 14365 50353 14368
rect 50387 14365 50399 14399
rect 50341 14359 50399 14365
rect 57885 14399 57943 14405
rect 57885 14365 57897 14399
rect 57931 14365 57943 14399
rect 57885 14359 57943 14365
rect 49697 14331 49755 14337
rect 49697 14297 49709 14331
rect 49743 14328 49755 14331
rect 50586 14331 50644 14337
rect 50586 14328 50598 14331
rect 49743 14300 50598 14328
rect 49743 14297 49755 14300
rect 49697 14291 49755 14297
rect 50586 14297 50598 14300
rect 50632 14297 50644 14331
rect 50586 14291 50644 14297
rect 50062 14260 50068 14272
rect 49620 14232 50068 14260
rect 35069 14223 35127 14229
rect 50062 14220 50068 14232
rect 50120 14220 50126 14272
rect 51718 14220 51724 14272
rect 51776 14260 51782 14272
rect 57900 14260 57928 14359
rect 58158 14288 58164 14340
rect 58216 14288 58222 14340
rect 51776 14232 57928 14260
rect 51776 14220 51782 14232
rect 1104 14170 58880 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 50294 14170
rect 50346 14118 50358 14170
rect 50410 14118 50422 14170
rect 50474 14118 50486 14170
rect 50538 14118 50550 14170
rect 50602 14118 58880 14170
rect 1104 14096 58880 14118
rect 15562 14016 15568 14068
rect 15620 14016 15626 14068
rect 20714 14016 20720 14068
rect 20772 14056 20778 14068
rect 21361 14059 21419 14065
rect 21361 14056 21373 14059
rect 20772 14028 21373 14056
rect 20772 14016 20778 14028
rect 21361 14025 21373 14028
rect 21407 14025 21419 14059
rect 21361 14019 21419 14025
rect 22278 14016 22284 14068
rect 22336 14056 22342 14068
rect 26326 14056 26332 14068
rect 22336 14028 26332 14056
rect 22336 14016 22342 14028
rect 26326 14016 26332 14028
rect 26384 14016 26390 14068
rect 26602 14016 26608 14068
rect 26660 14016 26666 14068
rect 27706 14016 27712 14068
rect 27764 14016 27770 14068
rect 29089 14059 29147 14065
rect 29089 14025 29101 14059
rect 29135 14056 29147 14059
rect 29178 14056 29184 14068
rect 29135 14028 29184 14056
rect 29135 14025 29147 14028
rect 29089 14019 29147 14025
rect 29178 14016 29184 14028
rect 29236 14016 29242 14068
rect 30190 14016 30196 14068
rect 30248 14056 30254 14068
rect 30653 14059 30711 14065
rect 30653 14056 30665 14059
rect 30248 14028 30665 14056
rect 30248 14016 30254 14028
rect 30653 14025 30665 14028
rect 30699 14025 30711 14059
rect 30653 14019 30711 14025
rect 31018 14016 31024 14068
rect 31076 14056 31082 14068
rect 31487 14059 31545 14065
rect 31487 14056 31499 14059
rect 31076 14028 31499 14056
rect 31076 14016 31082 14028
rect 31487 14025 31499 14028
rect 31533 14025 31545 14059
rect 31487 14019 31545 14025
rect 31573 14059 31631 14065
rect 31573 14025 31585 14059
rect 31619 14056 31631 14059
rect 31662 14056 31668 14068
rect 31619 14028 31668 14056
rect 31619 14025 31631 14028
rect 31573 14019 31631 14025
rect 31662 14016 31668 14028
rect 31720 14016 31726 14068
rect 32309 14059 32367 14065
rect 32309 14025 32321 14059
rect 32355 14056 32367 14059
rect 32355 14028 34376 14056
rect 32355 14025 32367 14028
rect 32309 14019 32367 14025
rect 15105 13991 15163 13997
rect 15105 13957 15117 13991
rect 15151 13988 15163 13991
rect 15470 13988 15476 14000
rect 15151 13960 15476 13988
rect 15151 13957 15163 13960
rect 15105 13951 15163 13957
rect 15470 13948 15476 13960
rect 15528 13948 15534 14000
rect 17310 13948 17316 14000
rect 17368 13988 17374 14000
rect 17368 13960 23060 13988
rect 17368 13948 17374 13960
rect 1581 13923 1639 13929
rect 1581 13889 1593 13923
rect 1627 13920 1639 13923
rect 21177 13923 21235 13929
rect 1627 13892 16574 13920
rect 1627 13889 1639 13892
rect 1581 13883 1639 13889
rect 934 13812 940 13864
rect 992 13852 998 13864
rect 1765 13855 1823 13861
rect 1765 13852 1777 13855
rect 992 13824 1777 13852
rect 992 13812 998 13824
rect 1765 13821 1777 13824
rect 1811 13821 1823 13855
rect 16546 13852 16574 13892
rect 21177 13889 21189 13923
rect 21223 13920 21235 13923
rect 22186 13920 22192 13932
rect 21223 13892 22192 13920
rect 21223 13889 21235 13892
rect 21177 13883 21235 13889
rect 22186 13880 22192 13892
rect 22244 13920 22250 13932
rect 22462 13920 22468 13932
rect 22244 13892 22468 13920
rect 22244 13880 22250 13892
rect 22462 13880 22468 13892
rect 22520 13880 22526 13932
rect 22094 13852 22100 13864
rect 16546 13824 22100 13852
rect 1765 13815 1823 13821
rect 22094 13812 22100 13824
rect 22152 13812 22158 13864
rect 23032 13852 23060 13960
rect 24118 13948 24124 14000
rect 24176 13988 24182 14000
rect 24314 13991 24372 13997
rect 24314 13988 24326 13991
rect 24176 13960 24326 13988
rect 24176 13948 24182 13960
rect 24314 13957 24326 13960
rect 24360 13988 24372 13991
rect 24854 13988 24860 14000
rect 24360 13960 24860 13988
rect 24360 13957 24372 13960
rect 24314 13951 24372 13957
rect 24854 13948 24860 13960
rect 24912 13948 24918 14000
rect 25958 13988 25964 14000
rect 25240 13960 25964 13988
rect 25240 13932 25268 13960
rect 25958 13948 25964 13960
rect 26016 13988 26022 14000
rect 29822 13988 29828 14000
rect 26016 13960 26372 13988
rect 26016 13948 26022 13960
rect 23934 13880 23940 13932
rect 23992 13880 23998 13932
rect 24486 13880 24492 13932
rect 24544 13920 24550 13932
rect 24581 13923 24639 13929
rect 24581 13920 24593 13923
rect 24544 13892 24593 13920
rect 24544 13880 24550 13892
rect 24581 13889 24593 13892
rect 24627 13889 24639 13923
rect 24581 13883 24639 13889
rect 25222 13880 25228 13932
rect 25280 13880 25286 13932
rect 25492 13923 25550 13929
rect 25492 13889 25504 13923
rect 25538 13920 25550 13923
rect 26234 13920 26240 13932
rect 25538 13892 26240 13920
rect 25538 13889 25550 13892
rect 25492 13883 25550 13889
rect 26234 13880 26240 13892
rect 26292 13880 26298 13932
rect 26344 13920 26372 13960
rect 26528 13960 29828 13988
rect 26528 13920 26556 13960
rect 29822 13948 29828 13960
rect 29880 13988 29886 14000
rect 29880 13960 34008 13988
rect 29880 13948 29886 13960
rect 26344 13892 26556 13920
rect 27525 13923 27583 13929
rect 27525 13889 27537 13923
rect 27571 13920 27583 13923
rect 28902 13920 28908 13932
rect 27571 13892 28908 13920
rect 27571 13889 27583 13892
rect 27525 13883 27583 13889
rect 28902 13880 28908 13892
rect 28960 13880 28966 13932
rect 29365 13923 29423 13929
rect 29365 13920 29377 13923
rect 29104 13892 29377 13920
rect 24302 13852 24308 13864
rect 23032 13824 24308 13852
rect 24302 13812 24308 13824
rect 24360 13812 24366 13864
rect 26326 13812 26332 13864
rect 26384 13852 26390 13864
rect 28718 13852 28724 13864
rect 26384 13824 28724 13852
rect 26384 13812 26390 13824
rect 28718 13812 28724 13824
rect 28776 13812 28782 13864
rect 15286 13744 15292 13796
rect 15344 13784 15350 13796
rect 15381 13787 15439 13793
rect 15381 13784 15393 13787
rect 15344 13756 15393 13784
rect 15344 13744 15350 13756
rect 15381 13753 15393 13756
rect 15427 13753 15439 13787
rect 15381 13747 15439 13753
rect 22738 13744 22744 13796
rect 22796 13784 22802 13796
rect 22796 13756 24440 13784
rect 22796 13744 22802 13756
rect 23566 13676 23572 13728
rect 23624 13716 23630 13728
rect 24210 13716 24216 13728
rect 23624 13688 24216 13716
rect 23624 13676 23630 13688
rect 24210 13676 24216 13688
rect 24268 13716 24274 13728
rect 24305 13719 24363 13725
rect 24305 13716 24317 13719
rect 24268 13688 24317 13716
rect 24268 13676 24274 13688
rect 24305 13685 24317 13688
rect 24351 13685 24363 13719
rect 24412 13716 24440 13756
rect 28810 13744 28816 13796
rect 28868 13784 28874 13796
rect 29104 13784 29132 13892
rect 29365 13889 29377 13892
rect 29411 13889 29423 13923
rect 29365 13883 29423 13889
rect 29457 13923 29515 13929
rect 29457 13889 29469 13923
rect 29503 13889 29515 13923
rect 29457 13883 29515 13889
rect 29472 13852 29500 13883
rect 29546 13880 29552 13932
rect 29604 13880 29610 13932
rect 29638 13880 29644 13932
rect 29696 13920 29702 13932
rect 29733 13923 29791 13929
rect 29733 13920 29745 13923
rect 29696 13892 29745 13920
rect 29696 13880 29702 13892
rect 29733 13889 29745 13892
rect 29779 13889 29791 13923
rect 29733 13883 29791 13889
rect 29914 13880 29920 13932
rect 29972 13920 29978 13932
rect 30469 13923 30527 13929
rect 30469 13920 30481 13923
rect 29972 13892 30481 13920
rect 29972 13880 29978 13892
rect 30469 13889 30481 13892
rect 30515 13889 30527 13923
rect 30469 13883 30527 13889
rect 31386 13880 31392 13932
rect 31444 13880 31450 13932
rect 31665 13923 31723 13929
rect 31665 13920 31677 13923
rect 31496 13892 31677 13920
rect 30098 13852 30104 13864
rect 29472 13824 30104 13852
rect 30098 13812 30104 13824
rect 30156 13812 30162 13864
rect 30650 13812 30656 13864
rect 30708 13852 30714 13864
rect 31496 13852 31524 13892
rect 31665 13889 31677 13892
rect 31711 13889 31723 13923
rect 31665 13883 31723 13889
rect 32493 13923 32551 13929
rect 32493 13889 32505 13923
rect 32539 13889 32551 13923
rect 32493 13883 32551 13889
rect 32508 13852 32536 13883
rect 32582 13880 32588 13932
rect 32640 13880 32646 13932
rect 32858 13880 32864 13932
rect 32916 13880 32922 13932
rect 33318 13880 33324 13932
rect 33376 13880 33382 13932
rect 33505 13923 33563 13929
rect 33505 13889 33517 13923
rect 33551 13920 33563 13923
rect 33778 13920 33784 13932
rect 33551 13892 33784 13920
rect 33551 13889 33563 13892
rect 33505 13883 33563 13889
rect 33778 13880 33784 13892
rect 33836 13880 33842 13932
rect 33980 13929 34008 13960
rect 33965 13923 34023 13929
rect 33965 13889 33977 13923
rect 34011 13889 34023 13923
rect 33965 13883 34023 13889
rect 34054 13880 34060 13932
rect 34112 13920 34118 13932
rect 34221 13923 34279 13929
rect 34221 13920 34233 13923
rect 34112 13892 34233 13920
rect 34112 13880 34118 13892
rect 34221 13889 34233 13892
rect 34267 13889 34279 13923
rect 34348 13920 34376 14028
rect 35342 14016 35348 14068
rect 35400 14016 35406 14068
rect 37829 14059 37887 14065
rect 37829 14025 37841 14059
rect 37875 14056 37887 14059
rect 38930 14056 38936 14068
rect 37875 14028 38936 14056
rect 37875 14025 37887 14028
rect 37829 14019 37887 14025
rect 38930 14016 38936 14028
rect 38988 14016 38994 14068
rect 50433 14059 50491 14065
rect 41386 14028 50384 14056
rect 34422 13948 34428 14000
rect 34480 13988 34486 14000
rect 41386 13988 41414 14028
rect 34480 13960 41414 13988
rect 34480 13948 34486 13960
rect 44910 13948 44916 14000
rect 44968 13988 44974 14000
rect 46658 13988 46664 14000
rect 44968 13960 46664 13988
rect 44968 13948 44974 13960
rect 46658 13948 46664 13960
rect 46716 13948 46722 14000
rect 49878 13948 49884 14000
rect 49936 13948 49942 14000
rect 50356 13988 50384 14028
rect 50433 14025 50445 14059
rect 50479 14056 50491 14059
rect 50890 14056 50896 14068
rect 50479 14028 50896 14056
rect 50479 14025 50491 14028
rect 50433 14019 50491 14025
rect 50890 14016 50896 14028
rect 50948 14016 50954 14068
rect 58250 13988 58256 14000
rect 50356 13960 58256 13988
rect 58250 13948 58256 13960
rect 58308 13948 58314 14000
rect 35802 13920 35808 13932
rect 34348 13892 35808 13920
rect 34221 13883 34279 13889
rect 35802 13880 35808 13892
rect 35860 13880 35866 13932
rect 42613 13923 42671 13929
rect 42613 13889 42625 13923
rect 42659 13920 42671 13923
rect 42702 13920 42708 13932
rect 42659 13892 42708 13920
rect 42659 13889 42671 13892
rect 42613 13883 42671 13889
rect 42702 13880 42708 13892
rect 42760 13880 42766 13932
rect 42880 13923 42938 13929
rect 42880 13889 42892 13923
rect 42926 13920 42938 13923
rect 43162 13920 43168 13932
rect 42926 13892 43168 13920
rect 42926 13889 42938 13892
rect 42880 13883 42938 13889
rect 43162 13880 43168 13892
rect 43220 13880 43226 13932
rect 49896 13920 49924 13948
rect 50430 13923 50488 13929
rect 49896 13892 50384 13920
rect 30708 13824 31524 13852
rect 31726 13824 32536 13852
rect 30708 13812 30714 13824
rect 28868 13756 29132 13784
rect 28868 13744 28874 13756
rect 30374 13744 30380 13796
rect 30432 13784 30438 13796
rect 31726 13784 31754 13824
rect 37918 13812 37924 13864
rect 37976 13812 37982 13864
rect 38102 13812 38108 13864
rect 38160 13852 38166 13864
rect 38470 13852 38476 13864
rect 38160 13824 38476 13852
rect 38160 13812 38166 13824
rect 38470 13812 38476 13824
rect 38528 13812 38534 13864
rect 50062 13812 50068 13864
rect 50120 13852 50126 13864
rect 50120 13824 50292 13852
rect 50120 13812 50126 13824
rect 30432 13756 31754 13784
rect 30432 13744 30438 13756
rect 32674 13744 32680 13796
rect 32732 13784 32738 13796
rect 50264 13793 50292 13824
rect 32769 13787 32827 13793
rect 32769 13784 32781 13787
rect 32732 13756 32781 13784
rect 32732 13744 32738 13756
rect 32769 13753 32781 13756
rect 32815 13753 32827 13787
rect 32769 13747 32827 13753
rect 50249 13787 50307 13793
rect 50249 13753 50261 13787
rect 50295 13753 50307 13787
rect 50356 13784 50384 13892
rect 50430 13889 50442 13923
rect 50476 13920 50488 13923
rect 51718 13920 51724 13932
rect 50476 13892 51724 13920
rect 50476 13889 50488 13892
rect 50430 13883 50488 13889
rect 51718 13880 51724 13892
rect 51776 13880 51782 13932
rect 56410 13880 56416 13932
rect 56468 13880 56474 13932
rect 57054 13880 57060 13932
rect 57112 13880 57118 13932
rect 58066 13880 58072 13932
rect 58124 13880 58130 13932
rect 50614 13812 50620 13864
rect 50672 13852 50678 13864
rect 50893 13855 50951 13861
rect 50893 13852 50905 13855
rect 50672 13824 50905 13852
rect 50672 13812 50678 13824
rect 50893 13821 50905 13824
rect 50939 13852 50951 13855
rect 51074 13852 51080 13864
rect 50939 13824 51080 13852
rect 50939 13821 50951 13824
rect 50893 13815 50951 13821
rect 51074 13812 51080 13824
rect 51132 13812 51138 13864
rect 56226 13812 56232 13864
rect 56284 13812 56290 13864
rect 57333 13855 57391 13861
rect 57333 13821 57345 13855
rect 57379 13852 57391 13855
rect 58986 13852 58992 13864
rect 57379 13824 58992 13852
rect 57379 13821 57391 13824
rect 57333 13815 57391 13821
rect 58986 13812 58992 13824
rect 59044 13812 59050 13864
rect 50801 13787 50859 13793
rect 50801 13784 50813 13787
rect 50356 13756 50813 13784
rect 50249 13747 50307 13753
rect 50801 13753 50813 13756
rect 50847 13753 50859 13787
rect 50801 13747 50859 13753
rect 58158 13744 58164 13796
rect 58216 13784 58222 13796
rect 58253 13787 58311 13793
rect 58253 13784 58265 13787
rect 58216 13756 58265 13784
rect 58216 13744 58222 13756
rect 58253 13753 58265 13756
rect 58299 13753 58311 13787
rect 58253 13747 58311 13753
rect 30006 13716 30012 13728
rect 24412 13688 30012 13716
rect 24305 13679 24363 13685
rect 30006 13676 30012 13688
rect 30064 13676 30070 13728
rect 31754 13676 31760 13728
rect 31812 13716 31818 13728
rect 32692 13716 32720 13744
rect 31812 13688 32720 13716
rect 33413 13719 33471 13725
rect 31812 13676 31818 13688
rect 33413 13685 33425 13719
rect 33459 13716 33471 13719
rect 34146 13716 34152 13728
rect 33459 13688 34152 13716
rect 33459 13685 33471 13688
rect 33413 13679 33471 13685
rect 34146 13676 34152 13688
rect 34204 13676 34210 13728
rect 37458 13676 37464 13728
rect 37516 13676 37522 13728
rect 43898 13676 43904 13728
rect 43956 13716 43962 13728
rect 43993 13719 44051 13725
rect 43993 13716 44005 13719
rect 43956 13688 44005 13716
rect 43956 13676 43962 13688
rect 43993 13685 44005 13688
rect 44039 13685 44051 13719
rect 43993 13679 44051 13685
rect 56594 13676 56600 13728
rect 56652 13676 56658 13728
rect 1104 13626 58880 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 58880 13626
rect 1104 13552 58880 13574
rect 16206 13472 16212 13524
rect 16264 13472 16270 13524
rect 21269 13515 21327 13521
rect 21269 13481 21281 13515
rect 21315 13512 21327 13515
rect 21358 13512 21364 13524
rect 21315 13484 21364 13512
rect 21315 13481 21327 13484
rect 21269 13475 21327 13481
rect 21358 13472 21364 13484
rect 21416 13472 21422 13524
rect 21450 13472 21456 13524
rect 21508 13512 21514 13524
rect 28166 13512 28172 13524
rect 21508 13484 28172 13512
rect 21508 13472 21514 13484
rect 28166 13472 28172 13484
rect 28224 13472 28230 13524
rect 29270 13472 29276 13524
rect 29328 13512 29334 13524
rect 30285 13515 30343 13521
rect 30285 13512 30297 13515
rect 29328 13484 30297 13512
rect 29328 13472 29334 13484
rect 30285 13481 30297 13484
rect 30331 13481 30343 13515
rect 30285 13475 30343 13481
rect 32582 13472 32588 13524
rect 32640 13512 32646 13524
rect 32861 13515 32919 13521
rect 32861 13512 32873 13515
rect 32640 13484 32873 13512
rect 32640 13472 32646 13484
rect 32861 13481 32873 13484
rect 32907 13481 32919 13515
rect 32861 13475 32919 13481
rect 33689 13515 33747 13521
rect 33689 13481 33701 13515
rect 33735 13512 33747 13515
rect 34054 13512 34060 13524
rect 33735 13484 34060 13512
rect 33735 13481 33747 13484
rect 33689 13475 33747 13481
rect 34054 13472 34060 13484
rect 34112 13472 34118 13524
rect 37553 13515 37611 13521
rect 37553 13512 37565 13515
rect 35728 13484 37565 13512
rect 16022 13404 16028 13456
rect 16080 13404 16086 13456
rect 23106 13404 23112 13456
rect 23164 13444 23170 13456
rect 24118 13444 24124 13456
rect 23164 13416 24124 13444
rect 23164 13404 23170 13416
rect 24118 13404 24124 13416
rect 24176 13404 24182 13456
rect 27065 13447 27123 13453
rect 27065 13444 27077 13447
rect 26252 13416 27077 13444
rect 15470 13336 15476 13388
rect 15528 13376 15534 13388
rect 15749 13379 15807 13385
rect 15749 13376 15761 13379
rect 15528 13348 15761 13376
rect 15528 13336 15534 13348
rect 15749 13345 15761 13348
rect 15795 13345 15807 13379
rect 23750 13376 23756 13388
rect 15749 13339 15807 13345
rect 16546 13348 23756 13376
rect 1581 13311 1639 13317
rect 1581 13277 1593 13311
rect 1627 13308 1639 13311
rect 4246 13308 4252 13320
rect 1627 13280 4252 13308
rect 1627 13277 1639 13280
rect 1581 13271 1639 13277
rect 4246 13268 4252 13280
rect 4304 13268 4310 13320
rect 8478 13268 8484 13320
rect 8536 13308 8542 13320
rect 16546 13308 16574 13348
rect 23750 13336 23756 13348
rect 23808 13336 23814 13388
rect 24578 13336 24584 13388
rect 24636 13376 24642 13388
rect 25222 13376 25228 13388
rect 24636 13348 25228 13376
rect 24636 13336 24642 13348
rect 25222 13336 25228 13348
rect 25280 13336 25286 13388
rect 8536 13280 16574 13308
rect 21085 13311 21143 13317
rect 8536 13268 8542 13280
rect 21085 13277 21097 13311
rect 21131 13308 21143 13311
rect 22554 13308 22560 13320
rect 21131 13280 22560 13308
rect 21131 13277 21143 13280
rect 21085 13271 21143 13277
rect 22554 13268 22560 13280
rect 22612 13268 22618 13320
rect 23658 13268 23664 13320
rect 23716 13268 23722 13320
rect 934 13200 940 13252
rect 992 13240 998 13252
rect 1857 13243 1915 13249
rect 1857 13240 1869 13243
rect 992 13212 1869 13240
rect 992 13200 998 13212
rect 1857 13209 1869 13212
rect 1903 13209 1915 13243
rect 1857 13203 1915 13209
rect 20530 13200 20536 13252
rect 20588 13240 20594 13252
rect 25492 13243 25550 13249
rect 20588 13212 25452 13240
rect 20588 13200 20594 13212
rect 23290 13132 23296 13184
rect 23348 13172 23354 13184
rect 23845 13175 23903 13181
rect 23845 13172 23857 13175
rect 23348 13144 23857 13172
rect 23348 13132 23354 13144
rect 23845 13141 23857 13144
rect 23891 13172 23903 13175
rect 25314 13172 25320 13184
rect 23891 13144 25320 13172
rect 23891 13141 23903 13144
rect 23845 13135 23903 13141
rect 25314 13132 25320 13144
rect 25372 13132 25378 13184
rect 25424 13172 25452 13212
rect 25492 13209 25504 13243
rect 25538 13240 25550 13243
rect 26252 13240 26280 13416
rect 27065 13413 27077 13416
rect 27111 13413 27123 13447
rect 27065 13407 27123 13413
rect 27154 13404 27160 13456
rect 27212 13444 27218 13456
rect 35728 13444 35756 13484
rect 37553 13481 37565 13484
rect 37599 13512 37611 13515
rect 37918 13512 37924 13524
rect 37599 13484 37924 13512
rect 37599 13481 37611 13484
rect 37553 13475 37611 13481
rect 37918 13472 37924 13484
rect 37976 13472 37982 13524
rect 48314 13472 48320 13524
rect 48372 13512 48378 13524
rect 55677 13515 55735 13521
rect 48372 13484 51074 13512
rect 48372 13472 48378 13484
rect 27212 13416 35756 13444
rect 27212 13404 27218 13416
rect 49878 13404 49884 13456
rect 49936 13444 49942 13456
rect 50341 13447 50399 13453
rect 50341 13444 50353 13447
rect 49936 13416 50353 13444
rect 49936 13404 49942 13416
rect 50341 13413 50353 13416
rect 50387 13413 50399 13447
rect 51046 13444 51074 13484
rect 55677 13481 55689 13515
rect 55723 13512 55735 13515
rect 56410 13512 56416 13524
rect 55723 13484 56416 13512
rect 55723 13481 55735 13484
rect 55677 13475 55735 13481
rect 56410 13472 56416 13484
rect 56468 13472 56474 13524
rect 57698 13472 57704 13524
rect 57756 13512 57762 13524
rect 58161 13515 58219 13521
rect 58161 13512 58173 13515
rect 57756 13484 58173 13512
rect 57756 13472 57762 13484
rect 58161 13481 58173 13484
rect 58207 13481 58219 13515
rect 58161 13475 58219 13481
rect 51046 13416 51672 13444
rect 50341 13407 50399 13413
rect 26878 13336 26884 13388
rect 26936 13376 26942 13388
rect 27617 13379 27675 13385
rect 27617 13376 27629 13379
rect 26936 13348 27629 13376
rect 26936 13336 26942 13348
rect 27617 13345 27629 13348
rect 27663 13345 27675 13379
rect 27617 13339 27675 13345
rect 27890 13336 27896 13388
rect 27948 13376 27954 13388
rect 34422 13376 34428 13388
rect 27948 13348 31754 13376
rect 27948 13336 27954 13348
rect 27525 13311 27583 13317
rect 27525 13308 27537 13311
rect 25538 13212 26280 13240
rect 26620 13280 27537 13308
rect 25538 13209 25550 13212
rect 25492 13203 25550 13209
rect 26620 13181 26648 13280
rect 27525 13277 27537 13280
rect 27571 13277 27583 13311
rect 27525 13271 27583 13277
rect 30101 13311 30159 13317
rect 30101 13277 30113 13311
rect 30147 13277 30159 13311
rect 30101 13271 30159 13277
rect 27433 13243 27491 13249
rect 27433 13209 27445 13243
rect 27479 13240 27491 13243
rect 28810 13240 28816 13252
rect 27479 13212 28816 13240
rect 27479 13209 27491 13212
rect 27433 13203 27491 13209
rect 28810 13200 28816 13212
rect 28868 13200 28874 13252
rect 30116 13240 30144 13271
rect 30282 13268 30288 13320
rect 30340 13308 30346 13320
rect 30650 13308 30656 13320
rect 30340 13280 30656 13308
rect 30340 13268 30346 13280
rect 30650 13268 30656 13280
rect 30708 13308 30714 13320
rect 30837 13311 30895 13317
rect 30837 13308 30849 13311
rect 30708 13280 30849 13308
rect 30708 13268 30714 13280
rect 30837 13277 30849 13280
rect 30883 13277 30895 13311
rect 30837 13271 30895 13277
rect 30116 13212 31064 13240
rect 26605 13175 26663 13181
rect 26605 13172 26617 13175
rect 25424 13144 26617 13172
rect 26605 13141 26617 13144
rect 26651 13141 26663 13175
rect 26605 13135 26663 13141
rect 28166 13132 28172 13184
rect 28224 13172 28230 13184
rect 30374 13172 30380 13184
rect 28224 13144 30380 13172
rect 28224 13132 28230 13144
rect 30374 13132 30380 13144
rect 30432 13132 30438 13184
rect 31036 13181 31064 13212
rect 31021 13175 31079 13181
rect 31021 13141 31033 13175
rect 31067 13141 31079 13175
rect 31726 13172 31754 13348
rect 33980 13348 34428 13376
rect 32677 13311 32735 13317
rect 32677 13277 32689 13311
rect 32723 13308 32735 13311
rect 33410 13308 33416 13320
rect 32723 13280 33416 13308
rect 32723 13277 32735 13280
rect 32677 13271 32735 13277
rect 33410 13268 33416 13280
rect 33468 13268 33474 13320
rect 33980 13317 34008 13348
rect 34422 13336 34428 13348
rect 34480 13336 34486 13388
rect 37182 13336 37188 13388
rect 37240 13376 37246 13388
rect 49786 13376 49792 13388
rect 37240 13348 49792 13376
rect 37240 13336 37246 13348
rect 49786 13336 49792 13348
rect 49844 13336 49850 13388
rect 51534 13376 51540 13388
rect 50080 13348 51540 13376
rect 33945 13311 34008 13317
rect 33945 13277 33957 13311
rect 33991 13280 34008 13311
rect 33991 13277 34003 13280
rect 33945 13271 34003 13277
rect 34054 13268 34060 13320
rect 34112 13268 34118 13320
rect 34146 13268 34152 13320
rect 34204 13268 34210 13320
rect 34238 13268 34244 13320
rect 34296 13308 34302 13320
rect 34333 13311 34391 13317
rect 34333 13308 34345 13311
rect 34296 13280 34345 13308
rect 34296 13268 34302 13280
rect 34333 13277 34345 13280
rect 34379 13277 34391 13311
rect 34333 13271 34391 13277
rect 36173 13311 36231 13317
rect 36173 13277 36185 13311
rect 36219 13308 36231 13311
rect 36262 13308 36268 13320
rect 36219 13280 36268 13308
rect 36219 13277 36231 13280
rect 36173 13271 36231 13277
rect 36262 13268 36268 13280
rect 36320 13268 36326 13320
rect 36440 13311 36498 13317
rect 36440 13277 36452 13311
rect 36486 13308 36498 13311
rect 37458 13308 37464 13320
rect 36486 13280 37464 13308
rect 36486 13277 36498 13280
rect 36440 13271 36498 13277
rect 37458 13268 37464 13280
rect 37516 13268 37522 13320
rect 41785 13311 41843 13317
rect 41785 13277 41797 13311
rect 41831 13308 41843 13311
rect 50080 13308 50108 13348
rect 51534 13336 51540 13348
rect 51592 13336 51598 13388
rect 41831 13280 50108 13308
rect 50525 13311 50583 13317
rect 41831 13277 41843 13280
rect 41785 13271 41843 13277
rect 50525 13277 50537 13311
rect 50571 13277 50583 13311
rect 50525 13271 50583 13277
rect 32306 13200 32312 13252
rect 32364 13240 32370 13252
rect 32493 13243 32551 13249
rect 32493 13240 32505 13243
rect 32364 13212 32505 13240
rect 32364 13200 32370 13212
rect 32493 13209 32505 13212
rect 32539 13209 32551 13243
rect 32493 13203 32551 13209
rect 41138 13200 41144 13252
rect 41196 13240 41202 13252
rect 43346 13240 43352 13252
rect 41196 13212 43352 13240
rect 41196 13200 41202 13212
rect 43346 13200 43352 13212
rect 43404 13200 43410 13252
rect 46845 13243 46903 13249
rect 46845 13240 46857 13243
rect 45526 13212 46857 13240
rect 36906 13172 36912 13184
rect 31726 13144 36912 13172
rect 31021 13135 31079 13141
rect 36906 13132 36912 13144
rect 36964 13132 36970 13184
rect 43070 13132 43076 13184
rect 43128 13172 43134 13184
rect 44174 13172 44180 13184
rect 43128 13144 44180 13172
rect 43128 13132 43134 13144
rect 44174 13132 44180 13144
rect 44232 13172 44238 13184
rect 45526 13172 45554 13212
rect 46845 13209 46857 13212
rect 46891 13240 46903 13243
rect 49418 13240 49424 13252
rect 46891 13212 49424 13240
rect 46891 13209 46903 13212
rect 46845 13203 46903 13209
rect 49418 13200 49424 13212
rect 49476 13200 49482 13252
rect 49786 13200 49792 13252
rect 49844 13240 49850 13252
rect 50540 13240 50568 13271
rect 50614 13268 50620 13320
rect 50672 13268 50678 13320
rect 51644 13308 51672 13416
rect 55784 13348 56088 13376
rect 55784 13308 55812 13348
rect 51644 13280 55812 13308
rect 55858 13268 55864 13320
rect 55916 13268 55922 13320
rect 49844 13212 50568 13240
rect 49844 13200 49850 13212
rect 44232 13144 45554 13172
rect 44232 13132 44238 13144
rect 47486 13132 47492 13184
rect 47544 13172 47550 13184
rect 48133 13175 48191 13181
rect 48133 13172 48145 13175
rect 47544 13144 48145 13172
rect 47544 13132 47550 13144
rect 48133 13141 48145 13144
rect 48179 13172 48191 13175
rect 50154 13172 50160 13184
rect 48179 13144 50160 13172
rect 48179 13141 48191 13144
rect 48133 13135 48191 13141
rect 50154 13132 50160 13144
rect 50212 13132 50218 13184
rect 50540 13172 50568 13212
rect 50890 13200 50896 13252
rect 50948 13200 50954 13252
rect 50985 13243 51043 13249
rect 50985 13209 50997 13243
rect 51031 13240 51043 13243
rect 51718 13240 51724 13252
rect 51031 13212 51724 13240
rect 51031 13209 51043 13212
rect 50985 13203 51043 13209
rect 51718 13200 51724 13212
rect 51776 13200 51782 13252
rect 55950 13200 55956 13252
rect 56008 13200 56014 13252
rect 56060 13249 56088 13348
rect 56778 13336 56784 13388
rect 56836 13336 56842 13388
rect 56321 13311 56379 13317
rect 56321 13277 56333 13311
rect 56367 13277 56379 13311
rect 56321 13271 56379 13277
rect 56045 13243 56103 13249
rect 56045 13209 56057 13243
rect 56091 13209 56103 13243
rect 56045 13203 56103 13209
rect 51261 13175 51319 13181
rect 51261 13172 51273 13175
rect 50540 13144 51273 13172
rect 51261 13141 51273 13144
rect 51307 13141 51319 13175
rect 56060 13172 56088 13203
rect 56134 13200 56140 13252
rect 56192 13249 56198 13252
rect 56192 13243 56221 13249
rect 56209 13209 56221 13243
rect 56336 13240 56364 13271
rect 56594 13268 56600 13320
rect 56652 13308 56658 13320
rect 57037 13311 57095 13317
rect 57037 13308 57049 13311
rect 56652 13280 57049 13308
rect 56652 13268 56658 13280
rect 57037 13277 57049 13280
rect 57083 13277 57095 13311
rect 57037 13271 57095 13277
rect 57698 13240 57704 13252
rect 56336 13212 57704 13240
rect 56192 13203 56221 13209
rect 56192 13200 56198 13203
rect 57698 13200 57704 13212
rect 57756 13200 57762 13252
rect 57146 13172 57152 13184
rect 56060 13144 57152 13172
rect 51261 13135 51319 13141
rect 57146 13132 57152 13144
rect 57204 13132 57210 13184
rect 1104 13082 58880 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 50294 13082
rect 50346 13030 50358 13082
rect 50410 13030 50422 13082
rect 50474 13030 50486 13082
rect 50538 13030 50550 13082
rect 50602 13030 58880 13082
rect 1104 13008 58880 13030
rect 6886 12940 22876 12968
rect 4246 12860 4252 12912
rect 4304 12900 4310 12912
rect 6886 12900 6914 12940
rect 4304 12872 6914 12900
rect 4304 12860 4310 12872
rect 1581 12835 1639 12841
rect 1581 12801 1593 12835
rect 1627 12832 1639 12835
rect 12342 12832 12348 12844
rect 1627 12804 12348 12832
rect 1627 12801 1639 12804
rect 1581 12795 1639 12801
rect 12342 12792 12348 12804
rect 12400 12792 12406 12844
rect 934 12724 940 12776
rect 992 12764 998 12776
rect 1765 12767 1823 12773
rect 1765 12764 1777 12767
rect 992 12736 1777 12764
rect 992 12724 998 12736
rect 1765 12733 1777 12736
rect 1811 12733 1823 12767
rect 1765 12727 1823 12733
rect 20806 12588 20812 12640
rect 20864 12628 20870 12640
rect 22738 12628 22744 12640
rect 20864 12600 22744 12628
rect 20864 12588 20870 12600
rect 22738 12588 22744 12600
rect 22796 12588 22802 12640
rect 22848 12628 22876 12940
rect 23290 12928 23296 12980
rect 23348 12928 23354 12980
rect 23658 12928 23664 12980
rect 23716 12968 23722 12980
rect 25501 12971 25559 12977
rect 25501 12968 25513 12971
rect 23716 12940 25513 12968
rect 23716 12928 23722 12940
rect 25501 12937 25513 12940
rect 25547 12937 25559 12971
rect 25501 12931 25559 12937
rect 26142 12928 26148 12980
rect 26200 12928 26206 12980
rect 26510 12928 26516 12980
rect 26568 12968 26574 12980
rect 26878 12968 26884 12980
rect 26568 12940 26884 12968
rect 26568 12928 26574 12940
rect 26878 12928 26884 12940
rect 26936 12928 26942 12980
rect 29454 12928 29460 12980
rect 29512 12968 29518 12980
rect 29825 12971 29883 12977
rect 29825 12968 29837 12971
rect 29512 12940 29837 12968
rect 29512 12928 29518 12940
rect 29825 12937 29837 12940
rect 29871 12937 29883 12971
rect 29825 12931 29883 12937
rect 30006 12928 30012 12980
rect 30064 12928 30070 12980
rect 35618 12928 35624 12980
rect 35676 12968 35682 12980
rect 58253 12971 58311 12977
rect 58253 12968 58265 12971
rect 35676 12940 58265 12968
rect 35676 12928 35682 12940
rect 58253 12937 58265 12940
rect 58299 12937 58311 12971
rect 58253 12931 58311 12937
rect 23014 12860 23020 12912
rect 23072 12900 23078 12912
rect 24578 12900 24584 12912
rect 23072 12872 23428 12900
rect 23072 12860 23078 12872
rect 23400 12832 23428 12872
rect 24136 12872 24584 12900
rect 24136 12841 24164 12872
rect 24578 12860 24584 12872
rect 24636 12860 24642 12912
rect 30024 12900 30052 12928
rect 30561 12903 30619 12909
rect 30561 12900 30573 12903
rect 30024 12872 30573 12900
rect 30561 12869 30573 12872
rect 30607 12869 30619 12903
rect 30561 12863 30619 12869
rect 30650 12860 30656 12912
rect 30708 12860 30714 12912
rect 31018 12860 31024 12912
rect 31076 12900 31082 12912
rect 31076 12872 31800 12900
rect 31076 12860 31082 12872
rect 24121 12835 24179 12841
rect 23400 12804 23520 12832
rect 23382 12724 23388 12776
rect 23440 12724 23446 12776
rect 23492 12773 23520 12804
rect 24121 12801 24133 12835
rect 24167 12801 24179 12835
rect 24377 12835 24435 12841
rect 24377 12832 24389 12835
rect 24121 12795 24179 12801
rect 24228 12804 24389 12832
rect 23477 12767 23535 12773
rect 23477 12733 23489 12767
rect 23523 12733 23535 12767
rect 24228 12764 24256 12804
rect 24377 12801 24389 12804
rect 24423 12801 24435 12835
rect 24377 12795 24435 12801
rect 25130 12792 25136 12844
rect 25188 12832 25194 12844
rect 25958 12832 25964 12844
rect 25188 12804 25964 12832
rect 25188 12792 25194 12804
rect 25958 12792 25964 12804
rect 26016 12792 26022 12844
rect 29641 12835 29699 12841
rect 29641 12801 29653 12835
rect 29687 12832 29699 12835
rect 29730 12832 29736 12844
rect 29687 12804 29736 12832
rect 29687 12801 29699 12804
rect 29641 12795 29699 12801
rect 29730 12792 29736 12804
rect 29788 12832 29794 12844
rect 30282 12832 30288 12844
rect 29788 12804 30288 12832
rect 29788 12792 29794 12804
rect 30282 12792 30288 12804
rect 30340 12792 30346 12844
rect 30374 12792 30380 12844
rect 30432 12792 30438 12844
rect 30797 12835 30855 12841
rect 30797 12801 30809 12835
rect 30843 12832 30855 12835
rect 31662 12832 31668 12844
rect 30843 12804 31668 12832
rect 30843 12801 30855 12804
rect 30797 12795 30855 12801
rect 31662 12792 31668 12804
rect 31720 12792 31726 12844
rect 31772 12832 31800 12872
rect 33778 12860 33784 12912
rect 33836 12900 33842 12912
rect 43070 12900 43076 12912
rect 33836 12872 43076 12900
rect 33836 12860 33842 12872
rect 43070 12860 43076 12872
rect 43128 12860 43134 12912
rect 49418 12860 49424 12912
rect 49476 12860 49482 12912
rect 51169 12903 51227 12909
rect 51169 12869 51181 12903
rect 51215 12900 51227 12903
rect 51810 12900 51816 12912
rect 51215 12872 51816 12900
rect 51215 12869 51227 12872
rect 51169 12863 51227 12869
rect 51810 12860 51816 12872
rect 51868 12860 51874 12912
rect 55766 12860 55772 12912
rect 55824 12860 55830 12912
rect 55861 12903 55919 12909
rect 55861 12869 55873 12903
rect 55907 12900 55919 12903
rect 57054 12900 57060 12912
rect 55907 12872 57060 12900
rect 55907 12869 55919 12872
rect 55861 12863 55919 12869
rect 57054 12860 57060 12872
rect 57112 12860 57118 12912
rect 57146 12860 57152 12912
rect 57204 12860 57210 12912
rect 37182 12832 37188 12844
rect 31772 12804 37188 12832
rect 37182 12792 37188 12804
rect 37240 12792 37246 12844
rect 37829 12835 37887 12841
rect 37829 12801 37841 12835
rect 37875 12832 37887 12835
rect 39298 12832 39304 12844
rect 37875 12804 39304 12832
rect 37875 12801 37887 12804
rect 37829 12795 37887 12801
rect 39298 12792 39304 12804
rect 39356 12792 39362 12844
rect 42978 12792 42984 12844
rect 43036 12792 43042 12844
rect 46934 12792 46940 12844
rect 46992 12832 46998 12844
rect 47946 12832 47952 12844
rect 46992 12804 47952 12832
rect 46992 12792 46998 12804
rect 47946 12792 47952 12804
rect 48004 12832 48010 12844
rect 51629 12835 51687 12841
rect 51629 12832 51641 12835
rect 48004 12804 51641 12832
rect 48004 12792 48010 12804
rect 51629 12801 51641 12804
rect 51675 12801 51687 12835
rect 51629 12795 51687 12801
rect 55582 12792 55588 12844
rect 55640 12792 55646 12844
rect 55953 12835 56011 12841
rect 55953 12801 55965 12835
rect 55999 12832 56011 12835
rect 56134 12832 56140 12844
rect 55999 12804 56140 12832
rect 55999 12801 56011 12804
rect 55953 12795 56011 12801
rect 23477 12727 23535 12733
rect 24136 12736 24256 12764
rect 22925 12699 22983 12705
rect 22925 12665 22937 12699
rect 22971 12696 22983 12699
rect 24136 12696 24164 12736
rect 25866 12724 25872 12776
rect 25924 12764 25930 12776
rect 34606 12764 34612 12776
rect 25924 12736 34612 12764
rect 25924 12724 25930 12736
rect 34606 12724 34612 12736
rect 34664 12724 34670 12776
rect 35529 12767 35587 12773
rect 35529 12733 35541 12767
rect 35575 12764 35587 12767
rect 36262 12764 36268 12776
rect 35575 12736 36268 12764
rect 35575 12733 35587 12736
rect 35529 12727 35587 12733
rect 36262 12724 36268 12736
rect 36320 12724 36326 12776
rect 37550 12724 37556 12776
rect 37608 12764 37614 12776
rect 37921 12767 37979 12773
rect 37921 12764 37933 12767
rect 37608 12736 37933 12764
rect 37608 12724 37614 12736
rect 37921 12733 37933 12736
rect 37967 12733 37979 12767
rect 37921 12727 37979 12733
rect 38102 12724 38108 12776
rect 38160 12724 38166 12776
rect 43073 12767 43131 12773
rect 43073 12733 43085 12767
rect 43119 12733 43131 12767
rect 43073 12727 43131 12733
rect 43257 12767 43315 12773
rect 43257 12733 43269 12767
rect 43303 12764 43315 12767
rect 43346 12764 43352 12776
rect 43303 12736 43352 12764
rect 43303 12733 43315 12736
rect 43257 12727 43315 12733
rect 29270 12696 29276 12708
rect 22971 12668 24164 12696
rect 25056 12668 29276 12696
rect 22971 12665 22983 12668
rect 22925 12659 22983 12665
rect 25056 12628 25084 12668
rect 29270 12656 29276 12668
rect 29328 12656 29334 12708
rect 30929 12699 30987 12705
rect 30929 12665 30941 12699
rect 30975 12696 30987 12699
rect 40034 12696 40040 12708
rect 30975 12668 40040 12696
rect 30975 12665 30987 12668
rect 30929 12659 30987 12665
rect 40034 12656 40040 12668
rect 40092 12656 40098 12708
rect 43088 12696 43116 12727
rect 43346 12724 43352 12736
rect 43404 12764 43410 12776
rect 45830 12764 45836 12776
rect 43404 12736 45836 12764
rect 43404 12724 43410 12736
rect 45830 12724 45836 12736
rect 45888 12724 45894 12776
rect 50890 12724 50896 12776
rect 50948 12764 50954 12776
rect 51905 12767 51963 12773
rect 51905 12764 51917 12767
rect 50948 12736 51917 12764
rect 50948 12724 50954 12736
rect 51905 12733 51917 12736
rect 51951 12764 51963 12767
rect 55968 12764 55996 12795
rect 56134 12792 56140 12804
rect 56192 12832 56198 12844
rect 56410 12832 56416 12844
rect 56192 12804 56416 12832
rect 56192 12792 56198 12804
rect 56410 12792 56416 12804
rect 56468 12792 56474 12844
rect 56502 12792 56508 12844
rect 56560 12832 56566 12844
rect 56689 12835 56747 12841
rect 56689 12832 56701 12835
rect 56560 12804 56701 12832
rect 56560 12792 56566 12804
rect 56689 12801 56701 12804
rect 56735 12801 56747 12835
rect 56689 12795 56747 12801
rect 58066 12792 58072 12844
rect 58124 12792 58130 12844
rect 51951 12736 55996 12764
rect 51951 12733 51963 12736
rect 51905 12727 51963 12733
rect 43898 12696 43904 12708
rect 43088 12668 43904 12696
rect 43898 12656 43904 12668
rect 43956 12656 43962 12708
rect 51534 12656 51540 12708
rect 51592 12696 51598 12708
rect 55858 12696 55864 12708
rect 51592 12668 55864 12696
rect 51592 12656 51598 12668
rect 55858 12656 55864 12668
rect 55916 12656 55922 12708
rect 22848 12600 25084 12628
rect 25866 12588 25872 12640
rect 25924 12628 25930 12640
rect 26050 12628 26056 12640
rect 25924 12600 26056 12628
rect 25924 12588 25930 12600
rect 26050 12588 26056 12600
rect 26108 12628 26114 12640
rect 32306 12628 32312 12640
rect 26108 12600 32312 12628
rect 26108 12588 26114 12600
rect 32306 12588 32312 12600
rect 32364 12588 32370 12640
rect 36630 12588 36636 12640
rect 36688 12628 36694 12640
rect 37461 12631 37519 12637
rect 37461 12628 37473 12631
rect 36688 12600 37473 12628
rect 36688 12588 36694 12600
rect 37461 12597 37473 12600
rect 37507 12597 37519 12631
rect 37461 12591 37519 12597
rect 38562 12588 38568 12640
rect 38620 12628 38626 12640
rect 41690 12628 41696 12640
rect 38620 12600 41696 12628
rect 38620 12588 38626 12600
rect 41690 12588 41696 12600
rect 41748 12588 41754 12640
rect 42613 12631 42671 12637
rect 42613 12597 42625 12631
rect 42659 12628 42671 12631
rect 43162 12628 43168 12640
rect 42659 12600 43168 12628
rect 42659 12597 42671 12600
rect 42613 12591 42671 12597
rect 43162 12588 43168 12600
rect 43220 12588 43226 12640
rect 56137 12631 56195 12637
rect 56137 12597 56149 12631
rect 56183 12628 56195 12631
rect 56502 12628 56508 12640
rect 56183 12600 56508 12628
rect 56183 12597 56195 12600
rect 56137 12591 56195 12597
rect 56502 12588 56508 12600
rect 56560 12588 56566 12640
rect 1104 12538 58880 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 58880 12538
rect 1104 12464 58880 12486
rect 12342 12384 12348 12436
rect 12400 12424 12406 12436
rect 13173 12427 13231 12433
rect 13173 12424 13185 12427
rect 12400 12396 13185 12424
rect 12400 12384 12406 12396
rect 13173 12393 13185 12396
rect 13219 12393 13231 12427
rect 13173 12387 13231 12393
rect 22554 12384 22560 12436
rect 22612 12424 22618 12436
rect 22741 12427 22799 12433
rect 22741 12424 22753 12427
rect 22612 12396 22753 12424
rect 22612 12384 22618 12396
rect 22741 12393 22753 12396
rect 22787 12393 22799 12427
rect 22741 12387 22799 12393
rect 23658 12384 23664 12436
rect 23716 12424 23722 12436
rect 23934 12424 23940 12436
rect 23716 12396 23940 12424
rect 23716 12384 23722 12396
rect 23934 12384 23940 12396
rect 23992 12384 23998 12436
rect 24762 12384 24768 12436
rect 24820 12424 24826 12436
rect 24820 12396 28488 12424
rect 24820 12384 24826 12396
rect 23014 12316 23020 12368
rect 23072 12356 23078 12368
rect 23072 12328 23888 12356
rect 23072 12316 23078 12328
rect 13538 12248 13544 12300
rect 13596 12288 13602 12300
rect 15470 12288 15476 12300
rect 13596 12260 15476 12288
rect 13596 12248 13602 12260
rect 15470 12248 15476 12260
rect 15528 12248 15534 12300
rect 23860 12297 23888 12328
rect 23845 12291 23903 12297
rect 22572 12260 23796 12288
rect 1581 12223 1639 12229
rect 1581 12189 1593 12223
rect 1627 12220 1639 12223
rect 13078 12220 13084 12232
rect 1627 12192 13084 12220
rect 1627 12189 1639 12192
rect 1581 12183 1639 12189
rect 13078 12180 13084 12192
rect 13136 12180 13142 12232
rect 13357 12223 13415 12229
rect 13357 12189 13369 12223
rect 13403 12189 13415 12223
rect 13357 12183 13415 12189
rect 934 12112 940 12164
rect 992 12152 998 12164
rect 1857 12155 1915 12161
rect 1857 12152 1869 12155
rect 992 12124 1869 12152
rect 992 12112 998 12124
rect 1857 12121 1869 12124
rect 1903 12121 1915 12155
rect 1857 12115 1915 12121
rect 13170 12112 13176 12164
rect 13228 12152 13234 12164
rect 13372 12152 13400 12183
rect 13446 12180 13452 12232
rect 13504 12180 13510 12232
rect 13630 12180 13636 12232
rect 13688 12180 13694 12232
rect 22572 12229 22600 12260
rect 22557 12223 22615 12229
rect 22557 12189 22569 12223
rect 22603 12189 22615 12223
rect 23474 12220 23480 12232
rect 22557 12183 22615 12189
rect 22756 12192 23480 12220
rect 22756 12152 22784 12192
rect 23474 12180 23480 12192
rect 23532 12180 23538 12232
rect 23658 12180 23664 12232
rect 23716 12180 23722 12232
rect 23768 12220 23796 12260
rect 23845 12257 23857 12291
rect 23891 12257 23903 12291
rect 23845 12251 23903 12257
rect 24578 12248 24584 12300
rect 24636 12248 24642 12300
rect 26142 12220 26148 12232
rect 23768 12192 26148 12220
rect 26142 12180 26148 12192
rect 26200 12180 26206 12232
rect 28460 12220 28488 12396
rect 28902 12384 28908 12436
rect 28960 12424 28966 12436
rect 29089 12427 29147 12433
rect 29089 12424 29101 12427
rect 28960 12396 29101 12424
rect 28960 12384 28966 12396
rect 29089 12393 29101 12396
rect 29135 12393 29147 12427
rect 29089 12387 29147 12393
rect 29178 12384 29184 12436
rect 29236 12424 29242 12436
rect 35710 12424 35716 12436
rect 29236 12396 35716 12424
rect 29236 12384 29242 12396
rect 35710 12384 35716 12396
rect 35768 12384 35774 12436
rect 38102 12384 38108 12436
rect 38160 12424 38166 12436
rect 56594 12424 56600 12436
rect 38160 12396 56600 12424
rect 38160 12384 38166 12396
rect 56594 12384 56600 12396
rect 56652 12384 56658 12436
rect 57054 12384 57060 12436
rect 57112 12424 57118 12436
rect 58161 12427 58219 12433
rect 58161 12424 58173 12427
rect 57112 12396 58173 12424
rect 57112 12384 57118 12396
rect 58161 12393 58173 12396
rect 58207 12393 58219 12427
rect 58161 12387 58219 12393
rect 32398 12356 32404 12368
rect 28920 12328 32404 12356
rect 28920 12229 28948 12328
rect 32398 12316 32404 12328
rect 32456 12316 32462 12368
rect 37366 12316 37372 12368
rect 37424 12356 37430 12368
rect 39758 12356 39764 12368
rect 37424 12328 39764 12356
rect 37424 12316 37430 12328
rect 39758 12316 39764 12328
rect 39816 12316 39822 12368
rect 30837 12291 30895 12297
rect 30837 12257 30849 12291
rect 30883 12288 30895 12291
rect 31018 12288 31024 12300
rect 30883 12260 31024 12288
rect 30883 12257 30895 12260
rect 30837 12251 30895 12257
rect 31018 12248 31024 12260
rect 31076 12248 31082 12300
rect 42153 12291 42211 12297
rect 42153 12257 42165 12291
rect 42199 12288 42211 12291
rect 42978 12288 42984 12300
rect 42199 12260 42984 12288
rect 42199 12257 42211 12260
rect 42153 12251 42211 12257
rect 42978 12248 42984 12260
rect 43036 12288 43042 12300
rect 43349 12291 43407 12297
rect 43349 12288 43361 12291
rect 43036 12260 43361 12288
rect 43036 12248 43042 12260
rect 43349 12257 43361 12260
rect 43395 12288 43407 12291
rect 44082 12288 44088 12300
rect 43395 12260 44088 12288
rect 43395 12257 43407 12260
rect 43349 12251 43407 12257
rect 44082 12248 44088 12260
rect 44140 12248 44146 12300
rect 50154 12248 50160 12300
rect 50212 12288 50218 12300
rect 50341 12291 50399 12297
rect 50341 12288 50353 12291
rect 50212 12260 50353 12288
rect 50212 12248 50218 12260
rect 50341 12257 50353 12260
rect 50387 12257 50399 12291
rect 50341 12251 50399 12257
rect 55766 12248 55772 12300
rect 55824 12288 55830 12300
rect 56045 12291 56103 12297
rect 56045 12288 56057 12291
rect 55824 12260 56057 12288
rect 55824 12248 55830 12260
rect 56045 12257 56057 12260
rect 56091 12257 56103 12291
rect 56045 12251 56103 12257
rect 56778 12248 56784 12300
rect 56836 12248 56842 12300
rect 28905 12223 28963 12229
rect 28905 12220 28917 12223
rect 28460 12192 28917 12220
rect 28905 12189 28917 12192
rect 28951 12189 28963 12223
rect 28905 12183 28963 12189
rect 30374 12180 30380 12232
rect 30432 12220 30438 12232
rect 30653 12223 30711 12229
rect 30653 12220 30665 12223
rect 30432 12192 30665 12220
rect 30432 12180 30438 12192
rect 30653 12189 30665 12192
rect 30699 12189 30711 12223
rect 30653 12183 30711 12189
rect 24826 12155 24884 12161
rect 24826 12152 24838 12155
rect 13228 12124 22784 12152
rect 23308 12124 24838 12152
rect 13228 12112 13234 12124
rect 23308 12093 23336 12124
rect 24826 12121 24838 12124
rect 24872 12121 24884 12155
rect 30668 12152 30696 12183
rect 30926 12180 30932 12232
rect 30984 12180 30990 12232
rect 31205 12223 31263 12229
rect 31205 12189 31217 12223
rect 31251 12189 31263 12223
rect 31205 12183 31263 12189
rect 31018 12152 31024 12164
rect 30668 12124 31024 12152
rect 24826 12115 24884 12121
rect 31018 12112 31024 12124
rect 31076 12112 31082 12164
rect 23293 12087 23351 12093
rect 23293 12053 23305 12087
rect 23339 12053 23351 12087
rect 23293 12047 23351 12053
rect 23750 12044 23756 12096
rect 23808 12044 23814 12096
rect 23934 12044 23940 12096
rect 23992 12084 23998 12096
rect 25961 12087 26019 12093
rect 25961 12084 25973 12087
rect 23992 12056 25973 12084
rect 23992 12044 23998 12056
rect 25961 12053 25973 12056
rect 26007 12053 26019 12087
rect 25961 12047 26019 12053
rect 30282 12044 30288 12096
rect 30340 12084 30346 12096
rect 31220 12084 31248 12183
rect 31754 12180 31760 12232
rect 31812 12220 31818 12232
rect 31849 12223 31907 12229
rect 31849 12220 31861 12223
rect 31812 12192 31861 12220
rect 31812 12180 31818 12192
rect 31849 12189 31861 12192
rect 31895 12220 31907 12223
rect 32674 12220 32680 12232
rect 31895 12192 32680 12220
rect 31895 12189 31907 12192
rect 31849 12183 31907 12189
rect 32674 12180 32680 12192
rect 32732 12220 32738 12232
rect 32950 12220 32956 12232
rect 32732 12192 32956 12220
rect 32732 12180 32738 12192
rect 32950 12180 32956 12192
rect 33008 12180 33014 12232
rect 36262 12180 36268 12232
rect 36320 12220 36326 12232
rect 36357 12223 36415 12229
rect 36357 12220 36369 12223
rect 36320 12192 36369 12220
rect 36320 12180 36326 12192
rect 36357 12189 36369 12192
rect 36403 12220 36415 12223
rect 37642 12220 37648 12232
rect 36403 12192 37648 12220
rect 36403 12189 36415 12192
rect 36357 12183 36415 12189
rect 37642 12180 37648 12192
rect 37700 12180 37706 12232
rect 41874 12180 41880 12232
rect 41932 12180 41938 12232
rect 43073 12223 43131 12229
rect 43073 12189 43085 12223
rect 43119 12220 43131 12223
rect 44266 12220 44272 12232
rect 43119 12192 44272 12220
rect 43119 12189 43131 12192
rect 43073 12183 43131 12189
rect 44266 12180 44272 12192
rect 44324 12180 44330 12232
rect 47118 12180 47124 12232
rect 47176 12220 47182 12232
rect 49326 12220 49332 12232
rect 47176 12192 49332 12220
rect 47176 12180 47182 12192
rect 49326 12180 49332 12192
rect 49384 12220 49390 12232
rect 49421 12223 49479 12229
rect 49421 12220 49433 12223
rect 49384 12192 49433 12220
rect 49384 12180 49390 12192
rect 49421 12189 49433 12192
rect 49467 12189 49479 12223
rect 49421 12183 49479 12189
rect 49605 12223 49663 12229
rect 49605 12189 49617 12223
rect 49651 12220 49663 12223
rect 49878 12220 49884 12232
rect 49651 12192 49884 12220
rect 49651 12189 49663 12192
rect 49605 12183 49663 12189
rect 36624 12155 36682 12161
rect 36624 12121 36636 12155
rect 36670 12152 36682 12155
rect 37458 12152 37464 12164
rect 36670 12124 37464 12152
rect 36670 12121 36682 12124
rect 36624 12115 36682 12121
rect 37458 12112 37464 12124
rect 37516 12112 37522 12164
rect 41322 12152 41328 12164
rect 37568 12124 41328 12152
rect 30340 12056 31248 12084
rect 30340 12044 30346 12056
rect 32490 12044 32496 12096
rect 32548 12084 32554 12096
rect 37568 12084 37596 12124
rect 41322 12112 41328 12124
rect 41380 12112 41386 12164
rect 32548 12056 37596 12084
rect 32548 12044 32554 12056
rect 37734 12044 37740 12096
rect 37792 12044 37798 12096
rect 41506 12044 41512 12096
rect 41564 12044 41570 12096
rect 41966 12044 41972 12096
rect 42024 12044 42030 12096
rect 42702 12044 42708 12096
rect 42760 12044 42766 12096
rect 43070 12044 43076 12096
rect 43128 12084 43134 12096
rect 43165 12087 43223 12093
rect 43165 12084 43177 12087
rect 43128 12056 43177 12084
rect 43128 12044 43134 12056
rect 43165 12053 43177 12056
rect 43211 12053 43223 12087
rect 49436 12084 49464 12183
rect 49878 12180 49884 12192
rect 49936 12180 49942 12232
rect 54938 12180 54944 12232
rect 54996 12220 55002 12232
rect 55861 12223 55919 12229
rect 55861 12220 55873 12223
rect 54996 12192 55873 12220
rect 54996 12180 55002 12192
rect 55861 12189 55873 12192
rect 55907 12189 55919 12223
rect 55861 12183 55919 12189
rect 49789 12155 49847 12161
rect 49789 12121 49801 12155
rect 49835 12152 49847 12155
rect 50586 12155 50644 12161
rect 50586 12152 50598 12155
rect 49835 12124 50598 12152
rect 49835 12121 49847 12124
rect 49789 12115 49847 12121
rect 50586 12121 50598 12124
rect 50632 12121 50644 12155
rect 56134 12152 56140 12164
rect 50586 12115 50644 12121
rect 51046 12124 56140 12152
rect 51046 12084 51074 12124
rect 56134 12112 56140 12124
rect 56192 12112 56198 12164
rect 56686 12112 56692 12164
rect 56744 12152 56750 12164
rect 57026 12155 57084 12161
rect 57026 12152 57038 12155
rect 56744 12124 57038 12152
rect 56744 12112 56750 12124
rect 57026 12121 57038 12124
rect 57072 12121 57084 12155
rect 57026 12115 57084 12121
rect 49436 12056 51074 12084
rect 43165 12047 43223 12053
rect 51718 12044 51724 12096
rect 51776 12044 51782 12096
rect 1104 11994 58880 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 50294 11994
rect 50346 11942 50358 11994
rect 50410 11942 50422 11994
rect 50474 11942 50486 11994
rect 50538 11942 50550 11994
rect 50602 11942 58880 11994
rect 1104 11920 58880 11942
rect 1578 11840 1584 11892
rect 1636 11880 1642 11892
rect 11698 11880 11704 11892
rect 1636 11852 11704 11880
rect 1636 11840 1642 11852
rect 11698 11840 11704 11852
rect 11756 11840 11762 11892
rect 13078 11840 13084 11892
rect 13136 11840 13142 11892
rect 13446 11840 13452 11892
rect 13504 11880 13510 11892
rect 23290 11880 23296 11892
rect 13504 11852 23296 11880
rect 13504 11840 13510 11852
rect 23290 11840 23296 11852
rect 23348 11840 23354 11892
rect 23658 11840 23664 11892
rect 23716 11880 23722 11892
rect 24029 11883 24087 11889
rect 24029 11880 24041 11883
rect 23716 11852 24041 11880
rect 23716 11840 23722 11852
rect 24029 11849 24041 11852
rect 24075 11849 24087 11883
rect 24029 11843 24087 11849
rect 24946 11840 24952 11892
rect 25004 11880 25010 11892
rect 25317 11883 25375 11889
rect 25317 11880 25329 11883
rect 25004 11852 25329 11880
rect 25004 11840 25010 11852
rect 25317 11849 25329 11852
rect 25363 11849 25375 11883
rect 25317 11843 25375 11849
rect 25406 11840 25412 11892
rect 25464 11880 25470 11892
rect 27341 11883 27399 11889
rect 27341 11880 27353 11883
rect 25464 11852 27353 11880
rect 25464 11840 25470 11852
rect 27341 11849 27353 11852
rect 27387 11849 27399 11883
rect 27341 11843 27399 11849
rect 30650 11840 30656 11892
rect 30708 11880 30714 11892
rect 30929 11883 30987 11889
rect 30929 11880 30941 11883
rect 30708 11852 30941 11880
rect 30708 11840 30714 11852
rect 30929 11849 30941 11852
rect 30975 11849 30987 11883
rect 30929 11843 30987 11849
rect 22738 11812 22744 11824
rect 17880 11784 22744 11812
rect 17880 11753 17908 11784
rect 22738 11772 22744 11784
rect 22796 11772 22802 11824
rect 23934 11772 23940 11824
rect 23992 11772 23998 11824
rect 29638 11812 29644 11824
rect 27172 11784 29644 11812
rect 1581 11747 1639 11753
rect 1581 11713 1593 11747
rect 1627 11744 1639 11747
rect 17865 11747 17923 11753
rect 1627 11716 17724 11744
rect 1627 11713 1639 11716
rect 1581 11707 1639 11713
rect 934 11636 940 11688
rect 992 11676 998 11688
rect 1765 11679 1823 11685
rect 1765 11676 1777 11679
rect 992 11648 1777 11676
rect 992 11636 998 11648
rect 1765 11645 1777 11648
rect 1811 11645 1823 11679
rect 1765 11639 1823 11645
rect 13170 11636 13176 11688
rect 13228 11676 13234 11688
rect 13265 11679 13323 11685
rect 13265 11676 13277 11679
rect 13228 11648 13277 11676
rect 13228 11636 13234 11648
rect 13265 11645 13277 11648
rect 13311 11645 13323 11679
rect 13265 11639 13323 11645
rect 13357 11679 13415 11685
rect 13357 11645 13369 11679
rect 13403 11645 13415 11679
rect 13357 11639 13415 11645
rect 13372 11608 13400 11639
rect 13446 11636 13452 11688
rect 13504 11636 13510 11688
rect 13538 11636 13544 11688
rect 13596 11636 13602 11688
rect 17696 11685 17724 11716
rect 17865 11713 17877 11747
rect 17911 11713 17923 11747
rect 17865 11707 17923 11713
rect 17957 11747 18015 11753
rect 17957 11713 17969 11747
rect 18003 11744 18015 11747
rect 18003 11716 22094 11744
rect 18003 11713 18015 11716
rect 17957 11707 18015 11713
rect 17681 11679 17739 11685
rect 17681 11645 17693 11679
rect 17727 11645 17739 11679
rect 17681 11639 17739 11645
rect 18046 11636 18052 11688
rect 18104 11636 18110 11688
rect 18138 11636 18144 11688
rect 18196 11636 18202 11688
rect 20714 11608 20720 11620
rect 13372 11580 20720 11608
rect 20714 11568 20720 11580
rect 20772 11568 20778 11620
rect 22066 11608 22094 11716
rect 25130 11704 25136 11756
rect 25188 11704 25194 11756
rect 27172 11753 27200 11784
rect 29638 11772 29644 11784
rect 29696 11772 29702 11824
rect 29822 11753 29828 11756
rect 27157 11747 27215 11753
rect 27157 11713 27169 11747
rect 27203 11713 27215 11747
rect 27157 11707 27215 11713
rect 29816 11707 29828 11753
rect 29822 11704 29828 11707
rect 29880 11704 29886 11756
rect 30944 11744 30972 11843
rect 31018 11840 31024 11892
rect 31076 11880 31082 11892
rect 32122 11880 32128 11892
rect 31076 11852 32128 11880
rect 31076 11840 31082 11852
rect 32122 11840 32128 11852
rect 32180 11880 32186 11892
rect 32401 11883 32459 11889
rect 32401 11880 32413 11883
rect 32180 11852 32413 11880
rect 32180 11840 32186 11852
rect 32401 11849 32413 11852
rect 32447 11849 32459 11883
rect 32401 11843 32459 11849
rect 37458 11840 37464 11892
rect 37516 11840 37522 11892
rect 37829 11883 37887 11889
rect 37829 11849 37841 11883
rect 37875 11880 37887 11883
rect 38838 11880 38844 11892
rect 37875 11852 38844 11880
rect 37875 11849 37887 11852
rect 37829 11843 37887 11849
rect 38838 11840 38844 11852
rect 38896 11840 38902 11892
rect 42978 11840 42984 11892
rect 43036 11840 43042 11892
rect 47762 11840 47768 11892
rect 47820 11880 47826 11892
rect 49050 11880 49056 11892
rect 47820 11852 49056 11880
rect 47820 11840 47826 11852
rect 49050 11840 49056 11852
rect 49108 11840 49114 11892
rect 56686 11840 56692 11892
rect 56744 11840 56750 11892
rect 31389 11815 31447 11821
rect 31389 11781 31401 11815
rect 31435 11812 31447 11815
rect 36262 11812 36268 11824
rect 31435 11784 31754 11812
rect 31435 11781 31447 11784
rect 31389 11775 31447 11781
rect 31573 11747 31631 11753
rect 31573 11744 31585 11747
rect 30944 11716 31585 11744
rect 31573 11713 31585 11716
rect 31619 11713 31631 11747
rect 31726 11744 31754 11784
rect 35544 11784 36268 11812
rect 32490 11744 32496 11756
rect 31726 11716 32496 11744
rect 31573 11707 31631 11713
rect 31864 11688 31892 11716
rect 32490 11704 32496 11716
rect 32548 11704 32554 11756
rect 32585 11747 32643 11753
rect 32585 11713 32597 11747
rect 32631 11744 32643 11747
rect 32674 11744 32680 11756
rect 32631 11716 32680 11744
rect 32631 11713 32643 11716
rect 32585 11707 32643 11713
rect 32674 11704 32680 11716
rect 32732 11704 32738 11756
rect 32766 11704 32772 11756
rect 32824 11704 32830 11756
rect 34790 11704 34796 11756
rect 34848 11744 34854 11756
rect 34885 11747 34943 11753
rect 34885 11744 34897 11747
rect 34848 11716 34897 11744
rect 34848 11704 34854 11716
rect 34885 11713 34897 11716
rect 34931 11713 34943 11747
rect 34885 11707 34943 11713
rect 35342 11704 35348 11756
rect 35400 11744 35406 11756
rect 35544 11753 35572 11784
rect 36262 11772 36268 11784
rect 36320 11772 36326 11824
rect 37734 11772 37740 11824
rect 37792 11812 37798 11824
rect 37921 11815 37979 11821
rect 37921 11812 37933 11815
rect 37792 11784 37933 11812
rect 37792 11772 37798 11784
rect 37921 11781 37933 11784
rect 37967 11781 37979 11815
rect 37921 11775 37979 11781
rect 40856 11815 40914 11821
rect 40856 11781 40868 11815
rect 40902 11812 40914 11815
rect 41506 11812 41512 11824
rect 40902 11784 41512 11812
rect 40902 11781 40914 11784
rect 40856 11775 40914 11781
rect 41506 11772 41512 11784
rect 41564 11772 41570 11824
rect 46201 11815 46259 11821
rect 46201 11812 46213 11815
rect 42812 11784 46213 11812
rect 42812 11756 42840 11784
rect 46201 11781 46213 11784
rect 46247 11812 46259 11815
rect 46474 11812 46480 11824
rect 46247 11784 46480 11812
rect 46247 11781 46259 11784
rect 46201 11775 46259 11781
rect 46474 11772 46480 11784
rect 46532 11772 46538 11824
rect 55950 11812 55956 11824
rect 48516 11784 55956 11812
rect 35529 11747 35587 11753
rect 35529 11744 35541 11747
rect 35400 11716 35541 11744
rect 35400 11704 35406 11716
rect 35529 11713 35541 11716
rect 35575 11713 35587 11747
rect 35529 11707 35587 11713
rect 35796 11747 35854 11753
rect 35796 11713 35808 11747
rect 35842 11744 35854 11747
rect 36630 11744 36636 11756
rect 35842 11716 36636 11744
rect 35842 11713 35854 11716
rect 35796 11707 35854 11713
rect 36630 11704 36636 11716
rect 36688 11704 36694 11756
rect 37642 11704 37648 11756
rect 37700 11744 37706 11756
rect 37700 11716 38240 11744
rect 37700 11704 37706 11716
rect 29546 11636 29552 11688
rect 29604 11636 29610 11688
rect 30926 11636 30932 11688
rect 30984 11676 30990 11688
rect 31757 11679 31815 11685
rect 31757 11676 31769 11679
rect 30984 11648 31769 11676
rect 30984 11636 30990 11648
rect 31757 11645 31769 11648
rect 31803 11645 31815 11679
rect 31757 11639 31815 11645
rect 31846 11636 31852 11688
rect 31904 11636 31910 11688
rect 32214 11636 32220 11688
rect 32272 11676 32278 11688
rect 32784 11676 32812 11704
rect 38212 11688 38240 11716
rect 42794 11704 42800 11756
rect 42852 11704 42858 11756
rect 44352 11747 44410 11753
rect 44352 11713 44364 11747
rect 44398 11744 44410 11747
rect 45186 11744 45192 11756
rect 44398 11716 45192 11744
rect 44398 11713 44410 11716
rect 44352 11707 44410 11713
rect 45186 11704 45192 11716
rect 45244 11704 45250 11756
rect 45925 11747 45983 11753
rect 45925 11713 45937 11747
rect 45971 11744 45983 11747
rect 46658 11744 46664 11756
rect 45971 11716 46664 11744
rect 45971 11713 45983 11716
rect 45925 11707 45983 11713
rect 46658 11704 46664 11716
rect 46716 11704 46722 11756
rect 32272 11648 32812 11676
rect 32272 11636 32278 11648
rect 34514 11636 34520 11688
rect 34572 11676 34578 11688
rect 34701 11679 34759 11685
rect 34701 11676 34713 11679
rect 34572 11648 34713 11676
rect 34572 11636 34578 11648
rect 34701 11645 34713 11648
rect 34747 11645 34759 11679
rect 34701 11639 34759 11645
rect 29086 11608 29092 11620
rect 22066 11580 29092 11608
rect 29086 11568 29092 11580
rect 29144 11568 29150 11620
rect 34716 11608 34744 11639
rect 38010 11636 38016 11688
rect 38068 11636 38074 11688
rect 38194 11636 38200 11688
rect 38252 11676 38258 11688
rect 40586 11676 40592 11688
rect 38252 11648 40592 11676
rect 38252 11636 38258 11648
rect 40586 11636 40592 11648
rect 40644 11636 40650 11688
rect 42886 11636 42892 11688
rect 42944 11676 42950 11688
rect 44082 11676 44088 11688
rect 42944 11648 44088 11676
rect 42944 11636 42950 11648
rect 44082 11636 44088 11648
rect 44140 11636 44146 11688
rect 39114 11608 39120 11620
rect 34716 11580 35572 11608
rect 23014 11500 23020 11552
rect 23072 11540 23078 11552
rect 28534 11540 28540 11552
rect 23072 11512 28540 11540
rect 23072 11500 23078 11512
rect 28534 11500 28540 11512
rect 28592 11500 28598 11552
rect 28810 11500 28816 11552
rect 28868 11540 28874 11552
rect 31846 11540 31852 11552
rect 28868 11512 31852 11540
rect 28868 11500 28874 11512
rect 31846 11500 31852 11512
rect 31904 11500 31910 11552
rect 35069 11543 35127 11549
rect 35069 11509 35081 11543
rect 35115 11540 35127 11543
rect 35434 11540 35440 11552
rect 35115 11512 35440 11540
rect 35115 11509 35127 11512
rect 35069 11503 35127 11509
rect 35434 11500 35440 11512
rect 35492 11500 35498 11552
rect 35544 11540 35572 11580
rect 36832 11580 39120 11608
rect 36832 11540 36860 11580
rect 39114 11568 39120 11580
rect 39172 11568 39178 11620
rect 48516 11608 48544 11784
rect 55950 11772 55956 11784
rect 56008 11772 56014 11824
rect 48774 11704 48780 11756
rect 48832 11744 48838 11756
rect 49145 11747 49203 11753
rect 49145 11744 49157 11747
rect 48832 11716 49157 11744
rect 48832 11704 48838 11716
rect 49145 11713 49157 11716
rect 49191 11713 49203 11747
rect 49145 11707 49203 11713
rect 49513 11747 49571 11753
rect 49513 11713 49525 11747
rect 49559 11744 49571 11747
rect 54202 11744 54208 11756
rect 49559 11716 54208 11744
rect 49559 11713 49571 11716
rect 49513 11707 49571 11713
rect 54202 11704 54208 11716
rect 54260 11704 54266 11756
rect 56502 11704 56508 11756
rect 56560 11704 56566 11756
rect 58066 11704 58072 11756
rect 58124 11704 58130 11756
rect 49050 11636 49056 11688
rect 49108 11636 49114 11688
rect 49605 11679 49663 11685
rect 49605 11645 49617 11679
rect 49651 11645 49663 11679
rect 49605 11639 49663 11645
rect 48593 11611 48651 11617
rect 48593 11608 48605 11611
rect 41892 11580 44128 11608
rect 35544 11512 36860 11540
rect 36909 11543 36967 11549
rect 36909 11509 36921 11543
rect 36955 11540 36967 11543
rect 37550 11540 37556 11552
rect 36955 11512 37556 11540
rect 36955 11509 36967 11512
rect 36909 11503 36967 11509
rect 37550 11500 37556 11512
rect 37608 11500 37614 11552
rect 37734 11500 37740 11552
rect 37792 11540 37798 11552
rect 41892 11540 41920 11580
rect 37792 11512 41920 11540
rect 37792 11500 37798 11512
rect 41966 11500 41972 11552
rect 42024 11500 42030 11552
rect 44100 11540 44128 11580
rect 45388 11580 48605 11608
rect 45388 11540 45416 11580
rect 48593 11577 48605 11580
rect 48639 11577 48651 11611
rect 48593 11571 48651 11577
rect 48866 11568 48872 11620
rect 48924 11608 48930 11620
rect 49620 11608 49648 11639
rect 56134 11636 56140 11688
rect 56192 11676 56198 11688
rect 56321 11679 56379 11685
rect 56321 11676 56333 11679
rect 56192 11648 56333 11676
rect 56192 11636 56198 11648
rect 56321 11645 56333 11648
rect 56367 11645 56379 11679
rect 56321 11639 56379 11645
rect 48924 11580 49648 11608
rect 48924 11568 48930 11580
rect 44100 11512 45416 11540
rect 45462 11500 45468 11552
rect 45520 11500 45526 11552
rect 48314 11500 48320 11552
rect 48372 11540 48378 11552
rect 58253 11543 58311 11549
rect 58253 11540 58265 11543
rect 48372 11512 58265 11540
rect 48372 11500 48378 11512
rect 58253 11509 58265 11512
rect 58299 11509 58311 11543
rect 58253 11503 58311 11509
rect 1104 11450 58880 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 58880 11450
rect 1104 11376 58880 11398
rect 13541 11339 13599 11345
rect 13541 11305 13553 11339
rect 13587 11336 13599 11339
rect 13630 11336 13636 11348
rect 13587 11308 13636 11336
rect 13587 11305 13599 11308
rect 13541 11299 13599 11305
rect 13630 11296 13636 11308
rect 13688 11296 13694 11348
rect 15470 11296 15476 11348
rect 15528 11296 15534 11348
rect 17221 11339 17279 11345
rect 17221 11305 17233 11339
rect 17267 11336 17279 11339
rect 18138 11336 18144 11348
rect 17267 11308 18144 11336
rect 17267 11305 17279 11308
rect 17221 11299 17279 11305
rect 18138 11296 18144 11308
rect 18196 11296 18202 11348
rect 19889 11339 19947 11345
rect 19889 11305 19901 11339
rect 19935 11336 19947 11339
rect 20622 11336 20628 11348
rect 19935 11308 20628 11336
rect 19935 11305 19947 11308
rect 19889 11299 19947 11305
rect 20622 11296 20628 11308
rect 20680 11296 20686 11348
rect 23293 11339 23351 11345
rect 23293 11305 23305 11339
rect 23339 11336 23351 11339
rect 23382 11336 23388 11348
rect 23339 11308 23388 11336
rect 23339 11305 23351 11308
rect 23293 11299 23351 11305
rect 23382 11296 23388 11308
rect 23440 11296 23446 11348
rect 29733 11339 29791 11345
rect 29733 11305 29745 11339
rect 29779 11336 29791 11339
rect 29822 11336 29828 11348
rect 29779 11308 29828 11336
rect 29779 11305 29791 11308
rect 29733 11299 29791 11305
rect 29822 11296 29828 11308
rect 29880 11296 29886 11348
rect 30466 11336 30472 11348
rect 30024 11308 30472 11336
rect 13170 11228 13176 11280
rect 13228 11268 13234 11280
rect 13357 11271 13415 11277
rect 13357 11268 13369 11271
rect 13228 11240 13369 11268
rect 13228 11228 13234 11240
rect 13357 11237 13369 11240
rect 13403 11237 13415 11271
rect 13357 11231 13415 11237
rect 14277 11203 14335 11209
rect 14277 11200 14289 11203
rect 6886 11172 14289 11200
rect 1581 11135 1639 11141
rect 1581 11101 1593 11135
rect 1627 11132 1639 11135
rect 6886 11132 6914 11172
rect 14277 11169 14289 11172
rect 14323 11169 14335 11203
rect 14277 11163 14335 11169
rect 14458 11160 14464 11212
rect 14516 11160 14522 11212
rect 14550 11160 14556 11212
rect 14608 11160 14614 11212
rect 14645 11203 14703 11209
rect 14645 11169 14657 11203
rect 14691 11200 14703 11203
rect 15488 11200 15516 11296
rect 15930 11228 15936 11280
rect 15988 11268 15994 11280
rect 17037 11271 17095 11277
rect 17037 11268 17049 11271
rect 15988 11240 17049 11268
rect 15988 11228 15994 11240
rect 17037 11237 17049 11240
rect 17083 11237 17095 11271
rect 17037 11231 17095 11237
rect 19705 11271 19763 11277
rect 19705 11237 19717 11271
rect 19751 11237 19763 11271
rect 19705 11231 19763 11237
rect 14691 11172 15516 11200
rect 14691 11169 14703 11172
rect 14645 11163 14703 11169
rect 16114 11160 16120 11212
rect 16172 11200 16178 11212
rect 19720 11200 19748 11231
rect 22186 11228 22192 11280
rect 22244 11268 22250 11280
rect 24765 11271 24823 11277
rect 24765 11268 24777 11271
rect 22244 11240 24777 11268
rect 22244 11228 22250 11240
rect 24765 11237 24777 11240
rect 24811 11237 24823 11271
rect 24765 11231 24823 11237
rect 28534 11228 28540 11280
rect 28592 11268 28598 11280
rect 30024 11268 30052 11308
rect 30466 11296 30472 11308
rect 30524 11296 30530 11348
rect 31404 11308 38700 11336
rect 28592 11240 30052 11268
rect 28592 11228 28598 11240
rect 30098 11228 30104 11280
rect 30156 11268 30162 11280
rect 31404 11277 31432 11308
rect 31389 11271 31447 11277
rect 30156 11240 31340 11268
rect 30156 11228 30162 11240
rect 16172 11172 19748 11200
rect 16172 11160 16178 11172
rect 23842 11160 23848 11212
rect 23900 11160 23906 11212
rect 29178 11200 29184 11212
rect 24504 11172 29184 11200
rect 1627 11104 6914 11132
rect 13081 11135 13139 11141
rect 1627 11101 1639 11104
rect 1581 11095 1639 11101
rect 13081 11101 13093 11135
rect 13127 11132 13139 11135
rect 13446 11132 13452 11144
rect 13127 11104 13452 11132
rect 13127 11101 13139 11104
rect 13081 11095 13139 11101
rect 13446 11092 13452 11104
rect 13504 11092 13510 11144
rect 14734 11092 14740 11144
rect 14792 11092 14798 11144
rect 15381 11135 15439 11141
rect 15381 11101 15393 11135
rect 15427 11132 15439 11135
rect 15838 11132 15844 11144
rect 15427 11104 15844 11132
rect 15427 11101 15439 11104
rect 15381 11095 15439 11101
rect 934 11024 940 11076
rect 992 11064 998 11076
rect 1857 11067 1915 11073
rect 1857 11064 1869 11067
rect 992 11036 1869 11064
rect 992 11024 998 11036
rect 1857 11033 1869 11036
rect 1903 11033 1915 11067
rect 1857 11027 1915 11033
rect 12434 11024 12440 11076
rect 12492 11064 12498 11076
rect 15396 11064 15424 11095
rect 15838 11092 15844 11104
rect 15896 11092 15902 11144
rect 23661 11135 23719 11141
rect 23661 11132 23673 11135
rect 15948 11104 23673 11132
rect 15948 11064 15976 11104
rect 23661 11101 23673 11104
rect 23707 11101 23719 11135
rect 23661 11095 23719 11101
rect 23753 11135 23811 11141
rect 23753 11101 23765 11135
rect 23799 11132 23811 11135
rect 24504 11132 24532 11172
rect 29178 11160 29184 11172
rect 29236 11160 29242 11212
rect 29822 11160 29828 11212
rect 29880 11200 29886 11212
rect 30926 11200 30932 11212
rect 29880 11172 30144 11200
rect 29880 11160 29886 11172
rect 23799 11104 24532 11132
rect 24581 11135 24639 11141
rect 23799 11101 23811 11104
rect 23753 11095 23811 11101
rect 24581 11101 24593 11135
rect 24627 11132 24639 11135
rect 27522 11132 27528 11144
rect 24627 11104 27528 11132
rect 24627 11101 24639 11104
rect 24581 11095 24639 11101
rect 27522 11092 27528 11104
rect 27580 11092 27586 11144
rect 28810 11092 28816 11144
rect 28868 11092 28874 11144
rect 28902 11092 28908 11144
rect 28960 11132 28966 11144
rect 29840 11132 29868 11160
rect 28960 11104 29868 11132
rect 28960 11092 28966 11104
rect 30006 11092 30012 11144
rect 30064 11092 30070 11144
rect 30116 11141 30144 11172
rect 30208 11172 30932 11200
rect 30101 11135 30159 11141
rect 30208 11138 30236 11172
rect 30926 11160 30932 11172
rect 30984 11160 30990 11212
rect 30101 11101 30113 11135
rect 30147 11101 30159 11135
rect 30101 11095 30159 11101
rect 30193 11132 30251 11138
rect 30193 11098 30205 11132
rect 30239 11098 30251 11132
rect 30193 11092 30251 11098
rect 30377 11135 30435 11141
rect 30377 11101 30389 11135
rect 30423 11132 30435 11135
rect 30466 11132 30472 11144
rect 30423 11104 30472 11132
rect 30423 11101 30435 11104
rect 30377 11095 30435 11101
rect 30466 11092 30472 11104
rect 30524 11092 30530 11144
rect 31312 11141 31340 11240
rect 31389 11237 31401 11271
rect 31435 11237 31447 11271
rect 36541 11271 36599 11277
rect 31389 11231 31447 11237
rect 31726 11240 35112 11268
rect 31297 11135 31355 11141
rect 31297 11101 31309 11135
rect 31343 11132 31355 11135
rect 31726 11132 31754 11240
rect 32122 11160 32128 11212
rect 32180 11160 32186 11212
rect 33226 11200 33232 11212
rect 32692 11172 33232 11200
rect 31343 11104 31754 11132
rect 31343 11101 31355 11104
rect 31297 11095 31355 11101
rect 31938 11092 31944 11144
rect 31996 11092 32002 11144
rect 32398 11092 32404 11144
rect 32456 11092 32462 11144
rect 12492 11036 15424 11064
rect 15488 11036 15976 11064
rect 16761 11067 16819 11073
rect 12492 11024 12498 11036
rect 15102 10956 15108 11008
rect 15160 10996 15166 11008
rect 15488 10996 15516 11036
rect 16761 11033 16773 11067
rect 16807 11064 16819 11067
rect 18046 11064 18052 11076
rect 16807 11036 18052 11064
rect 16807 11033 16819 11036
rect 16761 11027 16819 11033
rect 18046 11024 18052 11036
rect 18104 11064 18110 11076
rect 19429 11067 19487 11073
rect 19429 11064 19441 11067
rect 18104 11036 19441 11064
rect 18104 11024 18110 11036
rect 19429 11033 19441 11036
rect 19475 11064 19487 11067
rect 20438 11064 20444 11076
rect 19475 11036 20444 11064
rect 19475 11033 19487 11036
rect 19429 11027 19487 11033
rect 20438 11024 20444 11036
rect 20496 11064 20502 11076
rect 23842 11064 23848 11076
rect 20496 11036 23848 11064
rect 20496 11024 20502 11036
rect 23676 11008 23704 11036
rect 23842 11024 23848 11036
rect 23900 11024 23906 11076
rect 28997 11067 29055 11073
rect 28997 11033 29009 11067
rect 29043 11064 29055 11067
rect 29914 11064 29920 11076
rect 29043 11036 29920 11064
rect 29043 11033 29055 11036
rect 28997 11027 29055 11033
rect 29914 11024 29920 11036
rect 29972 11024 29978 11076
rect 30484 11064 30512 11092
rect 32692 11064 32720 11172
rect 33226 11160 33232 11172
rect 33284 11200 33290 11212
rect 33284 11172 34100 11200
rect 33284 11160 33290 11172
rect 32766 11092 32772 11144
rect 32824 11092 32830 11144
rect 33686 11092 33692 11144
rect 33744 11092 33750 11144
rect 34072 11141 34100 11172
rect 33781 11135 33839 11141
rect 33781 11101 33793 11135
rect 33827 11101 33839 11135
rect 33781 11095 33839 11101
rect 33873 11135 33931 11141
rect 33873 11101 33885 11135
rect 33919 11129 33931 11135
rect 34057 11135 34115 11141
rect 33919 11101 33988 11129
rect 33873 11095 33931 11101
rect 30484 11036 32720 11064
rect 32950 11024 32956 11076
rect 33008 11064 33014 11076
rect 33796 11064 33824 11095
rect 33960 11064 33988 11101
rect 34057 11101 34069 11135
rect 34103 11101 34115 11135
rect 34057 11095 34115 11101
rect 34146 11064 34152 11076
rect 33008 11036 33539 11064
rect 33796 11036 33916 11064
rect 33960 11036 34152 11064
rect 33008 11024 33014 11036
rect 15160 10968 15516 10996
rect 15160 10956 15166 10968
rect 23658 10956 23664 11008
rect 23716 10956 23722 11008
rect 27614 10956 27620 11008
rect 27672 10996 27678 11008
rect 27982 10996 27988 11008
rect 27672 10968 27988 10996
rect 27672 10956 27678 10968
rect 27982 10956 27988 10968
rect 28040 10956 28046 11008
rect 29086 10956 29092 11008
rect 29144 10996 29150 11008
rect 29181 10999 29239 11005
rect 29181 10996 29193 10999
rect 29144 10968 29193 10996
rect 29144 10956 29150 10968
rect 29181 10965 29193 10968
rect 29227 10965 29239 10999
rect 29181 10959 29239 10965
rect 33410 10956 33416 11008
rect 33468 10956 33474 11008
rect 33511 10996 33539 11036
rect 33888 10996 33916 11036
rect 34146 11024 34152 11036
rect 34204 11024 34210 11076
rect 35084 11064 35112 11240
rect 36541 11237 36553 11271
rect 36587 11268 36599 11271
rect 36587 11240 37412 11268
rect 36587 11237 36599 11240
rect 36541 11231 36599 11237
rect 35161 11135 35219 11141
rect 35161 11101 35173 11135
rect 35207 11132 35219 11135
rect 35250 11132 35256 11144
rect 35207 11104 35256 11132
rect 35207 11101 35219 11104
rect 35161 11095 35219 11101
rect 35250 11092 35256 11104
rect 35308 11092 35314 11144
rect 35434 11141 35440 11144
rect 35428 11132 35440 11141
rect 35395 11104 35440 11132
rect 35428 11095 35440 11104
rect 35434 11092 35440 11095
rect 35492 11092 35498 11144
rect 35710 11092 35716 11144
rect 35768 11132 35774 11144
rect 36556 11132 36584 11231
rect 37384 11141 37412 11240
rect 38102 11228 38108 11280
rect 38160 11228 38166 11280
rect 37461 11203 37519 11209
rect 37461 11169 37473 11203
rect 37507 11200 37519 11203
rect 37507 11172 38424 11200
rect 37507 11169 37519 11172
rect 37461 11163 37519 11169
rect 35768 11104 36584 11132
rect 37369 11135 37427 11141
rect 35768 11092 35774 11104
rect 37369 11101 37381 11135
rect 37415 11101 37427 11135
rect 38286 11132 38292 11144
rect 37369 11095 37427 11101
rect 37476 11104 38292 11132
rect 37476 11064 37504 11104
rect 38286 11092 38292 11104
rect 38344 11092 38350 11144
rect 38396 11141 38424 11172
rect 38672 11141 38700 11308
rect 45186 11296 45192 11348
rect 45244 11296 45250 11348
rect 48774 11296 48780 11348
rect 48832 11296 48838 11348
rect 43070 11228 43076 11280
rect 43128 11228 43134 11280
rect 46290 11228 46296 11280
rect 46348 11268 46354 11280
rect 49326 11268 49332 11280
rect 46348 11240 49332 11268
rect 46348 11228 46354 11240
rect 49326 11228 49332 11240
rect 49384 11228 49390 11280
rect 57241 11271 57299 11277
rect 57241 11268 57253 11271
rect 51046 11240 57253 11268
rect 40586 11160 40592 11212
rect 40644 11200 40650 11212
rect 41693 11203 41751 11209
rect 41693 11200 41705 11203
rect 40644 11172 41705 11200
rect 40644 11160 40650 11172
rect 41693 11169 41705 11172
rect 41739 11169 41751 11203
rect 41693 11163 41751 11169
rect 43990 11160 43996 11212
rect 44048 11200 44054 11212
rect 44048 11172 45784 11200
rect 44048 11160 44054 11172
rect 38381 11135 38439 11141
rect 38381 11101 38393 11135
rect 38427 11101 38439 11135
rect 38381 11095 38439 11101
rect 38565 11135 38623 11141
rect 38565 11101 38577 11135
rect 38611 11101 38623 11135
rect 38565 11095 38623 11101
rect 38657 11135 38715 11141
rect 38657 11101 38669 11135
rect 38703 11101 38715 11135
rect 38657 11095 38715 11101
rect 35084 11036 37504 11064
rect 38580 11064 38608 11095
rect 39114 11092 39120 11144
rect 39172 11092 39178 11144
rect 39298 11092 39304 11144
rect 39356 11092 39362 11144
rect 41960 11135 42018 11141
rect 41960 11101 41972 11135
rect 42006 11132 42018 11135
rect 42702 11132 42708 11144
rect 42006 11104 42708 11132
rect 42006 11101 42018 11104
rect 41960 11095 42018 11101
rect 42702 11092 42708 11104
rect 42760 11092 42766 11144
rect 45462 11132 45468 11144
rect 44928 11104 45468 11132
rect 39206 11064 39212 11076
rect 38580 11036 39212 11064
rect 39206 11024 39212 11036
rect 39264 11024 39270 11076
rect 39390 11024 39396 11076
rect 39448 11064 39454 11076
rect 44928 11064 44956 11104
rect 45462 11092 45468 11104
rect 45520 11132 45526 11144
rect 45649 11135 45707 11141
rect 45649 11132 45661 11135
rect 45520 11104 45661 11132
rect 45520 11092 45526 11104
rect 45649 11101 45661 11104
rect 45695 11101 45707 11135
rect 45756 11132 45784 11172
rect 45830 11160 45836 11212
rect 45888 11200 45894 11212
rect 46750 11200 46756 11212
rect 45888 11172 46756 11200
rect 45888 11160 45894 11172
rect 46750 11160 46756 11172
rect 46808 11160 46814 11212
rect 51046 11200 51074 11240
rect 57241 11237 57253 11240
rect 57287 11237 57299 11271
rect 57241 11231 57299 11237
rect 48332 11172 51074 11200
rect 45756 11104 45876 11132
rect 45649 11095 45707 11101
rect 39448 11036 44956 11064
rect 45557 11067 45615 11073
rect 39448 11024 39454 11036
rect 45557 11033 45569 11067
rect 45603 11064 45615 11067
rect 45738 11064 45744 11076
rect 45603 11036 45744 11064
rect 45603 11033 45615 11036
rect 45557 11027 45615 11033
rect 45738 11024 45744 11036
rect 45796 11024 45802 11076
rect 45848 11064 45876 11104
rect 46474 11092 46480 11144
rect 46532 11092 46538 11144
rect 46842 11092 46848 11144
rect 46900 11132 46906 11144
rect 48225 11135 48283 11141
rect 48225 11132 48237 11135
rect 46900 11104 48237 11132
rect 46900 11092 46906 11104
rect 48225 11101 48237 11104
rect 48271 11101 48283 11135
rect 48225 11095 48283 11101
rect 48332 11064 48360 11172
rect 58158 11160 58164 11212
rect 58216 11160 58222 11212
rect 48590 11092 48596 11144
rect 48648 11092 48654 11144
rect 51718 11092 51724 11144
rect 51776 11132 51782 11144
rect 57885 11135 57943 11141
rect 57885 11132 57897 11135
rect 51776 11104 57897 11132
rect 51776 11092 51782 11104
rect 57885 11101 57897 11104
rect 57931 11101 57943 11135
rect 57885 11095 57943 11101
rect 45848 11036 48360 11064
rect 48409 11067 48467 11073
rect 48409 11033 48421 11067
rect 48455 11033 48467 11067
rect 48409 11027 48467 11033
rect 48501 11067 48559 11073
rect 48501 11033 48513 11067
rect 48547 11064 48559 11067
rect 50798 11064 50804 11076
rect 48547 11036 50804 11064
rect 48547 11033 48559 11036
rect 48501 11027 48559 11033
rect 37366 10996 37372 11008
rect 33511 10968 37372 10996
rect 37366 10956 37372 10968
rect 37424 10956 37430 11008
rect 39482 10956 39488 11008
rect 39540 10956 39546 11008
rect 39574 10956 39580 11008
rect 39632 10996 39638 11008
rect 44450 10996 44456 11008
rect 39632 10968 44456 10996
rect 39632 10956 39638 10968
rect 44450 10956 44456 10968
rect 44508 10956 44514 11008
rect 48429 10996 48457 11027
rect 50798 11024 50804 11036
rect 50856 11024 50862 11076
rect 57057 11067 57115 11073
rect 57057 11033 57069 11067
rect 57103 11064 57115 11067
rect 58894 11064 58900 11076
rect 57103 11036 58900 11064
rect 57103 11033 57115 11036
rect 57057 11027 57115 11033
rect 58894 11024 58900 11036
rect 58952 11024 58958 11076
rect 49234 10996 49240 11008
rect 48429 10968 49240 10996
rect 49234 10956 49240 10968
rect 49292 10956 49298 11008
rect 1104 10906 58880 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 50294 10906
rect 50346 10854 50358 10906
rect 50410 10854 50422 10906
rect 50474 10854 50486 10906
rect 50538 10854 50550 10906
rect 50602 10854 58880 10906
rect 1104 10832 58880 10854
rect 12897 10795 12955 10801
rect 12897 10761 12909 10795
rect 12943 10792 12955 10795
rect 13538 10792 13544 10804
rect 12943 10764 13544 10792
rect 12943 10761 12955 10764
rect 12897 10755 12955 10761
rect 13538 10752 13544 10764
rect 13596 10752 13602 10804
rect 13817 10795 13875 10801
rect 13817 10761 13829 10795
rect 13863 10792 13875 10795
rect 14734 10792 14740 10804
rect 13863 10764 14740 10792
rect 13863 10761 13875 10764
rect 13817 10755 13875 10761
rect 14734 10752 14740 10764
rect 14792 10752 14798 10804
rect 23382 10792 23388 10804
rect 22066 10764 23388 10792
rect 2682 10684 2688 10736
rect 2740 10724 2746 10736
rect 22066 10724 22094 10764
rect 23382 10752 23388 10764
rect 23440 10752 23446 10804
rect 23477 10795 23535 10801
rect 23477 10761 23489 10795
rect 23523 10792 23535 10795
rect 23750 10792 23756 10804
rect 23523 10764 23756 10792
rect 23523 10761 23535 10764
rect 23477 10755 23535 10761
rect 23750 10752 23756 10764
rect 23808 10752 23814 10804
rect 25685 10795 25743 10801
rect 25685 10761 25697 10795
rect 25731 10792 25743 10795
rect 30006 10792 30012 10804
rect 25731 10764 30012 10792
rect 25731 10761 25743 10764
rect 25685 10755 25743 10761
rect 30006 10752 30012 10764
rect 30064 10752 30070 10804
rect 30282 10752 30288 10804
rect 30340 10792 30346 10804
rect 30377 10795 30435 10801
rect 30377 10792 30389 10795
rect 30340 10764 30389 10792
rect 30340 10752 30346 10764
rect 30377 10761 30389 10764
rect 30423 10761 30435 10795
rect 30377 10755 30435 10761
rect 30466 10752 30472 10804
rect 30524 10792 30530 10804
rect 30524 10764 34744 10792
rect 30524 10752 30530 10764
rect 28074 10724 28080 10736
rect 2740 10696 22094 10724
rect 23124 10696 28080 10724
rect 2740 10684 2746 10696
rect 1581 10659 1639 10665
rect 1581 10625 1593 10659
rect 1627 10656 1639 10659
rect 12342 10656 12348 10668
rect 1627 10628 12348 10656
rect 1627 10625 1639 10628
rect 1581 10619 1639 10625
rect 12342 10616 12348 10628
rect 12400 10616 12406 10668
rect 12434 10616 12440 10668
rect 12492 10616 12498 10668
rect 13357 10659 13415 10665
rect 13357 10625 13369 10659
rect 13403 10656 13415 10659
rect 13446 10656 13452 10668
rect 13403 10628 13452 10656
rect 13403 10625 13415 10628
rect 13357 10619 13415 10625
rect 13446 10616 13452 10628
rect 13504 10616 13510 10668
rect 18690 10616 18696 10668
rect 18748 10656 18754 10668
rect 23124 10656 23152 10696
rect 28074 10684 28080 10696
rect 28132 10684 28138 10736
rect 29086 10724 29092 10736
rect 28460 10696 29092 10724
rect 18748 10628 23152 10656
rect 23201 10659 23259 10665
rect 18748 10616 18754 10628
rect 23201 10625 23213 10659
rect 23247 10656 23259 10659
rect 23845 10659 23903 10665
rect 23845 10656 23857 10659
rect 23247 10628 23857 10656
rect 23247 10625 23259 10628
rect 23201 10619 23259 10625
rect 23845 10625 23857 10628
rect 23891 10625 23903 10659
rect 23845 10619 23903 10625
rect 934 10548 940 10600
rect 992 10588 998 10600
rect 1765 10591 1823 10597
rect 1765 10588 1777 10591
rect 992 10560 1777 10588
rect 992 10548 998 10560
rect 1765 10557 1777 10560
rect 1811 10557 1823 10591
rect 1765 10551 1823 10557
rect 12805 10523 12863 10529
rect 12805 10489 12817 10523
rect 12851 10489 12863 10523
rect 12805 10483 12863 10489
rect 12820 10452 12848 10483
rect 13078 10480 13084 10532
rect 13136 10520 13142 10532
rect 13633 10523 13691 10529
rect 13633 10520 13645 10523
rect 13136 10492 13645 10520
rect 13136 10480 13142 10492
rect 13633 10489 13645 10492
rect 13679 10489 13691 10523
rect 13633 10483 13691 10489
rect 13538 10452 13544 10464
rect 12820 10424 13544 10452
rect 13538 10412 13544 10424
rect 13596 10412 13602 10464
rect 17034 10412 17040 10464
rect 17092 10452 17098 10464
rect 23216 10452 23244 10619
rect 25406 10616 25412 10668
rect 25464 10656 25470 10668
rect 28169 10659 28227 10665
rect 28169 10656 28181 10659
rect 25464 10628 28181 10656
rect 25464 10616 25470 10628
rect 28169 10625 28181 10628
rect 28215 10625 28227 10659
rect 28169 10619 28227 10625
rect 28261 10659 28319 10665
rect 28261 10625 28273 10659
rect 28307 10625 28319 10659
rect 28261 10619 28319 10625
rect 28353 10659 28411 10665
rect 28460 10659 28488 10696
rect 29086 10684 29092 10696
rect 29144 10684 29150 10736
rect 30024 10724 30052 10752
rect 32944 10727 33002 10733
rect 30024 10696 32904 10724
rect 28353 10625 28365 10659
rect 28399 10631 28488 10659
rect 28399 10625 28411 10631
rect 28353 10619 28411 10625
rect 23934 10548 23940 10600
rect 23992 10548 23998 10600
rect 24029 10591 24087 10597
rect 24029 10557 24041 10591
rect 24075 10557 24087 10591
rect 24029 10551 24087 10557
rect 23658 10480 23664 10532
rect 23716 10520 23722 10532
rect 24044 10520 24072 10551
rect 25774 10548 25780 10600
rect 25832 10548 25838 10600
rect 25958 10548 25964 10600
rect 26016 10548 26022 10600
rect 27614 10520 27620 10532
rect 23716 10492 24072 10520
rect 24136 10492 27620 10520
rect 23716 10480 23722 10492
rect 17092 10424 23244 10452
rect 17092 10412 17098 10424
rect 23382 10412 23388 10464
rect 23440 10452 23446 10464
rect 24136 10452 24164 10492
rect 27614 10480 27620 10492
rect 27672 10480 27678 10532
rect 27706 10480 27712 10532
rect 27764 10520 27770 10532
rect 27893 10523 27951 10529
rect 27893 10520 27905 10523
rect 27764 10492 27905 10520
rect 27764 10480 27770 10492
rect 27893 10489 27905 10492
rect 27939 10489 27951 10523
rect 27893 10483 27951 10489
rect 23440 10424 24164 10452
rect 23440 10412 23446 10424
rect 25314 10412 25320 10464
rect 25372 10412 25378 10464
rect 28184 10452 28212 10619
rect 28276 10588 28304 10619
rect 28534 10616 28540 10668
rect 28592 10616 28598 10668
rect 28626 10616 28632 10668
rect 28684 10656 28690 10668
rect 29253 10659 29311 10665
rect 29253 10656 29265 10659
rect 28684 10628 29265 10656
rect 28684 10616 28690 10628
rect 29253 10625 29265 10628
rect 29299 10625 29311 10659
rect 29253 10619 29311 10625
rect 29546 10616 29552 10668
rect 29604 10656 29610 10668
rect 32876 10656 32904 10696
rect 32944 10693 32956 10727
rect 32990 10724 33002 10727
rect 33410 10724 33416 10736
rect 32990 10696 33416 10724
rect 32990 10693 33002 10696
rect 32944 10687 33002 10693
rect 33410 10684 33416 10696
rect 33468 10684 33474 10736
rect 34716 10724 34744 10764
rect 34790 10752 34796 10804
rect 34848 10792 34854 10804
rect 35437 10795 35495 10801
rect 35437 10792 35449 10795
rect 34848 10764 35449 10792
rect 34848 10752 34854 10764
rect 35437 10761 35449 10764
rect 35483 10761 35495 10795
rect 35437 10755 35495 10761
rect 35710 10752 35716 10804
rect 35768 10792 35774 10804
rect 35805 10795 35863 10801
rect 35805 10792 35817 10795
rect 35768 10764 35817 10792
rect 35768 10752 35774 10764
rect 35805 10761 35817 10764
rect 35851 10761 35863 10795
rect 35805 10755 35863 10761
rect 46385 10795 46443 10801
rect 46385 10761 46397 10795
rect 46431 10761 46443 10795
rect 46385 10755 46443 10761
rect 46753 10795 46811 10801
rect 46753 10761 46765 10795
rect 46799 10792 46811 10795
rect 59630 10792 59636 10804
rect 46799 10764 59636 10792
rect 46799 10761 46811 10764
rect 46753 10755 46811 10761
rect 38464 10727 38522 10733
rect 34716 10696 38424 10724
rect 35069 10659 35127 10665
rect 35069 10656 35081 10659
rect 29604 10628 31754 10656
rect 32876 10628 35081 10656
rect 29604 10616 29610 10628
rect 28276 10560 28488 10588
rect 28460 10520 28488 10560
rect 28994 10548 29000 10600
rect 29052 10548 29058 10600
rect 31726 10588 31754 10628
rect 35069 10625 35081 10628
rect 35115 10656 35127 10659
rect 35618 10656 35624 10668
rect 35115 10628 35624 10656
rect 35115 10625 35127 10628
rect 35069 10619 35127 10625
rect 35618 10616 35624 10628
rect 35676 10656 35682 10668
rect 35897 10659 35955 10665
rect 35897 10656 35909 10659
rect 35676 10628 35909 10656
rect 35676 10616 35682 10628
rect 35897 10625 35909 10628
rect 35943 10625 35955 10659
rect 35897 10619 35955 10625
rect 38194 10616 38200 10668
rect 38252 10616 38258 10668
rect 38396 10656 38424 10696
rect 38464 10693 38476 10727
rect 38510 10724 38522 10727
rect 39482 10724 39488 10736
rect 38510 10696 39488 10724
rect 38510 10693 38522 10696
rect 38464 10687 38522 10693
rect 39482 10684 39488 10696
rect 39540 10684 39546 10736
rect 44812 10727 44870 10733
rect 44812 10693 44824 10727
rect 44858 10724 44870 10727
rect 46400 10724 46428 10755
rect 59630 10752 59636 10764
rect 59688 10752 59694 10804
rect 44858 10696 46428 10724
rect 44858 10693 44870 10696
rect 44812 10687 44870 10693
rect 58069 10669 58127 10675
rect 39022 10656 39028 10668
rect 38396 10628 39028 10656
rect 39022 10616 39028 10628
rect 39080 10616 39086 10668
rect 40129 10659 40187 10665
rect 40129 10656 40141 10659
rect 39592 10628 40141 10656
rect 32674 10588 32680 10600
rect 31726 10560 32680 10588
rect 32674 10548 32680 10560
rect 32732 10548 32738 10600
rect 33686 10548 33692 10600
rect 33744 10588 33750 10600
rect 36081 10591 36139 10597
rect 36081 10588 36093 10591
rect 33744 10560 36093 10588
rect 33744 10548 33750 10560
rect 36081 10557 36093 10560
rect 36127 10588 36139 10591
rect 36127 10560 37596 10588
rect 36127 10557 36139 10560
rect 36081 10551 36139 10557
rect 28810 10520 28816 10532
rect 28460 10492 28816 10520
rect 28810 10480 28816 10492
rect 28868 10480 28874 10532
rect 30466 10452 30472 10464
rect 28184 10424 30472 10452
rect 30466 10412 30472 10424
rect 30524 10412 30530 10464
rect 32398 10412 32404 10464
rect 32456 10452 32462 10464
rect 34057 10455 34115 10461
rect 34057 10452 34069 10455
rect 32456 10424 34069 10452
rect 32456 10412 32462 10424
rect 34057 10421 34069 10424
rect 34103 10421 34115 10455
rect 37568 10452 37596 10560
rect 39592 10464 39620 10628
rect 40129 10625 40141 10628
rect 40175 10625 40187 10659
rect 40129 10619 40187 10625
rect 46750 10616 46756 10668
rect 46808 10656 46814 10668
rect 46808 10628 46980 10656
rect 46808 10616 46814 10628
rect 44082 10548 44088 10600
rect 44140 10588 44146 10600
rect 44542 10588 44548 10600
rect 44140 10560 44548 10588
rect 44140 10548 44146 10560
rect 44542 10548 44548 10560
rect 44600 10548 44606 10600
rect 46952 10597 46980 10628
rect 56042 10616 56048 10668
rect 56100 10656 56106 10668
rect 56321 10659 56379 10665
rect 56321 10656 56333 10659
rect 56100 10628 56333 10656
rect 56100 10616 56106 10628
rect 56321 10625 56333 10628
rect 56367 10625 56379 10659
rect 56321 10619 56379 10625
rect 56502 10616 56508 10668
rect 56560 10616 56566 10668
rect 56594 10616 56600 10668
rect 56652 10616 56658 10668
rect 57054 10616 57060 10668
rect 57112 10616 57118 10668
rect 58069 10666 58081 10669
rect 57946 10656 58081 10666
rect 57164 10638 58081 10656
rect 57164 10628 57974 10638
rect 58069 10635 58081 10638
rect 58115 10635 58127 10669
rect 58069 10629 58127 10635
rect 46845 10591 46903 10597
rect 46845 10557 46857 10591
rect 46891 10557 46903 10591
rect 46845 10551 46903 10557
rect 46937 10591 46995 10597
rect 46937 10557 46949 10591
rect 46983 10557 46995 10591
rect 46937 10551 46995 10557
rect 38378 10452 38384 10464
rect 37568 10424 38384 10452
rect 34057 10415 34115 10421
rect 38378 10412 38384 10424
rect 38436 10412 38442 10464
rect 39574 10412 39580 10464
rect 39632 10412 39638 10464
rect 40218 10412 40224 10464
rect 40276 10412 40282 10464
rect 44818 10412 44824 10464
rect 44876 10452 44882 10464
rect 45925 10455 45983 10461
rect 45925 10452 45937 10455
rect 44876 10424 45937 10452
rect 44876 10412 44882 10424
rect 45925 10421 45937 10424
rect 45971 10452 45983 10455
rect 46860 10452 46888 10551
rect 56410 10548 56416 10600
rect 56468 10588 56474 10600
rect 57164 10588 57192 10628
rect 58250 10616 58256 10668
rect 58308 10616 58314 10668
rect 56468 10560 57192 10588
rect 57333 10591 57391 10597
rect 56468 10548 56474 10560
rect 57333 10557 57345 10591
rect 57379 10588 57391 10591
rect 57882 10588 57888 10600
rect 57379 10560 57888 10588
rect 57379 10557 57391 10560
rect 57333 10551 57391 10557
rect 57882 10548 57888 10560
rect 57940 10548 57946 10600
rect 56502 10480 56508 10532
rect 56560 10520 56566 10532
rect 58161 10523 58219 10529
rect 58161 10520 58173 10523
rect 56560 10492 58173 10520
rect 56560 10480 56566 10492
rect 58161 10489 58173 10492
rect 58207 10489 58219 10523
rect 58161 10483 58219 10489
rect 45971 10424 46888 10452
rect 56321 10455 56379 10461
rect 45971 10421 45983 10424
rect 45925 10415 45983 10421
rect 56321 10421 56333 10455
rect 56367 10452 56379 10455
rect 56870 10452 56876 10464
rect 56367 10424 56876 10452
rect 56367 10421 56379 10424
rect 56321 10415 56379 10421
rect 56870 10412 56876 10424
rect 56928 10412 56934 10464
rect 57974 10412 57980 10464
rect 58032 10452 58038 10464
rect 58986 10452 58992 10464
rect 58032 10424 58992 10452
rect 58032 10412 58038 10424
rect 58986 10412 58992 10424
rect 59044 10412 59050 10464
rect 1104 10362 58880 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 58880 10362
rect 1104 10288 58880 10310
rect 12342 10208 12348 10260
rect 12400 10208 12406 10260
rect 23934 10208 23940 10260
rect 23992 10248 23998 10260
rect 23992 10220 31754 10248
rect 23992 10208 23998 10220
rect 23566 10140 23572 10192
rect 23624 10140 23630 10192
rect 26050 10140 26056 10192
rect 26108 10180 26114 10192
rect 27249 10183 27307 10189
rect 27249 10180 27261 10183
rect 26108 10152 27261 10180
rect 26108 10140 26114 10152
rect 27249 10149 27261 10152
rect 27295 10149 27307 10183
rect 27249 10143 27307 10149
rect 27522 10140 27528 10192
rect 27580 10180 27586 10192
rect 28261 10183 28319 10189
rect 28261 10180 28273 10183
rect 27580 10152 28273 10180
rect 27580 10140 27586 10152
rect 28261 10149 28273 10152
rect 28307 10149 28319 10183
rect 31726 10180 31754 10220
rect 32674 10208 32680 10260
rect 32732 10208 32738 10260
rect 38565 10251 38623 10257
rect 38565 10217 38577 10251
rect 38611 10248 38623 10251
rect 39298 10248 39304 10260
rect 38611 10220 39304 10248
rect 38611 10217 38623 10220
rect 38565 10211 38623 10217
rect 39298 10208 39304 10220
rect 39356 10208 39362 10260
rect 45830 10208 45836 10260
rect 45888 10248 45894 10260
rect 46569 10251 46627 10257
rect 46569 10248 46581 10251
rect 45888 10220 46581 10248
rect 45888 10208 45894 10220
rect 46569 10217 46581 10220
rect 46615 10217 46627 10251
rect 46569 10211 46627 10217
rect 57054 10208 57060 10260
rect 57112 10248 57118 10260
rect 58161 10251 58219 10257
rect 58161 10248 58173 10251
rect 57112 10220 58173 10248
rect 57112 10208 57118 10220
rect 58161 10217 58173 10220
rect 58207 10248 58219 10251
rect 58250 10248 58256 10260
rect 58207 10220 58256 10248
rect 58207 10217 58219 10220
rect 58161 10211 58219 10217
rect 58250 10208 58256 10220
rect 58308 10208 58314 10260
rect 39574 10180 39580 10192
rect 31726 10152 39580 10180
rect 28261 10143 28319 10149
rect 12526 10072 12532 10124
rect 12584 10072 12590 10124
rect 12618 10072 12624 10124
rect 12676 10072 12682 10124
rect 25958 10072 25964 10124
rect 26016 10112 26022 10124
rect 26016 10084 31754 10112
rect 26016 10072 26022 10084
rect 1581 10047 1639 10053
rect 1581 10013 1593 10047
rect 1627 10044 1639 10047
rect 12342 10044 12348 10056
rect 1627 10016 12348 10044
rect 1627 10013 1639 10016
rect 1581 10007 1639 10013
rect 12342 10004 12348 10016
rect 12400 10004 12406 10056
rect 12434 10004 12440 10056
rect 12492 10044 12498 10056
rect 12713 10047 12771 10053
rect 12713 10044 12725 10047
rect 12492 10016 12725 10044
rect 12492 10004 12498 10016
rect 12713 10013 12725 10016
rect 12759 10013 12771 10047
rect 12713 10007 12771 10013
rect 12805 10047 12863 10053
rect 12805 10013 12817 10047
rect 12851 10044 12863 10047
rect 13814 10044 13820 10056
rect 12851 10016 13820 10044
rect 12851 10013 12863 10016
rect 12805 10007 12863 10013
rect 934 9936 940 9988
rect 992 9976 998 9988
rect 1857 9979 1915 9985
rect 1857 9976 1869 9979
rect 992 9948 1869 9976
rect 992 9936 998 9948
rect 1857 9945 1869 9948
rect 1903 9945 1915 9979
rect 12728 9976 12756 10007
rect 13814 10004 13820 10016
rect 13872 10004 13878 10056
rect 24578 10004 24584 10056
rect 24636 10004 24642 10056
rect 24848 10047 24906 10053
rect 24848 10013 24860 10047
rect 24894 10044 24906 10047
rect 25314 10044 25320 10056
rect 24894 10016 25320 10044
rect 24894 10013 24906 10016
rect 24848 10007 24906 10013
rect 25314 10004 25320 10016
rect 25372 10004 25378 10056
rect 27065 10047 27123 10053
rect 27065 10013 27077 10047
rect 27111 10013 27123 10047
rect 27065 10007 27123 10013
rect 13354 9976 13360 9988
rect 12728 9948 13360 9976
rect 1857 9939 1915 9945
rect 13354 9936 13360 9948
rect 13412 9936 13418 9988
rect 23385 9979 23443 9985
rect 23385 9945 23397 9979
rect 23431 9976 23443 9979
rect 25222 9976 25228 9988
rect 23431 9948 25228 9976
rect 23431 9945 23443 9948
rect 23385 9939 23443 9945
rect 25222 9936 25228 9948
rect 25280 9936 25286 9988
rect 27080 9976 27108 10007
rect 28074 10004 28080 10056
rect 28132 10044 28138 10056
rect 30374 10044 30380 10056
rect 28132 10016 30380 10044
rect 28132 10004 28138 10016
rect 30374 10004 30380 10016
rect 30432 10004 30438 10056
rect 31726 10044 31754 10084
rect 33226 10072 33232 10124
rect 33284 10112 33290 10124
rect 35621 10115 35679 10121
rect 35621 10112 35633 10115
rect 33284 10084 35633 10112
rect 33284 10072 33290 10084
rect 35621 10081 35633 10084
rect 35667 10081 35679 10115
rect 35621 10075 35679 10081
rect 36357 10047 36415 10053
rect 36357 10044 36369 10047
rect 31726 10016 36369 10044
rect 36357 10013 36369 10016
rect 36403 10044 36415 10047
rect 38562 10044 38568 10056
rect 36403 10016 38568 10044
rect 36403 10013 36415 10016
rect 36357 10007 36415 10013
rect 38562 10004 38568 10016
rect 38620 10004 38626 10056
rect 38948 10053 38976 10152
rect 39574 10140 39580 10152
rect 39632 10140 39638 10192
rect 56045 10183 56103 10189
rect 56045 10149 56057 10183
rect 56091 10180 56103 10183
rect 56686 10180 56692 10192
rect 56091 10152 56692 10180
rect 56091 10149 56103 10152
rect 56045 10143 56103 10149
rect 56686 10140 56692 10152
rect 56744 10140 56750 10192
rect 39022 10072 39028 10124
rect 39080 10072 39086 10124
rect 39117 10115 39175 10121
rect 39117 10081 39129 10115
rect 39163 10081 39175 10115
rect 39117 10075 39175 10081
rect 38933 10047 38991 10053
rect 38933 10013 38945 10047
rect 38979 10013 38991 10047
rect 38933 10007 38991 10013
rect 28902 9976 28908 9988
rect 27080 9948 28908 9976
rect 28902 9936 28908 9948
rect 28960 9936 28966 9988
rect 31202 9936 31208 9988
rect 31260 9936 31266 9988
rect 32858 9936 32864 9988
rect 32916 9976 32922 9988
rect 34146 9976 34152 9988
rect 32916 9948 34152 9976
rect 32916 9936 32922 9948
rect 34146 9936 34152 9948
rect 34204 9936 34210 9988
rect 34330 9936 34336 9988
rect 34388 9976 34394 9988
rect 34885 9979 34943 9985
rect 34885 9976 34897 9979
rect 34388 9948 34897 9976
rect 34388 9936 34394 9948
rect 34885 9945 34897 9948
rect 34931 9976 34943 9979
rect 34931 9948 36400 9976
rect 34931 9945 34943 9948
rect 34885 9939 34943 9945
rect 23290 9868 23296 9920
rect 23348 9908 23354 9920
rect 25774 9908 25780 9920
rect 23348 9880 25780 9908
rect 23348 9868 23354 9880
rect 25774 9868 25780 9880
rect 25832 9908 25838 9920
rect 25961 9911 26019 9917
rect 25961 9908 25973 9911
rect 25832 9880 25973 9908
rect 25832 9868 25838 9880
rect 25961 9877 25973 9880
rect 26007 9877 26019 9911
rect 25961 9871 26019 9877
rect 29270 9868 29276 9920
rect 29328 9908 29334 9920
rect 36262 9908 36268 9920
rect 29328 9880 36268 9908
rect 29328 9868 29334 9880
rect 36262 9868 36268 9880
rect 36320 9868 36326 9920
rect 36372 9908 36400 9948
rect 36446 9936 36452 9988
rect 36504 9976 36510 9988
rect 36725 9979 36783 9985
rect 36725 9976 36737 9979
rect 36504 9948 36737 9976
rect 36504 9936 36510 9948
rect 36725 9945 36737 9948
rect 36771 9945 36783 9979
rect 36725 9939 36783 9945
rect 38378 9936 38384 9988
rect 38436 9976 38442 9988
rect 39132 9976 39160 10075
rect 56778 10072 56784 10124
rect 56836 10072 56842 10124
rect 44542 10004 44548 10056
rect 44600 10044 44606 10056
rect 45189 10047 45247 10053
rect 45189 10044 45201 10047
rect 44600 10016 45201 10044
rect 44600 10004 44606 10016
rect 45189 10013 45201 10016
rect 45235 10044 45247 10047
rect 47486 10044 47492 10056
rect 45235 10016 47492 10044
rect 45235 10013 45247 10016
rect 45189 10007 45247 10013
rect 47486 10004 47492 10016
rect 47544 10004 47550 10056
rect 56318 10004 56324 10056
rect 56376 10004 56382 10056
rect 56870 10004 56876 10056
rect 56928 10044 56934 10056
rect 57037 10047 57095 10053
rect 57037 10044 57049 10047
rect 56928 10016 57049 10044
rect 56928 10004 56934 10016
rect 57037 10013 57049 10016
rect 57083 10013 57095 10047
rect 57037 10007 57095 10013
rect 45462 9985 45468 9988
rect 38436 9948 39160 9976
rect 38436 9936 38442 9948
rect 45456 9939 45468 9985
rect 45462 9936 45468 9939
rect 45520 9936 45526 9988
rect 48314 9976 48320 9988
rect 46216 9948 48320 9976
rect 38010 9908 38016 9920
rect 36372 9880 38016 9908
rect 38010 9868 38016 9880
rect 38068 9868 38074 9920
rect 39022 9868 39028 9920
rect 39080 9908 39086 9920
rect 46216 9908 46244 9948
rect 48314 9936 48320 9948
rect 48372 9936 48378 9988
rect 56042 9936 56048 9988
rect 56100 9936 56106 9988
rect 39080 9880 46244 9908
rect 39080 9868 39086 9880
rect 56226 9868 56232 9920
rect 56284 9868 56290 9920
rect 1104 9818 58880 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 50294 9818
rect 50346 9766 50358 9818
rect 50410 9766 50422 9818
rect 50474 9766 50486 9818
rect 50538 9766 50550 9818
rect 50602 9766 58880 9818
rect 1104 9744 58880 9766
rect 17954 9664 17960 9716
rect 18012 9704 18018 9716
rect 18690 9704 18696 9716
rect 18012 9676 18696 9704
rect 18012 9664 18018 9676
rect 18690 9664 18696 9676
rect 18748 9664 18754 9716
rect 25222 9664 25228 9716
rect 25280 9704 25286 9716
rect 25317 9707 25375 9713
rect 25317 9704 25329 9707
rect 25280 9676 25329 9704
rect 25280 9664 25286 9676
rect 25317 9673 25329 9676
rect 25363 9673 25375 9707
rect 25317 9667 25375 9673
rect 28534 9664 28540 9716
rect 28592 9704 28598 9716
rect 30469 9707 30527 9713
rect 30469 9704 30481 9707
rect 28592 9676 29132 9704
rect 28592 9664 28598 9676
rect 23109 9639 23167 9645
rect 23109 9605 23121 9639
rect 23155 9636 23167 9639
rect 23566 9636 23572 9648
rect 23155 9608 23572 9636
rect 23155 9605 23167 9608
rect 23109 9599 23167 9605
rect 23566 9596 23572 9608
rect 23624 9596 23630 9648
rect 24578 9636 24584 9648
rect 23952 9608 24584 9636
rect 1581 9571 1639 9577
rect 1581 9537 1593 9571
rect 1627 9568 1639 9571
rect 12250 9568 12256 9580
rect 1627 9540 12256 9568
rect 1627 9537 1639 9540
rect 1581 9531 1639 9537
rect 12250 9528 12256 9540
rect 12308 9528 12314 9580
rect 12526 9528 12532 9580
rect 12584 9528 12590 9580
rect 12621 9571 12679 9577
rect 12621 9537 12633 9571
rect 12667 9568 12679 9571
rect 17310 9568 17316 9580
rect 12667 9540 17316 9568
rect 12667 9537 12679 9540
rect 12621 9531 12679 9537
rect 17310 9528 17316 9540
rect 17368 9528 17374 9580
rect 22738 9528 22744 9580
rect 22796 9568 22802 9580
rect 23014 9568 23020 9580
rect 22796 9540 23020 9568
rect 22796 9528 22802 9540
rect 23014 9528 23020 9540
rect 23072 9568 23078 9580
rect 23952 9577 23980 9608
rect 24578 9596 24584 9608
rect 24636 9636 24642 9648
rect 28994 9636 29000 9648
rect 24636 9608 29000 9636
rect 24636 9596 24642 9608
rect 27172 9580 27200 9608
rect 28994 9596 29000 9608
rect 29052 9596 29058 9648
rect 29104 9636 29132 9676
rect 30300 9676 30481 9704
rect 29454 9636 29460 9648
rect 29104 9608 29460 9636
rect 29454 9596 29460 9608
rect 29512 9596 29518 9648
rect 30190 9596 30196 9648
rect 30248 9636 30254 9648
rect 30300 9636 30328 9676
rect 30469 9673 30481 9676
rect 30515 9673 30527 9707
rect 30469 9667 30527 9673
rect 31018 9664 31024 9716
rect 31076 9704 31082 9716
rect 31076 9676 31432 9704
rect 31076 9664 31082 9676
rect 31404 9674 31432 9676
rect 31404 9646 31524 9674
rect 30248 9608 30328 9636
rect 30392 9608 31156 9636
rect 30248 9596 30254 9608
rect 23937 9571 23995 9577
rect 23072 9540 23336 9568
rect 23072 9528 23078 9540
rect 934 9460 940 9512
rect 992 9500 998 9512
rect 1765 9503 1823 9509
rect 1765 9500 1777 9503
rect 992 9472 1777 9500
rect 992 9460 998 9472
rect 1765 9469 1777 9472
rect 1811 9469 1823 9503
rect 1765 9463 1823 9469
rect 12342 9460 12348 9512
rect 12400 9460 12406 9512
rect 12713 9503 12771 9509
rect 12713 9500 12725 9503
rect 12636 9472 12725 9500
rect 12636 9444 12664 9472
rect 12713 9469 12725 9472
rect 12759 9469 12771 9503
rect 12713 9463 12771 9469
rect 12802 9460 12808 9512
rect 12860 9460 12866 9512
rect 13357 9503 13415 9509
rect 13357 9469 13369 9503
rect 13403 9469 13415 9503
rect 13357 9463 13415 9469
rect 12618 9392 12624 9444
rect 12676 9432 12682 9444
rect 13372 9432 13400 9463
rect 13814 9460 13820 9512
rect 13872 9460 13878 9512
rect 23198 9460 23204 9512
rect 23256 9460 23262 9512
rect 23308 9509 23336 9540
rect 23937 9537 23949 9571
rect 23983 9537 23995 9571
rect 24193 9571 24251 9577
rect 24193 9568 24205 9571
rect 23937 9531 23995 9537
rect 24044 9540 24205 9568
rect 23293 9503 23351 9509
rect 23293 9469 23305 9503
rect 23339 9469 23351 9503
rect 24044 9500 24072 9540
rect 24193 9537 24205 9540
rect 24239 9537 24251 9571
rect 24193 9531 24251 9537
rect 26326 9528 26332 9580
rect 26384 9528 26390 9580
rect 27154 9528 27160 9580
rect 27212 9528 27218 9580
rect 27424 9571 27482 9577
rect 27424 9537 27436 9571
rect 27470 9568 27482 9571
rect 27706 9568 27712 9580
rect 27470 9540 27712 9568
rect 27470 9537 27482 9540
rect 27424 9531 27482 9537
rect 27706 9528 27712 9540
rect 27764 9528 27770 9580
rect 27982 9528 27988 9580
rect 28040 9568 28046 9580
rect 29178 9568 29184 9580
rect 28040 9540 29184 9568
rect 28040 9528 28046 9540
rect 29178 9528 29184 9540
rect 29236 9528 29242 9580
rect 30282 9528 30288 9580
rect 30340 9528 30346 9580
rect 23293 9463 23351 9469
rect 23952 9472 24072 9500
rect 12676 9404 13400 9432
rect 13633 9435 13691 9441
rect 12676 9392 12682 9404
rect 13633 9401 13645 9435
rect 13679 9401 13691 9435
rect 13633 9395 13691 9401
rect 22741 9435 22799 9441
rect 22741 9401 22753 9435
rect 22787 9432 22799 9435
rect 23952 9432 23980 9472
rect 30006 9460 30012 9512
rect 30064 9500 30070 9512
rect 30392 9500 30420 9608
rect 30469 9571 30527 9577
rect 30469 9537 30481 9571
rect 30515 9568 30527 9571
rect 30515 9540 30880 9568
rect 30515 9537 30527 9540
rect 30469 9531 30527 9537
rect 30852 9512 30880 9540
rect 30926 9528 30932 9580
rect 30984 9570 30990 9580
rect 31128 9578 31156 9608
rect 31128 9577 31248 9578
rect 31025 9571 31083 9577
rect 31025 9570 31037 9571
rect 30984 9542 31037 9570
rect 30984 9528 30990 9542
rect 31025 9537 31037 9542
rect 31071 9537 31083 9571
rect 31128 9571 31263 9577
rect 31128 9550 31217 9571
rect 31025 9531 31083 9537
rect 31205 9537 31217 9550
rect 31251 9537 31263 9571
rect 31205 9531 31263 9537
rect 31297 9571 31355 9577
rect 31297 9537 31309 9571
rect 31343 9537 31355 9571
rect 31297 9531 31355 9537
rect 30064 9472 30420 9500
rect 30064 9460 30070 9472
rect 30834 9460 30840 9512
rect 30892 9460 30898 9512
rect 22787 9404 23980 9432
rect 22787 9401 22799 9404
rect 22741 9395 22799 9401
rect 12894 9324 12900 9376
rect 12952 9364 12958 9376
rect 13648 9364 13676 9395
rect 26142 9392 26148 9444
rect 26200 9432 26206 9444
rect 26513 9435 26571 9441
rect 26513 9432 26525 9435
rect 26200 9404 26525 9432
rect 26200 9392 26206 9404
rect 26513 9401 26525 9404
rect 26559 9401 26571 9435
rect 26513 9395 26571 9401
rect 28534 9392 28540 9444
rect 28592 9392 28598 9444
rect 28626 9392 28632 9444
rect 28684 9432 28690 9444
rect 29914 9432 29920 9444
rect 28684 9404 29920 9432
rect 28684 9392 28690 9404
rect 29914 9392 29920 9404
rect 29972 9392 29978 9444
rect 31110 9392 31116 9444
rect 31168 9432 31174 9444
rect 31312 9432 31340 9531
rect 31389 9503 31447 9509
rect 31389 9469 31401 9503
rect 31435 9500 31447 9503
rect 31496 9500 31524 9646
rect 31570 9634 31576 9686
rect 31628 9636 31634 9686
rect 32398 9664 32404 9716
rect 32456 9664 32462 9716
rect 45373 9707 45431 9713
rect 45373 9673 45385 9707
rect 45419 9704 45431 9707
rect 45462 9704 45468 9716
rect 45419 9676 45468 9704
rect 45419 9673 45431 9676
rect 45373 9667 45431 9673
rect 45462 9664 45468 9676
rect 45520 9664 45526 9716
rect 56226 9664 56232 9716
rect 56284 9704 56290 9716
rect 56505 9707 56563 9713
rect 56505 9704 56517 9707
rect 56284 9676 56517 9704
rect 56284 9664 56290 9676
rect 56505 9673 56517 9676
rect 56551 9673 56563 9707
rect 56505 9667 56563 9673
rect 32122 9636 32128 9648
rect 31628 9634 32128 9636
rect 31588 9608 32128 9634
rect 32122 9596 32128 9608
rect 32180 9596 32186 9648
rect 32416 9636 32444 9664
rect 32585 9639 32643 9645
rect 32585 9636 32597 9639
rect 32416 9608 32597 9636
rect 32585 9605 32597 9608
rect 32631 9605 32643 9639
rect 32585 9599 32643 9605
rect 32769 9639 32827 9645
rect 32769 9605 32781 9639
rect 32815 9636 32827 9639
rect 32858 9636 32864 9648
rect 32815 9608 32864 9636
rect 32815 9605 32827 9608
rect 32769 9599 32827 9605
rect 32858 9596 32864 9608
rect 32916 9596 32922 9648
rect 35618 9636 35624 9648
rect 34072 9608 35624 9636
rect 31570 9528 31576 9580
rect 31628 9528 31634 9580
rect 32401 9571 32459 9577
rect 32401 9537 32413 9571
rect 32447 9568 32459 9571
rect 32490 9568 32496 9580
rect 32447 9540 32496 9568
rect 32447 9537 32459 9540
rect 32401 9531 32459 9537
rect 32490 9528 32496 9540
rect 32548 9528 32554 9580
rect 33226 9528 33232 9580
rect 33284 9528 33290 9580
rect 33413 9571 33471 9577
rect 33413 9537 33425 9571
rect 33459 9568 33471 9571
rect 33686 9568 33692 9580
rect 33459 9540 33692 9568
rect 33459 9537 33471 9540
rect 33413 9531 33471 9537
rect 33686 9528 33692 9540
rect 33744 9528 33750 9580
rect 34072 9577 34100 9608
rect 35618 9596 35624 9608
rect 35676 9596 35682 9648
rect 35710 9596 35716 9648
rect 35768 9636 35774 9648
rect 36265 9639 36323 9645
rect 35768 9608 36032 9636
rect 35768 9596 35774 9608
rect 34057 9571 34115 9577
rect 34057 9537 34069 9571
rect 34103 9537 34115 9571
rect 34057 9531 34115 9537
rect 34324 9571 34382 9577
rect 34324 9537 34336 9571
rect 34370 9568 34382 9571
rect 36004 9568 36032 9608
rect 36265 9605 36277 9639
rect 36311 9636 36323 9639
rect 37090 9636 37096 9648
rect 36311 9608 37096 9636
rect 36311 9605 36323 9608
rect 36265 9599 36323 9605
rect 37090 9596 37096 9608
rect 37148 9596 37154 9648
rect 38838 9636 38844 9648
rect 37200 9608 38844 9636
rect 36357 9571 36415 9577
rect 36357 9568 36369 9571
rect 34370 9540 35940 9568
rect 36004 9540 36369 9568
rect 34370 9537 34382 9540
rect 34324 9531 34382 9537
rect 31435 9472 31524 9500
rect 31757 9503 31815 9509
rect 31435 9469 31447 9472
rect 31389 9463 31447 9469
rect 31757 9469 31769 9503
rect 31803 9500 31815 9503
rect 31803 9472 34100 9500
rect 31803 9469 31815 9472
rect 31757 9463 31815 9469
rect 31168 9404 31340 9432
rect 31404 9432 31432 9463
rect 31846 9432 31852 9444
rect 31404 9404 31852 9432
rect 31168 9392 31174 9404
rect 31846 9392 31852 9404
rect 31904 9392 31910 9444
rect 32398 9392 32404 9444
rect 32456 9432 32462 9444
rect 33597 9435 33655 9441
rect 33597 9432 33609 9435
rect 32456 9404 33609 9432
rect 32456 9392 32462 9404
rect 33597 9401 33609 9404
rect 33643 9401 33655 9435
rect 33597 9395 33655 9401
rect 12952 9336 13676 9364
rect 12952 9324 12958 9336
rect 24302 9324 24308 9376
rect 24360 9364 24366 9376
rect 26602 9364 26608 9376
rect 24360 9336 26608 9364
rect 24360 9324 24366 9336
rect 26602 9324 26608 9336
rect 26660 9324 26666 9376
rect 34072 9364 34100 9472
rect 35912 9441 35940 9540
rect 36357 9537 36369 9540
rect 36403 9537 36415 9571
rect 36357 9531 36415 9537
rect 36446 9460 36452 9512
rect 36504 9460 36510 9512
rect 35897 9435 35955 9441
rect 35176 9404 35848 9432
rect 35176 9364 35204 9404
rect 34072 9336 35204 9364
rect 35434 9324 35440 9376
rect 35492 9364 35498 9376
rect 35710 9364 35716 9376
rect 35492 9336 35716 9364
rect 35492 9324 35498 9336
rect 35710 9324 35716 9336
rect 35768 9324 35774 9376
rect 35820 9364 35848 9404
rect 35897 9401 35909 9435
rect 35943 9401 35955 9435
rect 35897 9395 35955 9401
rect 37200 9364 37228 9608
rect 38838 9596 38844 9608
rect 38896 9596 38902 9648
rect 40218 9636 40224 9648
rect 39132 9608 40224 9636
rect 38286 9528 38292 9580
rect 38344 9568 38350 9580
rect 39132 9577 39160 9608
rect 40218 9596 40224 9608
rect 40276 9596 40282 9648
rect 40862 9596 40868 9648
rect 40920 9636 40926 9648
rect 44634 9636 44640 9648
rect 40920 9608 44640 9636
rect 40920 9596 40926 9608
rect 44634 9596 44640 9608
rect 44692 9596 44698 9648
rect 45741 9639 45799 9645
rect 45741 9605 45753 9639
rect 45787 9636 45799 9639
rect 58802 9636 58808 9648
rect 45787 9608 58808 9636
rect 45787 9605 45799 9608
rect 45741 9599 45799 9605
rect 58802 9596 58808 9608
rect 58860 9596 58866 9648
rect 39025 9571 39083 9577
rect 39025 9568 39037 9571
rect 38344 9540 39037 9568
rect 38344 9528 38350 9540
rect 38856 9432 38884 9540
rect 39025 9537 39037 9540
rect 39071 9537 39083 9571
rect 39025 9531 39083 9537
rect 39117 9571 39175 9577
rect 39117 9537 39129 9571
rect 39163 9537 39175 9571
rect 39117 9531 39175 9537
rect 39298 9528 39304 9580
rect 39356 9528 39362 9580
rect 39393 9571 39451 9577
rect 39393 9537 39405 9571
rect 39439 9537 39451 9571
rect 39393 9531 39451 9537
rect 44177 9571 44235 9577
rect 44177 9537 44189 9571
rect 44223 9568 44235 9571
rect 44223 9540 51074 9568
rect 44223 9537 44235 9540
rect 44177 9531 44235 9537
rect 38930 9460 38936 9512
rect 38988 9500 38994 9512
rect 39408 9500 39436 9531
rect 43898 9500 43904 9512
rect 38988 9472 39436 9500
rect 41800 9472 43904 9500
rect 38988 9460 38994 9472
rect 41800 9432 41828 9472
rect 43898 9460 43904 9472
rect 43956 9500 43962 9512
rect 44453 9503 44511 9509
rect 44453 9500 44465 9503
rect 43956 9472 44465 9500
rect 43956 9460 43962 9472
rect 44453 9469 44465 9472
rect 44499 9469 44511 9503
rect 44453 9463 44511 9469
rect 45830 9460 45836 9512
rect 45888 9460 45894 9512
rect 46017 9503 46075 9509
rect 46017 9469 46029 9503
rect 46063 9500 46075 9503
rect 46750 9500 46756 9512
rect 46063 9472 46756 9500
rect 46063 9469 46075 9472
rect 46017 9463 46075 9469
rect 46750 9460 46756 9472
rect 46808 9460 46814 9512
rect 38856 9404 41828 9432
rect 41874 9392 41880 9444
rect 41932 9432 41938 9444
rect 45848 9432 45876 9460
rect 41932 9404 45876 9432
rect 51046 9432 51074 9540
rect 56410 9528 56416 9580
rect 56468 9528 56474 9580
rect 56597 9571 56655 9577
rect 56597 9537 56609 9571
rect 56643 9568 56655 9571
rect 57054 9568 57060 9580
rect 56643 9540 57060 9568
rect 56643 9537 56655 9540
rect 56597 9531 56655 9537
rect 57054 9528 57060 9540
rect 57112 9528 57118 9580
rect 57333 9503 57391 9509
rect 57333 9469 57345 9503
rect 57379 9500 57391 9503
rect 58986 9500 58992 9512
rect 57379 9472 58992 9500
rect 57379 9469 57391 9472
rect 57333 9463 57391 9469
rect 58986 9460 58992 9472
rect 59044 9460 59050 9512
rect 52086 9432 52092 9444
rect 51046 9404 52092 9432
rect 41932 9392 41938 9404
rect 52086 9392 52092 9404
rect 52144 9392 52150 9444
rect 35820 9336 37228 9364
rect 38841 9367 38899 9373
rect 38841 9333 38853 9367
rect 38887 9364 38899 9367
rect 56318 9364 56324 9376
rect 38887 9336 56324 9364
rect 38887 9333 38899 9336
rect 38841 9327 38899 9333
rect 56318 9324 56324 9336
rect 56376 9324 56382 9376
rect 1104 9274 58880 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 58880 9274
rect 1104 9200 58880 9222
rect 12250 9120 12256 9172
rect 12308 9120 12314 9172
rect 24302 9160 24308 9172
rect 12544 9132 24308 9160
rect 12544 9033 12572 9132
rect 24302 9120 24308 9132
rect 24360 9120 24366 9172
rect 25130 9120 25136 9172
rect 25188 9160 25194 9172
rect 26605 9163 26663 9169
rect 26605 9160 26617 9163
rect 25188 9132 26617 9160
rect 25188 9120 25194 9132
rect 26605 9129 26617 9132
rect 26651 9129 26663 9163
rect 26605 9123 26663 9129
rect 27338 9120 27344 9172
rect 27396 9160 27402 9172
rect 31021 9163 31079 9169
rect 27396 9132 28212 9160
rect 27396 9120 27402 9132
rect 25866 9092 25872 9104
rect 22066 9064 25872 9092
rect 12529 9027 12587 9033
rect 12529 8993 12541 9027
rect 12575 8993 12587 9027
rect 22066 9024 22094 9064
rect 25866 9052 25872 9064
rect 25924 9052 25930 9104
rect 23566 9024 23572 9036
rect 12529 8987 12587 8993
rect 15672 8996 22094 9024
rect 22940 8996 23572 9024
rect 1581 8959 1639 8965
rect 1581 8925 1593 8959
rect 1627 8956 1639 8959
rect 12158 8956 12164 8968
rect 1627 8928 12164 8956
rect 1627 8925 1639 8928
rect 1581 8919 1639 8925
rect 12158 8916 12164 8928
rect 12216 8916 12222 8968
rect 12437 8959 12495 8965
rect 12437 8925 12449 8959
rect 12483 8956 12495 8959
rect 12483 8928 12517 8956
rect 12483 8925 12495 8928
rect 12437 8919 12495 8925
rect 934 8848 940 8900
rect 992 8888 998 8900
rect 1857 8891 1915 8897
rect 1857 8888 1869 8891
rect 992 8860 1869 8888
rect 992 8848 998 8860
rect 1857 8857 1869 8860
rect 1903 8857 1915 8891
rect 1857 8851 1915 8857
rect 12342 8848 12348 8900
rect 12400 8888 12406 8900
rect 12452 8888 12480 8919
rect 12618 8916 12624 8968
rect 12676 8916 12682 8968
rect 12710 8916 12716 8968
rect 12768 8916 12774 8968
rect 15672 8888 15700 8996
rect 18414 8916 18420 8968
rect 18472 8956 18478 8968
rect 22830 8956 22836 8968
rect 18472 8928 22836 8956
rect 18472 8916 18478 8928
rect 22830 8916 22836 8928
rect 22888 8916 22894 8968
rect 22940 8965 22968 8996
rect 23566 8984 23572 8996
rect 23624 8984 23630 9036
rect 25682 8984 25688 9036
rect 25740 9024 25746 9036
rect 26970 9024 26976 9036
rect 25740 8996 26976 9024
rect 25740 8984 25746 8996
rect 26970 8984 26976 8996
rect 27028 8984 27034 9036
rect 27154 8984 27160 9036
rect 27212 8984 27218 9036
rect 28184 9024 28212 9132
rect 31021 9129 31033 9163
rect 31067 9129 31079 9163
rect 31021 9123 31079 9129
rect 28920 9064 29040 9092
rect 28920 9024 28948 9064
rect 28184 8996 28488 9024
rect 22925 8959 22983 8965
rect 22925 8925 22937 8959
rect 22971 8925 22983 8959
rect 22925 8919 22983 8925
rect 23014 8916 23020 8968
rect 23072 8916 23078 8968
rect 23106 8916 23112 8968
rect 23164 8956 23170 8968
rect 23201 8959 23259 8965
rect 23201 8956 23213 8959
rect 23164 8928 23213 8956
rect 23164 8916 23170 8928
rect 23201 8925 23213 8928
rect 23247 8925 23259 8959
rect 23201 8919 23259 8925
rect 25406 8916 25412 8968
rect 25464 8916 25470 8968
rect 26418 8916 26424 8968
rect 26476 8916 26482 8968
rect 28350 8956 28356 8968
rect 26528 8928 28356 8956
rect 12400 8860 15700 8888
rect 12400 8848 12406 8860
rect 17310 8848 17316 8900
rect 17368 8888 17374 8900
rect 26528 8888 26556 8928
rect 28350 8916 28356 8928
rect 28408 8916 28414 8968
rect 28460 8956 28488 8996
rect 28736 8996 28948 9024
rect 29012 9024 29040 9064
rect 29638 9052 29644 9104
rect 29696 9092 29702 9104
rect 31036 9092 31064 9123
rect 31478 9120 31484 9172
rect 31536 9160 31542 9172
rect 36446 9160 36452 9172
rect 31536 9132 36452 9160
rect 31536 9120 31542 9132
rect 36446 9120 36452 9132
rect 36504 9120 36510 9172
rect 36630 9120 36636 9172
rect 36688 9160 36694 9172
rect 39022 9160 39028 9172
rect 36688 9132 39028 9160
rect 36688 9120 36694 9132
rect 39022 9120 39028 9132
rect 39080 9160 39086 9172
rect 44085 9163 44143 9169
rect 44085 9160 44097 9163
rect 39080 9132 44097 9160
rect 39080 9120 39086 9132
rect 44085 9129 44097 9132
rect 44131 9160 44143 9163
rect 45186 9160 45192 9172
rect 44131 9132 45192 9160
rect 44131 9129 44143 9132
rect 44085 9123 44143 9129
rect 45186 9120 45192 9132
rect 45244 9120 45250 9172
rect 57054 9120 57060 9172
rect 57112 9160 57118 9172
rect 58161 9163 58219 9169
rect 58161 9160 58173 9163
rect 57112 9132 58173 9160
rect 57112 9120 57118 9132
rect 58161 9129 58173 9132
rect 58207 9129 58219 9163
rect 58161 9123 58219 9129
rect 44818 9092 44824 9104
rect 29696 9064 31064 9092
rect 35912 9064 44824 9092
rect 29696 9052 29702 9064
rect 29546 9024 29552 9036
rect 29012 8996 29552 9024
rect 28736 8956 28764 8996
rect 29012 8965 29040 8996
rect 29546 8984 29552 8996
rect 29604 8984 29610 9036
rect 29730 8984 29736 9036
rect 29788 9024 29794 9036
rect 30282 9024 30288 9036
rect 29788 8996 30288 9024
rect 29788 8984 29794 8996
rect 28460 8928 28764 8956
rect 28997 8959 29055 8965
rect 28997 8925 29009 8959
rect 29043 8925 29055 8959
rect 28997 8919 29055 8925
rect 29181 8959 29239 8965
rect 29181 8925 29193 8959
rect 29227 8956 29239 8959
rect 29638 8956 29644 8968
rect 29227 8928 29644 8956
rect 29227 8925 29239 8928
rect 29181 8919 29239 8925
rect 29638 8916 29644 8928
rect 29696 8916 29702 8968
rect 29822 8916 29828 8968
rect 29880 8956 29886 8968
rect 30116 8965 30144 8996
rect 30282 8984 30288 8996
rect 30340 8984 30346 9036
rect 34422 9024 34428 9036
rect 30392 8996 34428 9024
rect 30009 8959 30067 8965
rect 30009 8956 30021 8959
rect 29880 8928 30021 8956
rect 29880 8916 29886 8928
rect 30009 8925 30021 8928
rect 30055 8925 30067 8959
rect 30009 8919 30067 8925
rect 30101 8959 30159 8965
rect 30101 8925 30113 8959
rect 30147 8925 30159 8959
rect 30101 8919 30159 8925
rect 30190 8916 30196 8968
rect 30248 8916 30254 8968
rect 30392 8965 30420 8996
rect 34422 8984 34428 8996
rect 34480 8984 34486 9036
rect 30377 8959 30435 8965
rect 30377 8925 30389 8959
rect 30423 8925 30435 8959
rect 30377 8919 30435 8925
rect 30466 8916 30472 8968
rect 30524 8956 30530 8968
rect 30837 8959 30895 8965
rect 30837 8956 30849 8959
rect 30524 8928 30849 8956
rect 30524 8916 30530 8928
rect 30837 8925 30849 8928
rect 30883 8956 30895 8959
rect 31110 8956 31116 8968
rect 30883 8928 31116 8956
rect 30883 8925 30895 8928
rect 30837 8919 30895 8925
rect 31110 8916 31116 8928
rect 31168 8916 31174 8968
rect 31573 8959 31631 8965
rect 31573 8925 31585 8959
rect 31619 8925 31631 8959
rect 31573 8919 31631 8925
rect 17368 8860 26556 8888
rect 27424 8891 27482 8897
rect 17368 8848 17374 8860
rect 27424 8857 27436 8891
rect 27470 8888 27482 8891
rect 27798 8888 27804 8900
rect 27470 8860 27804 8888
rect 27470 8857 27482 8860
rect 27424 8851 27482 8857
rect 27798 8848 27804 8860
rect 27856 8848 27862 8900
rect 27982 8848 27988 8900
rect 28040 8888 28046 8900
rect 31478 8888 31484 8900
rect 28040 8860 31484 8888
rect 28040 8848 28046 8860
rect 31478 8848 31484 8860
rect 31536 8848 31542 8900
rect 31588 8832 31616 8919
rect 31662 8916 31668 8968
rect 31720 8916 31726 8968
rect 35342 8916 35348 8968
rect 35400 8956 35406 8968
rect 35529 8959 35587 8965
rect 35529 8956 35541 8959
rect 35400 8928 35541 8956
rect 35400 8916 35406 8928
rect 35529 8925 35541 8928
rect 35575 8925 35587 8959
rect 35529 8919 35587 8925
rect 35544 8888 35572 8919
rect 35802 8916 35808 8968
rect 35860 8916 35866 8968
rect 35912 8965 35940 9064
rect 44818 9052 44824 9064
rect 44876 9052 44882 9104
rect 35986 8984 35992 9036
rect 36044 9024 36050 9036
rect 36725 9027 36783 9033
rect 36725 9024 36737 9027
rect 36044 8996 36737 9024
rect 36044 8984 36050 8996
rect 36725 8993 36737 8996
rect 36771 8993 36783 9027
rect 36725 8987 36783 8993
rect 38562 8984 38568 9036
rect 38620 9024 38626 9036
rect 41233 9027 41291 9033
rect 41233 9024 41245 9027
rect 38620 8996 41245 9024
rect 38620 8984 38626 8996
rect 41233 8993 41245 8996
rect 41279 9024 41291 9027
rect 42794 9024 42800 9036
rect 41279 8996 42800 9024
rect 41279 8993 41291 8996
rect 41233 8987 41291 8993
rect 42794 8984 42800 8996
rect 42852 9024 42858 9036
rect 43254 9024 43260 9036
rect 42852 8996 43260 9024
rect 42852 8984 42858 8996
rect 43254 8984 43260 8996
rect 43312 8984 43318 9036
rect 48590 8984 48596 9036
rect 48648 9024 48654 9036
rect 48958 9024 48964 9036
rect 48648 8996 48964 9024
rect 48648 8984 48654 8996
rect 48958 8984 48964 8996
rect 49016 8984 49022 9036
rect 56778 8984 56784 9036
rect 56836 8984 56842 9036
rect 35897 8959 35955 8965
rect 35897 8925 35909 8959
rect 35943 8925 35955 8959
rect 37642 8956 37648 8968
rect 35897 8919 35955 8925
rect 36188 8928 37648 8956
rect 36188 8888 36216 8928
rect 37642 8916 37648 8928
rect 37700 8916 37706 8968
rect 41049 8959 41107 8965
rect 41049 8925 41061 8959
rect 41095 8956 41107 8959
rect 42334 8956 42340 8968
rect 41095 8928 42340 8956
rect 41095 8925 41107 8928
rect 41049 8919 41107 8925
rect 42334 8916 42340 8928
rect 42392 8916 42398 8968
rect 43898 8916 43904 8968
rect 43956 8956 43962 8968
rect 43993 8959 44051 8965
rect 43993 8956 44005 8959
rect 43956 8928 44005 8956
rect 43956 8916 43962 8928
rect 43993 8925 44005 8928
rect 44039 8956 44051 8959
rect 44358 8956 44364 8968
rect 44039 8928 44364 8956
rect 44039 8925 44051 8928
rect 43993 8919 44051 8925
rect 44358 8916 44364 8928
rect 44416 8916 44422 8968
rect 56686 8916 56692 8968
rect 56744 8956 56750 8968
rect 57037 8959 57095 8965
rect 57037 8956 57049 8959
rect 56744 8928 57049 8956
rect 56744 8916 56750 8928
rect 57037 8925 57049 8928
rect 57083 8925 57095 8959
rect 57037 8919 57095 8925
rect 35544 8860 36216 8888
rect 36262 8848 36268 8900
rect 36320 8848 36326 8900
rect 37918 8848 37924 8900
rect 37976 8888 37982 8900
rect 46198 8888 46204 8900
rect 37976 8860 46204 8888
rect 37976 8848 37982 8860
rect 46198 8848 46204 8860
rect 46256 8848 46262 8900
rect 48406 8848 48412 8900
rect 48464 8888 48470 8900
rect 48958 8888 48964 8900
rect 48464 8860 48964 8888
rect 48464 8848 48470 8860
rect 48958 8848 48964 8860
rect 49016 8848 49022 8900
rect 12434 8780 12440 8832
rect 12492 8820 12498 8832
rect 20530 8820 20536 8832
rect 12492 8792 20536 8820
rect 12492 8780 12498 8792
rect 20530 8780 20536 8792
rect 20588 8780 20594 8832
rect 25038 8780 25044 8832
rect 25096 8780 25102 8832
rect 25501 8823 25559 8829
rect 25501 8789 25513 8823
rect 25547 8820 25559 8823
rect 25590 8820 25596 8832
rect 25547 8792 25596 8820
rect 25547 8789 25559 8792
rect 25501 8783 25559 8789
rect 25590 8780 25596 8792
rect 25648 8780 25654 8832
rect 28258 8780 28264 8832
rect 28316 8820 28322 8832
rect 28537 8823 28595 8829
rect 28537 8820 28549 8823
rect 28316 8792 28549 8820
rect 28316 8780 28322 8792
rect 28537 8789 28549 8792
rect 28583 8789 28595 8823
rect 28537 8783 28595 8789
rect 29086 8780 29092 8832
rect 29144 8780 29150 8832
rect 29733 8823 29791 8829
rect 29733 8789 29745 8823
rect 29779 8820 29791 8823
rect 30282 8820 30288 8832
rect 29779 8792 30288 8820
rect 29779 8789 29791 8792
rect 29733 8783 29791 8789
rect 30282 8780 30288 8792
rect 30340 8780 30346 8832
rect 30374 8780 30380 8832
rect 30432 8820 30438 8832
rect 31570 8820 31576 8832
rect 30432 8792 31576 8820
rect 30432 8780 30438 8792
rect 31570 8780 31576 8792
rect 31628 8780 31634 8832
rect 33134 8780 33140 8832
rect 33192 8820 33198 8832
rect 33778 8820 33784 8832
rect 33192 8792 33784 8820
rect 33192 8780 33198 8792
rect 33778 8780 33784 8792
rect 33836 8780 33842 8832
rect 40678 8780 40684 8832
rect 40736 8780 40742 8832
rect 41138 8780 41144 8832
rect 41196 8780 41202 8832
rect 46106 8780 46112 8832
rect 46164 8820 46170 8832
rect 48774 8820 48780 8832
rect 46164 8792 48780 8820
rect 46164 8780 46170 8792
rect 48774 8780 48780 8792
rect 48832 8780 48838 8832
rect 1104 8730 58880 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 50294 8730
rect 50346 8678 50358 8730
rect 50410 8678 50422 8730
rect 50474 8678 50486 8730
rect 50538 8678 50550 8730
rect 50602 8678 58880 8730
rect 1104 8656 58880 8678
rect 11146 8616 11152 8628
rect 10796 8588 11152 8616
rect 10796 8489 10824 8588
rect 11146 8576 11152 8588
rect 11204 8616 11210 8628
rect 11330 8616 11336 8628
rect 11204 8588 11336 8616
rect 11204 8576 11210 8588
rect 11330 8576 11336 8588
rect 11388 8576 11394 8628
rect 12158 8576 12164 8628
rect 12216 8576 12222 8628
rect 23290 8616 23296 8628
rect 12360 8588 23296 8616
rect 12360 8548 12388 8588
rect 23290 8576 23296 8588
rect 23348 8576 23354 8628
rect 27706 8576 27712 8628
rect 27764 8616 27770 8628
rect 27893 8619 27951 8625
rect 27893 8616 27905 8619
rect 27764 8588 27905 8616
rect 27764 8576 27770 8588
rect 27893 8585 27905 8588
rect 27939 8585 27951 8619
rect 27893 8579 27951 8585
rect 28261 8619 28319 8625
rect 28261 8585 28273 8619
rect 28307 8616 28319 8619
rect 28442 8616 28448 8628
rect 28307 8588 28448 8616
rect 28307 8585 28319 8588
rect 28261 8579 28319 8585
rect 28442 8576 28448 8588
rect 28500 8576 28506 8628
rect 28902 8576 28908 8628
rect 28960 8616 28966 8628
rect 29457 8619 29515 8625
rect 29457 8616 29469 8619
rect 28960 8588 29469 8616
rect 28960 8576 28966 8588
rect 29457 8585 29469 8588
rect 29503 8585 29515 8619
rect 29457 8579 29515 8585
rect 29638 8576 29644 8628
rect 29696 8616 29702 8628
rect 30650 8616 30656 8628
rect 29696 8588 30656 8616
rect 29696 8576 29702 8588
rect 30650 8576 30656 8588
rect 30708 8576 30714 8628
rect 31570 8576 31576 8628
rect 31628 8576 31634 8628
rect 33042 8576 33048 8628
rect 33100 8616 33106 8628
rect 41138 8616 41144 8628
rect 33100 8588 34836 8616
rect 33100 8576 33106 8588
rect 10888 8520 12388 8548
rect 10888 8489 10916 8520
rect 12526 8508 12532 8560
rect 12584 8548 12590 8560
rect 13633 8551 13691 8557
rect 13633 8548 13645 8551
rect 12584 8520 13645 8548
rect 12584 8508 12590 8520
rect 13633 8517 13645 8520
rect 13679 8517 13691 8551
rect 24578 8548 24584 8560
rect 13633 8511 13691 8517
rect 24228 8520 24584 8548
rect 1581 8483 1639 8489
rect 1581 8449 1593 8483
rect 1627 8480 1639 8483
rect 10781 8483 10839 8489
rect 1627 8452 6914 8480
rect 1627 8449 1639 8452
rect 1581 8443 1639 8449
rect 934 8372 940 8424
rect 992 8412 998 8424
rect 1765 8415 1823 8421
rect 1765 8412 1777 8415
rect 992 8384 1777 8412
rect 992 8372 998 8384
rect 1765 8381 1777 8384
rect 1811 8381 1823 8415
rect 6886 8412 6914 8452
rect 10781 8449 10793 8483
rect 10827 8449 10839 8483
rect 10781 8443 10839 8449
rect 10873 8483 10931 8489
rect 10873 8449 10885 8483
rect 10919 8449 10931 8483
rect 10873 8443 10931 8449
rect 12342 8440 12348 8492
rect 12400 8440 12406 8492
rect 12434 8440 12440 8492
rect 12492 8440 12498 8492
rect 13265 8483 13323 8489
rect 13265 8449 13277 8483
rect 13311 8480 13323 8483
rect 13311 8452 13400 8480
rect 13311 8449 13323 8452
rect 13265 8443 13323 8449
rect 10597 8415 10655 8421
rect 10597 8412 10609 8415
rect 6886 8384 10609 8412
rect 1765 8375 1823 8381
rect 10597 8381 10609 8384
rect 10643 8381 10655 8415
rect 10597 8375 10655 8381
rect 10962 8372 10968 8424
rect 11020 8372 11026 8424
rect 11054 8372 11060 8424
rect 11112 8372 11118 8424
rect 12526 8372 12532 8424
rect 12584 8372 12590 8424
rect 12618 8372 12624 8424
rect 12676 8372 12682 8424
rect 10870 8304 10876 8356
rect 10928 8344 10934 8356
rect 13372 8344 13400 8452
rect 24118 8440 24124 8492
rect 24176 8480 24182 8492
rect 24228 8489 24256 8520
rect 24578 8508 24584 8520
rect 24636 8508 24642 8560
rect 24762 8508 24768 8560
rect 24820 8548 24826 8560
rect 27982 8548 27988 8560
rect 24820 8520 27988 8548
rect 24820 8508 24826 8520
rect 27982 8508 27988 8520
rect 28040 8508 28046 8560
rect 28966 8520 30144 8548
rect 24213 8483 24271 8489
rect 24213 8480 24225 8483
rect 24176 8452 24225 8480
rect 24176 8440 24182 8452
rect 24213 8449 24225 8452
rect 24259 8449 24271 8483
rect 24213 8443 24271 8449
rect 24480 8483 24538 8489
rect 24480 8449 24492 8483
rect 24526 8480 24538 8483
rect 25038 8480 25044 8492
rect 24526 8452 25044 8480
rect 24526 8449 24538 8452
rect 24480 8443 24538 8449
rect 25038 8440 25044 8452
rect 25096 8440 25102 8492
rect 27062 8440 27068 8492
rect 27120 8480 27126 8492
rect 28966 8480 28994 8520
rect 27120 8452 28994 8480
rect 27120 8440 27126 8452
rect 29270 8440 29276 8492
rect 29328 8440 29334 8492
rect 21174 8372 21180 8424
rect 21232 8412 21238 8424
rect 21542 8412 21548 8424
rect 21232 8384 21548 8412
rect 21232 8372 21238 8384
rect 21542 8372 21548 8384
rect 21600 8372 21606 8424
rect 28350 8372 28356 8424
rect 28408 8372 28414 8424
rect 28537 8415 28595 8421
rect 28537 8381 28549 8415
rect 28583 8412 28595 8415
rect 28626 8412 28632 8424
rect 28583 8384 28632 8412
rect 28583 8381 28595 8384
rect 28537 8375 28595 8381
rect 28626 8372 28632 8384
rect 28684 8372 28690 8424
rect 28994 8372 29000 8424
rect 29052 8412 29058 8424
rect 29914 8412 29920 8424
rect 29052 8384 29920 8412
rect 29052 8372 29058 8384
rect 29914 8372 29920 8384
rect 29972 8412 29978 8424
rect 30009 8415 30067 8421
rect 30009 8412 30021 8415
rect 29972 8384 30021 8412
rect 29972 8372 29978 8384
rect 30009 8381 30021 8384
rect 30055 8381 30067 8415
rect 30116 8412 30144 8520
rect 31846 8508 31852 8560
rect 31904 8548 31910 8560
rect 33597 8551 33655 8557
rect 33597 8548 33609 8551
rect 31904 8520 33609 8548
rect 31904 8508 31910 8520
rect 33597 8517 33609 8520
rect 33643 8517 33655 8551
rect 33597 8511 33655 8517
rect 33686 8508 33692 8560
rect 33744 8508 33750 8560
rect 30282 8440 30288 8492
rect 30340 8440 30346 8492
rect 30374 8440 30380 8492
rect 30432 8480 30438 8492
rect 31202 8480 31208 8492
rect 30432 8452 31208 8480
rect 30432 8440 30438 8452
rect 31202 8440 31208 8452
rect 31260 8480 31266 8492
rect 33134 8480 33140 8492
rect 31260 8452 33140 8480
rect 31260 8440 31266 8452
rect 33134 8440 33140 8452
rect 33192 8440 33198 8492
rect 33318 8440 33324 8492
rect 33376 8440 33382 8492
rect 33410 8440 33416 8492
rect 33468 8440 33474 8492
rect 33870 8489 33876 8492
rect 33827 8483 33876 8489
rect 33827 8449 33839 8483
rect 33873 8449 33876 8483
rect 33827 8443 33876 8449
rect 33870 8440 33876 8443
rect 33928 8440 33934 8492
rect 34606 8440 34612 8492
rect 34664 8480 34670 8492
rect 34808 8489 34836 8588
rect 35912 8588 41144 8616
rect 35526 8548 35532 8560
rect 34992 8520 35532 8548
rect 34992 8489 35020 8520
rect 35526 8508 35532 8520
rect 35584 8508 35590 8560
rect 35912 8557 35940 8588
rect 41138 8576 41144 8588
rect 41196 8616 41202 8628
rect 41417 8619 41475 8625
rect 41417 8616 41429 8619
rect 41196 8588 41429 8616
rect 41196 8576 41202 8588
rect 41417 8585 41429 8588
rect 41463 8585 41475 8619
rect 41417 8579 41475 8585
rect 46198 8576 46204 8628
rect 46256 8616 46262 8628
rect 58253 8619 58311 8625
rect 58253 8616 58265 8619
rect 46256 8588 58265 8616
rect 46256 8576 46262 8588
rect 58253 8585 58265 8588
rect 58299 8585 58311 8619
rect 58253 8579 58311 8585
rect 35897 8551 35955 8557
rect 35897 8517 35909 8551
rect 35943 8517 35955 8551
rect 35897 8511 35955 8517
rect 36170 8508 36176 8560
rect 36228 8548 36234 8560
rect 36265 8551 36323 8557
rect 36265 8548 36277 8551
rect 36228 8520 36277 8548
rect 36228 8508 36234 8520
rect 36265 8517 36277 8520
rect 36311 8517 36323 8551
rect 36265 8511 36323 8517
rect 40052 8520 41414 8548
rect 34701 8483 34759 8489
rect 34701 8480 34713 8483
rect 34664 8452 34713 8480
rect 34664 8440 34670 8452
rect 34701 8449 34713 8452
rect 34747 8449 34759 8483
rect 34701 8443 34759 8449
rect 34793 8483 34851 8489
rect 34793 8449 34805 8483
rect 34839 8449 34851 8483
rect 34793 8443 34851 8449
rect 34977 8483 35035 8489
rect 34977 8449 34989 8483
rect 35023 8449 35035 8483
rect 34977 8443 35035 8449
rect 35069 8483 35127 8489
rect 35069 8449 35081 8483
rect 35115 8449 35127 8483
rect 35069 8443 35127 8449
rect 35084 8412 35112 8443
rect 35802 8440 35808 8492
rect 35860 8440 35866 8492
rect 37461 8483 37519 8489
rect 37461 8449 37473 8483
rect 37507 8449 37519 8483
rect 37461 8443 37519 8449
rect 30116 8384 35112 8412
rect 30009 8375 30067 8381
rect 35342 8372 35348 8424
rect 35400 8412 35406 8424
rect 35529 8415 35587 8421
rect 35529 8412 35541 8415
rect 35400 8384 35541 8412
rect 35400 8372 35406 8384
rect 35529 8381 35541 8384
rect 35575 8381 35587 8415
rect 37476 8412 37504 8443
rect 39114 8440 39120 8492
rect 39172 8480 39178 8492
rect 40052 8489 40080 8520
rect 40037 8483 40095 8489
rect 40037 8480 40049 8483
rect 39172 8452 40049 8480
rect 39172 8440 39178 8452
rect 40037 8449 40049 8452
rect 40083 8449 40095 8483
rect 40037 8443 40095 8449
rect 40304 8483 40362 8489
rect 40304 8449 40316 8483
rect 40350 8480 40362 8483
rect 40678 8480 40684 8492
rect 40350 8452 40684 8480
rect 40350 8449 40362 8452
rect 40304 8443 40362 8449
rect 40678 8440 40684 8452
rect 40736 8440 40742 8492
rect 41386 8480 41414 8520
rect 47670 8508 47676 8560
rect 47728 8548 47734 8560
rect 47949 8551 48007 8557
rect 47949 8548 47961 8551
rect 47728 8520 47961 8548
rect 47728 8508 47734 8520
rect 47949 8517 47961 8520
rect 47995 8517 48007 8551
rect 47949 8511 48007 8517
rect 48041 8551 48099 8557
rect 48041 8517 48053 8551
rect 48087 8548 48099 8551
rect 53190 8548 53196 8560
rect 48087 8520 53196 8548
rect 48087 8517 48099 8520
rect 48041 8511 48099 8517
rect 53190 8508 53196 8520
rect 53248 8508 53254 8560
rect 42613 8483 42671 8489
rect 42613 8480 42625 8483
rect 41386 8452 42625 8480
rect 42613 8449 42625 8452
rect 42659 8480 42671 8483
rect 42702 8480 42708 8492
rect 42659 8452 42708 8480
rect 42659 8449 42671 8452
rect 42613 8443 42671 8449
rect 42702 8440 42708 8452
rect 42760 8440 42766 8492
rect 42886 8489 42892 8492
rect 42880 8443 42892 8489
rect 42886 8440 42892 8443
rect 42944 8440 42950 8492
rect 47765 8483 47823 8489
rect 47765 8449 47777 8483
rect 47811 8480 47823 8483
rect 47854 8480 47860 8492
rect 47811 8452 47860 8480
rect 47811 8449 47823 8452
rect 47765 8443 47823 8449
rect 47854 8440 47860 8452
rect 47912 8440 47918 8492
rect 48133 8483 48191 8489
rect 48133 8449 48145 8483
rect 48179 8449 48191 8483
rect 48133 8443 48191 8449
rect 35529 8375 35587 8381
rect 35636 8384 37504 8412
rect 22094 8344 22100 8356
rect 10928 8316 13400 8344
rect 20916 8316 22100 8344
rect 10928 8304 10934 8316
rect 17310 8236 17316 8288
rect 17368 8276 17374 8288
rect 18230 8276 18236 8288
rect 17368 8248 18236 8276
rect 17368 8236 17374 8248
rect 18230 8236 18236 8248
rect 18288 8276 18294 8288
rect 20916 8276 20944 8316
rect 22094 8304 22100 8316
rect 22152 8304 22158 8356
rect 25590 8304 25596 8356
rect 25648 8304 25654 8356
rect 28442 8304 28448 8356
rect 28500 8344 28506 8356
rect 29730 8344 29736 8356
rect 28500 8316 29736 8344
rect 28500 8304 28506 8316
rect 29730 8304 29736 8316
rect 29788 8304 29794 8356
rect 33134 8304 33140 8356
rect 33192 8344 33198 8356
rect 33192 8316 33824 8344
rect 33192 8304 33198 8316
rect 18288 8248 20944 8276
rect 18288 8236 18294 8248
rect 20990 8236 20996 8288
rect 21048 8276 21054 8288
rect 26602 8276 26608 8288
rect 21048 8248 26608 8276
rect 21048 8236 21054 8248
rect 26602 8236 26608 8248
rect 26660 8236 26666 8288
rect 26786 8236 26792 8288
rect 26844 8276 26850 8288
rect 31938 8276 31944 8288
rect 26844 8248 31944 8276
rect 26844 8236 26850 8248
rect 31938 8236 31944 8248
rect 31996 8236 32002 8288
rect 33796 8276 33824 8316
rect 34514 8304 34520 8356
rect 34572 8344 34578 8356
rect 35636 8344 35664 8384
rect 37642 8372 37648 8424
rect 37700 8372 37706 8424
rect 45094 8372 45100 8424
rect 45152 8412 45158 8424
rect 46474 8412 46480 8424
rect 45152 8384 46480 8412
rect 45152 8372 45158 8384
rect 46474 8372 46480 8384
rect 46532 8372 46538 8424
rect 47210 8372 47216 8424
rect 47268 8412 47274 8424
rect 48148 8412 48176 8443
rect 48314 8440 48320 8492
rect 48372 8480 48378 8492
rect 48372 8452 48728 8480
rect 48372 8440 48378 8452
rect 47268 8384 48176 8412
rect 48700 8412 48728 8452
rect 48958 8440 48964 8492
rect 49016 8440 49022 8492
rect 58066 8440 58072 8492
rect 58124 8440 58130 8492
rect 49050 8412 49056 8424
rect 48700 8384 49056 8412
rect 47268 8372 47274 8384
rect 49050 8372 49056 8384
rect 49108 8372 49114 8424
rect 34572 8316 35664 8344
rect 34572 8304 34578 8316
rect 36446 8304 36452 8356
rect 36504 8304 36510 8356
rect 37366 8304 37372 8356
rect 37424 8344 37430 8356
rect 37660 8344 37688 8372
rect 37424 8316 37688 8344
rect 37424 8304 37430 8316
rect 48130 8304 48136 8356
rect 48188 8344 48194 8356
rect 48317 8347 48375 8353
rect 48317 8344 48329 8347
rect 48188 8316 48329 8344
rect 48188 8304 48194 8316
rect 48317 8313 48329 8316
rect 48363 8313 48375 8347
rect 48317 8307 48375 8313
rect 48774 8304 48780 8356
rect 48832 8304 48838 8356
rect 53374 8304 53380 8356
rect 53432 8344 53438 8356
rect 55306 8344 55312 8356
rect 53432 8316 55312 8344
rect 53432 8304 53438 8316
rect 55306 8304 55312 8316
rect 55364 8304 55370 8356
rect 33965 8279 34023 8285
rect 33965 8276 33977 8279
rect 33796 8248 33977 8276
rect 33965 8245 33977 8248
rect 34011 8245 34023 8279
rect 33965 8239 34023 8245
rect 35434 8236 35440 8288
rect 35492 8276 35498 8288
rect 42610 8276 42616 8288
rect 35492 8248 42616 8276
rect 35492 8236 35498 8248
rect 42610 8236 42616 8248
rect 42668 8236 42674 8288
rect 43530 8236 43536 8288
rect 43588 8276 43594 8288
rect 43993 8279 44051 8285
rect 43993 8276 44005 8279
rect 43588 8248 44005 8276
rect 43588 8236 43594 8248
rect 43993 8245 44005 8248
rect 44039 8245 44051 8279
rect 43993 8239 44051 8245
rect 48958 8236 48964 8288
rect 49016 8276 49022 8288
rect 56594 8276 56600 8288
rect 49016 8248 56600 8276
rect 49016 8236 49022 8248
rect 56594 8236 56600 8248
rect 56652 8236 56658 8288
rect 1104 8186 58880 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 58880 8186
rect 1104 8112 58880 8134
rect 10505 8075 10563 8081
rect 10505 8041 10517 8075
rect 10551 8072 10563 8075
rect 11054 8072 11060 8084
rect 10551 8044 11060 8072
rect 10551 8041 10563 8044
rect 10505 8035 10563 8041
rect 11054 8032 11060 8044
rect 11112 8032 11118 8084
rect 12618 8032 12624 8084
rect 12676 8072 12682 8084
rect 13449 8075 13507 8081
rect 13449 8072 13461 8075
rect 12676 8044 13461 8072
rect 12676 8032 12682 8044
rect 13449 8041 13461 8044
rect 13495 8041 13507 8075
rect 13449 8035 13507 8041
rect 22833 8075 22891 8081
rect 22833 8041 22845 8075
rect 22879 8072 22891 8075
rect 23198 8072 23204 8084
rect 22879 8044 23204 8072
rect 22879 8041 22891 8044
rect 22833 8035 22891 8041
rect 23198 8032 23204 8044
rect 23256 8032 23262 8084
rect 26786 8072 26792 8084
rect 23308 8044 26792 8072
rect 8754 7964 8760 8016
rect 8812 8004 8818 8016
rect 10321 8007 10379 8013
rect 10321 8004 10333 8007
rect 8812 7976 10333 8004
rect 8812 7964 8818 7976
rect 10321 7973 10333 7976
rect 10367 7973 10379 8007
rect 10321 7967 10379 7973
rect 10594 7964 10600 8016
rect 10652 8004 10658 8016
rect 12345 8007 12403 8013
rect 12345 8004 12357 8007
rect 10652 7976 12357 8004
rect 10652 7964 10658 7976
rect 12345 7973 12357 7976
rect 12391 7973 12403 8007
rect 12345 7967 12403 7973
rect 12529 8007 12587 8013
rect 12529 7973 12541 8007
rect 12575 8004 12587 8007
rect 12802 8004 12808 8016
rect 12575 7976 12808 8004
rect 12575 7973 12587 7976
rect 12529 7967 12587 7973
rect 12802 7964 12808 7976
rect 12860 7964 12866 8016
rect 13265 8007 13323 8013
rect 13265 8004 13277 8007
rect 12912 7976 13277 8004
rect 10965 7939 11023 7945
rect 10965 7936 10977 7939
rect 6886 7908 10977 7936
rect 1581 7871 1639 7877
rect 1581 7837 1593 7871
rect 1627 7868 1639 7871
rect 6886 7868 6914 7908
rect 10965 7905 10977 7908
rect 11011 7905 11023 7939
rect 10965 7899 11023 7905
rect 11146 7896 11152 7948
rect 11204 7896 11210 7948
rect 11238 7896 11244 7948
rect 11296 7896 11302 7948
rect 12069 7939 12127 7945
rect 12069 7936 12081 7939
rect 11348 7908 12081 7936
rect 11348 7877 11376 7908
rect 12069 7905 12081 7908
rect 12115 7936 12127 7939
rect 12434 7936 12440 7948
rect 12115 7908 12440 7936
rect 12115 7905 12127 7908
rect 12069 7899 12127 7905
rect 12434 7896 12440 7908
rect 12492 7896 12498 7948
rect 1627 7840 6914 7868
rect 11333 7871 11391 7877
rect 1627 7837 1639 7840
rect 1581 7831 1639 7837
rect 11333 7837 11345 7871
rect 11379 7837 11391 7871
rect 11333 7831 11391 7837
rect 934 7760 940 7812
rect 992 7800 998 7812
rect 1857 7803 1915 7809
rect 1857 7800 1869 7803
rect 992 7772 1869 7800
rect 992 7760 998 7772
rect 1857 7769 1869 7772
rect 1903 7769 1915 7803
rect 1857 7763 1915 7769
rect 10045 7803 10103 7809
rect 10045 7769 10057 7803
rect 10091 7800 10103 7803
rect 10962 7800 10968 7812
rect 10091 7772 10968 7800
rect 10091 7769 10103 7772
rect 10045 7763 10103 7769
rect 10962 7760 10968 7772
rect 11020 7800 11026 7812
rect 11348 7800 11376 7831
rect 11422 7828 11428 7880
rect 11480 7828 11486 7880
rect 11514 7828 11520 7880
rect 11572 7868 11578 7880
rect 12912 7868 12940 7976
rect 13265 7973 13277 7976
rect 13311 7973 13323 8007
rect 13265 7967 13323 7973
rect 12989 7939 13047 7945
rect 12989 7905 13001 7939
rect 13035 7936 13047 7939
rect 13354 7936 13360 7948
rect 13035 7908 13360 7936
rect 13035 7905 13047 7908
rect 12989 7899 13047 7905
rect 13354 7896 13360 7908
rect 13412 7896 13418 7948
rect 19150 7896 19156 7948
rect 19208 7936 19214 7948
rect 23308 7936 23336 8044
rect 26786 8032 26792 8044
rect 26844 8032 26850 8084
rect 27798 8032 27804 8084
rect 27856 8072 27862 8084
rect 27893 8075 27951 8081
rect 27893 8072 27905 8075
rect 27856 8044 27905 8072
rect 27856 8032 27862 8044
rect 27893 8041 27905 8044
rect 27939 8041 27951 8075
rect 27893 8035 27951 8041
rect 30466 8032 30472 8084
rect 30524 8072 30530 8084
rect 31481 8075 31539 8081
rect 31481 8072 31493 8075
rect 30524 8044 31493 8072
rect 30524 8032 30530 8044
rect 31481 8041 31493 8044
rect 31527 8041 31539 8075
rect 31481 8035 31539 8041
rect 32398 8032 32404 8084
rect 32456 8072 32462 8084
rect 35434 8072 35440 8084
rect 32456 8044 35440 8072
rect 32456 8032 32462 8044
rect 35434 8032 35440 8044
rect 35492 8032 35498 8084
rect 35894 8032 35900 8084
rect 35952 8072 35958 8084
rect 39390 8072 39396 8084
rect 35952 8044 39396 8072
rect 35952 8032 35958 8044
rect 39390 8032 39396 8044
rect 39448 8032 39454 8084
rect 42886 8032 42892 8084
rect 42944 8072 42950 8084
rect 42981 8075 43039 8081
rect 42981 8072 42993 8075
rect 42944 8044 42993 8072
rect 42944 8032 42950 8044
rect 42981 8041 42993 8044
rect 43027 8041 43039 8075
rect 48869 8075 48927 8081
rect 48869 8072 48881 8075
rect 42981 8035 43039 8041
rect 46308 8044 48881 8072
rect 26602 7964 26608 8016
rect 26660 8004 26666 8016
rect 36630 8004 36636 8016
rect 26660 7976 36636 8004
rect 26660 7964 26666 7976
rect 36630 7964 36636 7976
rect 36688 7964 36694 8016
rect 36725 8007 36783 8013
rect 36725 7973 36737 8007
rect 36771 8004 36783 8007
rect 36906 8004 36912 8016
rect 36771 7976 36912 8004
rect 36771 7973 36783 7976
rect 36725 7967 36783 7973
rect 36906 7964 36912 7976
rect 36964 7964 36970 8016
rect 38102 7964 38108 8016
rect 38160 7964 38166 8016
rect 19208 7908 23336 7936
rect 23385 7939 23443 7945
rect 19208 7896 19214 7908
rect 23385 7905 23397 7939
rect 23431 7936 23443 7939
rect 23566 7936 23572 7948
rect 23431 7908 23572 7936
rect 23431 7905 23443 7908
rect 23385 7899 23443 7905
rect 23566 7896 23572 7908
rect 23624 7896 23630 7948
rect 27706 7936 27712 7948
rect 27080 7908 27712 7936
rect 11572 7840 12940 7868
rect 11572 7828 11578 7840
rect 25590 7800 25596 7812
rect 11020 7772 11376 7800
rect 12406 7772 12664 7800
rect 11020 7760 11026 7772
rect 11238 7692 11244 7744
rect 11296 7732 11302 7744
rect 12406 7732 12434 7772
rect 11296 7704 12434 7732
rect 12636 7732 12664 7772
rect 13372 7772 25596 7800
rect 13372 7732 13400 7772
rect 25590 7760 25596 7772
rect 25648 7760 25654 7812
rect 27080 7809 27108 7908
rect 27706 7896 27712 7908
rect 27764 7896 27770 7948
rect 28537 7939 28595 7945
rect 28537 7905 28549 7939
rect 28583 7936 28595 7939
rect 28626 7936 28632 7948
rect 28583 7908 28632 7936
rect 28583 7905 28595 7908
rect 28537 7899 28595 7905
rect 28626 7896 28632 7908
rect 28684 7896 28690 7948
rect 29086 7896 29092 7948
rect 29144 7936 29150 7948
rect 31846 7936 31852 7948
rect 29144 7908 30328 7936
rect 29144 7896 29150 7908
rect 27433 7871 27491 7877
rect 27433 7837 27445 7871
rect 27479 7868 27491 7871
rect 28810 7868 28816 7880
rect 27479 7840 28816 7868
rect 27479 7837 27491 7840
rect 27433 7831 27491 7837
rect 28810 7828 28816 7840
rect 28868 7828 28874 7880
rect 30098 7828 30104 7880
rect 30156 7868 30162 7880
rect 30300 7877 30328 7908
rect 30392 7908 31852 7936
rect 30193 7871 30251 7877
rect 30193 7868 30205 7871
rect 30156 7840 30205 7868
rect 30156 7828 30162 7840
rect 30193 7837 30205 7840
rect 30239 7837 30251 7871
rect 30193 7831 30251 7837
rect 30286 7871 30344 7877
rect 30286 7837 30298 7871
rect 30332 7837 30344 7871
rect 30286 7831 30344 7837
rect 27065 7803 27123 7809
rect 27065 7769 27077 7803
rect 27111 7769 27123 7803
rect 27065 7763 27123 7769
rect 27246 7760 27252 7812
rect 27304 7760 27310 7812
rect 28258 7760 28264 7812
rect 28316 7760 28322 7812
rect 29178 7760 29184 7812
rect 29236 7800 29242 7812
rect 30392 7800 30420 7908
rect 30650 7828 30656 7880
rect 30708 7877 30714 7880
rect 30708 7868 30716 7877
rect 31570 7868 31576 7880
rect 30708 7840 31576 7868
rect 30708 7831 30716 7840
rect 30708 7828 30714 7831
rect 31570 7828 31576 7840
rect 31628 7828 31634 7880
rect 31680 7877 31708 7908
rect 31846 7896 31852 7908
rect 31904 7896 31910 7948
rect 35986 7896 35992 7948
rect 36044 7936 36050 7948
rect 42978 7936 42984 7948
rect 36044 7908 42984 7936
rect 36044 7896 36050 7908
rect 42978 7896 42984 7908
rect 43036 7896 43042 7948
rect 43254 7896 43260 7948
rect 43312 7936 43318 7948
rect 43533 7939 43591 7945
rect 43533 7936 43545 7939
rect 43312 7908 43545 7936
rect 43312 7896 43318 7908
rect 43533 7905 43545 7908
rect 43579 7905 43591 7939
rect 43533 7899 43591 7905
rect 31665 7871 31723 7877
rect 31665 7837 31677 7871
rect 31711 7837 31723 7871
rect 31665 7831 31723 7837
rect 31754 7828 31760 7880
rect 31812 7828 31818 7880
rect 31938 7828 31944 7880
rect 31996 7828 32002 7880
rect 32033 7871 32091 7877
rect 32033 7837 32045 7871
rect 32079 7868 32091 7871
rect 32122 7868 32128 7880
rect 32079 7840 32128 7868
rect 32079 7837 32091 7840
rect 32033 7831 32091 7837
rect 32122 7828 32128 7840
rect 32180 7828 32186 7880
rect 33873 7871 33931 7877
rect 33873 7837 33885 7871
rect 33919 7868 33931 7871
rect 34514 7868 34520 7880
rect 33919 7840 34520 7868
rect 33919 7837 33931 7840
rect 33873 7831 33931 7837
rect 34514 7828 34520 7840
rect 34572 7828 34578 7880
rect 35434 7828 35440 7880
rect 35492 7868 35498 7880
rect 35529 7871 35587 7877
rect 35529 7868 35541 7871
rect 35492 7840 35541 7868
rect 35492 7828 35498 7840
rect 35529 7837 35541 7840
rect 35575 7837 35587 7871
rect 35529 7831 35587 7837
rect 35802 7828 35808 7880
rect 35860 7828 35866 7880
rect 37185 7871 37243 7877
rect 37185 7837 37197 7871
rect 37231 7868 37243 7871
rect 37366 7868 37372 7880
rect 37231 7840 37372 7868
rect 37231 7837 37243 7840
rect 37185 7831 37243 7837
rect 37366 7828 37372 7840
rect 37424 7828 37430 7880
rect 37458 7828 37464 7880
rect 37516 7828 37522 7880
rect 37550 7828 37556 7880
rect 37608 7828 37614 7880
rect 37826 7828 37832 7880
rect 37884 7868 37890 7880
rect 38838 7868 38844 7880
rect 37884 7840 38844 7868
rect 37884 7828 37890 7840
rect 38838 7828 38844 7840
rect 38896 7828 38902 7880
rect 43349 7871 43407 7877
rect 43349 7837 43361 7871
rect 43395 7868 43407 7871
rect 43622 7868 43628 7880
rect 43395 7840 43628 7868
rect 43395 7837 43407 7840
rect 43349 7831 43407 7837
rect 43622 7828 43628 7840
rect 43680 7828 43686 7880
rect 44818 7828 44824 7880
rect 44876 7868 44882 7880
rect 46308 7877 46336 8044
rect 48869 8041 48881 8044
rect 48915 8072 48927 8075
rect 48915 8044 51074 8072
rect 48915 8041 48927 8044
rect 48869 8035 48927 8041
rect 47486 7896 47492 7948
rect 47544 7896 47550 7948
rect 46017 7871 46075 7877
rect 46017 7868 46029 7871
rect 44876 7840 46029 7868
rect 44876 7828 44882 7840
rect 46017 7837 46029 7840
rect 46063 7837 46075 7871
rect 46017 7831 46075 7837
rect 46293 7871 46351 7877
rect 46293 7837 46305 7871
rect 46339 7837 46351 7871
rect 46293 7831 46351 7837
rect 46385 7871 46443 7877
rect 46385 7837 46397 7871
rect 46431 7868 46443 7871
rect 46934 7868 46940 7880
rect 46431 7840 46940 7868
rect 46431 7837 46443 7840
rect 46385 7831 46443 7837
rect 46934 7828 46940 7840
rect 46992 7828 46998 7880
rect 29236 7772 30420 7800
rect 29236 7760 29242 7772
rect 30466 7760 30472 7812
rect 30524 7760 30530 7812
rect 30561 7803 30619 7809
rect 30561 7769 30573 7803
rect 30607 7769 30619 7803
rect 30561 7763 30619 7769
rect 30852 7772 34100 7800
rect 12636 7704 13400 7732
rect 11296 7692 11302 7704
rect 22462 7692 22468 7744
rect 22520 7732 22526 7744
rect 23201 7735 23259 7741
rect 23201 7732 23213 7735
rect 22520 7704 23213 7732
rect 22520 7692 22526 7704
rect 23201 7701 23213 7704
rect 23247 7701 23259 7735
rect 23201 7695 23259 7701
rect 23293 7735 23351 7741
rect 23293 7701 23305 7735
rect 23339 7732 23351 7735
rect 27522 7732 27528 7744
rect 23339 7704 27528 7732
rect 23339 7701 23351 7704
rect 23293 7695 23351 7701
rect 27522 7692 27528 7704
rect 27580 7692 27586 7744
rect 28353 7735 28411 7741
rect 28353 7701 28365 7735
rect 28399 7732 28411 7735
rect 28442 7732 28448 7744
rect 28399 7704 28448 7732
rect 28399 7701 28411 7704
rect 28353 7695 28411 7701
rect 28442 7692 28448 7704
rect 28500 7692 28506 7744
rect 28994 7692 29000 7744
rect 29052 7732 29058 7744
rect 30576 7732 30604 7763
rect 30852 7741 30880 7772
rect 29052 7704 30604 7732
rect 30837 7735 30895 7741
rect 29052 7692 29058 7704
rect 30837 7701 30849 7735
rect 30883 7701 30895 7735
rect 34072 7732 34100 7772
rect 34146 7760 34152 7812
rect 34204 7760 34210 7812
rect 35894 7760 35900 7812
rect 35952 7760 35958 7812
rect 36262 7760 36268 7812
rect 36320 7760 36326 7812
rect 36630 7760 36636 7812
rect 36688 7800 36694 7812
rect 37921 7803 37979 7809
rect 37921 7800 37933 7803
rect 36688 7772 37933 7800
rect 36688 7760 36694 7772
rect 37921 7769 37933 7772
rect 37967 7769 37979 7803
rect 46201 7803 46259 7809
rect 46201 7800 46213 7803
rect 37921 7763 37979 7769
rect 41386 7772 46213 7800
rect 41386 7732 41414 7772
rect 46201 7769 46213 7772
rect 46247 7769 46259 7803
rect 46201 7763 46259 7769
rect 47756 7803 47814 7809
rect 47756 7769 47768 7803
rect 47802 7800 47814 7803
rect 48130 7800 48136 7812
rect 47802 7772 48136 7800
rect 47802 7769 47814 7772
rect 47756 7763 47814 7769
rect 48130 7760 48136 7772
rect 48188 7760 48194 7812
rect 51046 7800 51074 8044
rect 57974 7936 57980 7948
rect 57164 7908 57980 7936
rect 56410 7828 56416 7880
rect 56468 7868 56474 7880
rect 57164 7877 57192 7908
rect 57974 7896 57980 7908
rect 58032 7896 58038 7948
rect 58158 7896 58164 7948
rect 58216 7896 58222 7948
rect 56965 7871 57023 7877
rect 56965 7868 56977 7871
rect 56468 7840 56977 7868
rect 56468 7828 56474 7840
rect 56965 7837 56977 7840
rect 57011 7837 57023 7871
rect 56965 7831 57023 7837
rect 57149 7871 57207 7877
rect 57149 7837 57161 7871
rect 57195 7837 57207 7871
rect 57149 7831 57207 7837
rect 57885 7871 57943 7877
rect 57885 7837 57897 7871
rect 57931 7837 57943 7871
rect 57885 7831 57943 7837
rect 57900 7800 57928 7831
rect 51046 7772 57928 7800
rect 34072 7704 41414 7732
rect 30837 7695 30895 7701
rect 43438 7692 43444 7744
rect 43496 7692 43502 7744
rect 46569 7735 46627 7741
rect 46569 7701 46581 7735
rect 46615 7732 46627 7735
rect 47946 7732 47952 7744
rect 46615 7704 47952 7732
rect 46615 7701 46627 7704
rect 46569 7695 46627 7701
rect 47946 7692 47952 7704
rect 48004 7692 48010 7744
rect 56502 7692 56508 7744
rect 56560 7732 56566 7744
rect 57057 7735 57115 7741
rect 57057 7732 57069 7735
rect 56560 7704 57069 7732
rect 56560 7692 56566 7704
rect 57057 7701 57069 7704
rect 57103 7701 57115 7735
rect 57057 7695 57115 7701
rect 1104 7642 58880 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 50294 7642
rect 50346 7590 50358 7642
rect 50410 7590 50422 7642
rect 50474 7590 50486 7642
rect 50538 7590 50550 7642
rect 50602 7590 58880 7642
rect 1104 7568 58880 7590
rect 11149 7531 11207 7537
rect 11149 7497 11161 7531
rect 11195 7528 11207 7531
rect 11422 7528 11428 7540
rect 11195 7500 11428 7528
rect 11195 7497 11207 7500
rect 11149 7491 11207 7497
rect 11422 7488 11428 7500
rect 11480 7488 11486 7540
rect 12253 7531 12311 7537
rect 12253 7497 12265 7531
rect 12299 7528 12311 7531
rect 12710 7528 12716 7540
rect 12299 7500 12716 7528
rect 12299 7497 12311 7500
rect 12253 7491 12311 7497
rect 12710 7488 12716 7500
rect 12768 7488 12774 7540
rect 20533 7531 20591 7537
rect 20533 7497 20545 7531
rect 20579 7528 20591 7531
rect 20579 7500 26924 7528
rect 20579 7497 20591 7500
rect 20533 7491 20591 7497
rect 10689 7463 10747 7469
rect 10689 7429 10701 7463
rect 10735 7460 10747 7463
rect 10962 7460 10968 7472
rect 10735 7432 10968 7460
rect 10735 7429 10747 7432
rect 10689 7423 10747 7429
rect 10962 7420 10968 7432
rect 11020 7460 11026 7472
rect 11793 7463 11851 7469
rect 11793 7460 11805 7463
rect 11020 7432 11805 7460
rect 11020 7420 11026 7432
rect 11793 7429 11805 7432
rect 11839 7429 11851 7463
rect 11793 7423 11851 7429
rect 1581 7395 1639 7401
rect 1581 7361 1593 7395
rect 1627 7392 1639 7395
rect 12342 7392 12348 7404
rect 1627 7364 12348 7392
rect 1627 7361 1639 7364
rect 1581 7355 1639 7361
rect 12342 7352 12348 7364
rect 12400 7352 12406 7404
rect 24118 7352 24124 7404
rect 24176 7352 24182 7404
rect 24388 7395 24446 7401
rect 24388 7361 24400 7395
rect 24434 7392 24446 7395
rect 24946 7392 24952 7404
rect 24434 7364 24952 7392
rect 24434 7361 24446 7364
rect 24388 7355 24446 7361
rect 24946 7352 24952 7364
rect 25004 7352 25010 7404
rect 26896 7392 26924 7500
rect 29914 7488 29920 7540
rect 29972 7488 29978 7540
rect 30742 7488 30748 7540
rect 30800 7528 30806 7540
rect 31478 7528 31484 7540
rect 30800 7500 31484 7528
rect 30800 7488 30806 7500
rect 31478 7488 31484 7500
rect 31536 7488 31542 7540
rect 35342 7488 35348 7540
rect 35400 7528 35406 7540
rect 35802 7528 35808 7540
rect 35400 7500 35808 7528
rect 35400 7488 35406 7500
rect 35802 7488 35808 7500
rect 35860 7528 35866 7540
rect 37458 7528 37464 7540
rect 35860 7500 37464 7528
rect 35860 7488 35866 7500
rect 37458 7488 37464 7500
rect 37516 7488 37522 7540
rect 39301 7531 39359 7537
rect 39301 7497 39313 7531
rect 39347 7528 39359 7531
rect 39347 7500 44772 7528
rect 39347 7497 39359 7500
rect 39301 7491 39359 7497
rect 28629 7463 28687 7469
rect 28629 7429 28641 7463
rect 28675 7460 28687 7463
rect 30374 7460 30380 7472
rect 28675 7432 30380 7460
rect 28675 7429 28687 7432
rect 28629 7423 28687 7429
rect 30374 7420 30380 7432
rect 30432 7420 30438 7472
rect 30650 7420 30656 7472
rect 30708 7460 30714 7472
rect 30708 7432 31226 7460
rect 30708 7420 30714 7432
rect 30926 7392 30932 7404
rect 26896 7364 30932 7392
rect 30926 7352 30932 7364
rect 30984 7352 30990 7404
rect 31198 7401 31226 7432
rect 33778 7420 33784 7472
rect 33836 7420 33842 7472
rect 37476 7460 37504 7488
rect 37829 7463 37887 7469
rect 37476 7432 37780 7460
rect 31198 7395 31263 7401
rect 31198 7364 31217 7395
rect 31205 7361 31217 7364
rect 31251 7361 31263 7395
rect 31205 7355 31263 7361
rect 31389 7395 31447 7401
rect 31389 7361 31401 7395
rect 31435 7361 31447 7395
rect 31389 7358 31447 7361
rect 31389 7355 31524 7358
rect 934 7284 940 7336
rect 992 7324 998 7336
rect 1765 7327 1823 7333
rect 1765 7324 1777 7327
rect 992 7296 1777 7324
rect 992 7284 998 7296
rect 1765 7293 1777 7296
rect 1811 7293 1823 7327
rect 1765 7287 1823 7293
rect 20073 7327 20131 7333
rect 20073 7293 20085 7327
rect 20119 7324 20131 7327
rect 20438 7324 20444 7336
rect 20119 7296 20444 7324
rect 20119 7293 20131 7296
rect 20073 7287 20131 7293
rect 20438 7284 20444 7296
rect 20496 7284 20502 7336
rect 27522 7284 27528 7336
rect 27580 7324 27586 7336
rect 30742 7324 30748 7336
rect 27580 7296 30748 7324
rect 27580 7284 27586 7296
rect 30742 7284 30748 7296
rect 30800 7284 30806 7336
rect 31110 7284 31116 7336
rect 31168 7284 31174 7336
rect 31297 7327 31355 7333
rect 31405 7330 31524 7355
rect 32398 7352 32404 7404
rect 32456 7352 32462 7404
rect 32766 7352 32772 7404
rect 32824 7352 32830 7404
rect 37366 7352 37372 7404
rect 37424 7392 37430 7404
rect 37752 7401 37780 7432
rect 37829 7429 37841 7463
rect 37875 7460 37887 7463
rect 43438 7460 43444 7472
rect 37875 7432 43444 7460
rect 37875 7429 37887 7432
rect 37829 7423 37887 7429
rect 43438 7420 43444 7432
rect 43496 7420 43502 7472
rect 44744 7460 44772 7500
rect 44818 7488 44824 7540
rect 44876 7488 44882 7540
rect 46845 7531 46903 7537
rect 46845 7497 46857 7531
rect 46891 7528 46903 7531
rect 46934 7528 46940 7540
rect 46891 7500 46940 7528
rect 46891 7497 46903 7500
rect 46845 7491 46903 7497
rect 46934 7488 46940 7500
rect 46992 7488 46998 7540
rect 48130 7488 48136 7540
rect 48188 7488 48194 7540
rect 56502 7488 56508 7540
rect 56560 7488 56566 7540
rect 48958 7460 48964 7472
rect 44744 7432 48964 7460
rect 48958 7420 48964 7432
rect 49016 7420 49022 7472
rect 56042 7460 56048 7472
rect 55600 7432 56048 7460
rect 37461 7395 37519 7401
rect 37461 7392 37473 7395
rect 37424 7364 37473 7392
rect 37424 7352 37430 7364
rect 37461 7361 37473 7364
rect 37507 7361 37519 7395
rect 37461 7355 37519 7361
rect 37737 7395 37795 7401
rect 37737 7361 37749 7395
rect 37783 7361 37795 7395
rect 37737 7355 37795 7361
rect 38194 7352 38200 7404
rect 38252 7352 38258 7404
rect 44266 7352 44272 7404
rect 44324 7392 44330 7404
rect 45097 7395 45155 7401
rect 45097 7392 45109 7395
rect 44324 7364 45109 7392
rect 44324 7352 44330 7364
rect 45097 7361 45109 7364
rect 45143 7361 45155 7395
rect 45097 7355 45155 7361
rect 45186 7352 45192 7404
rect 45244 7352 45250 7404
rect 45281 7395 45339 7401
rect 45281 7361 45293 7395
rect 45327 7361 45339 7395
rect 45281 7355 45339 7361
rect 45465 7395 45523 7401
rect 45465 7361 45477 7395
rect 45511 7392 45523 7395
rect 46014 7392 46020 7404
rect 45511 7364 46020 7392
rect 45511 7361 45523 7364
rect 45465 7355 45523 7361
rect 31297 7293 31309 7327
rect 31343 7293 31355 7327
rect 31297 7287 31355 7293
rect 9122 7216 9128 7268
rect 9180 7256 9186 7268
rect 10965 7259 11023 7265
rect 10965 7256 10977 7259
rect 9180 7228 10977 7256
rect 9180 7216 9186 7228
rect 10965 7225 10977 7228
rect 11011 7225 11023 7259
rect 10965 7219 11023 7225
rect 12066 7216 12072 7268
rect 12124 7216 12130 7268
rect 13446 7216 13452 7268
rect 13504 7256 13510 7268
rect 20349 7259 20407 7265
rect 20349 7256 20361 7259
rect 13504 7228 20361 7256
rect 13504 7216 13510 7228
rect 20349 7225 20361 7228
rect 20395 7225 20407 7259
rect 30466 7256 30472 7268
rect 20349 7219 20407 7225
rect 25056 7228 30472 7256
rect 25056 7200 25084 7228
rect 30466 7216 30472 7228
rect 30524 7216 30530 7268
rect 30926 7216 30932 7268
rect 30984 7216 30990 7268
rect 31018 7216 31024 7268
rect 31076 7256 31082 7268
rect 31312 7256 31340 7287
rect 31076 7228 31340 7256
rect 31076 7216 31082 7228
rect 25038 7148 25044 7200
rect 25096 7148 25102 7200
rect 25130 7148 25136 7200
rect 25188 7188 25194 7200
rect 25501 7191 25559 7197
rect 25501 7188 25513 7191
rect 25188 7160 25513 7188
rect 25188 7148 25194 7160
rect 25501 7157 25513 7160
rect 25547 7157 25559 7191
rect 25501 7151 25559 7157
rect 27246 7148 27252 7200
rect 27304 7188 27310 7200
rect 28994 7188 29000 7200
rect 27304 7160 29000 7188
rect 27304 7148 27310 7160
rect 28994 7148 29000 7160
rect 29052 7148 29058 7200
rect 30006 7148 30012 7200
rect 30064 7188 30070 7200
rect 31496 7188 31524 7330
rect 35529 7327 35587 7333
rect 35529 7293 35541 7327
rect 35575 7324 35587 7327
rect 35618 7324 35624 7336
rect 35575 7296 35624 7324
rect 35575 7293 35587 7296
rect 35529 7287 35587 7293
rect 35618 7284 35624 7296
rect 35676 7284 35682 7336
rect 39117 7327 39175 7333
rect 39117 7324 39129 7327
rect 35728 7296 39129 7324
rect 34790 7216 34796 7268
rect 34848 7256 34854 7268
rect 35728 7256 35756 7296
rect 39117 7293 39129 7296
rect 39163 7293 39175 7327
rect 39117 7287 39175 7293
rect 39482 7284 39488 7336
rect 39540 7284 39546 7336
rect 44450 7284 44456 7336
rect 44508 7324 44514 7336
rect 44818 7324 44824 7336
rect 44508 7296 44824 7324
rect 44508 7284 44514 7296
rect 44818 7284 44824 7296
rect 44876 7284 44882 7336
rect 45002 7284 45008 7336
rect 45060 7324 45066 7336
rect 45296 7324 45324 7355
rect 46014 7352 46020 7364
rect 46072 7352 46078 7404
rect 46566 7352 46572 7404
rect 46624 7352 46630 7404
rect 47946 7352 47952 7404
rect 48004 7352 48010 7404
rect 55490 7352 55496 7404
rect 55548 7392 55554 7404
rect 55600 7401 55628 7432
rect 56042 7420 56048 7432
rect 56100 7460 56106 7472
rect 56318 7460 56324 7472
rect 56100 7432 56324 7460
rect 56100 7420 56106 7432
rect 56318 7420 56324 7432
rect 56376 7420 56382 7472
rect 55585 7395 55643 7401
rect 55585 7392 55597 7395
rect 55548 7364 55597 7392
rect 55548 7352 55554 7364
rect 55585 7361 55597 7364
rect 55631 7361 55643 7395
rect 55585 7355 55643 7361
rect 55766 7352 55772 7404
rect 55824 7352 55830 7404
rect 55861 7395 55919 7401
rect 55861 7361 55873 7395
rect 55907 7361 55919 7395
rect 55861 7355 55919 7361
rect 45060 7296 45324 7324
rect 45060 7284 45066 7296
rect 47118 7284 47124 7336
rect 47176 7324 47182 7336
rect 47486 7324 47492 7336
rect 47176 7296 47492 7324
rect 47176 7284 47182 7296
rect 47486 7284 47492 7296
rect 47544 7324 47550 7336
rect 47765 7327 47823 7333
rect 47765 7324 47777 7327
rect 47544 7296 47777 7324
rect 47544 7284 47550 7296
rect 47765 7293 47777 7296
rect 47811 7293 47823 7327
rect 47765 7287 47823 7293
rect 34848 7228 35756 7256
rect 34848 7216 34854 7228
rect 38378 7216 38384 7268
rect 38436 7216 38442 7268
rect 39592 7228 41414 7256
rect 30064 7160 31524 7188
rect 30064 7148 30070 7160
rect 31754 7148 31760 7200
rect 31812 7188 31818 7200
rect 39592 7188 39620 7228
rect 31812 7160 39620 7188
rect 31812 7148 31818 7160
rect 39666 7148 39672 7200
rect 39724 7148 39730 7200
rect 41386 7188 41414 7228
rect 42702 7216 42708 7268
rect 42760 7256 42766 7268
rect 55876 7256 55904 7355
rect 56594 7352 56600 7404
rect 56652 7352 56658 7404
rect 57057 7395 57115 7401
rect 57057 7361 57069 7395
rect 57103 7392 57115 7395
rect 57974 7392 57980 7404
rect 57103 7364 57980 7392
rect 57103 7361 57115 7364
rect 57057 7355 57115 7361
rect 57974 7352 57980 7364
rect 58032 7352 58038 7404
rect 58066 7352 58072 7404
rect 58124 7352 58130 7404
rect 57333 7327 57391 7333
rect 57333 7293 57345 7327
rect 57379 7324 57391 7327
rect 58986 7324 58992 7336
rect 57379 7296 58992 7324
rect 57379 7293 57391 7296
rect 57333 7287 57391 7293
rect 58986 7284 58992 7296
rect 59044 7284 59050 7336
rect 42760 7228 55904 7256
rect 42760 7216 42766 7228
rect 58250 7216 58256 7268
rect 58308 7216 58314 7268
rect 42978 7188 42984 7200
rect 41386 7160 42984 7188
rect 42978 7148 42984 7160
rect 43036 7148 43042 7200
rect 47670 7148 47676 7200
rect 47728 7188 47734 7200
rect 48130 7188 48136 7200
rect 47728 7160 48136 7188
rect 47728 7148 47734 7160
rect 48130 7148 48136 7160
rect 48188 7148 48194 7200
rect 55585 7191 55643 7197
rect 55585 7157 55597 7191
rect 55631 7188 55643 7191
rect 56042 7188 56048 7200
rect 55631 7160 56048 7188
rect 55631 7157 55643 7160
rect 55585 7151 55643 7157
rect 56042 7148 56048 7160
rect 56100 7148 56106 7200
rect 56321 7191 56379 7197
rect 56321 7157 56333 7191
rect 56367 7188 56379 7191
rect 56962 7188 56968 7200
rect 56367 7160 56968 7188
rect 56367 7157 56379 7160
rect 56321 7151 56379 7157
rect 56962 7148 56968 7160
rect 57020 7148 57026 7200
rect 1104 7098 58880 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 58880 7098
rect 1104 7024 58880 7046
rect 20901 6987 20959 6993
rect 20901 6953 20913 6987
rect 20947 6984 20959 6987
rect 20990 6984 20996 6996
rect 20947 6956 20996 6984
rect 20947 6953 20959 6956
rect 20901 6947 20959 6953
rect 20990 6944 20996 6956
rect 21048 6944 21054 6996
rect 24946 6944 24952 6996
rect 25004 6944 25010 6996
rect 26896 6956 28488 6984
rect 19797 6919 19855 6925
rect 19797 6885 19809 6919
rect 19843 6885 19855 6919
rect 19797 6879 19855 6885
rect 20717 6919 20775 6925
rect 20717 6885 20729 6919
rect 20763 6885 20775 6919
rect 20717 6879 20775 6885
rect 14458 6808 14464 6860
rect 14516 6848 14522 6860
rect 19812 6848 19840 6879
rect 14516 6820 19840 6848
rect 14516 6808 14522 6820
rect 1581 6783 1639 6789
rect 1581 6749 1593 6783
rect 1627 6780 1639 6783
rect 10410 6780 10416 6792
rect 1627 6752 10416 6780
rect 1627 6749 1639 6752
rect 1581 6743 1639 6749
rect 10410 6740 10416 6752
rect 10468 6740 10474 6792
rect 13906 6740 13912 6792
rect 13964 6780 13970 6792
rect 20732 6780 20760 6879
rect 21174 6876 21180 6928
rect 21232 6916 21238 6928
rect 26896 6916 26924 6956
rect 21232 6888 26924 6916
rect 28460 6916 28488 6956
rect 31386 6944 31392 6996
rect 31444 6944 31450 6996
rect 38194 6984 38200 6996
rect 31496 6956 38200 6984
rect 31496 6916 31524 6956
rect 38194 6944 38200 6956
rect 38252 6944 38258 6996
rect 39209 6987 39267 6993
rect 39209 6953 39221 6987
rect 39255 6984 39267 6987
rect 39666 6984 39672 6996
rect 39255 6956 39672 6984
rect 39255 6953 39267 6956
rect 39209 6947 39267 6953
rect 39666 6944 39672 6956
rect 39724 6984 39730 6996
rect 40957 6987 41015 6993
rect 40957 6984 40969 6987
rect 39724 6956 40969 6984
rect 39724 6944 39730 6956
rect 40957 6953 40969 6956
rect 41003 6984 41015 6987
rect 41414 6984 41420 6996
rect 41003 6956 41420 6984
rect 41003 6953 41015 6956
rect 40957 6947 41015 6953
rect 41414 6944 41420 6956
rect 41472 6984 41478 6996
rect 46934 6984 46940 6996
rect 41472 6956 46940 6984
rect 41472 6944 41478 6956
rect 46934 6944 46940 6956
rect 46992 6944 46998 6996
rect 47210 6944 47216 6996
rect 47268 6984 47274 6996
rect 47673 6987 47731 6993
rect 47673 6984 47685 6987
rect 47268 6956 47685 6984
rect 47268 6944 47274 6956
rect 47673 6953 47685 6956
rect 47719 6953 47731 6987
rect 47673 6947 47731 6953
rect 28460 6888 31524 6916
rect 21232 6876 21238 6888
rect 31570 6876 31576 6928
rect 31628 6916 31634 6928
rect 31938 6916 31944 6928
rect 31628 6888 31944 6916
rect 31628 6876 31634 6888
rect 31938 6876 31944 6888
rect 31996 6916 32002 6928
rect 32766 6916 32772 6928
rect 31996 6888 32772 6916
rect 31996 6876 32002 6888
rect 32766 6876 32772 6888
rect 32824 6876 32830 6928
rect 38286 6916 38292 6928
rect 37844 6888 38292 6916
rect 25593 6851 25651 6857
rect 25593 6817 25605 6851
rect 25639 6848 25651 6851
rect 25682 6848 25688 6860
rect 25639 6820 25688 6848
rect 25639 6817 25651 6820
rect 25593 6811 25651 6817
rect 25682 6808 25688 6820
rect 25740 6808 25746 6860
rect 27154 6808 27160 6860
rect 27212 6848 27218 6860
rect 27522 6848 27528 6860
rect 27212 6820 27528 6848
rect 27212 6808 27218 6820
rect 27522 6808 27528 6820
rect 27580 6808 27586 6860
rect 28166 6848 28172 6860
rect 27816 6820 28172 6848
rect 27614 6780 27620 6792
rect 13964 6752 20760 6780
rect 22066 6752 27620 6780
rect 13964 6740 13970 6752
rect 934 6672 940 6724
rect 992 6712 998 6724
rect 1857 6715 1915 6721
rect 1857 6712 1869 6715
rect 992 6684 1869 6712
rect 992 6672 998 6684
rect 1857 6681 1869 6684
rect 1903 6681 1915 6715
rect 1857 6675 1915 6681
rect 19521 6715 19579 6721
rect 19521 6681 19533 6715
rect 19567 6712 19579 6715
rect 20438 6712 20444 6724
rect 19567 6684 20444 6712
rect 19567 6681 19579 6684
rect 19521 6675 19579 6681
rect 20438 6672 20444 6684
rect 20496 6672 20502 6724
rect 19981 6647 20039 6653
rect 19981 6613 19993 6647
rect 20027 6644 20039 6647
rect 22066 6644 22094 6752
rect 27614 6740 27620 6752
rect 27672 6740 27678 6792
rect 27816 6789 27844 6820
rect 28166 6808 28172 6820
rect 28224 6808 28230 6860
rect 28994 6808 29000 6860
rect 29052 6808 29058 6860
rect 29270 6808 29276 6860
rect 29328 6848 29334 6860
rect 30466 6848 30472 6860
rect 29328 6820 30472 6848
rect 29328 6808 29334 6820
rect 30466 6808 30472 6820
rect 30524 6808 30530 6860
rect 30650 6808 30656 6860
rect 30708 6808 30714 6860
rect 30837 6851 30895 6857
rect 30837 6817 30849 6851
rect 30883 6848 30895 6851
rect 32309 6851 32367 6857
rect 32309 6848 32321 6851
rect 30883 6820 32321 6848
rect 30883 6817 30895 6820
rect 30837 6811 30895 6817
rect 32309 6817 32321 6820
rect 32355 6817 32367 6851
rect 32309 6811 32367 6817
rect 32416 6820 34008 6848
rect 27801 6783 27859 6789
rect 27801 6749 27813 6783
rect 27847 6749 27859 6783
rect 27801 6743 27859 6749
rect 27890 6740 27896 6792
rect 27948 6780 27954 6792
rect 30561 6783 30619 6789
rect 30561 6780 30573 6783
rect 27948 6752 30573 6780
rect 27948 6740 27954 6752
rect 30561 6749 30573 6752
rect 30607 6749 30619 6783
rect 30561 6743 30619 6749
rect 30742 6740 30748 6792
rect 30800 6780 30806 6792
rect 31018 6780 31024 6792
rect 30800 6752 31024 6780
rect 30800 6740 30806 6752
rect 31018 6740 31024 6752
rect 31076 6740 31082 6792
rect 31389 6783 31447 6789
rect 31389 6749 31401 6783
rect 31435 6749 31447 6783
rect 31389 6743 31447 6749
rect 25130 6672 25136 6724
rect 25188 6712 25194 6724
rect 25409 6715 25467 6721
rect 25409 6712 25421 6715
rect 25188 6684 25421 6712
rect 25188 6672 25194 6684
rect 25409 6681 25421 6684
rect 25455 6681 25467 6715
rect 29822 6712 29828 6724
rect 25409 6675 25467 6681
rect 28828 6684 29828 6712
rect 20027 6616 22094 6644
rect 25317 6647 25375 6653
rect 20027 6613 20039 6616
rect 19981 6607 20039 6613
rect 25317 6613 25329 6647
rect 25363 6644 25375 6647
rect 28828 6644 28856 6684
rect 29822 6672 29828 6684
rect 29880 6672 29886 6724
rect 31404 6712 31432 6743
rect 31570 6740 31576 6792
rect 31628 6740 31634 6792
rect 32030 6740 32036 6792
rect 32088 6780 32094 6792
rect 32416 6780 32444 6820
rect 32088 6752 32444 6780
rect 32088 6740 32094 6752
rect 32490 6740 32496 6792
rect 32548 6740 32554 6792
rect 32766 6740 32772 6792
rect 32824 6740 32830 6792
rect 33980 6789 34008 6820
rect 37274 6808 37280 6860
rect 37332 6848 37338 6860
rect 37844 6848 37872 6888
rect 37332 6820 37872 6848
rect 37332 6808 37338 6820
rect 37918 6808 37924 6860
rect 37976 6808 37982 6860
rect 38028 6857 38056 6888
rect 38286 6876 38292 6888
rect 38344 6876 38350 6928
rect 40678 6876 40684 6928
rect 40736 6916 40742 6928
rect 45189 6919 45247 6925
rect 40736 6888 43852 6916
rect 40736 6876 40742 6888
rect 38013 6851 38071 6857
rect 38013 6817 38025 6851
rect 38059 6817 38071 6851
rect 38013 6811 38071 6817
rect 38102 6808 38108 6860
rect 38160 6848 38166 6860
rect 43824 6857 43852 6888
rect 45189 6885 45201 6919
rect 45235 6916 45247 6919
rect 46014 6916 46020 6928
rect 45235 6888 46020 6916
rect 45235 6885 45247 6888
rect 45189 6879 45247 6885
rect 46014 6876 46020 6888
rect 46072 6876 46078 6928
rect 47688 6916 47716 6947
rect 57974 6944 57980 6996
rect 58032 6984 58038 6996
rect 58069 6987 58127 6993
rect 58069 6984 58081 6987
rect 58032 6956 58081 6984
rect 58032 6944 58038 6956
rect 58069 6953 58081 6956
rect 58115 6953 58127 6987
rect 58069 6947 58127 6953
rect 47688 6888 47808 6916
rect 43809 6851 43867 6857
rect 38160 6820 40908 6848
rect 38160 6808 38166 6820
rect 33965 6783 34023 6789
rect 33965 6749 33977 6783
rect 34011 6749 34023 6783
rect 33965 6743 34023 6749
rect 35618 6740 35624 6792
rect 35676 6740 35682 6792
rect 35710 6740 35716 6792
rect 35768 6780 35774 6792
rect 38657 6783 38715 6789
rect 38657 6780 38669 6783
rect 35768 6752 38669 6780
rect 35768 6740 35774 6752
rect 38657 6749 38669 6752
rect 38703 6749 38715 6783
rect 38657 6743 38715 6749
rect 39025 6783 39083 6789
rect 39025 6749 39037 6783
rect 39071 6780 39083 6783
rect 39850 6780 39856 6792
rect 39071 6752 39856 6780
rect 39071 6749 39083 6752
rect 39025 6743 39083 6749
rect 39850 6740 39856 6752
rect 39908 6740 39914 6792
rect 39942 6740 39948 6792
rect 40000 6780 40006 6792
rect 40405 6783 40463 6789
rect 40405 6780 40417 6783
rect 40000 6752 40417 6780
rect 40000 6740 40006 6752
rect 40405 6749 40417 6752
rect 40451 6749 40463 6783
rect 40405 6743 40463 6749
rect 40494 6740 40500 6792
rect 40552 6780 40558 6792
rect 40773 6783 40831 6789
rect 40773 6780 40785 6783
rect 40552 6752 40785 6780
rect 40552 6740 40558 6752
rect 40773 6749 40785 6752
rect 40819 6749 40831 6783
rect 40880 6780 40908 6820
rect 43809 6817 43821 6851
rect 43855 6848 43867 6851
rect 43898 6848 43904 6860
rect 43855 6820 43904 6848
rect 43855 6817 43867 6820
rect 43809 6811 43867 6817
rect 43898 6808 43904 6820
rect 43956 6808 43962 6860
rect 44468 6820 47716 6848
rect 44468 6792 44496 6820
rect 43625 6783 43683 6789
rect 43625 6780 43637 6783
rect 40880 6752 43637 6780
rect 40773 6743 40831 6749
rect 43625 6749 43637 6752
rect 43671 6780 43683 6783
rect 44266 6780 44272 6792
rect 43671 6752 44272 6780
rect 43671 6749 43683 6752
rect 43625 6743 43683 6749
rect 44266 6740 44272 6752
rect 44324 6740 44330 6792
rect 44450 6740 44456 6792
rect 44508 6740 44514 6792
rect 44637 6783 44695 6789
rect 44637 6749 44649 6783
rect 44683 6780 44695 6783
rect 44910 6780 44916 6792
rect 44683 6752 44916 6780
rect 44683 6749 44695 6752
rect 44637 6743 44695 6749
rect 44910 6740 44916 6752
rect 44968 6740 44974 6792
rect 45457 6783 45515 6789
rect 45365 6761 45423 6767
rect 45365 6758 45377 6761
rect 45296 6730 45377 6758
rect 33134 6712 33140 6724
rect 31404 6684 33140 6712
rect 33134 6672 33140 6684
rect 33192 6672 33198 6724
rect 33781 6715 33839 6721
rect 33781 6681 33793 6715
rect 33827 6712 33839 6715
rect 34146 6712 34152 6724
rect 33827 6684 34152 6712
rect 33827 6681 33839 6684
rect 33781 6675 33839 6681
rect 34146 6672 34152 6684
rect 34204 6672 34210 6724
rect 34698 6672 34704 6724
rect 34756 6712 34762 6724
rect 35866 6715 35924 6721
rect 35866 6712 35878 6715
rect 34756 6684 35878 6712
rect 34756 6672 34762 6684
rect 35866 6681 35878 6684
rect 35912 6681 35924 6715
rect 37829 6715 37887 6721
rect 37829 6712 37841 6715
rect 35866 6675 35924 6681
rect 37016 6684 37841 6712
rect 25363 6616 28856 6644
rect 30377 6647 30435 6653
rect 25363 6613 25375 6616
rect 25317 6607 25375 6613
rect 30377 6613 30389 6647
rect 30423 6644 30435 6647
rect 31018 6644 31024 6656
rect 30423 6616 31024 6644
rect 30423 6613 30435 6616
rect 30377 6607 30435 6613
rect 31018 6604 31024 6616
rect 31076 6604 31082 6656
rect 31754 6604 31760 6656
rect 31812 6604 31818 6656
rect 32677 6647 32735 6653
rect 32677 6613 32689 6647
rect 32723 6644 32735 6647
rect 32766 6644 32772 6656
rect 32723 6616 32772 6644
rect 32723 6613 32735 6616
rect 32677 6607 32735 6613
rect 32766 6604 32772 6616
rect 32824 6604 32830 6656
rect 34054 6604 34060 6656
rect 34112 6604 34118 6656
rect 34606 6604 34612 6656
rect 34664 6644 34670 6656
rect 37016 6653 37044 6684
rect 37829 6681 37841 6684
rect 37875 6712 37887 6715
rect 39298 6712 39304 6724
rect 37875 6684 39304 6712
rect 37875 6681 37887 6684
rect 37829 6675 37887 6681
rect 39298 6672 39304 6684
rect 39356 6672 39362 6724
rect 43717 6715 43775 6721
rect 43717 6681 43729 6715
rect 43763 6712 43775 6715
rect 43990 6712 43996 6724
rect 43763 6684 43996 6712
rect 43763 6681 43775 6684
rect 43717 6675 43775 6681
rect 43990 6672 43996 6684
rect 44048 6672 44054 6724
rect 45002 6672 45008 6724
rect 45060 6712 45066 6724
rect 45296 6712 45324 6730
rect 45365 6727 45377 6730
rect 45411 6727 45423 6761
rect 45457 6749 45469 6783
rect 45503 6749 45515 6783
rect 45457 6743 45515 6749
rect 45634 6783 45692 6789
rect 45634 6749 45646 6783
rect 45680 6749 45692 6783
rect 45634 6743 45692 6749
rect 45365 6721 45423 6727
rect 45060 6684 45324 6712
rect 45060 6672 45066 6684
rect 37001 6647 37059 6653
rect 37001 6644 37013 6647
rect 34664 6616 37013 6644
rect 34664 6604 34670 6616
rect 37001 6613 37013 6616
rect 37047 6613 37059 6647
rect 37001 6607 37059 6613
rect 37090 6604 37096 6656
rect 37148 6644 37154 6656
rect 37461 6647 37519 6653
rect 37461 6644 37473 6647
rect 37148 6616 37473 6644
rect 37148 6604 37154 6616
rect 37461 6613 37473 6616
rect 37507 6613 37519 6647
rect 37461 6607 37519 6613
rect 38841 6647 38899 6653
rect 38841 6613 38853 6647
rect 38887 6644 38899 6647
rect 40218 6644 40224 6656
rect 38887 6616 40224 6644
rect 38887 6613 38899 6616
rect 38841 6607 38899 6613
rect 40218 6604 40224 6616
rect 40276 6604 40282 6656
rect 40589 6647 40647 6653
rect 40589 6613 40601 6647
rect 40635 6644 40647 6647
rect 42702 6644 42708 6656
rect 40635 6616 42708 6644
rect 40635 6613 40647 6616
rect 40589 6607 40647 6613
rect 42702 6604 42708 6616
rect 42760 6604 42766 6656
rect 43254 6604 43260 6656
rect 43312 6604 43318 6656
rect 44542 6604 44548 6656
rect 44600 6604 44606 6656
rect 45370 6604 45376 6656
rect 45428 6644 45434 6656
rect 45471 6644 45499 6743
rect 45428 6616 45499 6644
rect 45664 6644 45692 6743
rect 45738 6740 45744 6792
rect 45796 6740 45802 6792
rect 46106 6740 46112 6792
rect 46164 6740 46170 6792
rect 46658 6740 46664 6792
rect 46716 6780 46722 6792
rect 46716 6752 47624 6780
rect 46716 6740 46722 6752
rect 46845 6715 46903 6721
rect 46845 6681 46857 6715
rect 46891 6681 46903 6715
rect 46845 6675 46903 6681
rect 45830 6644 45836 6656
rect 45664 6616 45836 6644
rect 45428 6604 45434 6616
rect 45830 6604 45836 6616
rect 45888 6644 45894 6656
rect 46382 6644 46388 6656
rect 45888 6616 46388 6644
rect 45888 6604 45894 6616
rect 46382 6604 46388 6616
rect 46440 6604 46446 6656
rect 46658 6604 46664 6656
rect 46716 6644 46722 6656
rect 46860 6644 46888 6675
rect 46716 6616 46888 6644
rect 46716 6604 46722 6616
rect 47210 6604 47216 6656
rect 47268 6644 47274 6656
rect 47305 6647 47363 6653
rect 47305 6644 47317 6647
rect 47268 6616 47317 6644
rect 47268 6604 47274 6616
rect 47305 6613 47317 6616
rect 47351 6613 47363 6647
rect 47596 6644 47624 6752
rect 47688 6724 47716 6820
rect 47670 6672 47676 6724
rect 47728 6672 47734 6724
rect 47780 6712 47808 6888
rect 55876 6820 56272 6848
rect 47854 6740 47860 6792
rect 47912 6740 47918 6792
rect 47949 6783 48007 6789
rect 47949 6749 47961 6783
rect 47995 6780 48007 6783
rect 48590 6780 48596 6792
rect 47995 6752 48596 6780
rect 47995 6749 48007 6752
rect 47949 6743 48007 6749
rect 48590 6740 48596 6752
rect 48648 6740 48654 6792
rect 55398 6712 55404 6724
rect 47780 6684 55404 6712
rect 55398 6672 55404 6684
rect 55456 6672 55462 6724
rect 55876 6721 55904 6820
rect 55861 6715 55919 6721
rect 55861 6681 55873 6715
rect 55907 6681 55919 6715
rect 56244 6712 56272 6820
rect 56689 6783 56747 6789
rect 56689 6749 56701 6783
rect 56735 6780 56747 6783
rect 56778 6780 56784 6792
rect 56735 6752 56784 6780
rect 56735 6749 56747 6752
rect 56689 6743 56747 6749
rect 56778 6740 56784 6752
rect 56836 6740 56842 6792
rect 56962 6789 56968 6792
rect 56956 6780 56968 6789
rect 56923 6752 56968 6780
rect 56956 6743 56968 6752
rect 56962 6740 56968 6743
rect 57020 6740 57026 6792
rect 58986 6712 58992 6724
rect 56244 6684 58992 6712
rect 55861 6675 55919 6681
rect 58986 6672 58992 6684
rect 59044 6672 59050 6724
rect 48133 6647 48191 6653
rect 48133 6644 48145 6647
rect 47596 6616 48145 6644
rect 47305 6607 47363 6613
rect 48133 6613 48145 6616
rect 48179 6613 48191 6647
rect 48133 6607 48191 6613
rect 48222 6604 48228 6656
rect 48280 6644 48286 6656
rect 55953 6647 56011 6653
rect 55953 6644 55965 6647
rect 48280 6616 55965 6644
rect 48280 6604 48286 6616
rect 55953 6613 55965 6616
rect 55999 6613 56011 6647
rect 55953 6607 56011 6613
rect 1104 6554 58880 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 50294 6554
rect 50346 6502 50358 6554
rect 50410 6502 50422 6554
rect 50474 6502 50486 6554
rect 50538 6502 50550 6554
rect 50602 6502 58880 6554
rect 1104 6480 58880 6502
rect 10410 6400 10416 6452
rect 10468 6400 10474 6452
rect 18322 6400 18328 6452
rect 18380 6440 18386 6452
rect 18380 6412 27844 6440
rect 18380 6400 18386 6412
rect 10686 6332 10692 6384
rect 10744 6372 10750 6384
rect 25130 6372 25136 6384
rect 10744 6344 25136 6372
rect 10744 6332 10750 6344
rect 25130 6332 25136 6344
rect 25188 6332 25194 6384
rect 25222 6332 25228 6384
rect 25280 6332 25286 6384
rect 27525 6375 27583 6381
rect 27525 6341 27537 6375
rect 27571 6372 27583 6375
rect 27816 6372 27844 6412
rect 28166 6400 28172 6452
rect 28224 6440 28230 6452
rect 28353 6443 28411 6449
rect 28353 6440 28365 6443
rect 28224 6412 28365 6440
rect 28224 6400 28230 6412
rect 28353 6409 28365 6412
rect 28399 6409 28411 6443
rect 28353 6403 28411 6409
rect 29178 6400 29184 6452
rect 29236 6440 29242 6452
rect 29638 6440 29644 6452
rect 29236 6412 29644 6440
rect 29236 6400 29242 6412
rect 29638 6400 29644 6412
rect 29696 6400 29702 6452
rect 29840 6412 30788 6440
rect 29840 6372 29868 6412
rect 27571 6344 27752 6372
rect 27816 6344 29868 6372
rect 29917 6375 29975 6381
rect 27571 6341 27583 6344
rect 27525 6335 27583 6341
rect 1581 6307 1639 6313
rect 1581 6273 1593 6307
rect 1627 6304 1639 6307
rect 26050 6304 26056 6316
rect 1627 6276 26056 6304
rect 1627 6273 1639 6276
rect 1581 6267 1639 6273
rect 26050 6264 26056 6276
rect 26108 6264 26114 6316
rect 27617 6307 27675 6313
rect 27540 6279 27629 6307
rect 934 6196 940 6248
rect 992 6236 998 6248
rect 1765 6239 1823 6245
rect 1765 6236 1777 6239
rect 992 6208 1777 6236
rect 992 6196 998 6208
rect 1765 6205 1777 6208
rect 1811 6205 1823 6239
rect 1765 6199 1823 6205
rect 10502 6196 10508 6248
rect 10560 6236 10566 6248
rect 10597 6239 10655 6245
rect 10597 6236 10609 6239
rect 10560 6208 10609 6236
rect 10560 6196 10566 6208
rect 10597 6205 10609 6208
rect 10643 6205 10655 6239
rect 10597 6199 10655 6205
rect 10612 6168 10640 6199
rect 10686 6196 10692 6248
rect 10744 6196 10750 6248
rect 10778 6196 10784 6248
rect 10836 6196 10842 6248
rect 10873 6239 10931 6245
rect 10873 6205 10885 6239
rect 10919 6236 10931 6239
rect 11054 6236 11060 6248
rect 10919 6208 11060 6236
rect 10919 6205 10931 6208
rect 10873 6199 10931 6205
rect 11054 6196 11060 6208
rect 11112 6196 11118 6248
rect 20438 6196 20444 6248
rect 20496 6236 20502 6248
rect 20717 6239 20775 6245
rect 20717 6236 20729 6239
rect 20496 6208 20729 6236
rect 20496 6196 20502 6208
rect 20717 6205 20729 6208
rect 20763 6205 20775 6239
rect 20717 6199 20775 6205
rect 25314 6196 25320 6248
rect 25372 6196 25378 6248
rect 25501 6239 25559 6245
rect 25501 6205 25513 6239
rect 25547 6236 25559 6239
rect 25682 6236 25688 6248
rect 25547 6208 25688 6236
rect 25547 6205 25559 6208
rect 25501 6199 25559 6205
rect 25682 6196 25688 6208
rect 25740 6196 25746 6248
rect 26326 6196 26332 6248
rect 26384 6236 26390 6248
rect 26786 6236 26792 6248
rect 26384 6208 26792 6236
rect 26384 6196 26390 6208
rect 26786 6196 26792 6208
rect 26844 6236 26850 6248
rect 27540 6236 27568 6279
rect 27617 6273 27629 6279
rect 27663 6273 27675 6307
rect 27724 6304 27752 6344
rect 29917 6341 29929 6375
rect 29963 6372 29975 6375
rect 30760 6372 30788 6412
rect 30834 6400 30840 6452
rect 30892 6440 30898 6452
rect 34606 6440 34612 6452
rect 30892 6412 34612 6440
rect 30892 6400 30898 6412
rect 34606 6400 34612 6412
rect 34664 6400 34670 6452
rect 34698 6400 34704 6452
rect 34756 6400 34762 6452
rect 39209 6443 39267 6449
rect 39209 6409 39221 6443
rect 39255 6440 39267 6443
rect 39482 6440 39488 6452
rect 39255 6412 39488 6440
rect 39255 6409 39267 6412
rect 39209 6403 39267 6409
rect 39482 6400 39488 6412
rect 39540 6400 39546 6452
rect 39850 6400 39856 6452
rect 39908 6400 39914 6452
rect 40494 6400 40500 6452
rect 40552 6400 40558 6452
rect 44266 6400 44272 6452
rect 44324 6400 44330 6452
rect 45186 6400 45192 6452
rect 45244 6440 45250 6452
rect 45462 6440 45468 6452
rect 45244 6412 45468 6440
rect 45244 6400 45250 6412
rect 45462 6400 45468 6412
rect 45520 6400 45526 6452
rect 45646 6400 45652 6452
rect 45704 6440 45710 6452
rect 46201 6443 46259 6449
rect 46201 6440 46213 6443
rect 45704 6412 46213 6440
rect 45704 6400 45710 6412
rect 46201 6409 46213 6412
rect 46247 6409 46259 6443
rect 46201 6403 46259 6409
rect 46382 6400 46388 6452
rect 46440 6440 46446 6452
rect 48406 6440 48412 6452
rect 46440 6412 48412 6440
rect 46440 6400 46446 6412
rect 48406 6400 48412 6412
rect 48464 6400 48470 6452
rect 55309 6443 55367 6449
rect 55309 6409 55321 6443
rect 55355 6440 55367 6443
rect 58253 6443 58311 6449
rect 58253 6440 58265 6443
rect 55355 6412 58265 6440
rect 55355 6409 55367 6412
rect 55309 6403 55367 6409
rect 58253 6409 58265 6412
rect 58299 6409 58311 6443
rect 58253 6403 58311 6409
rect 31110 6372 31116 6384
rect 29963 6344 30696 6372
rect 30760 6344 31116 6372
rect 29963 6341 29975 6344
rect 29917 6335 29975 6341
rect 30668 6316 30696 6344
rect 31110 6332 31116 6344
rect 31168 6372 31174 6384
rect 31754 6372 31760 6384
rect 31168 6344 31760 6372
rect 31168 6332 31174 6344
rect 31754 6332 31760 6344
rect 31812 6332 31818 6384
rect 37090 6372 37096 6384
rect 34532 6344 37096 6372
rect 28350 6304 28356 6316
rect 27724 6276 28356 6304
rect 27617 6267 27675 6273
rect 28350 6264 28356 6276
rect 28408 6304 28414 6316
rect 28629 6307 28687 6313
rect 28629 6304 28641 6307
rect 28408 6276 28641 6304
rect 28408 6264 28414 6276
rect 28629 6273 28641 6276
rect 28675 6273 28687 6307
rect 28629 6267 28687 6273
rect 28721 6307 28779 6313
rect 28721 6273 28733 6307
rect 28767 6273 28779 6307
rect 28721 6267 28779 6273
rect 26844 6208 27568 6236
rect 26844 6196 26850 6208
rect 27798 6196 27804 6248
rect 27856 6196 27862 6248
rect 28074 6196 28080 6248
rect 28132 6236 28138 6248
rect 28534 6236 28540 6248
rect 28132 6208 28540 6236
rect 28132 6196 28138 6208
rect 28534 6196 28540 6208
rect 28592 6236 28598 6248
rect 28736 6236 28764 6267
rect 28810 6264 28816 6316
rect 28868 6264 28874 6316
rect 28997 6307 29055 6313
rect 28997 6273 29009 6307
rect 29043 6304 29055 6307
rect 29454 6304 29460 6316
rect 29043 6276 29460 6304
rect 29043 6273 29055 6276
rect 28997 6267 29055 6273
rect 29454 6264 29460 6276
rect 29512 6264 29518 6316
rect 29638 6264 29644 6316
rect 29696 6264 29702 6316
rect 29822 6264 29828 6316
rect 29880 6264 29886 6316
rect 30650 6264 30656 6316
rect 30708 6264 30714 6316
rect 30742 6264 30748 6316
rect 30800 6264 30806 6316
rect 32582 6264 32588 6316
rect 32640 6264 32646 6316
rect 32766 6264 32772 6316
rect 32824 6264 32830 6316
rect 34532 6313 34560 6344
rect 37090 6332 37096 6344
rect 37148 6332 37154 6384
rect 43346 6372 43352 6384
rect 37200 6344 43352 6372
rect 34517 6307 34575 6313
rect 34517 6273 34529 6307
rect 34563 6273 34575 6307
rect 34517 6267 34575 6273
rect 35342 6264 35348 6316
rect 35400 6304 35406 6316
rect 35437 6307 35495 6313
rect 35437 6304 35449 6307
rect 35400 6276 35449 6304
rect 35400 6264 35406 6276
rect 35437 6273 35449 6276
rect 35483 6273 35495 6307
rect 35437 6267 35495 6273
rect 35526 6264 35532 6316
rect 35584 6264 35590 6316
rect 35894 6264 35900 6316
rect 35952 6264 35958 6316
rect 36354 6264 36360 6316
rect 36412 6304 36418 6316
rect 37200 6304 37228 6344
rect 43346 6332 43352 6344
rect 43404 6332 43410 6384
rect 45738 6372 45744 6384
rect 44836 6344 45744 6372
rect 36412 6276 37228 6304
rect 36412 6264 36418 6276
rect 37458 6264 37464 6316
rect 37516 6264 37522 6316
rect 38473 6307 38531 6313
rect 38473 6273 38485 6307
rect 38519 6273 38531 6307
rect 38473 6267 38531 6273
rect 28592 6208 28764 6236
rect 28592 6196 28598 6208
rect 30558 6196 30564 6248
rect 30616 6196 30622 6248
rect 30837 6239 30895 6245
rect 30837 6205 30849 6239
rect 30883 6236 30895 6239
rect 30926 6236 30932 6248
rect 30883 6208 30932 6236
rect 30883 6205 30895 6208
rect 30837 6199 30895 6205
rect 30926 6196 30932 6208
rect 30984 6196 30990 6248
rect 33134 6196 33140 6248
rect 33192 6236 33198 6248
rect 34333 6239 34391 6245
rect 34333 6236 34345 6239
rect 33192 6208 34345 6236
rect 33192 6196 33198 6208
rect 34333 6205 34345 6208
rect 34379 6205 34391 6239
rect 34333 6199 34391 6205
rect 10612 6140 12434 6168
rect 12406 6100 12434 6140
rect 16574 6128 16580 6180
rect 16632 6168 16638 6180
rect 20993 6171 21051 6177
rect 20993 6168 21005 6171
rect 16632 6140 21005 6168
rect 16632 6128 16638 6140
rect 20993 6137 21005 6140
rect 21039 6137 21051 6171
rect 20993 6131 21051 6137
rect 21177 6171 21235 6177
rect 21177 6137 21189 6171
rect 21223 6168 21235 6171
rect 28994 6168 29000 6180
rect 21223 6140 29000 6168
rect 21223 6137 21235 6140
rect 21177 6131 21235 6137
rect 28994 6128 29000 6140
rect 29052 6128 29058 6180
rect 30282 6128 30288 6180
rect 30340 6168 30346 6180
rect 30377 6171 30435 6177
rect 30377 6168 30389 6171
rect 30340 6140 30389 6168
rect 30340 6128 30346 6140
rect 30377 6137 30389 6140
rect 30423 6137 30435 6171
rect 34054 6168 34060 6180
rect 30377 6131 30435 6137
rect 32876 6140 34060 6168
rect 24578 6100 24584 6112
rect 12406 6072 24584 6100
rect 24578 6060 24584 6072
rect 24636 6060 24642 6112
rect 24670 6060 24676 6112
rect 24728 6100 24734 6112
rect 24857 6103 24915 6109
rect 24857 6100 24869 6103
rect 24728 6072 24869 6100
rect 24728 6060 24734 6072
rect 24857 6069 24869 6072
rect 24903 6069 24915 6103
rect 24857 6063 24915 6069
rect 25682 6060 25688 6112
rect 25740 6100 25746 6112
rect 27157 6103 27215 6109
rect 27157 6100 27169 6103
rect 25740 6072 27169 6100
rect 25740 6060 25746 6072
rect 27157 6069 27169 6072
rect 27203 6069 27215 6103
rect 27157 6063 27215 6069
rect 28718 6060 28724 6112
rect 28776 6100 28782 6112
rect 32876 6100 32904 6140
rect 34054 6128 34060 6140
rect 34112 6128 34118 6180
rect 34348 6168 34376 6199
rect 34606 6196 34612 6248
rect 34664 6236 34670 6248
rect 35161 6239 35219 6245
rect 35161 6236 35173 6239
rect 34664 6208 35173 6236
rect 34664 6196 34670 6208
rect 35161 6205 35173 6208
rect 35207 6236 35219 6239
rect 35207 6208 37504 6236
rect 35207 6205 35219 6208
rect 35161 6199 35219 6205
rect 34422 6168 34428 6180
rect 34348 6140 34428 6168
rect 34422 6128 34428 6140
rect 34480 6168 34486 6180
rect 35710 6168 35716 6180
rect 34480 6140 35716 6168
rect 34480 6128 34486 6140
rect 35710 6128 35716 6140
rect 35768 6128 35774 6180
rect 36262 6128 36268 6180
rect 36320 6128 36326 6180
rect 37476 6168 37504 6208
rect 37550 6196 37556 6248
rect 37608 6236 37614 6248
rect 37645 6239 37703 6245
rect 37645 6236 37657 6239
rect 37608 6208 37657 6236
rect 37608 6196 37614 6208
rect 37645 6205 37657 6208
rect 37691 6205 37703 6239
rect 37645 6199 37703 6205
rect 38194 6168 38200 6180
rect 37476 6140 38200 6168
rect 38194 6128 38200 6140
rect 38252 6168 38258 6180
rect 38488 6168 38516 6267
rect 39022 6264 39028 6316
rect 39080 6304 39086 6316
rect 39117 6307 39175 6313
rect 39117 6304 39129 6307
rect 39080 6276 39129 6304
rect 39080 6264 39086 6276
rect 39117 6273 39129 6276
rect 39163 6273 39175 6307
rect 39117 6267 39175 6273
rect 39132 6236 39160 6267
rect 39298 6264 39304 6316
rect 39356 6264 39362 6316
rect 39761 6307 39819 6313
rect 39761 6273 39773 6307
rect 39807 6273 39819 6307
rect 39761 6267 39819 6273
rect 39945 6310 40003 6313
rect 40034 6310 40040 6316
rect 39945 6307 40040 6310
rect 39945 6273 39957 6307
rect 39991 6282 40040 6307
rect 39991 6273 40003 6282
rect 39945 6267 40003 6273
rect 39776 6236 39804 6267
rect 40034 6264 40040 6282
rect 40092 6264 40098 6316
rect 40405 6307 40463 6313
rect 40405 6273 40417 6307
rect 40451 6273 40463 6307
rect 40405 6267 40463 6273
rect 39132 6208 39896 6236
rect 38252 6140 38516 6168
rect 38657 6171 38715 6177
rect 38252 6128 38258 6140
rect 38657 6137 38669 6171
rect 38703 6168 38715 6171
rect 39298 6168 39304 6180
rect 38703 6140 39304 6168
rect 38703 6137 38715 6140
rect 38657 6131 38715 6137
rect 39298 6128 39304 6140
rect 39356 6128 39362 6180
rect 39868 6168 39896 6208
rect 40420 6168 40448 6267
rect 40494 6264 40500 6316
rect 40552 6304 40558 6316
rect 40589 6307 40647 6313
rect 40589 6304 40601 6307
rect 40552 6276 40601 6304
rect 40552 6264 40558 6276
rect 40589 6273 40601 6276
rect 40635 6273 40647 6307
rect 40589 6267 40647 6273
rect 42794 6264 42800 6316
rect 42852 6304 42858 6316
rect 42889 6307 42947 6313
rect 42889 6304 42901 6307
rect 42852 6276 42901 6304
rect 42852 6264 42858 6276
rect 42889 6273 42901 6276
rect 42935 6273 42947 6307
rect 42889 6267 42947 6273
rect 43156 6307 43214 6313
rect 43156 6273 43168 6307
rect 43202 6304 43214 6307
rect 43438 6304 43444 6316
rect 43202 6276 43444 6304
rect 43202 6273 43214 6276
rect 43156 6267 43214 6273
rect 43438 6264 43444 6276
rect 43496 6264 43502 6316
rect 44358 6264 44364 6316
rect 44416 6304 44422 6316
rect 44836 6313 44864 6344
rect 45738 6332 45744 6344
rect 45796 6332 45802 6384
rect 44821 6307 44879 6313
rect 44821 6304 44833 6307
rect 44416 6276 44833 6304
rect 44416 6264 44422 6276
rect 44821 6273 44833 6276
rect 44867 6273 44879 6307
rect 44821 6267 44879 6273
rect 45005 6307 45063 6313
rect 45005 6273 45017 6307
rect 45051 6273 45063 6307
rect 45005 6267 45063 6273
rect 45020 6236 45048 6267
rect 45094 6264 45100 6316
rect 45152 6264 45158 6316
rect 45186 6264 45192 6316
rect 45244 6304 45250 6316
rect 46400 6313 46428 6400
rect 54662 6372 54668 6384
rect 51046 6344 54668 6372
rect 46017 6307 46075 6313
rect 46017 6304 46029 6307
rect 45244 6276 46029 6304
rect 45244 6264 45250 6276
rect 46017 6273 46029 6276
rect 46063 6273 46075 6307
rect 46017 6267 46075 6273
rect 46385 6307 46443 6313
rect 46385 6273 46397 6307
rect 46431 6273 46443 6307
rect 46385 6267 46443 6273
rect 46661 6307 46719 6313
rect 46661 6273 46673 6307
rect 46707 6304 46719 6307
rect 47670 6304 47676 6316
rect 46707 6276 47676 6304
rect 46707 6273 46719 6276
rect 46661 6267 46719 6273
rect 45462 6236 45468 6248
rect 45020 6208 45468 6236
rect 45462 6196 45468 6208
rect 45520 6196 45526 6248
rect 45557 6239 45615 6245
rect 45557 6205 45569 6239
rect 45603 6205 45615 6239
rect 46032 6236 46060 6267
rect 47670 6264 47676 6276
rect 47728 6264 47734 6316
rect 51046 6236 51074 6344
rect 54662 6332 54668 6344
rect 54720 6332 54726 6384
rect 56778 6372 56784 6384
rect 55784 6344 56784 6372
rect 55125 6307 55183 6313
rect 55125 6273 55137 6307
rect 55171 6273 55183 6307
rect 55125 6267 55183 6273
rect 55309 6307 55367 6313
rect 55309 6273 55321 6307
rect 55355 6304 55367 6307
rect 55674 6304 55680 6316
rect 55355 6276 55680 6304
rect 55355 6273 55367 6276
rect 55309 6267 55367 6273
rect 46032 6208 51074 6236
rect 45557 6199 45615 6205
rect 39868 6140 40448 6168
rect 43898 6128 43904 6180
rect 43956 6168 43962 6180
rect 45572 6168 45600 6199
rect 43956 6140 45600 6168
rect 43956 6128 43962 6140
rect 46658 6128 46664 6180
rect 46716 6168 46722 6180
rect 48590 6168 48596 6180
rect 46716 6140 48596 6168
rect 46716 6128 46722 6140
rect 48590 6128 48596 6140
rect 48648 6128 48654 6180
rect 28776 6072 32904 6100
rect 28776 6060 28782 6072
rect 32950 6060 32956 6112
rect 33008 6060 33014 6112
rect 35802 6060 35808 6112
rect 35860 6100 35866 6112
rect 37550 6100 37556 6112
rect 35860 6072 37556 6100
rect 35860 6060 35866 6072
rect 37550 6060 37556 6072
rect 37608 6060 37614 6112
rect 37826 6060 37832 6112
rect 37884 6100 37890 6112
rect 40034 6100 40040 6112
rect 37884 6072 40040 6100
rect 37884 6060 37890 6072
rect 40034 6060 40040 6072
rect 40092 6060 40098 6112
rect 44082 6060 44088 6112
rect 44140 6100 44146 6112
rect 46382 6100 46388 6112
rect 44140 6072 46388 6100
rect 44140 6060 44146 6072
rect 46382 6060 46388 6072
rect 46440 6060 46446 6112
rect 46477 6103 46535 6109
rect 46477 6069 46489 6103
rect 46523 6100 46535 6103
rect 47854 6100 47860 6112
rect 46523 6072 47860 6100
rect 46523 6069 46535 6072
rect 46477 6063 46535 6069
rect 47854 6060 47860 6072
rect 47912 6100 47918 6112
rect 54754 6100 54760 6112
rect 47912 6072 54760 6100
rect 47912 6060 47918 6072
rect 54754 6060 54760 6072
rect 54812 6060 54818 6112
rect 55140 6100 55168 6267
rect 55674 6264 55680 6276
rect 55732 6264 55738 6316
rect 55784 6313 55812 6344
rect 56778 6332 56784 6344
rect 56836 6332 56842 6384
rect 56042 6313 56048 6316
rect 55769 6307 55827 6313
rect 55769 6273 55781 6307
rect 55815 6273 55827 6307
rect 56036 6304 56048 6313
rect 56003 6276 56048 6304
rect 55769 6267 55827 6273
rect 56036 6267 56048 6276
rect 56042 6264 56048 6267
rect 56100 6264 56106 6316
rect 56318 6264 56324 6316
rect 56376 6304 56382 6316
rect 58069 6307 58127 6313
rect 58069 6304 58081 6307
rect 56376 6276 58081 6304
rect 56376 6264 56382 6276
rect 58069 6273 58081 6276
rect 58115 6273 58127 6307
rect 58069 6267 58127 6273
rect 58345 6307 58403 6313
rect 58345 6273 58357 6307
rect 58391 6273 58403 6307
rect 58345 6267 58403 6273
rect 57146 6196 57152 6248
rect 57204 6236 57210 6248
rect 58360 6236 58388 6267
rect 57204 6208 58388 6236
rect 57204 6196 57210 6208
rect 56410 6100 56416 6112
rect 55140 6072 56416 6100
rect 56410 6060 56416 6072
rect 56468 6060 56474 6112
rect 57054 6060 57060 6112
rect 57112 6100 57118 6112
rect 57149 6103 57207 6109
rect 57149 6100 57161 6103
rect 57112 6072 57161 6100
rect 57112 6060 57118 6072
rect 57149 6069 57161 6072
rect 57195 6069 57207 6103
rect 57149 6063 57207 6069
rect 58066 6060 58072 6112
rect 58124 6060 58130 6112
rect 1104 6010 58880 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 58880 6010
rect 1104 5936 58880 5958
rect 11054 5856 11060 5908
rect 11112 5856 11118 5908
rect 12342 5856 12348 5908
rect 12400 5896 12406 5908
rect 17773 5899 17831 5905
rect 17773 5896 17785 5899
rect 12400 5868 17785 5896
rect 12400 5856 12406 5868
rect 17773 5865 17785 5868
rect 17819 5865 17831 5899
rect 17773 5859 17831 5865
rect 23106 5856 23112 5908
rect 23164 5856 23170 5908
rect 24578 5856 24584 5908
rect 24636 5896 24642 5908
rect 24636 5868 26372 5896
rect 24636 5856 24642 5868
rect 8386 5788 8392 5840
rect 8444 5828 8450 5840
rect 10873 5831 10931 5837
rect 10873 5828 10885 5831
rect 8444 5800 10885 5828
rect 8444 5788 8450 5800
rect 10873 5797 10885 5800
rect 10919 5797 10931 5831
rect 10873 5791 10931 5797
rect 13814 5788 13820 5840
rect 13872 5828 13878 5840
rect 20257 5831 20315 5837
rect 20257 5828 20269 5831
rect 13872 5800 20269 5828
rect 13872 5788 13878 5800
rect 20257 5797 20269 5800
rect 20303 5797 20315 5831
rect 20257 5791 20315 5797
rect 20441 5831 20499 5837
rect 20441 5797 20453 5831
rect 20487 5828 20499 5831
rect 24762 5828 24768 5840
rect 20487 5800 24768 5828
rect 20487 5797 20499 5800
rect 20441 5791 20499 5797
rect 24762 5788 24768 5800
rect 24820 5788 24826 5840
rect 26344 5828 26372 5868
rect 26786 5856 26792 5908
rect 26844 5856 26850 5908
rect 29914 5896 29920 5908
rect 26896 5868 29920 5896
rect 26896 5828 26924 5868
rect 29914 5856 29920 5868
rect 29972 5896 29978 5908
rect 30834 5896 30840 5908
rect 29972 5868 30840 5896
rect 29972 5856 29978 5868
rect 30834 5856 30840 5868
rect 30892 5856 30898 5908
rect 30926 5856 30932 5908
rect 30984 5856 30990 5908
rect 31018 5856 31024 5908
rect 31076 5896 31082 5908
rect 39942 5896 39948 5908
rect 31076 5868 39948 5896
rect 31076 5856 31082 5868
rect 39942 5856 39948 5868
rect 40000 5856 40006 5908
rect 40221 5899 40279 5905
rect 40221 5865 40233 5899
rect 40267 5896 40279 5899
rect 40310 5896 40316 5908
rect 40267 5868 40316 5896
rect 40267 5865 40279 5868
rect 40221 5859 40279 5865
rect 40310 5856 40316 5868
rect 40368 5856 40374 5908
rect 45094 5856 45100 5908
rect 45152 5896 45158 5908
rect 45373 5899 45431 5905
rect 45373 5896 45385 5899
rect 45152 5868 45385 5896
rect 45152 5856 45158 5868
rect 45373 5865 45385 5868
rect 45419 5865 45431 5899
rect 45373 5859 45431 5865
rect 26344 5800 26924 5828
rect 27706 5788 27712 5840
rect 27764 5828 27770 5840
rect 31386 5828 31392 5840
rect 27764 5800 31392 5828
rect 27764 5788 27770 5800
rect 31386 5788 31392 5800
rect 31444 5828 31450 5840
rect 32582 5828 32588 5840
rect 31444 5800 32588 5828
rect 31444 5788 31450 5800
rect 32582 5788 32588 5800
rect 32640 5788 32646 5840
rect 43806 5828 43812 5840
rect 35912 5800 43812 5828
rect 10134 5720 10140 5772
rect 10192 5720 10198 5772
rect 10597 5763 10655 5769
rect 10597 5729 10609 5763
rect 10643 5760 10655 5763
rect 10778 5760 10784 5772
rect 10643 5732 10784 5760
rect 10643 5729 10655 5732
rect 10597 5723 10655 5729
rect 1581 5695 1639 5701
rect 1581 5661 1593 5695
rect 1627 5692 1639 5695
rect 4614 5692 4620 5704
rect 1627 5664 4620 5692
rect 1627 5661 1639 5664
rect 1581 5655 1639 5661
rect 4614 5652 4620 5664
rect 4672 5652 4678 5704
rect 9398 5652 9404 5704
rect 9456 5652 9462 5704
rect 9490 5652 9496 5704
rect 9548 5652 9554 5704
rect 9677 5695 9735 5701
rect 9677 5661 9689 5695
rect 9723 5692 9735 5695
rect 10612 5692 10640 5723
rect 10778 5720 10784 5732
rect 10836 5720 10842 5772
rect 18049 5763 18107 5769
rect 18049 5729 18061 5763
rect 18095 5760 18107 5763
rect 25314 5760 25320 5772
rect 18095 5732 25320 5760
rect 18095 5729 18107 5732
rect 18049 5723 18107 5729
rect 25314 5720 25320 5732
rect 25372 5720 25378 5772
rect 30006 5720 30012 5772
rect 30064 5720 30070 5772
rect 30098 5720 30104 5772
rect 30156 5760 30162 5772
rect 32490 5760 32496 5772
rect 30156 5732 32496 5760
rect 30156 5720 30162 5732
rect 9723 5664 10640 5692
rect 17957 5695 18015 5701
rect 9723 5661 9735 5664
rect 9677 5655 9735 5661
rect 10152 5636 10180 5664
rect 17957 5661 17969 5695
rect 18003 5661 18015 5695
rect 17957 5655 18015 5661
rect 934 5584 940 5636
rect 992 5624 998 5636
rect 1857 5627 1915 5633
rect 1857 5624 1869 5627
rect 992 5596 1869 5624
rect 992 5584 998 5596
rect 1857 5593 1869 5596
rect 1903 5593 1915 5627
rect 1857 5587 1915 5593
rect 10134 5584 10140 5636
rect 10192 5584 10198 5636
rect 17972 5556 18000 5655
rect 18138 5652 18144 5704
rect 18196 5652 18202 5704
rect 18230 5652 18236 5704
rect 18288 5652 18294 5704
rect 19981 5695 20039 5701
rect 19981 5692 19993 5695
rect 19306 5664 19993 5692
rect 18156 5624 18184 5652
rect 19306 5624 19334 5664
rect 19981 5661 19993 5664
rect 20027 5692 20039 5695
rect 20438 5692 20444 5704
rect 20027 5664 20444 5692
rect 20027 5661 20039 5664
rect 19981 5655 20039 5661
rect 20438 5652 20444 5664
rect 20496 5652 20502 5704
rect 25409 5695 25467 5701
rect 25409 5661 25421 5695
rect 25455 5692 25467 5695
rect 27522 5692 27528 5704
rect 25455 5664 27528 5692
rect 25455 5661 25467 5664
rect 25409 5655 25467 5661
rect 25884 5636 25912 5664
rect 27522 5652 27528 5664
rect 27580 5652 27586 5704
rect 27706 5652 27712 5704
rect 27764 5652 27770 5704
rect 29178 5692 29184 5704
rect 27908 5664 29184 5692
rect 22833 5627 22891 5633
rect 18156 5596 19334 5624
rect 20364 5596 20576 5624
rect 20364 5556 20392 5596
rect 17972 5528 20392 5556
rect 20548 5556 20576 5596
rect 22833 5593 22845 5627
rect 22879 5624 22891 5627
rect 24762 5624 24768 5636
rect 22879 5596 24768 5624
rect 22879 5593 22891 5596
rect 22833 5587 22891 5593
rect 24762 5584 24768 5596
rect 24820 5584 24826 5636
rect 25682 5633 25688 5636
rect 25676 5624 25688 5633
rect 25643 5596 25688 5624
rect 25676 5587 25688 5596
rect 25682 5584 25688 5587
rect 25740 5584 25746 5636
rect 25866 5584 25872 5636
rect 25924 5584 25930 5636
rect 26418 5584 26424 5636
rect 26476 5624 26482 5636
rect 27908 5633 27936 5664
rect 29178 5652 29184 5664
rect 29236 5652 29242 5704
rect 30208 5701 30236 5732
rect 31128 5701 31156 5732
rect 32490 5720 32496 5732
rect 32548 5720 32554 5772
rect 33042 5760 33048 5772
rect 32876 5732 33048 5760
rect 30193 5695 30251 5701
rect 30193 5661 30205 5695
rect 30239 5692 30251 5695
rect 30469 5695 30527 5701
rect 30239 5664 30273 5692
rect 30239 5661 30251 5664
rect 30193 5655 30251 5661
rect 30469 5661 30481 5695
rect 30515 5692 30527 5695
rect 31113 5695 31171 5701
rect 30515 5664 31064 5692
rect 30515 5661 30527 5664
rect 30469 5655 30527 5661
rect 27893 5627 27951 5633
rect 27893 5624 27905 5627
rect 26476 5596 27905 5624
rect 26476 5584 26482 5596
rect 27893 5593 27905 5596
rect 27939 5593 27951 5627
rect 30098 5624 30104 5636
rect 27893 5587 27951 5593
rect 28000 5596 30104 5624
rect 28000 5556 28028 5596
rect 30098 5584 30104 5596
rect 30156 5584 30162 5636
rect 31036 5624 31064 5664
rect 31113 5661 31125 5695
rect 31159 5692 31171 5695
rect 31389 5695 31447 5701
rect 31159 5664 31193 5692
rect 31159 5661 31171 5664
rect 31113 5655 31171 5661
rect 31389 5661 31401 5695
rect 31435 5692 31447 5695
rect 31938 5692 31944 5704
rect 31435 5664 31944 5692
rect 31435 5661 31447 5664
rect 31389 5655 31447 5661
rect 31404 5624 31432 5655
rect 31938 5652 31944 5664
rect 31996 5652 32002 5704
rect 32030 5652 32036 5704
rect 32088 5692 32094 5704
rect 32674 5692 32680 5704
rect 32088 5664 32680 5692
rect 32088 5652 32094 5664
rect 32674 5652 32680 5664
rect 32732 5692 32738 5704
rect 32876 5701 32904 5732
rect 33042 5720 33048 5732
rect 33100 5720 33106 5772
rect 32769 5695 32827 5701
rect 32769 5692 32781 5695
rect 32732 5664 32781 5692
rect 32732 5652 32738 5664
rect 32769 5661 32781 5664
rect 32815 5661 32827 5695
rect 32769 5655 32827 5661
rect 32861 5695 32919 5701
rect 32861 5661 32873 5695
rect 32907 5661 32919 5695
rect 32861 5655 32919 5661
rect 30208 5596 30512 5624
rect 31036 5596 31432 5624
rect 20548 5528 28028 5556
rect 28077 5559 28135 5565
rect 28077 5525 28089 5559
rect 28123 5556 28135 5559
rect 28166 5556 28172 5568
rect 28123 5528 28172 5556
rect 28123 5525 28135 5528
rect 28077 5519 28135 5525
rect 28166 5516 28172 5528
rect 28224 5516 28230 5568
rect 29178 5516 29184 5568
rect 29236 5556 29242 5568
rect 30208 5556 30236 5596
rect 29236 5528 30236 5556
rect 29236 5516 29242 5528
rect 30374 5516 30380 5568
rect 30432 5516 30438 5568
rect 30484 5556 30512 5596
rect 32122 5584 32128 5636
rect 32180 5624 32186 5636
rect 32876 5624 32904 5655
rect 32950 5652 32956 5704
rect 33008 5652 33014 5704
rect 33134 5652 33140 5704
rect 33192 5652 33198 5704
rect 34146 5652 34152 5704
rect 34204 5692 34210 5704
rect 34606 5692 34612 5704
rect 34204 5664 34612 5692
rect 34204 5652 34210 5664
rect 34606 5652 34612 5664
rect 34664 5652 34670 5704
rect 35526 5652 35532 5704
rect 35584 5652 35590 5704
rect 35802 5652 35808 5704
rect 35860 5652 35866 5704
rect 35912 5701 35940 5800
rect 43806 5788 43812 5800
rect 43864 5788 43870 5840
rect 45388 5828 45416 5859
rect 45554 5856 45560 5908
rect 45612 5856 45618 5908
rect 46109 5899 46167 5905
rect 46109 5865 46121 5899
rect 46155 5896 46167 5899
rect 46566 5896 46572 5908
rect 46155 5868 46572 5896
rect 46155 5865 46167 5868
rect 46109 5859 46167 5865
rect 46566 5856 46572 5868
rect 46624 5856 46630 5908
rect 46750 5856 46756 5908
rect 46808 5856 46814 5908
rect 55766 5856 55772 5908
rect 55824 5896 55830 5908
rect 56229 5899 56287 5905
rect 56229 5896 56241 5899
rect 55824 5868 56241 5896
rect 55824 5856 55830 5868
rect 56229 5865 56241 5868
rect 56275 5865 56287 5899
rect 58434 5896 58440 5908
rect 56229 5859 56287 5865
rect 56336 5868 58440 5896
rect 45388 5800 46244 5828
rect 36078 5720 36084 5772
rect 36136 5760 36142 5772
rect 36725 5763 36783 5769
rect 36725 5760 36737 5763
rect 36136 5732 36737 5760
rect 36136 5720 36142 5732
rect 36725 5729 36737 5732
rect 36771 5729 36783 5763
rect 36725 5723 36783 5729
rect 37200 5732 40172 5760
rect 37200 5701 37228 5732
rect 35897 5695 35955 5701
rect 35897 5661 35909 5695
rect 35943 5661 35955 5695
rect 35897 5655 35955 5661
rect 37185 5695 37243 5701
rect 37185 5661 37197 5695
rect 37231 5661 37243 5695
rect 39117 5695 39175 5701
rect 39117 5692 39129 5695
rect 37185 5655 37243 5661
rect 37292 5664 39129 5692
rect 32180 5596 32904 5624
rect 34333 5627 34391 5633
rect 32180 5584 32186 5596
rect 34333 5593 34345 5627
rect 34379 5624 34391 5627
rect 35434 5624 35440 5636
rect 34379 5596 35440 5624
rect 34379 5593 34391 5596
rect 34333 5587 34391 5593
rect 35434 5584 35440 5596
rect 35492 5584 35498 5636
rect 36262 5584 36268 5636
rect 36320 5584 36326 5636
rect 31297 5559 31355 5565
rect 31297 5556 31309 5559
rect 30484 5528 31309 5556
rect 31297 5525 31309 5528
rect 31343 5525 31355 5559
rect 31297 5519 31355 5525
rect 32493 5559 32551 5565
rect 32493 5525 32505 5559
rect 32539 5556 32551 5559
rect 32582 5556 32588 5568
rect 32539 5528 32588 5556
rect 32539 5525 32551 5528
rect 32493 5519 32551 5525
rect 32582 5516 32588 5528
rect 32640 5516 32646 5568
rect 33410 5516 33416 5568
rect 33468 5556 33474 5568
rect 37292 5556 37320 5664
rect 39117 5661 39129 5664
rect 39163 5661 39175 5695
rect 39117 5655 39175 5661
rect 39574 5652 39580 5704
rect 39632 5692 39638 5704
rect 40037 5695 40095 5701
rect 40037 5692 40049 5695
rect 39632 5664 40049 5692
rect 39632 5652 39638 5664
rect 40037 5661 40049 5664
rect 40083 5661 40095 5695
rect 40144 5692 40172 5732
rect 40218 5720 40224 5772
rect 40276 5760 40282 5772
rect 46216 5760 46244 5800
rect 46382 5788 46388 5840
rect 46440 5828 46446 5840
rect 47486 5828 47492 5840
rect 46440 5800 47492 5828
rect 46440 5788 46446 5800
rect 47486 5788 47492 5800
rect 47544 5788 47550 5840
rect 54662 5788 54668 5840
rect 54720 5828 54726 5840
rect 56336 5828 56364 5868
rect 58434 5856 58440 5868
rect 58492 5856 58498 5908
rect 54720 5800 56364 5828
rect 54720 5788 54726 5800
rect 53650 5760 53656 5772
rect 40276 5732 46152 5760
rect 40276 5720 40282 5732
rect 43073 5695 43131 5701
rect 43073 5692 43085 5695
rect 40144 5664 43085 5692
rect 40037 5655 40095 5661
rect 43073 5661 43085 5664
rect 43119 5692 43131 5695
rect 43162 5692 43168 5704
rect 43119 5664 43168 5692
rect 43119 5661 43131 5664
rect 43073 5655 43131 5661
rect 43162 5652 43168 5664
rect 43220 5652 43226 5704
rect 44542 5652 44548 5704
rect 44600 5692 44606 5704
rect 44600 5664 45324 5692
rect 44600 5652 44606 5664
rect 37461 5627 37519 5633
rect 37461 5593 37473 5627
rect 37507 5593 37519 5627
rect 37461 5587 37519 5593
rect 33468 5528 37320 5556
rect 37476 5556 37504 5587
rect 38194 5584 38200 5636
rect 38252 5584 38258 5636
rect 38286 5584 38292 5636
rect 38344 5624 38350 5636
rect 38381 5627 38439 5633
rect 38381 5624 38393 5627
rect 38344 5596 38393 5624
rect 38344 5584 38350 5596
rect 38381 5593 38393 5596
rect 38427 5593 38439 5627
rect 38381 5587 38439 5593
rect 38930 5584 38936 5636
rect 38988 5584 38994 5636
rect 42886 5584 42892 5636
rect 42944 5624 42950 5636
rect 43809 5627 43867 5633
rect 43809 5624 43821 5627
rect 42944 5596 43821 5624
rect 42944 5584 42950 5596
rect 43809 5593 43821 5596
rect 43855 5624 43867 5627
rect 44082 5624 44088 5636
rect 43855 5596 44088 5624
rect 43855 5593 43867 5596
rect 43809 5587 43867 5593
rect 44082 5584 44088 5596
rect 44140 5584 44146 5636
rect 45186 5584 45192 5636
rect 45244 5584 45250 5636
rect 45296 5624 45324 5664
rect 46014 5652 46020 5704
rect 46072 5652 46078 5704
rect 45389 5627 45447 5633
rect 45389 5624 45401 5627
rect 45296 5596 45401 5624
rect 45389 5593 45401 5596
rect 45435 5593 45447 5627
rect 46124 5624 46152 5732
rect 46216 5732 53656 5760
rect 46216 5701 46244 5732
rect 53650 5720 53656 5732
rect 53708 5720 53714 5772
rect 56410 5760 56416 5772
rect 56152 5732 56416 5760
rect 46201 5695 46259 5701
rect 46201 5661 46213 5695
rect 46247 5661 46259 5695
rect 46201 5655 46259 5661
rect 46658 5652 46664 5704
rect 46716 5652 46722 5704
rect 56152 5701 56180 5732
rect 56410 5720 56416 5732
rect 56468 5720 56474 5772
rect 56778 5720 56784 5772
rect 56836 5720 56842 5772
rect 56137 5695 56195 5701
rect 56137 5661 56149 5695
rect 56183 5661 56195 5695
rect 56137 5655 56195 5661
rect 56321 5695 56379 5701
rect 56321 5661 56333 5695
rect 56367 5692 56379 5695
rect 56870 5692 56876 5704
rect 56367 5664 56876 5692
rect 56367 5661 56379 5664
rect 56321 5655 56379 5661
rect 56870 5652 56876 5664
rect 56928 5652 56934 5704
rect 57048 5695 57106 5701
rect 57048 5661 57060 5695
rect 57094 5692 57106 5695
rect 58066 5692 58072 5704
rect 57094 5664 58072 5692
rect 57094 5661 57106 5664
rect 57048 5655 57106 5661
rect 58066 5652 58072 5664
rect 58124 5652 58130 5704
rect 57146 5624 57152 5636
rect 46124 5596 57152 5624
rect 45389 5587 45447 5593
rect 57146 5584 57152 5596
rect 57204 5584 57210 5636
rect 57330 5584 57336 5636
rect 57388 5624 57394 5636
rect 58986 5624 58992 5636
rect 57388 5596 58992 5624
rect 57388 5584 57394 5596
rect 58986 5584 58992 5596
rect 59044 5584 59050 5636
rect 38010 5556 38016 5568
rect 37476 5528 38016 5556
rect 33468 5516 33474 5528
rect 38010 5516 38016 5528
rect 38068 5556 38074 5568
rect 40034 5556 40040 5568
rect 38068 5528 40040 5556
rect 38068 5516 38074 5528
rect 40034 5516 40040 5528
rect 40092 5516 40098 5568
rect 43346 5516 43352 5568
rect 43404 5556 43410 5568
rect 47210 5556 47216 5568
rect 43404 5528 47216 5556
rect 43404 5516 43410 5528
rect 47210 5516 47216 5528
rect 47268 5516 47274 5568
rect 55674 5516 55680 5568
rect 55732 5556 55738 5568
rect 58161 5559 58219 5565
rect 58161 5556 58173 5559
rect 55732 5528 58173 5556
rect 55732 5516 55738 5528
rect 58161 5525 58173 5528
rect 58207 5525 58219 5559
rect 58161 5519 58219 5525
rect 1104 5466 58880 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 50294 5466
rect 50346 5414 50358 5466
rect 50410 5414 50422 5466
rect 50474 5414 50486 5466
rect 50538 5414 50550 5466
rect 50602 5414 58880 5466
rect 1104 5392 58880 5414
rect 22649 5355 22707 5361
rect 22649 5321 22661 5355
rect 22695 5352 22707 5355
rect 23106 5352 23112 5364
rect 22695 5324 23112 5352
rect 22695 5321 22707 5324
rect 22649 5315 22707 5321
rect 23106 5312 23112 5324
rect 23164 5312 23170 5364
rect 24302 5312 24308 5364
rect 24360 5352 24366 5364
rect 25038 5352 25044 5364
rect 24360 5324 25044 5352
rect 24360 5312 24366 5324
rect 25038 5312 25044 5324
rect 25096 5312 25102 5364
rect 25314 5312 25320 5364
rect 25372 5352 25378 5364
rect 25501 5355 25559 5361
rect 25501 5352 25513 5355
rect 25372 5324 25513 5352
rect 25372 5312 25378 5324
rect 25501 5321 25513 5324
rect 25547 5321 25559 5355
rect 25501 5315 25559 5321
rect 26326 5312 26332 5364
rect 26384 5312 26390 5364
rect 26418 5312 26424 5364
rect 26476 5312 26482 5364
rect 27632 5324 28994 5352
rect 24388 5287 24446 5293
rect 24388 5253 24400 5287
rect 24434 5284 24446 5287
rect 24670 5284 24676 5296
rect 24434 5256 24676 5284
rect 24434 5253 24446 5256
rect 24388 5247 24446 5253
rect 24670 5244 24676 5256
rect 24728 5244 24734 5296
rect 26050 5244 26056 5296
rect 26108 5244 26114 5296
rect 26237 5287 26295 5293
rect 26237 5253 26249 5287
rect 26283 5284 26295 5287
rect 27632 5284 27660 5324
rect 26283 5256 27660 5284
rect 28966 5284 28994 5324
rect 29178 5312 29184 5364
rect 29236 5312 29242 5364
rect 40218 5352 40224 5364
rect 35452 5324 40224 5352
rect 29822 5284 29828 5296
rect 28966 5256 29828 5284
rect 26283 5253 26295 5256
rect 26237 5247 26295 5253
rect 29822 5244 29828 5256
rect 29880 5244 29886 5296
rect 31113 5287 31171 5293
rect 31113 5253 31125 5287
rect 31159 5284 31171 5287
rect 31159 5256 31432 5284
rect 31159 5253 31171 5256
rect 31113 5247 31171 5253
rect 1581 5219 1639 5225
rect 1581 5185 1593 5219
rect 1627 5216 1639 5219
rect 9582 5216 9588 5228
rect 1627 5188 9588 5216
rect 1627 5185 1639 5188
rect 1581 5179 1639 5185
rect 9582 5176 9588 5188
rect 9640 5176 9646 5228
rect 19794 5176 19800 5228
rect 19852 5176 19858 5228
rect 20806 5176 20812 5228
rect 20864 5216 20870 5228
rect 20993 5219 21051 5225
rect 20993 5216 21005 5219
rect 20864 5188 21005 5216
rect 20864 5176 20870 5188
rect 20993 5185 21005 5188
rect 21039 5185 21051 5219
rect 20993 5179 21051 5185
rect 24118 5176 24124 5228
rect 24176 5176 24182 5228
rect 26602 5176 26608 5228
rect 26660 5176 26666 5228
rect 27614 5176 27620 5228
rect 27672 5216 27678 5228
rect 27801 5219 27859 5225
rect 27801 5216 27813 5219
rect 27672 5188 27813 5216
rect 27672 5176 27678 5188
rect 27801 5185 27813 5188
rect 27847 5216 27859 5219
rect 29178 5216 29184 5228
rect 27847 5188 29184 5216
rect 27847 5185 27859 5188
rect 27801 5179 27859 5185
rect 29178 5176 29184 5188
rect 29236 5176 29242 5228
rect 30285 5219 30343 5225
rect 30285 5185 30297 5219
rect 30331 5216 30343 5219
rect 30650 5216 30656 5228
rect 30331 5188 30656 5216
rect 30331 5185 30343 5188
rect 30285 5179 30343 5185
rect 30650 5176 30656 5188
rect 30708 5176 30714 5228
rect 31294 5176 31300 5228
rect 31352 5176 31358 5228
rect 31404 5216 31432 5256
rect 34606 5244 34612 5296
rect 34664 5244 34670 5296
rect 31754 5216 31760 5228
rect 31404 5188 31760 5216
rect 31754 5176 31760 5188
rect 31812 5216 31818 5228
rect 32214 5216 32220 5228
rect 31812 5188 32220 5216
rect 31812 5176 31818 5188
rect 32214 5176 32220 5188
rect 32272 5176 32278 5228
rect 32582 5176 32588 5228
rect 32640 5176 32646 5228
rect 32674 5176 32680 5228
rect 32732 5216 32738 5228
rect 35452 5216 35480 5324
rect 40218 5312 40224 5324
rect 40276 5312 40282 5364
rect 40494 5312 40500 5364
rect 40552 5312 40558 5364
rect 41230 5312 41236 5364
rect 41288 5312 41294 5364
rect 58253 5355 58311 5361
rect 58253 5352 58265 5355
rect 41386 5324 58265 5352
rect 35618 5244 35624 5296
rect 35676 5284 35682 5296
rect 36170 5284 36176 5296
rect 35676 5256 36176 5284
rect 35676 5244 35682 5256
rect 36170 5244 36176 5256
rect 36228 5284 36234 5296
rect 40236 5284 40264 5312
rect 41386 5284 41414 5324
rect 58253 5321 58265 5324
rect 58299 5321 58311 5355
rect 58253 5315 58311 5321
rect 36228 5256 39160 5284
rect 40236 5256 41414 5284
rect 36228 5244 36234 5256
rect 39132 5228 39160 5256
rect 43438 5244 43444 5296
rect 43496 5244 43502 5296
rect 44450 5244 44456 5296
rect 44508 5284 44514 5296
rect 45189 5287 45247 5293
rect 45189 5284 45201 5287
rect 44508 5256 45201 5284
rect 44508 5244 44514 5256
rect 45189 5253 45201 5256
rect 45235 5253 45247 5287
rect 45189 5247 45247 5253
rect 47946 5244 47952 5296
rect 48004 5284 48010 5296
rect 49602 5284 49608 5296
rect 48004 5256 49608 5284
rect 48004 5244 48010 5256
rect 49602 5244 49608 5256
rect 49660 5244 49666 5296
rect 57330 5244 57336 5296
rect 57388 5244 57394 5296
rect 32732 5188 35480 5216
rect 32732 5176 32738 5188
rect 35526 5176 35532 5228
rect 35584 5176 35590 5228
rect 35802 5176 35808 5228
rect 35860 5176 35866 5228
rect 35897 5219 35955 5225
rect 35897 5185 35909 5219
rect 35943 5185 35955 5219
rect 35897 5179 35955 5185
rect 934 5108 940 5160
rect 992 5148 998 5160
rect 1765 5151 1823 5157
rect 1765 5148 1777 5151
rect 992 5120 1777 5148
rect 992 5108 998 5120
rect 1765 5117 1777 5120
rect 1811 5117 1823 5151
rect 1765 5111 1823 5117
rect 19978 5108 19984 5160
rect 20036 5108 20042 5160
rect 21266 5108 21272 5160
rect 21324 5108 21330 5160
rect 21726 5108 21732 5160
rect 21784 5148 21790 5160
rect 22741 5151 22799 5157
rect 22741 5148 22753 5151
rect 21784 5120 22753 5148
rect 21784 5108 21790 5120
rect 22741 5117 22753 5120
rect 22787 5117 22799 5151
rect 22741 5111 22799 5117
rect 22830 5108 22836 5160
rect 22888 5108 22894 5160
rect 27706 5108 27712 5160
rect 27764 5148 27770 5160
rect 28077 5151 28135 5157
rect 28077 5148 28089 5151
rect 27764 5120 28089 5148
rect 27764 5108 27770 5120
rect 28077 5117 28089 5120
rect 28123 5117 28135 5151
rect 28077 5111 28135 5117
rect 30098 5108 30104 5160
rect 30156 5148 30162 5160
rect 31481 5151 31539 5157
rect 31481 5148 31493 5151
rect 30156 5120 31493 5148
rect 30156 5108 30162 5120
rect 31481 5117 31493 5120
rect 31527 5148 31539 5151
rect 31938 5148 31944 5160
rect 31527 5120 31944 5148
rect 31527 5117 31539 5120
rect 31481 5111 31539 5117
rect 31938 5108 31944 5120
rect 31996 5108 32002 5160
rect 32306 5108 32312 5160
rect 32364 5108 32370 5160
rect 35912 5148 35940 5179
rect 36262 5176 36268 5228
rect 36320 5176 36326 5228
rect 36722 5176 36728 5228
rect 36780 5176 36786 5228
rect 37550 5176 37556 5228
rect 37608 5176 37614 5228
rect 39114 5176 39120 5228
rect 39172 5176 39178 5228
rect 39390 5225 39396 5228
rect 39384 5179 39396 5225
rect 39390 5176 39396 5179
rect 39448 5176 39454 5228
rect 41046 5176 41052 5228
rect 41104 5176 41110 5228
rect 41230 5176 41236 5228
rect 41288 5216 41294 5228
rect 41785 5219 41843 5225
rect 41785 5216 41797 5219
rect 41288 5188 41797 5216
rect 41288 5176 41294 5188
rect 41785 5185 41797 5188
rect 41831 5185 41843 5219
rect 41785 5179 41843 5185
rect 43254 5176 43260 5228
rect 43312 5176 43318 5228
rect 44542 5176 44548 5228
rect 44600 5216 44606 5228
rect 44818 5216 44824 5228
rect 44600 5188 44824 5216
rect 44600 5176 44606 5188
rect 44818 5176 44824 5188
rect 44876 5176 44882 5228
rect 45097 5219 45155 5225
rect 45097 5185 45109 5219
rect 45143 5185 45155 5219
rect 45097 5179 45155 5185
rect 45281 5219 45339 5225
rect 45281 5185 45293 5219
rect 45327 5216 45339 5219
rect 45370 5216 45376 5228
rect 45327 5188 45376 5216
rect 45327 5185 45339 5188
rect 45281 5179 45339 5185
rect 35912 5120 37780 5148
rect 1578 5040 1584 5092
rect 1636 5080 1642 5092
rect 1636 5052 6914 5080
rect 1636 5040 1642 5052
rect 6886 5012 6914 5052
rect 20346 5040 20352 5092
rect 20404 5080 20410 5092
rect 23474 5080 23480 5092
rect 20404 5052 23480 5080
rect 20404 5040 20410 5052
rect 23474 5040 23480 5052
rect 23532 5040 23538 5092
rect 30116 5052 31754 5080
rect 22094 5012 22100 5024
rect 6886 4984 22100 5012
rect 22094 4972 22100 4984
rect 22152 4972 22158 5024
rect 22281 5015 22339 5021
rect 22281 4981 22293 5015
rect 22327 5012 22339 5015
rect 24854 5012 24860 5024
rect 22327 4984 24860 5012
rect 22327 4981 22339 4984
rect 22281 4975 22339 4981
rect 24854 4972 24860 4984
rect 24912 4972 24918 5024
rect 25038 4972 25044 5024
rect 25096 5012 25102 5024
rect 26602 5012 26608 5024
rect 25096 4984 26608 5012
rect 25096 4972 25102 4984
rect 26602 4972 26608 4984
rect 26660 4972 26666 5024
rect 26694 4972 26700 5024
rect 26752 5012 26758 5024
rect 30116 5012 30144 5052
rect 26752 4984 30144 5012
rect 26752 4972 26758 4984
rect 30190 4972 30196 5024
rect 30248 5012 30254 5024
rect 30377 5015 30435 5021
rect 30377 5012 30389 5015
rect 30248 4984 30389 5012
rect 30248 4972 30254 4984
rect 30377 4981 30389 4984
rect 30423 4981 30435 5015
rect 31726 5012 31754 5052
rect 33686 5040 33692 5092
rect 33744 5040 33750 5092
rect 35342 5080 35348 5092
rect 34624 5052 35348 5080
rect 34624 5012 34652 5052
rect 35342 5040 35348 5052
rect 35400 5040 35406 5092
rect 31726 4984 34652 5012
rect 30377 4975 30435 4981
rect 34698 4972 34704 5024
rect 34756 4972 34762 5024
rect 37752 5012 37780 5120
rect 37826 5108 37832 5160
rect 37884 5108 37890 5160
rect 42886 5108 42892 5160
rect 42944 5148 42950 5160
rect 43073 5151 43131 5157
rect 43073 5148 43085 5151
rect 42944 5120 43085 5148
rect 42944 5108 42950 5120
rect 43073 5117 43085 5120
rect 43119 5117 43131 5151
rect 45112 5148 45140 5179
rect 45370 5176 45376 5188
rect 45428 5176 45434 5228
rect 46198 5176 46204 5228
rect 46256 5216 46262 5228
rect 46293 5219 46351 5225
rect 46293 5216 46305 5219
rect 46256 5188 46305 5216
rect 46256 5176 46262 5188
rect 46293 5185 46305 5188
rect 46339 5185 46351 5219
rect 46293 5179 46351 5185
rect 55493 5219 55551 5225
rect 55493 5185 55505 5219
rect 55539 5216 55551 5219
rect 55539 5188 55628 5216
rect 55539 5185 55551 5188
rect 55493 5179 55551 5185
rect 45462 5148 45468 5160
rect 45112 5120 45468 5148
rect 43073 5111 43131 5117
rect 45462 5108 45468 5120
rect 45520 5148 45526 5160
rect 46658 5148 46664 5160
rect 45520 5120 46664 5148
rect 45520 5108 45526 5120
rect 46658 5108 46664 5120
rect 46716 5108 46722 5160
rect 41874 5080 41880 5092
rect 40052 5052 41880 5080
rect 40052 5012 40080 5052
rect 41874 5040 41880 5052
rect 41932 5040 41938 5092
rect 41966 5040 41972 5092
rect 42024 5040 42030 5092
rect 42426 5040 42432 5092
rect 42484 5080 42490 5092
rect 45370 5080 45376 5092
rect 42484 5052 45376 5080
rect 42484 5040 42490 5052
rect 45370 5040 45376 5052
rect 45428 5040 45434 5092
rect 46474 5040 46480 5092
rect 46532 5040 46538 5092
rect 37752 4984 40080 5012
rect 55600 5012 55628 5188
rect 55674 5176 55680 5228
rect 55732 5216 55738 5228
rect 56137 5219 56195 5225
rect 56137 5216 56149 5219
rect 55732 5188 56149 5216
rect 55732 5176 55738 5188
rect 56137 5185 56149 5188
rect 56183 5185 56195 5219
rect 56137 5179 56195 5185
rect 57054 5176 57060 5228
rect 57112 5176 57118 5228
rect 58066 5176 58072 5228
rect 58124 5176 58130 5228
rect 56413 5151 56471 5157
rect 56413 5117 56425 5151
rect 56459 5148 56471 5151
rect 58986 5148 58992 5160
rect 56459 5120 58992 5148
rect 56459 5117 56471 5120
rect 56413 5111 56471 5117
rect 58986 5108 58992 5120
rect 59044 5108 59050 5160
rect 55677 5083 55735 5089
rect 55677 5049 55689 5083
rect 55723 5080 55735 5083
rect 57330 5080 57336 5092
rect 55723 5052 57336 5080
rect 55723 5049 55735 5052
rect 55677 5043 55735 5049
rect 57330 5040 57336 5052
rect 57388 5040 57394 5092
rect 58894 5012 58900 5024
rect 55600 4984 58900 5012
rect 58894 4972 58900 4984
rect 58952 4972 58958 5024
rect 1104 4922 58880 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 58880 4922
rect 1104 4848 58880 4870
rect 15838 4768 15844 4820
rect 15896 4808 15902 4820
rect 17865 4811 17923 4817
rect 15896 4780 17816 4808
rect 15896 4768 15902 4780
rect 11793 4743 11851 4749
rect 11793 4709 11805 4743
rect 11839 4740 11851 4743
rect 12066 4740 12072 4752
rect 11839 4712 12072 4740
rect 11839 4709 11851 4712
rect 11793 4703 11851 4709
rect 12066 4700 12072 4712
rect 12124 4700 12130 4752
rect 17681 4743 17739 4749
rect 17681 4740 17693 4743
rect 12406 4712 17693 4740
rect 10689 4675 10747 4681
rect 10689 4641 10701 4675
rect 10735 4672 10747 4675
rect 12406 4672 12434 4712
rect 17681 4709 17693 4712
rect 17727 4709 17739 4743
rect 17788 4740 17816 4780
rect 17865 4777 17877 4811
rect 17911 4808 17923 4811
rect 18230 4808 18236 4820
rect 17911 4780 18236 4808
rect 17911 4777 17923 4780
rect 17865 4771 17923 4777
rect 18230 4768 18236 4780
rect 18288 4768 18294 4820
rect 21726 4768 21732 4820
rect 21784 4808 21790 4820
rect 22189 4811 22247 4817
rect 22189 4808 22201 4811
rect 21784 4780 22201 4808
rect 21784 4768 21790 4780
rect 22189 4777 22201 4780
rect 22235 4777 22247 4811
rect 22189 4771 22247 4777
rect 27706 4768 27712 4820
rect 27764 4768 27770 4820
rect 27798 4768 27804 4820
rect 27856 4808 27862 4820
rect 38102 4808 38108 4820
rect 27856 4780 38108 4808
rect 27856 4768 27862 4780
rect 38102 4768 38108 4780
rect 38160 4768 38166 4820
rect 39390 4768 39396 4820
rect 39448 4808 39454 4820
rect 39485 4811 39543 4817
rect 39485 4808 39497 4811
rect 39448 4780 39497 4808
rect 39448 4768 39454 4780
rect 39485 4777 39497 4780
rect 39531 4777 39543 4811
rect 39485 4771 39543 4777
rect 39960 4780 41414 4808
rect 22002 4740 22008 4752
rect 17788 4712 22008 4740
rect 17681 4703 17739 4709
rect 22002 4700 22008 4712
rect 22060 4700 22066 4752
rect 24302 4740 24308 4752
rect 22204 4712 24308 4740
rect 10735 4644 12434 4672
rect 17405 4675 17463 4681
rect 10735 4641 10747 4644
rect 10689 4635 10747 4641
rect 17405 4641 17417 4675
rect 17451 4672 17463 4675
rect 18138 4672 18144 4684
rect 17451 4644 18144 4672
rect 17451 4641 17463 4644
rect 17405 4635 17463 4641
rect 18138 4632 18144 4644
rect 18196 4632 18202 4684
rect 22204 4672 22232 4712
rect 24302 4700 24308 4712
rect 24360 4700 24366 4752
rect 25590 4700 25596 4752
rect 25648 4740 25654 4752
rect 31202 4740 31208 4752
rect 25648 4712 31208 4740
rect 25648 4700 25654 4712
rect 31202 4700 31208 4712
rect 31260 4740 31266 4752
rect 32766 4740 32772 4752
rect 31260 4712 32772 4740
rect 31260 4700 31266 4712
rect 32766 4700 32772 4712
rect 32824 4740 32830 4752
rect 33686 4740 33692 4752
rect 32824 4712 33692 4740
rect 32824 4700 32830 4712
rect 33686 4700 33692 4712
rect 33744 4700 33750 4752
rect 35342 4700 35348 4752
rect 35400 4740 35406 4752
rect 37826 4740 37832 4752
rect 35400 4712 37832 4740
rect 35400 4700 35406 4712
rect 19444 4644 22232 4672
rect 1578 4564 1584 4616
rect 1636 4564 1642 4616
rect 18046 4564 18052 4616
rect 18104 4604 18110 4616
rect 19444 4613 19472 4644
rect 22278 4632 22284 4684
rect 22336 4672 22342 4684
rect 22833 4675 22891 4681
rect 22833 4672 22845 4675
rect 22336 4644 22845 4672
rect 22336 4632 22342 4644
rect 22833 4641 22845 4644
rect 22879 4672 22891 4675
rect 23290 4672 23296 4684
rect 22879 4644 23296 4672
rect 22879 4641 22891 4644
rect 22833 4635 22891 4641
rect 23290 4632 23296 4644
rect 23348 4632 23354 4684
rect 24118 4632 24124 4684
rect 24176 4672 24182 4684
rect 24176 4644 24624 4672
rect 24176 4632 24182 4644
rect 24596 4616 24624 4644
rect 27890 4632 27896 4684
rect 27948 4672 27954 4684
rect 28442 4672 28448 4684
rect 27948 4644 28448 4672
rect 27948 4632 27954 4644
rect 28442 4632 28448 4644
rect 28500 4672 28506 4684
rect 36354 4672 36360 4684
rect 28500 4644 36360 4672
rect 28500 4632 28506 4644
rect 18509 4607 18567 4613
rect 18509 4604 18521 4607
rect 18104 4576 18521 4604
rect 18104 4564 18110 4576
rect 18509 4573 18521 4576
rect 18555 4573 18567 4607
rect 18509 4567 18567 4573
rect 19429 4607 19487 4613
rect 19429 4573 19441 4607
rect 19475 4573 19487 4607
rect 19429 4567 19487 4573
rect 20346 4564 20352 4616
rect 20404 4564 20410 4616
rect 20898 4564 20904 4616
rect 20956 4604 20962 4616
rect 21085 4607 21143 4613
rect 21085 4604 21097 4607
rect 20956 4576 21097 4604
rect 20956 4564 20962 4576
rect 21085 4573 21097 4576
rect 21131 4573 21143 4607
rect 22649 4607 22707 4613
rect 22649 4604 22661 4607
rect 21085 4567 21143 4573
rect 22066 4576 22661 4604
rect 934 4496 940 4548
rect 992 4536 998 4548
rect 1857 4539 1915 4545
rect 1857 4536 1869 4539
rect 992 4508 1869 4536
rect 992 4496 998 4508
rect 1857 4505 1869 4508
rect 1903 4505 1915 4539
rect 1857 4499 1915 4505
rect 10318 4496 10324 4548
rect 10376 4536 10382 4548
rect 10505 4539 10563 4545
rect 10505 4536 10517 4539
rect 10376 4508 10517 4536
rect 10376 4496 10382 4508
rect 10505 4505 10517 4508
rect 10551 4505 10563 4539
rect 10505 4499 10563 4505
rect 11422 4496 11428 4548
rect 11480 4536 11486 4548
rect 11609 4539 11667 4545
rect 11609 4536 11621 4539
rect 11480 4508 11621 4536
rect 11480 4496 11486 4508
rect 11609 4505 11621 4508
rect 11655 4505 11667 4539
rect 11609 4499 11667 4505
rect 19705 4539 19763 4545
rect 19705 4505 19717 4539
rect 19751 4536 19763 4539
rect 20254 4536 20260 4548
rect 19751 4508 20260 4536
rect 19751 4505 19763 4508
rect 19705 4499 19763 4505
rect 20254 4496 20260 4508
rect 20312 4496 20318 4548
rect 20625 4539 20683 4545
rect 20625 4505 20637 4539
rect 20671 4536 20683 4539
rect 20806 4536 20812 4548
rect 20671 4508 20812 4536
rect 20671 4505 20683 4508
rect 20625 4499 20683 4505
rect 20806 4496 20812 4508
rect 20864 4496 20870 4548
rect 21358 4496 21364 4548
rect 21416 4496 21422 4548
rect 21913 4539 21971 4545
rect 21913 4505 21925 4539
rect 21959 4536 21971 4539
rect 22066 4536 22094 4576
rect 22649 4573 22661 4576
rect 22695 4604 22707 4607
rect 22695 4576 24532 4604
rect 22695 4573 22707 4576
rect 22649 4567 22707 4573
rect 21959 4508 22094 4536
rect 23477 4539 23535 4545
rect 21959 4505 21971 4508
rect 21913 4499 21971 4505
rect 23477 4505 23489 4539
rect 23523 4536 23535 4539
rect 23566 4536 23572 4548
rect 23523 4508 23572 4536
rect 23523 4505 23535 4508
rect 23477 4499 23535 4505
rect 23566 4496 23572 4508
rect 23624 4496 23630 4548
rect 24504 4536 24532 4576
rect 24578 4564 24584 4616
rect 24636 4564 24642 4616
rect 24854 4613 24860 4616
rect 24848 4604 24860 4613
rect 24815 4576 24860 4604
rect 24848 4567 24860 4576
rect 24854 4564 24860 4567
rect 24912 4564 24918 4616
rect 26605 4607 26663 4613
rect 26605 4573 26617 4607
rect 26651 4604 26663 4607
rect 27062 4604 27068 4616
rect 26651 4576 27068 4604
rect 26651 4573 26663 4576
rect 26605 4567 26663 4573
rect 27062 4564 27068 4576
rect 27120 4564 27126 4616
rect 27249 4607 27307 4613
rect 27249 4573 27261 4607
rect 27295 4604 27307 4607
rect 27706 4604 27712 4616
rect 27295 4576 27712 4604
rect 27295 4573 27307 4576
rect 27249 4567 27307 4573
rect 27706 4564 27712 4576
rect 27764 4564 27770 4616
rect 27982 4564 27988 4616
rect 28040 4564 28046 4616
rect 28074 4564 28080 4616
rect 28132 4564 28138 4616
rect 28166 4564 28172 4616
rect 28224 4564 28230 4616
rect 28353 4607 28411 4613
rect 28353 4573 28365 4607
rect 28399 4604 28411 4607
rect 29454 4604 29460 4616
rect 28399 4576 29460 4604
rect 28399 4573 28411 4576
rect 28353 4567 28411 4573
rect 29454 4564 29460 4576
rect 29512 4564 29518 4616
rect 31021 4607 31079 4613
rect 31021 4573 31033 4607
rect 31067 4604 31079 4607
rect 31754 4604 31760 4616
rect 31067 4576 31760 4604
rect 31067 4573 31079 4576
rect 31021 4567 31079 4573
rect 31754 4564 31760 4576
rect 31812 4564 31818 4616
rect 31956 4613 31984 4644
rect 36354 4632 36360 4644
rect 36412 4632 36418 4684
rect 31941 4607 31999 4613
rect 31941 4573 31953 4607
rect 31987 4573 31999 4607
rect 31941 4567 31999 4573
rect 32033 4607 32091 4613
rect 32033 4573 32045 4607
rect 32079 4573 32091 4607
rect 32033 4567 32091 4573
rect 27798 4536 27804 4548
rect 24504 4508 27804 4536
rect 27798 4496 27804 4508
rect 27856 4496 27862 4548
rect 29546 4536 29552 4548
rect 28092 4508 29552 4536
rect 17126 4428 17132 4480
rect 17184 4468 17190 4480
rect 20898 4468 20904 4480
rect 17184 4440 20904 4468
rect 17184 4428 17190 4440
rect 20898 4428 20904 4440
rect 20956 4428 20962 4480
rect 22554 4428 22560 4480
rect 22612 4428 22618 4480
rect 23290 4428 23296 4480
rect 23348 4468 23354 4480
rect 23753 4471 23811 4477
rect 23753 4468 23765 4471
rect 23348 4440 23765 4468
rect 23348 4428 23354 4440
rect 23753 4437 23765 4440
rect 23799 4437 23811 4471
rect 23753 4431 23811 4437
rect 24762 4428 24768 4480
rect 24820 4468 24826 4480
rect 25961 4471 26019 4477
rect 25961 4468 25973 4471
rect 24820 4440 25973 4468
rect 24820 4428 24826 4440
rect 25961 4437 25973 4440
rect 26007 4437 26019 4471
rect 25961 4431 26019 4437
rect 27982 4428 27988 4480
rect 28040 4468 28046 4480
rect 28092 4468 28120 4508
rect 29546 4496 29552 4508
rect 29604 4496 29610 4548
rect 31205 4539 31263 4545
rect 31205 4505 31217 4539
rect 31251 4536 31263 4539
rect 31846 4536 31852 4548
rect 31251 4508 31852 4536
rect 31251 4505 31263 4508
rect 31205 4499 31263 4505
rect 31846 4496 31852 4508
rect 31904 4496 31910 4548
rect 32048 4536 32076 4567
rect 32122 4564 32128 4616
rect 32180 4564 32186 4616
rect 32309 4607 32367 4613
rect 32309 4573 32321 4607
rect 32355 4573 32367 4607
rect 32309 4567 32367 4573
rect 32214 4536 32220 4548
rect 32048 4508 32220 4536
rect 32214 4496 32220 4508
rect 32272 4496 32278 4548
rect 32324 4536 32352 4567
rect 32398 4564 32404 4616
rect 32456 4604 32462 4616
rect 32861 4607 32919 4613
rect 32861 4604 32873 4607
rect 32456 4576 32873 4604
rect 32456 4564 32462 4576
rect 32861 4573 32873 4576
rect 32907 4604 32919 4607
rect 32950 4604 32956 4616
rect 32907 4576 32956 4604
rect 32907 4573 32919 4576
rect 32861 4567 32919 4573
rect 32950 4564 32956 4576
rect 33008 4564 33014 4616
rect 33502 4564 33508 4616
rect 33560 4604 33566 4616
rect 33597 4607 33655 4613
rect 33597 4604 33609 4607
rect 33560 4576 33609 4604
rect 33560 4564 33566 4576
rect 33597 4573 33609 4576
rect 33643 4604 33655 4607
rect 33686 4604 33692 4616
rect 33643 4576 33692 4604
rect 33643 4573 33655 4576
rect 33597 4567 33655 4573
rect 33686 4564 33692 4576
rect 33744 4564 33750 4616
rect 34054 4564 34060 4616
rect 34112 4604 34118 4616
rect 35158 4604 35164 4616
rect 34112 4576 35164 4604
rect 34112 4564 34118 4576
rect 35158 4564 35164 4576
rect 35216 4564 35222 4616
rect 35710 4564 35716 4616
rect 35768 4604 35774 4616
rect 35894 4604 35900 4616
rect 35768 4576 35900 4604
rect 35768 4564 35774 4576
rect 35894 4564 35900 4576
rect 35952 4564 35958 4616
rect 35986 4564 35992 4616
rect 36044 4564 36050 4616
rect 36648 4604 36676 4712
rect 37826 4700 37832 4712
rect 37884 4700 37890 4752
rect 37182 4632 37188 4684
rect 37240 4632 37246 4684
rect 38013 4675 38071 4681
rect 38013 4672 38025 4675
rect 37292 4644 38025 4672
rect 37001 4607 37059 4613
rect 37001 4604 37013 4607
rect 36648 4576 37013 4604
rect 37001 4573 37013 4576
rect 37047 4573 37059 4607
rect 37001 4567 37059 4573
rect 37090 4564 37096 4616
rect 37148 4604 37154 4616
rect 37292 4604 37320 4644
rect 38013 4641 38025 4644
rect 38059 4641 38071 4675
rect 38013 4635 38071 4641
rect 39117 4675 39175 4681
rect 39117 4641 39129 4675
rect 39163 4672 39175 4675
rect 39960 4672 39988 4780
rect 40037 4743 40095 4749
rect 40037 4709 40049 4743
rect 40083 4709 40095 4743
rect 40037 4703 40095 4709
rect 39163 4644 39988 4672
rect 39163 4641 39175 4644
rect 39117 4635 39175 4641
rect 37148 4576 37320 4604
rect 37148 4564 37154 4576
rect 37734 4564 37740 4616
rect 37792 4604 37798 4616
rect 37829 4607 37887 4613
rect 37829 4604 37841 4607
rect 37792 4576 37841 4604
rect 37792 4564 37798 4576
rect 37829 4573 37841 4576
rect 37875 4573 37887 4607
rect 37829 4567 37887 4573
rect 39301 4607 39359 4613
rect 39301 4573 39313 4607
rect 39347 4604 39359 4607
rect 40052 4604 40080 4703
rect 40126 4700 40132 4752
rect 40184 4740 40190 4752
rect 40862 4740 40868 4752
rect 40184 4712 40868 4740
rect 40184 4700 40190 4712
rect 40862 4700 40868 4712
rect 40920 4700 40926 4752
rect 41386 4740 41414 4780
rect 42150 4768 42156 4820
rect 42208 4768 42214 4820
rect 43162 4768 43168 4820
rect 43220 4808 43226 4820
rect 43533 4811 43591 4817
rect 43533 4808 43545 4811
rect 43220 4780 43545 4808
rect 43220 4768 43226 4780
rect 43533 4777 43545 4780
rect 43579 4777 43591 4811
rect 43533 4771 43591 4777
rect 45925 4811 45983 4817
rect 45925 4777 45937 4811
rect 45971 4808 45983 4811
rect 46842 4808 46848 4820
rect 45971 4780 46848 4808
rect 45971 4777 45983 4780
rect 45925 4771 45983 4777
rect 46842 4768 46848 4780
rect 46900 4768 46906 4820
rect 48682 4768 48688 4820
rect 48740 4768 48746 4820
rect 42886 4740 42892 4752
rect 41386 4712 42892 4740
rect 42886 4700 42892 4712
rect 42944 4700 42950 4752
rect 46753 4743 46811 4749
rect 46753 4709 46765 4743
rect 46799 4740 46811 4743
rect 48222 4740 48228 4752
rect 46799 4712 48228 4740
rect 46799 4709 46811 4712
rect 46753 4703 46811 4709
rect 48222 4700 48228 4712
rect 48280 4700 48286 4752
rect 48406 4700 48412 4752
rect 48464 4740 48470 4752
rect 48464 4712 48590 4740
rect 48464 4700 48470 4712
rect 40218 4632 40224 4684
rect 40276 4672 40282 4684
rect 40497 4675 40555 4681
rect 40497 4672 40509 4675
rect 40276 4644 40509 4672
rect 40276 4632 40282 4644
rect 40497 4641 40509 4644
rect 40543 4641 40555 4675
rect 40497 4635 40555 4641
rect 40678 4632 40684 4684
rect 40736 4632 40742 4684
rect 46382 4632 46388 4684
rect 46440 4672 46446 4684
rect 46440 4644 48452 4672
rect 46440 4632 46446 4644
rect 39347 4576 40080 4604
rect 39347 4573 39359 4576
rect 39301 4567 39359 4573
rect 32324 4508 32904 4536
rect 28040 4440 28120 4468
rect 28040 4428 28046 4440
rect 28258 4428 28264 4480
rect 28316 4468 28322 4480
rect 28813 4471 28871 4477
rect 28813 4468 28825 4471
rect 28316 4440 28825 4468
rect 28316 4428 28322 4440
rect 28813 4437 28825 4440
rect 28859 4437 28871 4471
rect 28813 4431 28871 4437
rect 31665 4471 31723 4477
rect 31665 4437 31677 4471
rect 31711 4468 31723 4471
rect 32582 4468 32588 4480
rect 31711 4440 32588 4468
rect 31711 4437 31723 4440
rect 31665 4431 31723 4437
rect 32582 4428 32588 4440
rect 32640 4428 32646 4480
rect 32876 4468 32904 4508
rect 33042 4496 33048 4548
rect 33100 4496 33106 4548
rect 33781 4539 33839 4545
rect 33781 4505 33793 4539
rect 33827 4536 33839 4539
rect 34146 4536 34152 4548
rect 33827 4508 34152 4536
rect 33827 4505 33839 4508
rect 33781 4499 33839 4505
rect 34146 4496 34152 4508
rect 34204 4496 34210 4548
rect 35345 4539 35403 4545
rect 35345 4505 35357 4539
rect 35391 4536 35403 4539
rect 37550 4536 37556 4548
rect 35391 4508 37556 4536
rect 35391 4505 35403 4508
rect 35345 4499 35403 4505
rect 37550 4496 37556 4508
rect 37608 4496 37614 4548
rect 33134 4468 33140 4480
rect 32876 4440 33140 4468
rect 33134 4428 33140 4440
rect 33192 4428 33198 4480
rect 36173 4471 36231 4477
rect 36173 4437 36185 4471
rect 36219 4468 36231 4471
rect 36354 4468 36360 4480
rect 36219 4440 36360 4468
rect 36219 4437 36231 4440
rect 36173 4431 36231 4437
rect 36354 4428 36360 4440
rect 36412 4428 36418 4480
rect 36630 4428 36636 4480
rect 36688 4428 36694 4480
rect 37093 4471 37151 4477
rect 37093 4437 37105 4471
rect 37139 4468 37151 4471
rect 37182 4468 37188 4480
rect 37139 4440 37188 4468
rect 37139 4437 37151 4440
rect 37093 4431 37151 4437
rect 37182 4428 37188 4440
rect 37240 4428 37246 4480
rect 37844 4468 37872 4567
rect 40402 4564 40408 4616
rect 40460 4604 40466 4616
rect 41969 4607 42027 4613
rect 41969 4604 41981 4607
rect 40460 4576 41981 4604
rect 40460 4564 40466 4576
rect 41969 4573 41981 4576
rect 42015 4573 42027 4607
rect 41969 4567 42027 4573
rect 43346 4564 43352 4616
rect 43404 4604 43410 4616
rect 43441 4607 43499 4613
rect 43441 4604 43453 4607
rect 43404 4576 43453 4604
rect 43404 4564 43410 4576
rect 43441 4573 43453 4576
rect 43487 4573 43499 4607
rect 43441 4567 43499 4573
rect 46474 4564 46480 4616
rect 46532 4604 46538 4616
rect 47213 4607 47271 4613
rect 47213 4604 47225 4607
rect 46532 4576 47225 4604
rect 46532 4564 46538 4576
rect 47213 4573 47225 4576
rect 47259 4573 47271 4607
rect 47213 4567 47271 4573
rect 48038 4564 48044 4616
rect 48096 4564 48102 4616
rect 48189 4607 48247 4613
rect 48189 4573 48201 4607
rect 48235 4604 48247 4607
rect 48235 4573 48268 4604
rect 48189 4567 48268 4573
rect 38654 4496 38660 4548
rect 38712 4536 38718 4548
rect 38712 4508 40632 4536
rect 38712 4496 38718 4508
rect 40126 4468 40132 4480
rect 37844 4440 40132 4468
rect 40126 4428 40132 4440
rect 40184 4428 40190 4480
rect 40310 4428 40316 4480
rect 40368 4468 40374 4480
rect 40405 4471 40463 4477
rect 40405 4468 40417 4471
rect 40368 4440 40417 4468
rect 40368 4428 40374 4440
rect 40405 4437 40417 4440
rect 40451 4437 40463 4471
rect 40604 4468 40632 4508
rect 41322 4496 41328 4548
rect 41380 4496 41386 4548
rect 42058 4496 42064 4548
rect 42116 4536 42122 4548
rect 42797 4539 42855 4545
rect 42797 4536 42809 4539
rect 42116 4508 42809 4536
rect 42116 4496 42122 4508
rect 42797 4505 42809 4508
rect 42843 4505 42855 4539
rect 42797 4499 42855 4505
rect 45646 4496 45652 4548
rect 45704 4536 45710 4548
rect 45833 4539 45891 4545
rect 45833 4536 45845 4539
rect 45704 4508 45845 4536
rect 45704 4496 45710 4508
rect 45833 4505 45845 4508
rect 45879 4505 45891 4539
rect 45833 4499 45891 4505
rect 46014 4496 46020 4548
rect 46072 4536 46078 4548
rect 46569 4539 46627 4545
rect 46569 4536 46581 4539
rect 46072 4508 46581 4536
rect 46072 4496 46078 4508
rect 46569 4505 46581 4508
rect 46615 4505 46627 4539
rect 46569 4499 46627 4505
rect 41417 4471 41475 4477
rect 41417 4468 41429 4471
rect 40604 4440 41429 4468
rect 40405 4431 40463 4437
rect 41417 4437 41429 4440
rect 41463 4437 41475 4471
rect 41417 4431 41475 4437
rect 42886 4428 42892 4480
rect 42944 4428 42950 4480
rect 47394 4428 47400 4480
rect 47452 4428 47458 4480
rect 48240 4468 48268 4567
rect 48314 4564 48320 4616
rect 48372 4564 48378 4616
rect 48424 4613 48452 4644
rect 48562 4613 48590 4712
rect 56410 4632 56416 4684
rect 56468 4672 56474 4684
rect 56778 4672 56784 4684
rect 56468 4644 56784 4672
rect 56468 4632 56474 4644
rect 56778 4632 56784 4644
rect 56836 4672 56842 4684
rect 56873 4675 56931 4681
rect 56873 4672 56885 4675
rect 56836 4644 56885 4672
rect 56836 4632 56842 4644
rect 56873 4641 56885 4644
rect 56919 4641 56931 4675
rect 56873 4635 56931 4641
rect 48409 4607 48467 4613
rect 48409 4573 48421 4607
rect 48455 4573 48467 4607
rect 48409 4567 48467 4573
rect 48545 4607 48603 4613
rect 48545 4573 48557 4607
rect 48591 4604 48603 4607
rect 49234 4604 49240 4616
rect 48591 4576 49240 4604
rect 48591 4573 48603 4576
rect 48545 4567 48603 4573
rect 49234 4564 49240 4576
rect 49292 4564 49298 4616
rect 55398 4564 55404 4616
rect 55456 4604 55462 4616
rect 55953 4607 56011 4613
rect 55953 4604 55965 4607
rect 55456 4576 55965 4604
rect 55456 4564 55462 4576
rect 55953 4573 55965 4576
rect 55999 4604 56011 4607
rect 56318 4604 56324 4616
rect 55999 4576 56324 4604
rect 55999 4573 56011 4576
rect 55953 4567 56011 4573
rect 56318 4564 56324 4576
rect 56376 4564 56382 4616
rect 48332 4536 48360 4564
rect 48774 4536 48780 4548
rect 48332 4508 48780 4536
rect 48774 4496 48780 4508
rect 48832 4496 48838 4548
rect 55490 4496 55496 4548
rect 55548 4536 55554 4548
rect 56229 4539 56287 4545
rect 56229 4536 56241 4539
rect 55548 4508 56241 4536
rect 55548 4496 55554 4508
rect 56229 4505 56241 4508
rect 56275 4505 56287 4539
rect 56229 4499 56287 4505
rect 56962 4496 56968 4548
rect 57020 4536 57026 4548
rect 57118 4539 57176 4545
rect 57118 4536 57130 4539
rect 57020 4508 57130 4536
rect 57020 4496 57026 4508
rect 57118 4505 57130 4508
rect 57164 4505 57176 4539
rect 57118 4499 57176 4505
rect 53466 4468 53472 4480
rect 48240 4440 53472 4468
rect 53466 4428 53472 4440
rect 53524 4428 53530 4480
rect 58250 4428 58256 4480
rect 58308 4428 58314 4480
rect 1104 4378 58880 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 50294 4378
rect 50346 4326 50358 4378
rect 50410 4326 50422 4378
rect 50474 4326 50486 4378
rect 50538 4326 50550 4378
rect 50602 4326 58880 4378
rect 1104 4304 58880 4326
rect 12161 4267 12219 4273
rect 10244 4236 11652 4264
rect 8938 4156 8944 4208
rect 8996 4196 9002 4208
rect 9125 4199 9183 4205
rect 9125 4196 9137 4199
rect 8996 4168 9137 4196
rect 8996 4156 9002 4168
rect 9125 4165 9137 4168
rect 9171 4165 9183 4199
rect 10244 4196 10272 4236
rect 9125 4159 9183 4165
rect 10060 4168 10272 4196
rect 10965 4199 11023 4205
rect 8110 4088 8116 4140
rect 8168 4128 8174 4140
rect 8297 4131 8355 4137
rect 8297 4128 8309 4131
rect 8168 4100 8309 4128
rect 8168 4088 8174 4100
rect 8297 4097 8309 4100
rect 8343 4097 8355 4131
rect 8297 4091 8355 4097
rect 8481 4131 8539 4137
rect 8481 4097 8493 4131
rect 8527 4128 8539 4131
rect 10060 4128 10088 4168
rect 10965 4165 10977 4199
rect 11011 4196 11023 4199
rect 11054 4196 11060 4208
rect 11011 4168 11060 4196
rect 11011 4165 11023 4168
rect 10965 4159 11023 4165
rect 11054 4156 11060 4168
rect 11112 4156 11118 4208
rect 8527 4100 10088 4128
rect 8527 4097 8539 4100
rect 8481 4091 8539 4097
rect 10134 4088 10140 4140
rect 10192 4128 10198 4140
rect 11149 4131 11207 4137
rect 10192 4100 10732 4128
rect 10192 4088 10198 4100
rect 9674 4020 9680 4072
rect 9732 4060 9738 4072
rect 9953 4063 10011 4069
rect 9953 4060 9965 4063
rect 9732 4032 9965 4060
rect 9732 4020 9738 4032
rect 9953 4029 9965 4032
rect 9999 4029 10011 4063
rect 9953 4023 10011 4029
rect 4614 3952 4620 4004
rect 4672 3992 4678 4004
rect 9769 3995 9827 4001
rect 9769 3992 9781 3995
rect 4672 3964 9781 3992
rect 4672 3952 4678 3964
rect 9769 3961 9781 3964
rect 9815 3961 9827 3995
rect 9968 3992 9996 4023
rect 10042 4020 10048 4072
rect 10100 4020 10106 4072
rect 10226 4020 10232 4072
rect 10284 4020 10290 4072
rect 10704 4060 10732 4100
rect 11149 4097 11161 4131
rect 11195 4128 11207 4131
rect 11514 4128 11520 4140
rect 11195 4100 11520 4128
rect 11195 4097 11207 4100
rect 11149 4091 11207 4097
rect 11514 4088 11520 4100
rect 11572 4088 11578 4140
rect 11624 4128 11652 4236
rect 12161 4233 12173 4267
rect 12207 4264 12219 4267
rect 25038 4264 25044 4276
rect 12207 4236 25044 4264
rect 12207 4233 12219 4236
rect 12161 4227 12219 4233
rect 25038 4224 25044 4236
rect 25096 4224 25102 4276
rect 25222 4224 25228 4276
rect 25280 4224 25286 4276
rect 25593 4267 25651 4273
rect 25593 4233 25605 4267
rect 25639 4264 25651 4267
rect 27982 4264 27988 4276
rect 25639 4236 27988 4264
rect 25639 4233 25651 4236
rect 25593 4227 25651 4233
rect 27982 4224 27988 4236
rect 28040 4224 28046 4276
rect 30466 4264 30472 4276
rect 29380 4236 30472 4264
rect 12544 4168 12756 4196
rect 12544 4128 12572 4168
rect 11624 4100 12572 4128
rect 12621 4131 12679 4137
rect 12621 4097 12633 4131
rect 12667 4097 12679 4131
rect 12728 4128 12756 4168
rect 15562 4156 15568 4208
rect 15620 4196 15626 4208
rect 15749 4199 15807 4205
rect 15749 4196 15761 4199
rect 15620 4168 15761 4196
rect 15620 4156 15626 4168
rect 15749 4165 15761 4168
rect 15795 4165 15807 4199
rect 15749 4159 15807 4165
rect 21358 4156 21364 4208
rect 21416 4196 21422 4208
rect 22922 4196 22928 4208
rect 21416 4168 22928 4196
rect 21416 4156 21422 4168
rect 22922 4156 22928 4168
rect 22980 4156 22986 4208
rect 23400 4168 24808 4196
rect 15102 4128 15108 4140
rect 12728 4100 15108 4128
rect 12621 4091 12679 4097
rect 11701 4063 11759 4069
rect 11701 4060 11713 4063
rect 10704 4032 11713 4060
rect 11701 4029 11713 4032
rect 11747 4029 11759 4063
rect 11701 4023 11759 4029
rect 11808 4032 12112 4060
rect 11808 3992 11836 4032
rect 9968 3964 11836 3992
rect 9769 3955 9827 3961
rect 11974 3952 11980 4004
rect 12032 3952 12038 4004
rect 9217 3927 9275 3933
rect 9217 3893 9229 3927
rect 9263 3924 9275 3927
rect 11882 3924 11888 3936
rect 9263 3896 11888 3924
rect 9263 3893 9275 3896
rect 9217 3887 9275 3893
rect 11882 3884 11888 3896
rect 11940 3884 11946 3936
rect 12084 3924 12112 4032
rect 12636 3992 12664 4091
rect 15102 4088 15108 4100
rect 15160 4088 15166 4140
rect 15654 4088 15660 4140
rect 15712 4128 15718 4140
rect 17034 4128 17040 4140
rect 15712 4100 17040 4128
rect 15712 4088 15718 4100
rect 17034 4088 17040 4100
rect 17092 4088 17098 4140
rect 17310 4088 17316 4140
rect 17368 4088 17374 4140
rect 19150 4088 19156 4140
rect 19208 4088 19214 4140
rect 19426 4088 19432 4140
rect 19484 4088 19490 4140
rect 20073 4131 20131 4137
rect 20073 4097 20085 4131
rect 20119 4128 20131 4131
rect 20438 4128 20444 4140
rect 20119 4100 20444 4128
rect 20119 4097 20131 4100
rect 20073 4091 20131 4097
rect 20438 4088 20444 4100
rect 20496 4128 20502 4140
rect 22278 4128 22284 4140
rect 20496 4100 22284 4128
rect 20496 4088 20502 4100
rect 22278 4088 22284 4100
rect 22336 4088 22342 4140
rect 22465 4131 22523 4137
rect 22465 4097 22477 4131
rect 22511 4097 22523 4131
rect 22465 4091 22523 4097
rect 12710 4020 12716 4072
rect 12768 4060 12774 4072
rect 16114 4060 16120 4072
rect 12768 4032 16120 4060
rect 12768 4020 12774 4032
rect 16114 4020 16120 4032
rect 16172 4020 16178 4072
rect 17218 4020 17224 4072
rect 17276 4060 17282 4072
rect 17497 4063 17555 4069
rect 17497 4060 17509 4063
rect 17276 4032 17509 4060
rect 17276 4020 17282 4032
rect 17497 4029 17509 4032
rect 17543 4029 17555 4063
rect 17497 4023 17555 4029
rect 19886 3992 19892 4004
rect 12636 3964 19892 3992
rect 19886 3952 19892 3964
rect 19944 3952 19950 4004
rect 20349 3995 20407 4001
rect 20349 3961 20361 3995
rect 20395 3961 20407 3995
rect 20349 3955 20407 3961
rect 12710 3924 12716 3936
rect 12084 3896 12716 3924
rect 12710 3884 12716 3896
rect 12768 3884 12774 3936
rect 12805 3927 12863 3933
rect 12805 3893 12817 3927
rect 12851 3924 12863 3927
rect 12986 3924 12992 3936
rect 12851 3896 12992 3924
rect 12851 3893 12863 3896
rect 12805 3887 12863 3893
rect 12986 3884 12992 3896
rect 13044 3924 13050 3936
rect 13354 3924 13360 3936
rect 13044 3896 13360 3924
rect 13044 3884 13050 3896
rect 13354 3884 13360 3896
rect 13412 3884 13418 3936
rect 15841 3927 15899 3933
rect 15841 3893 15853 3927
rect 15887 3924 15899 3927
rect 18138 3924 18144 3936
rect 15887 3896 18144 3924
rect 15887 3893 15899 3896
rect 15841 3887 15899 3893
rect 18138 3884 18144 3896
rect 18196 3884 18202 3936
rect 18322 3884 18328 3936
rect 18380 3924 18386 3936
rect 18601 3927 18659 3933
rect 18601 3924 18613 3927
rect 18380 3896 18613 3924
rect 18380 3884 18386 3896
rect 18601 3893 18613 3896
rect 18647 3893 18659 3927
rect 18601 3887 18659 3893
rect 18690 3884 18696 3936
rect 18748 3924 18754 3936
rect 20364 3924 20392 3955
rect 20438 3952 20444 4004
rect 20496 3992 20502 4004
rect 21542 3992 21548 4004
rect 20496 3964 21548 3992
rect 20496 3952 20502 3964
rect 21542 3952 21548 3964
rect 21600 3952 21606 4004
rect 22490 3992 22518 4091
rect 22554 4088 22560 4140
rect 22612 4128 22618 4140
rect 23400 4137 23428 4168
rect 23385 4131 23443 4137
rect 23385 4128 23397 4131
rect 22612 4100 23397 4128
rect 22612 4088 22618 4100
rect 23385 4097 23397 4100
rect 23431 4097 23443 4131
rect 23385 4091 23443 4097
rect 24305 4131 24363 4137
rect 24305 4097 24317 4131
rect 24351 4128 24363 4131
rect 24486 4128 24492 4140
rect 24351 4100 24492 4128
rect 24351 4097 24363 4100
rect 24305 4091 24363 4097
rect 24486 4088 24492 4100
rect 24544 4088 24550 4140
rect 24581 4131 24639 4137
rect 24581 4097 24593 4131
rect 24627 4128 24639 4131
rect 24670 4128 24676 4140
rect 24627 4100 24676 4128
rect 24627 4097 24639 4100
rect 24581 4091 24639 4097
rect 24670 4088 24676 4100
rect 24728 4088 24734 4140
rect 24780 4128 24808 4168
rect 25774 4156 25780 4208
rect 25832 4196 25838 4208
rect 27525 4199 27583 4205
rect 25832 4168 27476 4196
rect 25832 4156 25838 4168
rect 27448 4128 27476 4168
rect 27525 4165 27537 4199
rect 27571 4196 27583 4199
rect 27890 4196 27896 4208
rect 27571 4168 27896 4196
rect 27571 4165 27583 4168
rect 27525 4159 27583 4165
rect 27890 4156 27896 4168
rect 27948 4156 27954 4208
rect 28534 4156 28540 4208
rect 28592 4156 28598 4208
rect 24780 4100 25912 4128
rect 27448 4100 27752 4128
rect 22741 4063 22799 4069
rect 22741 4029 22753 4063
rect 22787 4060 22799 4063
rect 23198 4060 23204 4072
rect 22787 4032 23204 4060
rect 22787 4029 22799 4032
rect 22741 4023 22799 4029
rect 23198 4020 23204 4032
rect 23256 4020 23262 4072
rect 23566 4020 23572 4072
rect 23624 4020 23630 4072
rect 25682 4020 25688 4072
rect 25740 4020 25746 4072
rect 25774 4020 25780 4072
rect 25832 4020 25838 4072
rect 25884 4060 25912 4100
rect 25884 4032 27568 4060
rect 24026 3992 24032 4004
rect 22490 3964 24032 3992
rect 24026 3952 24032 3964
rect 24084 3952 24090 4004
rect 24578 3952 24584 4004
rect 24636 3992 24642 4004
rect 25866 3992 25872 4004
rect 24636 3964 25872 3992
rect 24636 3952 24642 3964
rect 25866 3952 25872 3964
rect 25924 3952 25930 4004
rect 26605 3995 26663 4001
rect 26605 3961 26617 3995
rect 26651 3992 26663 3995
rect 27430 3992 27436 4004
rect 26651 3964 27436 3992
rect 26651 3961 26663 3964
rect 26605 3955 26663 3961
rect 27430 3952 27436 3964
rect 27488 3952 27494 4004
rect 27540 3992 27568 4032
rect 27614 4020 27620 4072
rect 27672 4020 27678 4072
rect 27724 4069 27752 4100
rect 29178 4088 29184 4140
rect 29236 4088 29242 4140
rect 29380 4128 29408 4236
rect 30466 4224 30472 4236
rect 30524 4224 30530 4276
rect 31757 4267 31815 4273
rect 31757 4233 31769 4267
rect 31803 4264 31815 4267
rect 32122 4264 32128 4276
rect 31803 4236 32128 4264
rect 31803 4233 31815 4236
rect 31757 4227 31815 4233
rect 32122 4224 32128 4236
rect 32180 4224 32186 4276
rect 37182 4264 37188 4276
rect 32416 4236 37188 4264
rect 29546 4156 29552 4208
rect 29604 4196 29610 4208
rect 32416 4196 32444 4236
rect 37182 4224 37188 4236
rect 37240 4224 37246 4276
rect 37274 4224 37280 4276
rect 37332 4264 37338 4276
rect 37332 4236 37688 4264
rect 37332 4224 37338 4236
rect 36170 4196 36176 4208
rect 29604 4168 32444 4196
rect 33244 4168 36176 4196
rect 29604 4156 29610 4168
rect 29288 4100 29408 4128
rect 29448 4131 29506 4137
rect 27709 4063 27767 4069
rect 27709 4029 27721 4063
rect 27755 4060 27767 4063
rect 29288 4060 29316 4100
rect 29448 4097 29460 4131
rect 29494 4128 29506 4131
rect 30006 4128 30012 4140
rect 29494 4100 30012 4128
rect 29494 4097 29506 4100
rect 29448 4091 29506 4097
rect 30006 4088 30012 4100
rect 30064 4088 30070 4140
rect 31386 4088 31392 4140
rect 31444 4088 31450 4140
rect 31573 4131 31631 4137
rect 31573 4097 31585 4131
rect 31619 4128 31631 4131
rect 31619 4100 31653 4128
rect 31619 4097 31631 4100
rect 31573 4091 31631 4097
rect 27755 4032 29316 4060
rect 27755 4029 27767 4032
rect 27709 4023 27767 4029
rect 30374 4020 30380 4072
rect 30432 4060 30438 4072
rect 31588 4060 31616 4091
rect 32306 4088 32312 4140
rect 32364 4128 32370 4140
rect 33244 4128 33272 4168
rect 36170 4156 36176 4168
rect 36228 4156 36234 4208
rect 36538 4156 36544 4208
rect 36596 4196 36602 4208
rect 36633 4199 36691 4205
rect 36633 4196 36645 4199
rect 36596 4168 36645 4196
rect 36596 4156 36602 4168
rect 36633 4165 36645 4168
rect 36679 4165 36691 4199
rect 37660 4196 37688 4236
rect 39206 4224 39212 4276
rect 39264 4264 39270 4276
rect 39264 4236 39344 4264
rect 39264 4224 39270 4236
rect 39114 4196 39120 4208
rect 36633 4159 36691 4165
rect 37384 4168 37596 4196
rect 37660 4168 39120 4196
rect 32364 4100 33272 4128
rect 32364 4088 32370 4100
rect 34698 4088 34704 4140
rect 34756 4088 34762 4140
rect 35434 4088 35440 4140
rect 35492 4128 35498 4140
rect 35621 4131 35679 4137
rect 35621 4128 35633 4131
rect 35492 4100 35633 4128
rect 35492 4088 35498 4100
rect 35621 4097 35633 4100
rect 35667 4097 35679 4131
rect 35621 4091 35679 4097
rect 30432 4032 32352 4060
rect 30432 4020 30438 4032
rect 32214 3992 32220 4004
rect 27540 3964 28994 3992
rect 18748 3896 20392 3924
rect 20533 3927 20591 3933
rect 18748 3884 18754 3896
rect 20533 3893 20545 3927
rect 20579 3924 20591 3927
rect 22830 3924 22836 3936
rect 20579 3896 22836 3924
rect 20579 3893 20591 3896
rect 20533 3887 20591 3893
rect 22830 3884 22836 3896
rect 22888 3884 22894 3936
rect 23750 3884 23756 3936
rect 23808 3924 23814 3936
rect 26970 3924 26976 3936
rect 23808 3896 26976 3924
rect 23808 3884 23814 3896
rect 26970 3884 26976 3896
rect 27028 3884 27034 3936
rect 27154 3884 27160 3936
rect 27212 3884 27218 3936
rect 28966 3924 28994 3964
rect 30116 3964 32220 3992
rect 30116 3924 30144 3964
rect 32214 3952 32220 3964
rect 32272 3952 32278 4004
rect 28966 3896 30144 3924
rect 30282 3884 30288 3936
rect 30340 3924 30346 3936
rect 30561 3927 30619 3933
rect 30561 3924 30573 3927
rect 30340 3896 30573 3924
rect 30340 3884 30346 3896
rect 30561 3893 30573 3896
rect 30607 3893 30619 3927
rect 32324 3924 32352 4032
rect 32582 4020 32588 4072
rect 32640 4020 32646 4072
rect 34606 4020 34612 4072
rect 34664 4060 34670 4072
rect 34885 4063 34943 4069
rect 34885 4060 34897 4063
rect 34664 4032 34897 4060
rect 34664 4020 34670 4032
rect 34885 4029 34897 4032
rect 34931 4029 34943 4063
rect 34885 4023 34943 4029
rect 35342 4020 35348 4072
rect 35400 4060 35406 4072
rect 35805 4063 35863 4069
rect 35805 4060 35817 4063
rect 35400 4032 35817 4060
rect 35400 4020 35406 4032
rect 35805 4029 35817 4032
rect 35851 4029 35863 4063
rect 35805 4023 35863 4029
rect 36078 4020 36084 4072
rect 36136 4060 36142 4072
rect 37384 4060 37412 4168
rect 37461 4131 37519 4137
rect 37461 4097 37473 4131
rect 37507 4097 37519 4131
rect 37568 4128 37596 4168
rect 39114 4156 39120 4168
rect 39172 4156 39178 4208
rect 37737 4131 37795 4137
rect 37737 4128 37749 4131
rect 37568 4100 37749 4128
rect 37461 4091 37519 4097
rect 37737 4097 37749 4100
rect 37783 4097 37795 4131
rect 37737 4091 37795 4097
rect 36136 4032 37412 4060
rect 36136 4020 36142 4032
rect 37476 3992 37504 4091
rect 38194 4088 38200 4140
rect 38252 4128 38258 4140
rect 38381 4131 38439 4137
rect 38381 4128 38393 4131
rect 38252 4100 38393 4128
rect 38252 4088 38258 4100
rect 38381 4097 38393 4100
rect 38427 4097 38439 4131
rect 38381 4091 38439 4097
rect 38562 4088 38568 4140
rect 38620 4128 38626 4140
rect 39022 4128 39028 4140
rect 38620 4100 39028 4128
rect 38620 4088 38626 4100
rect 39022 4088 39028 4100
rect 39080 4088 39086 4140
rect 39316 4137 39344 4236
rect 40126 4224 40132 4276
rect 40184 4264 40190 4276
rect 41046 4264 41052 4276
rect 40184 4236 41052 4264
rect 40184 4224 40190 4236
rect 41046 4224 41052 4236
rect 41104 4224 41110 4276
rect 44634 4224 44640 4276
rect 44692 4264 44698 4276
rect 45005 4267 45063 4273
rect 45005 4264 45017 4267
rect 44692 4236 45017 4264
rect 44692 4224 44698 4236
rect 45005 4233 45017 4236
rect 45051 4233 45063 4267
rect 45005 4227 45063 4233
rect 45186 4224 45192 4276
rect 45244 4264 45250 4276
rect 45244 4236 46428 4264
rect 45244 4224 45250 4236
rect 44358 4156 44364 4208
rect 44416 4196 44422 4208
rect 46400 4205 46428 4236
rect 48038 4224 48044 4276
rect 48096 4264 48102 4276
rect 48096 4236 49832 4264
rect 48096 4224 48102 4236
rect 45649 4199 45707 4205
rect 45649 4196 45661 4199
rect 44416 4168 45661 4196
rect 44416 4156 44422 4168
rect 45649 4165 45661 4168
rect 45695 4165 45707 4199
rect 45649 4159 45707 4165
rect 46385 4199 46443 4205
rect 46385 4165 46397 4199
rect 46431 4165 46443 4199
rect 46385 4159 46443 4165
rect 39301 4131 39359 4137
rect 39301 4097 39313 4131
rect 39347 4097 39359 4131
rect 39301 4091 39359 4097
rect 40034 4088 40040 4140
rect 40092 4128 40098 4140
rect 40221 4131 40279 4137
rect 40221 4128 40233 4131
rect 40092 4100 40233 4128
rect 40092 4088 40098 4100
rect 40221 4097 40233 4100
rect 40267 4097 40279 4131
rect 40221 4091 40279 4097
rect 41046 4088 41052 4140
rect 41104 4088 41110 4140
rect 41782 4088 41788 4140
rect 41840 4088 41846 4140
rect 42702 4088 42708 4140
rect 42760 4088 42766 4140
rect 42889 4131 42947 4137
rect 42889 4097 42901 4131
rect 42935 4128 42947 4131
rect 42978 4128 42984 4140
rect 42935 4100 42984 4128
rect 42935 4097 42947 4100
rect 42889 4091 42947 4097
rect 42978 4088 42984 4100
rect 43036 4088 43042 4140
rect 43346 4088 43352 4140
rect 43404 4088 43410 4140
rect 44085 4131 44143 4137
rect 44085 4097 44097 4131
rect 44131 4097 44143 4131
rect 44085 4091 44143 4097
rect 44913 4131 44971 4137
rect 44913 4097 44925 4131
rect 44959 4097 44971 4131
rect 44913 4091 44971 4097
rect 45833 4131 45891 4137
rect 45833 4097 45845 4131
rect 45879 4128 45891 4131
rect 47486 4128 47492 4140
rect 45879 4100 47492 4128
rect 45879 4097 45891 4100
rect 45833 4091 45891 4097
rect 38657 4063 38715 4069
rect 38657 4029 38669 4063
rect 38703 4060 38715 4063
rect 38746 4060 38752 4072
rect 38703 4032 38752 4060
rect 38703 4029 38715 4032
rect 38657 4023 38715 4029
rect 38746 4020 38752 4032
rect 38804 4020 38810 4072
rect 39114 4020 39120 4072
rect 39172 4060 39178 4072
rect 39485 4063 39543 4069
rect 39485 4060 39497 4063
rect 39172 4032 39497 4060
rect 39172 4020 39178 4032
rect 39485 4029 39497 4032
rect 39531 4029 39543 4063
rect 39485 4023 39543 4029
rect 40770 4020 40776 4072
rect 40828 4060 40834 4072
rect 41969 4063 42027 4069
rect 41969 4060 41981 4063
rect 40828 4032 41981 4060
rect 40828 4020 40834 4032
rect 41969 4029 41981 4032
rect 42015 4029 42027 4063
rect 41969 4023 42027 4029
rect 42610 4020 42616 4072
rect 42668 4060 42674 4072
rect 44100 4060 44128 4091
rect 42668 4032 44128 4060
rect 42668 4020 42674 4032
rect 41233 3995 41291 4001
rect 41233 3992 41245 3995
rect 37476 3964 41245 3992
rect 41233 3961 41245 3964
rect 41279 3961 41291 3995
rect 41233 3955 41291 3961
rect 43530 3952 43536 4004
rect 43588 3952 43594 4004
rect 44266 3952 44272 4004
rect 44324 3952 44330 4004
rect 33689 3927 33747 3933
rect 33689 3924 33701 3927
rect 32324 3896 33701 3924
rect 30561 3887 30619 3893
rect 33689 3893 33701 3896
rect 33735 3893 33747 3927
rect 33689 3887 33747 3893
rect 36722 3884 36728 3936
rect 36780 3884 36786 3936
rect 38194 3884 38200 3936
rect 38252 3924 38258 3936
rect 40034 3924 40040 3936
rect 38252 3896 40040 3924
rect 38252 3884 38258 3896
rect 40034 3884 40040 3896
rect 40092 3884 40098 3936
rect 40218 3884 40224 3936
rect 40276 3924 40282 3936
rect 40405 3927 40463 3933
rect 40405 3924 40417 3927
rect 40276 3896 40417 3924
rect 40276 3884 40282 3896
rect 40405 3893 40417 3896
rect 40451 3893 40463 3927
rect 40405 3887 40463 3893
rect 43162 3884 43168 3936
rect 43220 3924 43226 3936
rect 44928 3924 44956 4091
rect 47486 4088 47492 4100
rect 47544 4088 47550 4140
rect 47762 4088 47768 4140
rect 47820 4088 47826 4140
rect 48225 4129 48283 4135
rect 48225 4095 48237 4129
rect 48271 4126 48283 4129
rect 48314 4126 48320 4140
rect 48271 4098 48320 4126
rect 48271 4095 48283 4098
rect 48225 4089 48283 4095
rect 48314 4088 48320 4098
rect 48372 4088 48378 4140
rect 48501 4131 48559 4137
rect 48501 4097 48513 4131
rect 48547 4097 48559 4131
rect 48501 4091 48559 4097
rect 47118 4020 47124 4072
rect 47176 4060 47182 4072
rect 48516 4060 48544 4091
rect 48590 4088 48596 4140
rect 48648 4088 48654 4140
rect 48866 4088 48872 4140
rect 48924 4088 48930 4140
rect 49804 4137 49832 4236
rect 51166 4224 51172 4276
rect 51224 4264 51230 4276
rect 51224 4236 52040 4264
rect 51224 4224 51230 4236
rect 50522 4156 50528 4208
rect 50580 4156 50586 4208
rect 50706 4156 50712 4208
rect 50764 4196 50770 4208
rect 52012 4205 52040 4236
rect 51261 4199 51319 4205
rect 51261 4196 51273 4199
rect 50764 4168 51273 4196
rect 50764 4156 50770 4168
rect 51261 4165 51273 4168
rect 51307 4165 51319 4199
rect 51261 4159 51319 4165
rect 51997 4199 52055 4205
rect 51997 4165 52009 4199
rect 52043 4165 52055 4199
rect 51997 4159 52055 4165
rect 54573 4199 54631 4205
rect 54573 4165 54585 4199
rect 54619 4196 54631 4199
rect 55214 4196 55220 4208
rect 54619 4168 55220 4196
rect 54619 4165 54631 4168
rect 54573 4159 54631 4165
rect 55214 4156 55220 4168
rect 55272 4156 55278 4208
rect 55309 4199 55367 4205
rect 55309 4165 55321 4199
rect 55355 4196 55367 4199
rect 58802 4196 58808 4208
rect 55355 4168 58808 4196
rect 55355 4165 55367 4168
rect 55309 4159 55367 4165
rect 58802 4156 58808 4168
rect 58860 4156 58866 4208
rect 49145 4131 49203 4137
rect 49145 4097 49157 4131
rect 49191 4097 49203 4131
rect 49145 4091 49203 4097
rect 49789 4131 49847 4137
rect 49789 4097 49801 4131
rect 49835 4097 49847 4131
rect 49789 4091 49847 4097
rect 47176 4032 48544 4060
rect 49160 4060 49188 4091
rect 51350 4088 51356 4140
rect 51408 4128 51414 4140
rect 51445 4131 51503 4137
rect 51445 4128 51457 4131
rect 51408 4100 51457 4128
rect 51408 4088 51414 4100
rect 51445 4097 51457 4100
rect 51491 4097 51503 4131
rect 51445 4091 51503 4097
rect 52270 4088 52276 4140
rect 52328 4128 52334 4140
rect 53009 4131 53067 4137
rect 53009 4128 53021 4131
rect 52328 4100 53021 4128
rect 52328 4088 52334 4100
rect 53009 4097 53021 4100
rect 53055 4097 53067 4131
rect 53009 4091 53067 4097
rect 55493 4131 55551 4137
rect 55493 4097 55505 4131
rect 55539 4128 55551 4131
rect 56045 4131 56103 4137
rect 56045 4128 56057 4131
rect 55539 4100 56057 4128
rect 55539 4097 55551 4100
rect 55493 4091 55551 4097
rect 56045 4097 56057 4100
rect 56091 4097 56103 4131
rect 56045 4091 56103 4097
rect 56870 4088 56876 4140
rect 56928 4128 56934 4140
rect 57149 4131 57207 4137
rect 57149 4128 57161 4131
rect 56928 4100 57161 4128
rect 56928 4088 56934 4100
rect 57149 4097 57161 4100
rect 57195 4097 57207 4131
rect 57149 4091 57207 4097
rect 57330 4088 57336 4140
rect 57388 4088 57394 4140
rect 58066 4088 58072 4140
rect 58124 4088 58130 4140
rect 49973 4063 50031 4069
rect 49973 4060 49985 4063
rect 49160 4032 49985 4060
rect 47176 4020 47182 4032
rect 49973 4029 49985 4032
rect 50019 4029 50031 4063
rect 49973 4023 50031 4029
rect 52914 4020 52920 4072
rect 52972 4060 52978 4072
rect 53193 4063 53251 4069
rect 53193 4060 53205 4063
rect 52972 4032 53205 4060
rect 52972 4020 52978 4032
rect 53193 4029 53205 4032
rect 53239 4029 53251 4063
rect 53193 4023 53251 4029
rect 53742 4020 53748 4072
rect 53800 4060 53806 4072
rect 53800 4032 54892 4060
rect 53800 4020 53806 4032
rect 46569 3995 46627 4001
rect 46569 3961 46581 3995
rect 46615 3992 46627 3995
rect 48314 3992 48320 4004
rect 46615 3964 48320 3992
rect 46615 3961 46627 3964
rect 46569 3955 46627 3961
rect 48314 3952 48320 3964
rect 48372 3952 48378 4004
rect 54757 3995 54815 4001
rect 54757 3992 54769 3995
rect 48424 3964 54769 3992
rect 43220 3896 44956 3924
rect 43220 3884 43226 3896
rect 46658 3884 46664 3936
rect 46716 3924 46722 3936
rect 48424 3924 48452 3964
rect 54757 3961 54769 3964
rect 54803 3961 54815 3995
rect 54864 3992 54892 4032
rect 56318 4020 56324 4072
rect 56376 4020 56382 4072
rect 58253 3995 58311 4001
rect 58253 3992 58265 3995
rect 54864 3964 58265 3992
rect 54757 3955 54815 3961
rect 58253 3961 58265 3964
rect 58299 3961 58311 3995
rect 58253 3955 58311 3961
rect 46716 3896 48452 3924
rect 46716 3884 46722 3896
rect 49510 3884 49516 3936
rect 49568 3924 49574 3936
rect 50522 3924 50528 3936
rect 49568 3896 50528 3924
rect 49568 3884 49574 3896
rect 50522 3884 50528 3896
rect 50580 3884 50586 3936
rect 50614 3884 50620 3936
rect 50672 3884 50678 3936
rect 51442 3884 51448 3936
rect 51500 3924 51506 3936
rect 52089 3927 52147 3933
rect 52089 3924 52101 3927
rect 51500 3896 52101 3924
rect 51500 3884 51506 3896
rect 52089 3893 52101 3896
rect 52135 3893 52147 3927
rect 52089 3887 52147 3893
rect 54846 3884 54852 3936
rect 54904 3924 54910 3936
rect 57241 3927 57299 3933
rect 57241 3924 57253 3927
rect 54904 3896 57253 3924
rect 54904 3884 54910 3896
rect 57241 3893 57253 3896
rect 57287 3893 57299 3927
rect 57241 3887 57299 3893
rect 1104 3834 58880 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 58880 3834
rect 1104 3760 58880 3782
rect 8478 3680 8484 3732
rect 8536 3680 8542 3732
rect 9582 3680 9588 3732
rect 9640 3720 9646 3732
rect 9677 3723 9735 3729
rect 9677 3720 9689 3723
rect 9640 3692 9689 3720
rect 9640 3680 9646 3692
rect 9677 3689 9689 3692
rect 9723 3689 9735 3723
rect 9677 3683 9735 3689
rect 9766 3680 9772 3732
rect 9824 3720 9830 3732
rect 12897 3723 12955 3729
rect 9824 3692 12434 3720
rect 9824 3680 9830 3692
rect 7837 3655 7895 3661
rect 7837 3621 7849 3655
rect 7883 3652 7895 3655
rect 9398 3652 9404 3664
rect 7883 3624 9404 3652
rect 7883 3621 7895 3624
rect 7837 3615 7895 3621
rect 9398 3612 9404 3624
rect 9456 3612 9462 3664
rect 10965 3655 11023 3661
rect 10965 3652 10977 3655
rect 9508 3624 10977 3652
rect 7650 3544 7656 3596
rect 7708 3584 7714 3596
rect 9508 3584 9536 3624
rect 10965 3621 10977 3624
rect 11011 3621 11023 3655
rect 12406 3652 12434 3692
rect 12897 3689 12909 3723
rect 12943 3720 12955 3723
rect 13538 3720 13544 3732
rect 12943 3692 13544 3720
rect 12943 3689 12955 3692
rect 12897 3683 12955 3689
rect 13538 3680 13544 3692
rect 13596 3680 13602 3732
rect 14458 3680 14464 3732
rect 14516 3680 14522 3732
rect 15286 3680 15292 3732
rect 15344 3680 15350 3732
rect 16022 3680 16028 3732
rect 16080 3680 16086 3732
rect 16666 3680 16672 3732
rect 16724 3720 16730 3732
rect 20438 3720 20444 3732
rect 16724 3692 20444 3720
rect 16724 3680 16730 3692
rect 20438 3680 20444 3692
rect 20496 3680 20502 3732
rect 20714 3680 20720 3732
rect 20772 3720 20778 3732
rect 27249 3723 27307 3729
rect 27249 3720 27261 3723
rect 20772 3692 27261 3720
rect 20772 3680 20778 3692
rect 27249 3689 27261 3692
rect 27295 3720 27307 3723
rect 27614 3720 27620 3732
rect 27295 3692 27620 3720
rect 27295 3689 27307 3692
rect 27249 3683 27307 3689
rect 27614 3680 27620 3692
rect 27672 3680 27678 3732
rect 27890 3680 27896 3732
rect 27948 3720 27954 3732
rect 27948 3692 31248 3720
rect 27948 3680 27954 3692
rect 17126 3652 17132 3664
rect 12406 3624 17132 3652
rect 10965 3615 11023 3621
rect 17126 3612 17132 3624
rect 17184 3612 17190 3664
rect 17310 3612 17316 3664
rect 17368 3652 17374 3664
rect 20625 3655 20683 3661
rect 20625 3652 20637 3655
rect 17368 3624 20637 3652
rect 17368 3612 17374 3624
rect 20625 3621 20637 3624
rect 20671 3621 20683 3655
rect 20625 3615 20683 3621
rect 20809 3655 20867 3661
rect 20809 3621 20821 3655
rect 20855 3652 20867 3655
rect 21174 3652 21180 3664
rect 20855 3624 21180 3652
rect 20855 3621 20867 3624
rect 20809 3615 20867 3621
rect 21174 3612 21180 3624
rect 21232 3612 21238 3664
rect 22094 3612 22100 3664
rect 22152 3652 22158 3664
rect 22833 3655 22891 3661
rect 22833 3652 22845 3655
rect 22152 3624 22845 3652
rect 22152 3612 22158 3624
rect 22833 3621 22845 3624
rect 22879 3621 22891 3655
rect 22833 3615 22891 3621
rect 23014 3612 23020 3664
rect 23072 3652 23078 3664
rect 23072 3624 23796 3652
rect 23072 3612 23078 3624
rect 7708 3556 9536 3584
rect 7708 3544 7714 3556
rect 9674 3544 9680 3596
rect 9732 3584 9738 3596
rect 9861 3587 9919 3593
rect 9861 3584 9873 3587
rect 9732 3556 9873 3584
rect 9732 3544 9738 3556
rect 9861 3553 9873 3556
rect 9907 3553 9919 3587
rect 9861 3547 9919 3553
rect 10042 3544 10048 3596
rect 10100 3544 10106 3596
rect 10137 3587 10195 3593
rect 10137 3553 10149 3587
rect 10183 3584 10195 3587
rect 11149 3587 11207 3593
rect 11149 3584 11161 3587
rect 10183 3556 11161 3584
rect 10183 3553 10195 3556
rect 10137 3547 10195 3553
rect 11149 3553 11161 3556
rect 11195 3553 11207 3587
rect 11149 3547 11207 3553
rect 12710 3544 12716 3596
rect 12768 3584 12774 3596
rect 22189 3587 22247 3593
rect 12768 3556 16804 3584
rect 12768 3544 12774 3556
rect 7101 3519 7159 3525
rect 7101 3485 7113 3519
rect 7147 3516 7159 3519
rect 9766 3516 9772 3528
rect 7147 3488 9772 3516
rect 7147 3485 7159 3488
rect 7101 3479 7159 3485
rect 9766 3476 9772 3488
rect 9824 3476 9830 3528
rect 9942 3519 10000 3525
rect 9942 3485 9954 3519
rect 9988 3516 10000 3519
rect 16577 3519 16635 3525
rect 9988 3488 16528 3516
rect 9988 3485 10000 3488
rect 9942 3479 10000 3485
rect 6917 3451 6975 3457
rect 6917 3417 6929 3451
rect 6963 3448 6975 3451
rect 7558 3448 7564 3460
rect 6963 3420 7564 3448
rect 6963 3417 6975 3420
rect 6917 3411 6975 3417
rect 7558 3408 7564 3420
rect 7616 3408 7622 3460
rect 7653 3451 7711 3457
rect 7653 3417 7665 3451
rect 7699 3448 7711 3451
rect 8202 3448 8208 3460
rect 7699 3420 8208 3448
rect 7699 3417 7711 3420
rect 7653 3411 7711 3417
rect 8202 3408 8208 3420
rect 8260 3408 8266 3460
rect 8389 3451 8447 3457
rect 8389 3417 8401 3451
rect 8435 3448 8447 3451
rect 8662 3448 8668 3460
rect 8435 3420 8668 3448
rect 8435 3417 8447 3420
rect 8389 3411 8447 3417
rect 8662 3408 8668 3420
rect 8720 3408 8726 3460
rect 10689 3451 10747 3457
rect 10689 3417 10701 3451
rect 10735 3417 10747 3451
rect 10689 3411 10747 3417
rect 11701 3451 11759 3457
rect 11701 3417 11713 3451
rect 11747 3448 11759 3451
rect 11747 3420 12756 3448
rect 11747 3417 11759 3420
rect 11701 3411 11759 3417
rect 10042 3340 10048 3392
rect 10100 3380 10106 3392
rect 10704 3380 10732 3411
rect 10870 3380 10876 3392
rect 10100 3352 10876 3380
rect 10100 3340 10106 3352
rect 10870 3340 10876 3352
rect 10928 3380 10934 3392
rect 11793 3383 11851 3389
rect 11793 3380 11805 3383
rect 10928 3352 11805 3380
rect 10928 3340 10934 3352
rect 11793 3349 11805 3352
rect 11839 3349 11851 3383
rect 11793 3343 11851 3349
rect 12066 3340 12072 3392
rect 12124 3380 12130 3392
rect 12618 3380 12624 3392
rect 12124 3352 12624 3380
rect 12124 3340 12130 3352
rect 12618 3340 12624 3352
rect 12676 3340 12682 3392
rect 12728 3380 12756 3420
rect 12802 3408 12808 3460
rect 12860 3408 12866 3460
rect 13354 3408 13360 3460
rect 13412 3448 13418 3460
rect 13541 3451 13599 3457
rect 13541 3448 13553 3451
rect 13412 3420 13553 3448
rect 13412 3408 13418 3420
rect 13541 3417 13553 3420
rect 13587 3417 13599 3451
rect 13541 3411 13599 3417
rect 14182 3408 14188 3460
rect 14240 3448 14246 3460
rect 14369 3451 14427 3457
rect 14369 3448 14381 3451
rect 14240 3420 14381 3448
rect 14240 3408 14246 3420
rect 14369 3417 14381 3420
rect 14415 3417 14427 3451
rect 14369 3411 14427 3417
rect 15197 3451 15255 3457
rect 15197 3417 15209 3451
rect 15243 3448 15255 3451
rect 15286 3448 15292 3460
rect 15243 3420 15292 3448
rect 15243 3417 15255 3420
rect 15197 3411 15255 3417
rect 15286 3408 15292 3420
rect 15344 3408 15350 3460
rect 15933 3451 15991 3457
rect 15933 3417 15945 3451
rect 15979 3448 15991 3451
rect 16114 3448 16120 3460
rect 15979 3420 16120 3448
rect 15979 3417 15991 3420
rect 15933 3411 15991 3417
rect 16114 3408 16120 3420
rect 16172 3408 16178 3460
rect 16500 3448 16528 3488
rect 16577 3485 16589 3519
rect 16623 3516 16635 3519
rect 16666 3516 16672 3528
rect 16623 3488 16672 3516
rect 16623 3485 16635 3488
rect 16577 3479 16635 3485
rect 16666 3476 16672 3488
rect 16724 3476 16730 3528
rect 16776 3516 16804 3556
rect 17328 3556 22048 3584
rect 17328 3516 17356 3556
rect 16776 3488 17356 3516
rect 17497 3519 17555 3525
rect 17497 3485 17509 3519
rect 17543 3516 17555 3519
rect 17954 3516 17960 3528
rect 17543 3488 17960 3516
rect 17543 3485 17555 3488
rect 17497 3479 17555 3485
rect 17954 3476 17960 3488
rect 18012 3476 18018 3528
rect 18417 3519 18475 3525
rect 18417 3485 18429 3519
rect 18463 3516 18475 3519
rect 18506 3516 18512 3528
rect 18463 3488 18512 3516
rect 18463 3485 18475 3488
rect 18417 3479 18475 3485
rect 18506 3476 18512 3488
rect 18564 3476 18570 3528
rect 19429 3519 19487 3525
rect 19429 3485 19441 3519
rect 19475 3485 19487 3519
rect 19429 3479 19487 3485
rect 19705 3519 19763 3525
rect 19705 3485 19717 3519
rect 19751 3516 19763 3519
rect 20530 3516 20536 3528
rect 19751 3488 20536 3516
rect 19751 3485 19763 3488
rect 19705 3479 19763 3485
rect 16758 3448 16764 3460
rect 16500 3420 16764 3448
rect 16758 3408 16764 3420
rect 16816 3408 16822 3460
rect 16853 3451 16911 3457
rect 16853 3417 16865 3451
rect 16899 3448 16911 3451
rect 16942 3448 16948 3460
rect 16899 3420 16948 3448
rect 16899 3417 16911 3420
rect 16853 3411 16911 3417
rect 16942 3408 16948 3420
rect 17000 3408 17006 3460
rect 17586 3408 17592 3460
rect 17644 3448 17650 3460
rect 17773 3451 17831 3457
rect 17773 3448 17785 3451
rect 17644 3420 17785 3448
rect 17644 3408 17650 3420
rect 17773 3417 17785 3420
rect 17819 3417 17831 3451
rect 17773 3411 17831 3417
rect 18690 3408 18696 3460
rect 18748 3408 18754 3460
rect 19444 3448 19472 3479
rect 20530 3476 20536 3488
rect 20588 3476 20594 3528
rect 21910 3476 21916 3528
rect 21968 3476 21974 3528
rect 20162 3448 20168 3460
rect 19444 3420 20168 3448
rect 20162 3408 20168 3420
rect 20220 3408 20226 3460
rect 20346 3408 20352 3460
rect 20404 3408 20410 3460
rect 22020 3448 22048 3556
rect 22189 3553 22201 3587
rect 22235 3584 22247 3587
rect 23474 3584 23480 3596
rect 22235 3556 23480 3584
rect 22235 3553 22247 3556
rect 22189 3547 22247 3553
rect 23474 3544 23480 3556
rect 23532 3544 23538 3596
rect 23768 3584 23796 3624
rect 23842 3612 23848 3664
rect 23900 3652 23906 3664
rect 25314 3652 25320 3664
rect 23900 3624 25320 3652
rect 23900 3612 23906 3624
rect 25314 3612 25320 3624
rect 25372 3612 25378 3664
rect 29362 3612 29368 3664
rect 29420 3652 29426 3664
rect 31220 3652 31248 3692
rect 31570 3680 31576 3732
rect 31628 3720 31634 3732
rect 32033 3723 32091 3729
rect 32033 3720 32045 3723
rect 31628 3692 32045 3720
rect 31628 3680 31634 3692
rect 32033 3689 32045 3692
rect 32079 3689 32091 3723
rect 32033 3683 32091 3689
rect 32214 3680 32220 3732
rect 32272 3720 32278 3732
rect 35802 3720 35808 3732
rect 32272 3692 35808 3720
rect 32272 3680 32278 3692
rect 35802 3680 35808 3692
rect 35860 3680 35866 3732
rect 36538 3720 36544 3732
rect 36004 3692 36544 3720
rect 32122 3652 32128 3664
rect 29420 3624 31156 3652
rect 31220 3624 32128 3652
rect 29420 3612 29426 3624
rect 23768 3556 25820 3584
rect 22554 3476 22560 3528
rect 22612 3516 22618 3528
rect 23385 3519 23443 3525
rect 23385 3516 23397 3519
rect 22612 3488 23397 3516
rect 22612 3476 22618 3488
rect 23385 3485 23397 3488
rect 23431 3485 23443 3519
rect 23385 3479 23443 3485
rect 23845 3519 23903 3525
rect 23845 3485 23857 3519
rect 23891 3485 23903 3519
rect 23845 3479 23903 3485
rect 22738 3448 22744 3460
rect 22020 3420 22744 3448
rect 22738 3408 22744 3420
rect 22796 3408 22802 3460
rect 23014 3408 23020 3460
rect 23072 3408 23078 3460
rect 23106 3408 23112 3460
rect 23164 3457 23170 3460
rect 23164 3451 23177 3457
rect 23165 3417 23177 3451
rect 23860 3448 23888 3479
rect 24946 3476 24952 3528
rect 25004 3476 25010 3528
rect 25792 3516 25820 3556
rect 25866 3544 25872 3596
rect 25924 3544 25930 3596
rect 26970 3544 26976 3596
rect 27028 3584 27034 3596
rect 30374 3584 30380 3596
rect 27028 3556 30380 3584
rect 27028 3544 27034 3556
rect 30374 3544 30380 3556
rect 30432 3544 30438 3596
rect 30466 3544 30472 3596
rect 30524 3544 30530 3596
rect 25958 3516 25964 3528
rect 25792 3488 25964 3516
rect 25958 3476 25964 3488
rect 26016 3476 26022 3528
rect 26136 3519 26194 3525
rect 26136 3485 26148 3519
rect 26182 3516 26194 3519
rect 27154 3516 27160 3528
rect 26182 3488 27160 3516
rect 26182 3485 26194 3488
rect 26136 3479 26194 3485
rect 27154 3476 27160 3488
rect 27212 3476 27218 3528
rect 28902 3476 28908 3528
rect 28960 3516 28966 3528
rect 30282 3516 30288 3528
rect 28960 3488 30288 3516
rect 28960 3476 28966 3488
rect 30282 3476 30288 3488
rect 30340 3476 30346 3528
rect 31018 3476 31024 3528
rect 31076 3476 31082 3528
rect 31128 3516 31156 3624
rect 32122 3612 32128 3624
rect 32180 3612 32186 3664
rect 31478 3584 31484 3596
rect 31404 3556 31484 3584
rect 31205 3519 31263 3525
rect 31205 3516 31217 3519
rect 31128 3488 31217 3516
rect 31205 3485 31217 3488
rect 31251 3485 31263 3519
rect 31205 3479 31263 3485
rect 31294 3476 31300 3528
rect 31352 3476 31358 3528
rect 31404 3525 31432 3556
rect 31478 3544 31484 3556
rect 31536 3544 31542 3596
rect 32398 3544 32404 3596
rect 32456 3584 32462 3596
rect 33137 3587 33195 3593
rect 33137 3584 33149 3587
rect 32456 3556 33149 3584
rect 32456 3544 32462 3556
rect 33137 3553 33149 3556
rect 33183 3553 33195 3587
rect 33137 3547 33195 3553
rect 34054 3544 34060 3596
rect 34112 3584 34118 3596
rect 35069 3587 35127 3593
rect 35069 3584 35081 3587
rect 34112 3556 35081 3584
rect 34112 3544 34118 3556
rect 35069 3553 35081 3556
rect 35115 3553 35127 3587
rect 35069 3547 35127 3553
rect 31389 3519 31447 3525
rect 31389 3485 31401 3519
rect 31435 3485 31447 3519
rect 32030 3516 32036 3528
rect 31389 3479 31447 3485
rect 31496 3488 32036 3516
rect 25225 3451 25283 3457
rect 23860 3420 25176 3448
rect 23164 3411 23177 3417
rect 23164 3408 23170 3411
rect 12986 3380 12992 3392
rect 12728 3352 12992 3380
rect 12986 3340 12992 3352
rect 13044 3340 13050 3392
rect 13633 3383 13691 3389
rect 13633 3349 13645 3383
rect 13679 3380 13691 3383
rect 16574 3380 16580 3392
rect 13679 3352 16580 3380
rect 13679 3349 13691 3352
rect 13633 3343 13691 3349
rect 16574 3340 16580 3352
rect 16632 3340 16638 3392
rect 19426 3340 19432 3392
rect 19484 3380 19490 3392
rect 20438 3380 20444 3392
rect 19484 3352 20444 3380
rect 19484 3340 19490 3352
rect 20438 3340 20444 3352
rect 20496 3340 20502 3392
rect 23201 3383 23259 3389
rect 23201 3349 23213 3383
rect 23247 3380 23259 3383
rect 23290 3380 23296 3392
rect 23247 3352 23296 3380
rect 23247 3349 23259 3352
rect 23201 3343 23259 3349
rect 23290 3340 23296 3352
rect 23348 3340 23354 3392
rect 23934 3340 23940 3392
rect 23992 3340 23998 3392
rect 25148 3380 25176 3420
rect 25225 3417 25237 3451
rect 25271 3448 25283 3451
rect 25774 3448 25780 3460
rect 25271 3420 25780 3448
rect 25271 3417 25283 3420
rect 25225 3411 25283 3417
rect 25774 3408 25780 3420
rect 25832 3408 25838 3460
rect 26234 3408 26240 3460
rect 26292 3448 26298 3460
rect 28997 3451 29055 3457
rect 28997 3448 29009 3451
rect 26292 3420 29009 3448
rect 26292 3408 26298 3420
rect 28997 3417 29009 3420
rect 29043 3448 29055 3451
rect 30193 3451 30251 3457
rect 29043 3420 30144 3448
rect 29043 3417 29055 3420
rect 28997 3411 29055 3417
rect 27154 3380 27160 3392
rect 25148 3352 27160 3380
rect 27154 3340 27160 3352
rect 27212 3340 27218 3392
rect 28261 3383 28319 3389
rect 28261 3349 28273 3383
rect 28307 3380 28319 3383
rect 28810 3380 28816 3392
rect 28307 3352 28816 3380
rect 28307 3349 28319 3352
rect 28261 3343 28319 3349
rect 28810 3340 28816 3352
rect 28868 3340 28874 3392
rect 29089 3383 29147 3389
rect 29089 3349 29101 3383
rect 29135 3380 29147 3383
rect 29730 3380 29736 3392
rect 29135 3352 29736 3380
rect 29135 3349 29147 3352
rect 29089 3343 29147 3349
rect 29730 3340 29736 3352
rect 29788 3340 29794 3392
rect 29825 3383 29883 3389
rect 29825 3349 29837 3383
rect 29871 3380 29883 3383
rect 30006 3380 30012 3392
rect 29871 3352 30012 3380
rect 29871 3349 29883 3352
rect 29825 3343 29883 3349
rect 30006 3340 30012 3352
rect 30064 3340 30070 3392
rect 30116 3380 30144 3420
rect 30193 3417 30205 3451
rect 30239 3448 30251 3451
rect 30239 3420 30972 3448
rect 30239 3417 30251 3420
rect 30193 3411 30251 3417
rect 30282 3380 30288 3392
rect 30116 3352 30288 3380
rect 30282 3340 30288 3352
rect 30340 3340 30346 3392
rect 30944 3380 30972 3420
rect 31496 3380 31524 3488
rect 32030 3476 32036 3488
rect 32088 3476 32094 3528
rect 32217 3519 32275 3525
rect 32217 3485 32229 3519
rect 32263 3485 32275 3519
rect 32493 3519 32551 3525
rect 32493 3516 32505 3519
rect 32217 3479 32275 3485
rect 32324 3488 32505 3516
rect 32232 3448 32260 3479
rect 31726 3420 32260 3448
rect 30944 3352 31524 3380
rect 31573 3383 31631 3389
rect 31573 3349 31585 3383
rect 31619 3380 31631 3383
rect 31726 3380 31754 3420
rect 31619 3352 31754 3380
rect 31619 3349 31631 3352
rect 31573 3343 31631 3349
rect 32122 3340 32128 3392
rect 32180 3380 32186 3392
rect 32324 3380 32352 3488
rect 32493 3485 32505 3488
rect 32539 3485 32551 3519
rect 32493 3479 32551 3485
rect 32950 3476 32956 3528
rect 33008 3476 33014 3528
rect 33873 3519 33931 3525
rect 33873 3485 33885 3519
rect 33919 3516 33931 3519
rect 33962 3516 33968 3528
rect 33919 3488 33968 3516
rect 33919 3485 33931 3488
rect 33873 3479 33931 3485
rect 33962 3476 33968 3488
rect 34020 3476 34026 3528
rect 34885 3519 34943 3525
rect 34885 3485 34897 3519
rect 34931 3516 34943 3519
rect 36004 3516 36032 3692
rect 36538 3680 36544 3692
rect 36596 3680 36602 3732
rect 37458 3680 37464 3732
rect 37516 3720 37522 3732
rect 37645 3723 37703 3729
rect 37645 3720 37657 3723
rect 37516 3692 37657 3720
rect 37516 3680 37522 3692
rect 37645 3689 37657 3692
rect 37691 3689 37703 3723
rect 37645 3683 37703 3689
rect 37918 3680 37924 3732
rect 37976 3720 37982 3732
rect 38930 3720 38936 3732
rect 37976 3692 38936 3720
rect 37976 3680 37982 3692
rect 38930 3680 38936 3692
rect 38988 3680 38994 3732
rect 42702 3720 42708 3732
rect 39040 3692 42708 3720
rect 38194 3612 38200 3664
rect 38252 3652 38258 3664
rect 39040 3652 39068 3692
rect 42702 3680 42708 3692
rect 42760 3680 42766 3732
rect 42978 3680 42984 3732
rect 43036 3720 43042 3732
rect 44082 3720 44088 3732
rect 43036 3692 44088 3720
rect 43036 3680 43042 3692
rect 44082 3680 44088 3692
rect 44140 3680 44146 3732
rect 44174 3680 44180 3732
rect 44232 3680 44238 3732
rect 44284 3692 47440 3720
rect 41782 3652 41788 3664
rect 38252 3624 39068 3652
rect 39132 3624 41788 3652
rect 38252 3612 38258 3624
rect 36170 3544 36176 3596
rect 36228 3584 36234 3596
rect 36265 3587 36323 3593
rect 36265 3584 36277 3587
rect 36228 3556 36277 3584
rect 36228 3544 36234 3556
rect 36265 3553 36277 3556
rect 36311 3553 36323 3587
rect 36265 3547 36323 3553
rect 37366 3544 37372 3596
rect 37424 3584 37430 3596
rect 39132 3584 39160 3624
rect 41782 3612 41788 3624
rect 41840 3612 41846 3664
rect 44284 3652 44312 3692
rect 47302 3652 47308 3664
rect 42628 3624 44312 3652
rect 46952 3624 47308 3652
rect 42628 3593 42656 3624
rect 42613 3587 42671 3593
rect 37424 3556 39160 3584
rect 39316 3556 42564 3584
rect 37424 3544 37430 3556
rect 34931 3488 36032 3516
rect 34931 3485 34943 3488
rect 34885 3479 34943 3485
rect 36354 3476 36360 3528
rect 36412 3516 36418 3528
rect 36521 3519 36579 3525
rect 36521 3516 36533 3519
rect 36412 3488 36533 3516
rect 36412 3476 36418 3488
rect 36521 3485 36533 3488
rect 36567 3485 36579 3519
rect 39206 3516 39212 3528
rect 36521 3479 36579 3485
rect 36648 3488 39212 3516
rect 32401 3451 32459 3457
rect 32401 3417 32413 3451
rect 32447 3448 32459 3451
rect 32858 3448 32864 3460
rect 32447 3420 32864 3448
rect 32447 3417 32459 3420
rect 32401 3411 32459 3417
rect 32858 3408 32864 3420
rect 32916 3408 32922 3460
rect 33226 3408 33232 3460
rect 33284 3448 33290 3460
rect 34149 3451 34207 3457
rect 34149 3448 34161 3451
rect 33284 3420 34161 3448
rect 33284 3408 33290 3420
rect 34149 3417 34161 3420
rect 34195 3417 34207 3451
rect 36648 3448 36676 3488
rect 39206 3476 39212 3488
rect 39264 3476 39270 3528
rect 34149 3411 34207 3417
rect 34256 3420 36676 3448
rect 34256 3380 34284 3420
rect 38470 3408 38476 3460
rect 38528 3448 38534 3460
rect 38565 3451 38623 3457
rect 38565 3448 38577 3451
rect 38528 3420 38577 3448
rect 38528 3408 38534 3420
rect 38565 3417 38577 3420
rect 38611 3417 38623 3451
rect 38565 3411 38623 3417
rect 39114 3408 39120 3460
rect 39172 3448 39178 3460
rect 39316 3448 39344 3556
rect 39390 3476 39396 3528
rect 39448 3516 39454 3528
rect 42536 3525 42564 3556
rect 42613 3553 42625 3587
rect 42659 3553 42671 3587
rect 42613 3547 42671 3553
rect 43438 3544 43444 3596
rect 43496 3584 43502 3596
rect 43496 3556 45324 3584
rect 43496 3544 43502 3556
rect 42521 3519 42579 3525
rect 39448 3488 41828 3516
rect 39448 3476 39454 3488
rect 39172 3420 39344 3448
rect 39172 3408 39178 3420
rect 40034 3408 40040 3460
rect 40092 3448 40098 3460
rect 40129 3451 40187 3457
rect 40129 3448 40141 3451
rect 40092 3420 40141 3448
rect 40092 3408 40098 3420
rect 40129 3417 40141 3420
rect 40175 3448 40187 3451
rect 40865 3451 40923 3457
rect 40865 3448 40877 3451
rect 40175 3420 40877 3448
rect 40175 3417 40187 3420
rect 40129 3411 40187 3417
rect 40865 3417 40877 3420
rect 40911 3448 40923 3451
rect 41046 3448 41052 3460
rect 40911 3420 41052 3448
rect 40911 3417 40923 3420
rect 40865 3411 40923 3417
rect 41046 3408 41052 3420
rect 41104 3408 41110 3460
rect 32180 3352 34284 3380
rect 32180 3340 32186 3352
rect 35986 3340 35992 3392
rect 36044 3380 36050 3392
rect 40221 3383 40279 3389
rect 40221 3380 40233 3383
rect 36044 3352 40233 3380
rect 36044 3340 36050 3352
rect 40221 3349 40233 3352
rect 40267 3349 40279 3383
rect 40221 3343 40279 3349
rect 40954 3340 40960 3392
rect 41012 3340 41018 3392
rect 41800 3380 41828 3488
rect 42521 3485 42533 3519
rect 42567 3516 42579 3519
rect 42794 3516 42800 3528
rect 42567 3488 42800 3516
rect 42567 3485 42579 3488
rect 42521 3479 42579 3485
rect 42794 3476 42800 3488
rect 42852 3476 42858 3528
rect 42886 3476 42892 3528
rect 42944 3476 42950 3528
rect 42978 3476 42984 3528
rect 43036 3476 43042 3528
rect 43070 3476 43076 3528
rect 43128 3516 43134 3528
rect 43714 3525 43720 3528
rect 43533 3519 43591 3525
rect 43533 3516 43545 3519
rect 43128 3488 43545 3516
rect 43128 3476 43134 3488
rect 43533 3485 43545 3488
rect 43579 3485 43591 3519
rect 43533 3479 43591 3485
rect 43681 3519 43720 3525
rect 43681 3485 43693 3519
rect 43681 3479 43720 3485
rect 43714 3476 43720 3479
rect 43772 3476 43778 3528
rect 43898 3476 43904 3528
rect 43956 3476 43962 3528
rect 44039 3519 44097 3525
rect 44039 3485 44051 3519
rect 44085 3516 44097 3519
rect 44174 3516 44180 3528
rect 44085 3488 44180 3516
rect 44085 3485 44097 3488
rect 44039 3479 44097 3485
rect 44174 3476 44180 3488
rect 44232 3476 44238 3528
rect 45296 3525 45324 3556
rect 46952 3525 46980 3624
rect 47302 3612 47308 3624
rect 47360 3612 47366 3664
rect 47412 3652 47440 3692
rect 47578 3680 47584 3732
rect 47636 3680 47642 3732
rect 49970 3680 49976 3732
rect 50028 3720 50034 3732
rect 50525 3723 50583 3729
rect 50525 3720 50537 3723
rect 50028 3692 50537 3720
rect 50028 3680 50034 3692
rect 50525 3689 50537 3692
rect 50571 3689 50583 3723
rect 50525 3683 50583 3689
rect 53466 3680 53472 3732
rect 53524 3680 53530 3732
rect 54202 3680 54208 3732
rect 54260 3680 54266 3732
rect 57793 3723 57851 3729
rect 57793 3720 57805 3723
rect 54404 3692 57805 3720
rect 50614 3652 50620 3664
rect 47412 3624 50620 3652
rect 50614 3612 50620 3624
rect 50672 3612 50678 3664
rect 52089 3655 52147 3661
rect 52089 3621 52101 3655
rect 52135 3652 52147 3655
rect 52178 3652 52184 3664
rect 52135 3624 52184 3652
rect 52135 3621 52147 3624
rect 52089 3615 52147 3621
rect 52178 3612 52184 3624
rect 52236 3612 52242 3664
rect 53650 3612 53656 3664
rect 53708 3652 53714 3664
rect 54404 3652 54432 3692
rect 57793 3689 57805 3692
rect 57839 3689 57851 3723
rect 57793 3683 57851 3689
rect 53708 3624 54432 3652
rect 53708 3612 53714 3624
rect 52825 3587 52883 3593
rect 52825 3584 52837 3587
rect 47320 3556 52837 3584
rect 45281 3519 45339 3525
rect 45281 3485 45293 3519
rect 45327 3485 45339 3519
rect 46937 3519 46995 3525
rect 45281 3479 45339 3485
rect 45388 3488 46428 3516
rect 41874 3408 41880 3460
rect 41932 3408 41938 3460
rect 42812 3448 42840 3476
rect 43809 3451 43867 3457
rect 43809 3448 43821 3451
rect 42812 3420 43821 3448
rect 43640 3392 43668 3420
rect 43809 3417 43821 3420
rect 43855 3417 43867 3451
rect 43809 3411 43867 3417
rect 44450 3408 44456 3460
rect 44508 3448 44514 3460
rect 45388 3448 45416 3488
rect 44508 3420 45416 3448
rect 44508 3408 44514 3420
rect 45462 3408 45468 3460
rect 45520 3448 45526 3460
rect 46293 3451 46351 3457
rect 46293 3448 46305 3451
rect 45520 3420 46305 3448
rect 45520 3408 45526 3420
rect 46293 3417 46305 3420
rect 46339 3417 46351 3451
rect 46400 3448 46428 3488
rect 46937 3485 46949 3519
rect 46983 3485 46995 3519
rect 46937 3479 46995 3485
rect 47085 3519 47143 3525
rect 47085 3485 47097 3519
rect 47131 3516 47143 3519
rect 47320 3516 47348 3556
rect 52825 3553 52837 3556
rect 52871 3553 52883 3587
rect 52825 3547 52883 3553
rect 57330 3544 57336 3596
rect 57388 3584 57394 3596
rect 57425 3587 57483 3593
rect 57425 3584 57437 3587
rect 57388 3556 57437 3584
rect 57388 3544 57394 3556
rect 57425 3553 57437 3556
rect 57471 3553 57483 3587
rect 57425 3547 57483 3553
rect 47131 3488 47348 3516
rect 47131 3485 47143 3488
rect 47085 3479 47143 3485
rect 47394 3476 47400 3528
rect 47452 3525 47458 3528
rect 47452 3516 47460 3525
rect 47452 3488 47497 3516
rect 47452 3479 47460 3488
rect 47452 3476 47458 3479
rect 47946 3476 47952 3528
rect 48004 3516 48010 3528
rect 48133 3519 48191 3525
rect 48133 3516 48145 3519
rect 48004 3488 48145 3516
rect 48004 3476 48010 3488
rect 48133 3485 48145 3488
rect 48179 3485 48191 3519
rect 48133 3479 48191 3485
rect 48590 3476 48596 3528
rect 48648 3476 48654 3528
rect 48774 3476 48780 3528
rect 48832 3476 48838 3528
rect 49145 3519 49203 3525
rect 49145 3485 49157 3519
rect 49191 3485 49203 3519
rect 49145 3479 49203 3485
rect 47210 3448 47216 3460
rect 46400 3420 47216 3448
rect 46293 3411 46351 3417
rect 47210 3408 47216 3420
rect 47268 3408 47274 3460
rect 47302 3408 47308 3460
rect 47360 3408 47366 3460
rect 49160 3448 49188 3479
rect 49234 3476 49240 3528
rect 49292 3476 49298 3528
rect 49970 3476 49976 3528
rect 50028 3516 50034 3528
rect 50341 3519 50399 3525
rect 50341 3516 50353 3519
rect 50028 3488 50353 3516
rect 50028 3476 50034 3488
rect 50341 3485 50353 3488
rect 50387 3485 50399 3519
rect 50341 3479 50399 3485
rect 50430 3476 50436 3528
rect 50488 3516 50494 3528
rect 51353 3519 51411 3525
rect 51353 3516 51365 3519
rect 50488 3488 51365 3516
rect 50488 3476 50494 3488
rect 51353 3485 51365 3488
rect 51399 3485 51411 3519
rect 51353 3479 51411 3485
rect 51442 3476 51448 3528
rect 51500 3516 51506 3528
rect 52641 3519 52699 3525
rect 52641 3516 52653 3519
rect 51500 3488 52653 3516
rect 51500 3476 51506 3488
rect 52641 3485 52653 3488
rect 52687 3485 52699 3519
rect 52641 3479 52699 3485
rect 53098 3476 53104 3528
rect 53156 3516 53162 3528
rect 54113 3519 54171 3525
rect 54113 3516 54125 3519
rect 53156 3488 54125 3516
rect 53156 3476 53162 3488
rect 54113 3485 54125 3488
rect 54159 3485 54171 3519
rect 54113 3479 54171 3485
rect 54754 3476 54760 3528
rect 54812 3476 54818 3528
rect 54941 3519 54999 3525
rect 54941 3485 54953 3519
rect 54987 3516 54999 3519
rect 55490 3516 55496 3528
rect 54987 3488 55496 3516
rect 54987 3485 54999 3488
rect 54941 3479 54999 3485
rect 55490 3476 55496 3488
rect 55548 3476 55554 3528
rect 55585 3519 55643 3525
rect 55585 3485 55597 3519
rect 55631 3516 55643 3519
rect 56410 3516 56416 3528
rect 55631 3488 56416 3516
rect 55631 3485 55643 3488
rect 55585 3479 55643 3485
rect 56410 3476 56416 3488
rect 56468 3476 56474 3528
rect 57609 3519 57667 3525
rect 57609 3485 57621 3519
rect 57655 3485 57667 3519
rect 57609 3479 57667 3485
rect 48148 3420 49188 3448
rect 42978 3380 42984 3392
rect 41800 3352 42984 3380
rect 42978 3340 42984 3352
rect 43036 3340 43042 3392
rect 43622 3340 43628 3392
rect 43680 3340 43686 3392
rect 44082 3340 44088 3392
rect 44140 3380 44146 3392
rect 45373 3383 45431 3389
rect 45373 3380 45385 3383
rect 44140 3352 45385 3380
rect 44140 3340 44146 3352
rect 45373 3349 45385 3352
rect 45419 3349 45431 3383
rect 45373 3343 45431 3349
rect 46385 3383 46443 3389
rect 46385 3349 46397 3383
rect 46431 3380 46443 3383
rect 48148 3380 48176 3420
rect 49786 3408 49792 3460
rect 49844 3448 49850 3460
rect 51169 3451 51227 3457
rect 51169 3448 51181 3451
rect 49844 3420 51181 3448
rect 49844 3408 49850 3420
rect 51169 3417 51181 3420
rect 51215 3417 51227 3451
rect 51169 3411 51227 3417
rect 51905 3451 51963 3457
rect 51905 3417 51917 3451
rect 51951 3417 51963 3451
rect 51905 3411 51963 3417
rect 46431 3352 48176 3380
rect 46431 3349 46443 3352
rect 46385 3343 46443 3349
rect 50062 3340 50068 3392
rect 50120 3380 50126 3392
rect 51920 3380 51948 3411
rect 51994 3408 52000 3460
rect 52052 3448 52058 3460
rect 53377 3451 53435 3457
rect 53377 3448 53389 3451
rect 52052 3420 53389 3448
rect 52052 3408 52058 3420
rect 53377 3417 53389 3420
rect 53423 3417 53435 3451
rect 53377 3411 53435 3417
rect 54849 3451 54907 3457
rect 54849 3417 54861 3451
rect 54895 3448 54907 3451
rect 55830 3451 55888 3457
rect 55830 3448 55842 3451
rect 54895 3420 55842 3448
rect 54895 3417 54907 3420
rect 54849 3411 54907 3417
rect 55830 3417 55842 3420
rect 55876 3417 55888 3451
rect 55830 3411 55888 3417
rect 56870 3408 56876 3460
rect 56928 3448 56934 3460
rect 57624 3448 57652 3479
rect 56928 3420 57652 3448
rect 56928 3408 56934 3420
rect 50120 3352 51948 3380
rect 50120 3340 50126 3352
rect 56778 3340 56784 3392
rect 56836 3380 56842 3392
rect 56965 3383 57023 3389
rect 56965 3380 56977 3383
rect 56836 3352 56977 3380
rect 56836 3340 56842 3352
rect 56965 3349 56977 3352
rect 57011 3349 57023 3383
rect 56965 3343 57023 3349
rect 1104 3290 58880 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 50294 3290
rect 50346 3238 50358 3290
rect 50410 3238 50422 3290
rect 50474 3238 50486 3290
rect 50538 3238 50550 3290
rect 50602 3238 58880 3290
rect 1104 3216 58880 3238
rect 7650 3136 7656 3188
rect 7708 3136 7714 3188
rect 12066 3176 12072 3188
rect 8220 3148 12072 3176
rect 5997 3111 6055 3117
rect 5997 3077 6009 3111
rect 6043 3108 6055 3111
rect 8220 3108 8248 3148
rect 12066 3136 12072 3148
rect 12124 3136 12130 3188
rect 12161 3179 12219 3185
rect 12161 3145 12173 3179
rect 12207 3145 12219 3179
rect 12161 3139 12219 3145
rect 6043 3080 8248 3108
rect 8297 3111 8355 3117
rect 6043 3077 6055 3080
rect 5997 3071 6055 3077
rect 8297 3077 8309 3111
rect 8343 3108 8355 3111
rect 9582 3108 9588 3120
rect 8343 3080 9588 3108
rect 8343 3077 8355 3080
rect 8297 3071 8355 3077
rect 9582 3068 9588 3080
rect 9640 3068 9646 3120
rect 9677 3111 9735 3117
rect 9677 3077 9689 3111
rect 9723 3108 9735 3111
rect 10042 3108 10048 3120
rect 9723 3080 10048 3108
rect 9723 3077 9735 3080
rect 9677 3071 9735 3077
rect 10042 3068 10048 3080
rect 10100 3068 10106 3120
rect 11974 3108 11980 3120
rect 10152 3080 11980 3108
rect 5813 3043 5871 3049
rect 5813 3009 5825 3043
rect 5859 3040 5871 3043
rect 5902 3040 5908 3052
rect 5859 3012 5908 3040
rect 5859 3009 5871 3012
rect 5813 3003 5871 3009
rect 5902 3000 5908 3012
rect 5960 3000 5966 3052
rect 6822 3000 6828 3052
rect 6880 3000 6886 3052
rect 7561 3043 7619 3049
rect 7561 3009 7573 3043
rect 7607 3040 7619 3043
rect 7926 3040 7932 3052
rect 7607 3012 7932 3040
rect 7607 3009 7619 3012
rect 7561 3003 7619 3009
rect 7926 3000 7932 3012
rect 7984 3000 7990 3052
rect 9030 3000 9036 3052
rect 9088 3000 9094 3052
rect 9122 3000 9128 3052
rect 9180 3040 9186 3052
rect 9217 3043 9275 3049
rect 9217 3040 9229 3043
rect 9180 3012 9229 3040
rect 9180 3000 9186 3012
rect 9217 3009 9229 3012
rect 9263 3009 9275 3043
rect 10152 3040 10180 3080
rect 11974 3068 11980 3080
rect 12032 3068 12038 3120
rect 12176 3108 12204 3139
rect 13814 3136 13820 3188
rect 13872 3136 13878 3188
rect 15289 3179 15347 3185
rect 15289 3145 15301 3179
rect 15335 3176 15347 3179
rect 18598 3176 18604 3188
rect 15335 3148 18604 3176
rect 15335 3145 15347 3148
rect 15289 3139 15347 3145
rect 18598 3136 18604 3148
rect 18656 3136 18662 3188
rect 21910 3176 21916 3188
rect 18708 3148 21916 3176
rect 17954 3108 17960 3120
rect 12176 3080 17960 3108
rect 17954 3068 17960 3080
rect 18012 3068 18018 3120
rect 18708 3117 18736 3148
rect 21910 3136 21916 3148
rect 21968 3136 21974 3188
rect 23750 3176 23756 3188
rect 22204 3148 23756 3176
rect 18693 3111 18751 3117
rect 18693 3077 18705 3111
rect 18739 3077 18751 3111
rect 22094 3108 22100 3120
rect 18693 3071 18751 3077
rect 19352 3080 22100 3108
rect 9217 3003 9275 3009
rect 9600 3012 10180 3040
rect 8481 2975 8539 2981
rect 8481 2941 8493 2975
rect 8527 2972 8539 2975
rect 9600 2972 9628 3012
rect 10962 3000 10968 3052
rect 11020 3000 11026 3052
rect 11149 3043 11207 3049
rect 11149 3009 11161 3043
rect 11195 3040 11207 3043
rect 12989 3043 13047 3049
rect 11195 3012 12296 3040
rect 11195 3009 11207 3012
rect 11149 3003 11207 3009
rect 8527 2944 9628 2972
rect 10137 2975 10195 2981
rect 8527 2941 8539 2944
rect 8481 2935 8539 2941
rect 10137 2941 10149 2975
rect 10183 2972 10195 2975
rect 10226 2972 10232 2984
rect 10183 2944 10232 2972
rect 10183 2941 10195 2944
rect 10137 2935 10195 2941
rect 10226 2932 10232 2944
rect 10284 2932 10290 2984
rect 10870 2932 10876 2984
rect 10928 2972 10934 2984
rect 11701 2975 11759 2981
rect 11701 2972 11713 2975
rect 10928 2944 11713 2972
rect 10928 2932 10934 2944
rect 11701 2941 11713 2944
rect 11747 2941 11759 2975
rect 12268 2972 12296 3012
rect 12989 3009 13001 3043
rect 13035 3040 13047 3043
rect 13630 3040 13636 3052
rect 13035 3012 13636 3040
rect 13035 3009 13047 3012
rect 12989 3003 13047 3009
rect 13630 3000 13636 3012
rect 13688 3000 13694 3052
rect 13722 3000 13728 3052
rect 13780 3000 13786 3052
rect 14461 3043 14519 3049
rect 14461 3009 14473 3043
rect 14507 3040 14519 3043
rect 15010 3040 15016 3052
rect 14507 3012 15016 3040
rect 14507 3009 14519 3012
rect 14461 3003 14519 3009
rect 15010 3000 15016 3012
rect 15068 3000 15074 3052
rect 15197 3043 15255 3049
rect 15197 3009 15209 3043
rect 15243 3040 15255 3043
rect 15746 3040 15752 3052
rect 15243 3012 15752 3040
rect 15243 3009 15255 3012
rect 15197 3003 15255 3009
rect 15746 3000 15752 3012
rect 15804 3000 15810 3052
rect 15838 3000 15844 3052
rect 15896 3000 15902 3052
rect 17497 3043 17555 3049
rect 17497 3009 17509 3043
rect 17543 3040 17555 3043
rect 18230 3040 18236 3052
rect 17543 3012 18236 3040
rect 17543 3009 17555 3012
rect 17497 3003 17555 3009
rect 18230 3000 18236 3012
rect 18288 3000 18294 3052
rect 19352 3049 19380 3080
rect 22094 3068 22100 3080
rect 22152 3068 22158 3120
rect 18417 3043 18475 3049
rect 18417 3009 18429 3043
rect 18463 3040 18475 3043
rect 19337 3043 19395 3049
rect 18463 3012 19288 3040
rect 18463 3009 18475 3012
rect 18417 3003 18475 3009
rect 13078 2972 13084 2984
rect 12268 2944 13084 2972
rect 11701 2935 11759 2941
rect 13078 2932 13084 2944
rect 13136 2932 13142 2984
rect 13173 2975 13231 2981
rect 13173 2941 13185 2975
rect 13219 2972 13231 2975
rect 13906 2972 13912 2984
rect 13219 2944 13912 2972
rect 13219 2941 13231 2944
rect 13173 2935 13231 2941
rect 13906 2932 13912 2944
rect 13964 2932 13970 2984
rect 14645 2975 14703 2981
rect 14645 2941 14657 2975
rect 14691 2941 14703 2975
rect 14645 2935 14703 2941
rect 16117 2975 16175 2981
rect 16117 2941 16129 2975
rect 16163 2972 16175 2975
rect 16482 2972 16488 2984
rect 16163 2944 16488 2972
rect 16163 2941 16175 2944
rect 16117 2935 16175 2941
rect 8294 2864 8300 2916
rect 8352 2904 8358 2916
rect 9953 2907 10011 2913
rect 9953 2904 9965 2907
rect 8352 2876 9965 2904
rect 8352 2864 8358 2876
rect 9953 2873 9965 2876
rect 9999 2873 10011 2907
rect 9953 2867 10011 2873
rect 11882 2864 11888 2916
rect 11940 2904 11946 2916
rect 11977 2907 12035 2913
rect 11977 2904 11989 2907
rect 11940 2876 11989 2904
rect 11940 2864 11946 2876
rect 11977 2873 11989 2876
rect 12023 2873 12035 2907
rect 14660 2904 14688 2935
rect 16482 2932 16488 2944
rect 16540 2932 16546 2984
rect 17773 2975 17831 2981
rect 17773 2941 17785 2975
rect 17819 2972 17831 2975
rect 17862 2972 17868 2984
rect 17819 2944 17868 2972
rect 17819 2941 17831 2944
rect 17773 2935 17831 2941
rect 17862 2932 17868 2944
rect 17920 2932 17926 2984
rect 19260 2972 19288 3012
rect 19337 3009 19349 3043
rect 19383 3009 19395 3043
rect 19337 3003 19395 3009
rect 19613 3043 19671 3049
rect 19613 3009 19625 3043
rect 19659 3040 19671 3043
rect 21174 3040 21180 3052
rect 19659 3012 21180 3040
rect 19659 3009 19671 3012
rect 19613 3003 19671 3009
rect 21174 3000 21180 3012
rect 21232 3000 21238 3052
rect 21269 3043 21327 3049
rect 21269 3009 21281 3043
rect 21315 3040 21327 3043
rect 21450 3040 21456 3052
rect 21315 3012 21456 3040
rect 21315 3009 21327 3012
rect 21269 3003 21327 3009
rect 21450 3000 21456 3012
rect 21508 3000 21514 3052
rect 19426 2972 19432 2984
rect 19260 2944 19432 2972
rect 19426 2932 19432 2944
rect 19484 2932 19490 2984
rect 20257 2975 20315 2981
rect 20257 2941 20269 2975
rect 20303 2972 20315 2975
rect 20346 2972 20352 2984
rect 20303 2944 20352 2972
rect 20303 2941 20315 2944
rect 20257 2935 20315 2941
rect 20346 2932 20352 2944
rect 20404 2972 20410 2984
rect 22204 2972 22232 3148
rect 23750 3136 23756 3148
rect 23808 3136 23814 3188
rect 25682 3136 25688 3188
rect 25740 3176 25746 3188
rect 25777 3179 25835 3185
rect 25777 3176 25789 3179
rect 25740 3148 25789 3176
rect 25740 3136 25746 3148
rect 25777 3145 25789 3148
rect 25823 3145 25835 3179
rect 25777 3139 25835 3145
rect 25958 3136 25964 3188
rect 26016 3176 26022 3188
rect 26605 3179 26663 3185
rect 26605 3176 26617 3179
rect 26016 3148 26617 3176
rect 26016 3136 26022 3148
rect 26605 3145 26617 3148
rect 26651 3145 26663 3179
rect 26605 3139 26663 3145
rect 27154 3136 27160 3188
rect 27212 3176 27218 3188
rect 33594 3176 33600 3188
rect 27212 3148 33600 3176
rect 27212 3136 27218 3148
rect 33594 3136 33600 3148
rect 33652 3136 33658 3188
rect 38470 3136 38476 3188
rect 38528 3176 38534 3188
rect 41322 3176 41328 3188
rect 38528 3148 41328 3176
rect 38528 3136 38534 3148
rect 41322 3136 41328 3148
rect 41380 3136 41386 3188
rect 41690 3136 41696 3188
rect 41748 3176 41754 3188
rect 41785 3179 41843 3185
rect 41785 3176 41797 3179
rect 41748 3148 41797 3176
rect 41748 3136 41754 3148
rect 41785 3145 41797 3148
rect 41831 3145 41843 3179
rect 41785 3139 41843 3145
rect 43898 3136 43904 3188
rect 43956 3136 43962 3188
rect 44634 3136 44640 3188
rect 44692 3136 44698 3188
rect 46106 3176 46112 3188
rect 44836 3148 46112 3176
rect 22370 3068 22376 3120
rect 22428 3108 22434 3120
rect 23934 3108 23940 3120
rect 22428 3080 23940 3108
rect 22428 3068 22434 3080
rect 23934 3068 23940 3080
rect 23992 3068 23998 3120
rect 24664 3111 24722 3117
rect 24664 3077 24676 3111
rect 24710 3108 24722 3111
rect 25222 3108 25228 3120
rect 24710 3080 25228 3108
rect 24710 3077 24722 3080
rect 24664 3071 24722 3077
rect 25222 3068 25228 3080
rect 25280 3068 25286 3120
rect 25314 3068 25320 3120
rect 25372 3108 25378 3120
rect 27890 3108 27896 3120
rect 25372 3080 27896 3108
rect 25372 3068 25378 3080
rect 27890 3068 27896 3080
rect 27948 3068 27954 3120
rect 29822 3068 29828 3120
rect 29880 3108 29886 3120
rect 29880 3080 30880 3108
rect 29880 3068 29886 3080
rect 22281 3043 22339 3049
rect 22281 3009 22293 3043
rect 22327 3040 22339 3043
rect 22557 3043 22615 3049
rect 22557 3040 22569 3043
rect 22327 3012 22569 3040
rect 22327 3009 22339 3012
rect 22281 3003 22339 3009
rect 22557 3009 22569 3012
rect 22603 3040 22615 3043
rect 23382 3040 23388 3052
rect 22603 3012 23388 3040
rect 22603 3009 22615 3012
rect 22557 3003 22615 3009
rect 23382 3000 23388 3012
rect 23440 3000 23446 3052
rect 23477 3043 23535 3049
rect 23477 3009 23489 3043
rect 23523 3009 23535 3043
rect 23477 3003 23535 3009
rect 24397 3043 24455 3049
rect 24397 3009 24409 3043
rect 24443 3040 24455 3043
rect 24486 3040 24492 3052
rect 24443 3012 24492 3040
rect 24443 3009 24455 3012
rect 24397 3003 24455 3009
rect 20404 2944 21496 2972
rect 20404 2932 20410 2944
rect 17310 2904 17316 2916
rect 14660 2876 17316 2904
rect 11977 2867 12035 2873
rect 17310 2864 17316 2876
rect 17368 2864 17374 2916
rect 18138 2864 18144 2916
rect 18196 2904 18202 2916
rect 20533 2907 20591 2913
rect 20533 2904 20545 2907
rect 18196 2876 20545 2904
rect 18196 2864 18202 2876
rect 20533 2873 20545 2876
rect 20579 2873 20591 2907
rect 20533 2867 20591 2873
rect 20717 2907 20775 2913
rect 20717 2873 20729 2907
rect 20763 2904 20775 2907
rect 20990 2904 20996 2916
rect 20763 2876 20996 2904
rect 20763 2873 20775 2876
rect 20717 2867 20775 2873
rect 20990 2864 20996 2876
rect 21048 2864 21054 2916
rect 6917 2839 6975 2845
rect 6917 2805 6929 2839
rect 6963 2836 6975 2839
rect 15654 2836 15660 2848
rect 6963 2808 15660 2836
rect 6963 2805 6975 2808
rect 6917 2799 6975 2805
rect 15654 2796 15660 2808
rect 15712 2796 15718 2848
rect 17034 2796 17040 2848
rect 17092 2796 17098 2848
rect 20806 2796 20812 2848
rect 20864 2836 20870 2848
rect 21361 2839 21419 2845
rect 21361 2836 21373 2839
rect 20864 2808 21373 2836
rect 20864 2796 20870 2808
rect 21361 2805 21373 2808
rect 21407 2805 21419 2839
rect 21468 2836 21496 2944
rect 22066 2944 22232 2972
rect 21542 2864 21548 2916
rect 21600 2904 21606 2916
rect 22066 2904 22094 2944
rect 22830 2932 22836 2984
rect 22888 2932 22894 2984
rect 23492 2972 23520 3003
rect 24486 3000 24492 3012
rect 24544 3000 24550 3052
rect 26234 3040 26240 3052
rect 25424 3012 26240 3040
rect 23492 2944 23704 2972
rect 21600 2876 22094 2904
rect 23676 2904 23704 2944
rect 23750 2932 23756 2984
rect 23808 2932 23814 2984
rect 24210 2904 24216 2916
rect 23676 2876 24216 2904
rect 21600 2864 21606 2876
rect 24210 2864 24216 2876
rect 24268 2864 24274 2916
rect 22646 2836 22652 2848
rect 21468 2808 22652 2836
rect 21361 2799 21419 2805
rect 22646 2796 22652 2808
rect 22704 2796 22710 2848
rect 22738 2796 22744 2848
rect 22796 2836 22802 2848
rect 25424 2836 25452 3012
rect 26234 3000 26240 3012
rect 26292 3000 26298 3052
rect 26421 3043 26479 3049
rect 26421 3009 26433 3043
rect 26467 3009 26479 3043
rect 26421 3003 26479 3009
rect 27157 3043 27215 3049
rect 27157 3009 27169 3043
rect 27203 3040 27215 3043
rect 28629 3043 28687 3049
rect 27203 3012 28580 3040
rect 27203 3009 27215 3012
rect 27157 3003 27215 3009
rect 26436 2904 26464 3003
rect 26510 2932 26516 2984
rect 26568 2972 26574 2984
rect 27341 2975 27399 2981
rect 27341 2972 27353 2975
rect 26568 2944 27353 2972
rect 26568 2932 26574 2944
rect 27341 2941 27353 2944
rect 27387 2941 27399 2975
rect 28552 2972 28580 3012
rect 28629 3009 28641 3043
rect 28675 3040 28687 3043
rect 29362 3040 29368 3052
rect 28675 3012 29368 3040
rect 28675 3009 28687 3012
rect 28629 3003 28687 3009
rect 29362 3000 29368 3012
rect 29420 3000 29426 3052
rect 29730 3000 29736 3052
rect 29788 3040 29794 3052
rect 30852 3049 30880 3080
rect 32674 3068 32680 3120
rect 32732 3108 32738 3120
rect 34425 3111 34483 3117
rect 34425 3108 34437 3111
rect 32732 3080 34437 3108
rect 32732 3068 32738 3080
rect 34425 3077 34437 3080
rect 34471 3077 34483 3111
rect 34425 3071 34483 3077
rect 38565 3111 38623 3117
rect 38565 3077 38577 3111
rect 38611 3108 38623 3111
rect 39114 3108 39120 3120
rect 38611 3080 39120 3108
rect 38611 3077 38623 3080
rect 38565 3071 38623 3077
rect 39114 3068 39120 3080
rect 39172 3068 39178 3120
rect 40681 3111 40739 3117
rect 40681 3108 40693 3111
rect 39500 3080 40693 3108
rect 29917 3043 29975 3049
rect 29917 3040 29929 3043
rect 29788 3012 29929 3040
rect 29788 3000 29794 3012
rect 29917 3009 29929 3012
rect 29963 3009 29975 3043
rect 29917 3003 29975 3009
rect 30837 3043 30895 3049
rect 30837 3009 30849 3043
rect 30883 3009 30895 3043
rect 30837 3003 30895 3009
rect 31846 3000 31852 3052
rect 31904 3040 31910 3052
rect 32309 3043 32367 3049
rect 32309 3040 32321 3043
rect 31904 3012 32321 3040
rect 31904 3000 31910 3012
rect 32309 3009 32321 3012
rect 32355 3009 32367 3043
rect 32309 3003 32367 3009
rect 33042 3000 33048 3052
rect 33100 3040 33106 3052
rect 33229 3043 33287 3049
rect 33229 3040 33241 3043
rect 33100 3012 33241 3040
rect 33100 3000 33106 3012
rect 33229 3009 33241 3012
rect 33275 3009 33287 3043
rect 33229 3003 33287 3009
rect 34146 3000 34152 3052
rect 34204 3000 34210 3052
rect 34238 3000 34244 3052
rect 34296 3040 34302 3052
rect 35069 3043 35127 3049
rect 35069 3040 35081 3043
rect 34296 3012 35081 3040
rect 34296 3000 34302 3012
rect 35069 3009 35081 3012
rect 35115 3009 35127 3043
rect 35069 3003 35127 3009
rect 35986 3000 35992 3052
rect 36044 3000 36050 3052
rect 37461 3043 37519 3049
rect 37461 3009 37473 3043
rect 37507 3040 37519 3043
rect 38286 3040 38292 3052
rect 37507 3012 38292 3040
rect 37507 3009 37519 3012
rect 37461 3003 37519 3009
rect 38286 3000 38292 3012
rect 38344 3000 38350 3052
rect 38378 3000 38384 3052
rect 38436 3000 38442 3052
rect 38654 3000 38660 3052
rect 38712 3000 38718 3052
rect 38801 3043 38859 3049
rect 38801 3009 38813 3043
rect 38847 3040 38859 3043
rect 39390 3040 39396 3052
rect 38847 3012 39396 3040
rect 38847 3009 38859 3012
rect 38801 3003 38859 3009
rect 39390 3000 39396 3012
rect 39448 3000 39454 3052
rect 39500 3049 39528 3080
rect 40681 3077 40693 3080
rect 40727 3077 40739 3111
rect 40681 3071 40739 3077
rect 42794 3068 42800 3120
rect 42852 3068 42858 3120
rect 42889 3111 42947 3117
rect 42889 3077 42901 3111
rect 42935 3108 42947 3111
rect 44836 3108 44864 3148
rect 46106 3136 46112 3148
rect 46164 3136 46170 3188
rect 46290 3136 46296 3188
rect 46348 3176 46354 3188
rect 46845 3179 46903 3185
rect 46845 3176 46857 3179
rect 46348 3148 46857 3176
rect 46348 3136 46354 3148
rect 46845 3145 46857 3148
rect 46891 3145 46903 3179
rect 48406 3176 48412 3188
rect 46845 3139 46903 3145
rect 46952 3148 48412 3176
rect 42935 3080 44864 3108
rect 42935 3077 42947 3080
rect 42889 3071 42947 3077
rect 44910 3068 44916 3120
rect 44968 3108 44974 3120
rect 46017 3111 46075 3117
rect 46017 3108 46029 3111
rect 44968 3080 46029 3108
rect 44968 3068 44974 3080
rect 46017 3077 46029 3080
rect 46063 3077 46075 3111
rect 46017 3071 46075 3077
rect 46201 3111 46259 3117
rect 46201 3077 46213 3111
rect 46247 3108 46259 3111
rect 46382 3108 46388 3120
rect 46247 3080 46388 3108
rect 46247 3077 46259 3080
rect 46201 3071 46259 3077
rect 46382 3068 46388 3080
rect 46440 3068 46446 3120
rect 39485 3043 39543 3049
rect 39485 3009 39497 3043
rect 39531 3009 39543 3043
rect 39485 3003 39543 3009
rect 40497 3043 40555 3049
rect 40497 3009 40509 3043
rect 40543 3040 40555 3043
rect 40862 3040 40868 3052
rect 40543 3012 40868 3040
rect 40543 3009 40555 3012
rect 40497 3003 40555 3009
rect 40862 3000 40868 3012
rect 40920 3000 40926 3052
rect 41506 3000 41512 3052
rect 41564 3040 41570 3052
rect 41693 3043 41751 3049
rect 41693 3040 41705 3043
rect 41564 3012 41705 3040
rect 41564 3000 41570 3012
rect 41693 3009 41705 3012
rect 41739 3009 41751 3043
rect 41693 3003 41751 3009
rect 42613 3043 42671 3049
rect 42613 3009 42625 3043
rect 42659 3040 42671 3043
rect 42702 3040 42708 3052
rect 42659 3012 42708 3040
rect 42659 3009 42671 3012
rect 42613 3003 42671 3009
rect 42702 3000 42708 3012
rect 42760 3000 42766 3052
rect 43033 3043 43091 3049
rect 43033 3009 43045 3043
rect 43079 3040 43091 3043
rect 43079 3012 43199 3040
rect 43079 3009 43091 3012
rect 43033 3003 43091 3009
rect 29086 2972 29092 2984
rect 28552 2944 29092 2972
rect 27341 2935 27399 2941
rect 29086 2932 29092 2944
rect 29144 2932 29150 2984
rect 29273 2975 29331 2981
rect 29273 2941 29285 2975
rect 29319 2972 29331 2975
rect 29638 2972 29644 2984
rect 29319 2944 29644 2972
rect 29319 2941 29331 2944
rect 29273 2935 29331 2941
rect 29638 2932 29644 2944
rect 29696 2932 29702 2984
rect 30190 2932 30196 2984
rect 30248 2932 30254 2984
rect 30742 2932 30748 2984
rect 30800 2972 30806 2984
rect 31021 2975 31079 2981
rect 31021 2972 31033 2975
rect 30800 2944 31033 2972
rect 30800 2932 30806 2944
rect 31021 2941 31033 2944
rect 31067 2941 31079 2975
rect 31021 2935 31079 2941
rect 31570 2932 31576 2984
rect 31628 2972 31634 2984
rect 32493 2975 32551 2981
rect 32493 2972 32505 2975
rect 31628 2944 32505 2972
rect 31628 2932 31634 2944
rect 32493 2941 32505 2944
rect 32539 2941 32551 2975
rect 32493 2935 32551 2941
rect 33413 2975 33471 2981
rect 33413 2941 33425 2975
rect 33459 2941 33471 2975
rect 33413 2935 33471 2941
rect 35253 2975 35311 2981
rect 35253 2941 35265 2975
rect 35299 2941 35311 2975
rect 35253 2935 35311 2941
rect 31478 2904 31484 2916
rect 26436 2876 31484 2904
rect 31478 2864 31484 2876
rect 31536 2864 31542 2916
rect 32122 2864 32128 2916
rect 32180 2904 32186 2916
rect 33428 2904 33456 2935
rect 32180 2876 33456 2904
rect 32180 2864 32186 2876
rect 33502 2864 33508 2916
rect 33560 2904 33566 2916
rect 35268 2904 35296 2935
rect 36170 2932 36176 2984
rect 36228 2932 36234 2984
rect 37274 2932 37280 2984
rect 37332 2972 37338 2984
rect 37645 2975 37703 2981
rect 37645 2972 37657 2975
rect 37332 2944 37657 2972
rect 37332 2932 37338 2944
rect 37645 2941 37657 2944
rect 37691 2941 37703 2975
rect 37645 2935 37703 2941
rect 39666 2932 39672 2984
rect 39724 2932 39730 2984
rect 43171 2972 43199 3012
rect 43254 3000 43260 3052
rect 43312 3040 43318 3052
rect 43809 3043 43867 3049
rect 43809 3040 43821 3043
rect 43312 3012 43821 3040
rect 43312 3000 43318 3012
rect 43809 3009 43821 3012
rect 43855 3009 43867 3043
rect 43809 3003 43867 3009
rect 44082 3000 44088 3052
rect 44140 3040 44146 3052
rect 44453 3043 44511 3049
rect 44453 3040 44465 3043
rect 44140 3012 44465 3040
rect 44140 3000 44146 3012
rect 44453 3009 44465 3012
rect 44499 3009 44511 3043
rect 44453 3003 44511 3009
rect 45278 3000 45284 3052
rect 45336 3000 45342 3052
rect 45370 3000 45376 3052
rect 45428 3040 45434 3052
rect 45465 3043 45523 3049
rect 45465 3040 45477 3043
rect 45428 3012 45477 3040
rect 45428 3000 45434 3012
rect 45465 3009 45477 3012
rect 45511 3009 45523 3043
rect 45465 3003 45523 3009
rect 46290 3000 46296 3052
rect 46348 3040 46354 3052
rect 46753 3043 46811 3049
rect 46753 3040 46765 3043
rect 46348 3012 46765 3040
rect 46348 3000 46354 3012
rect 46753 3009 46765 3012
rect 46799 3009 46811 3043
rect 46753 3003 46811 3009
rect 44174 2972 44180 2984
rect 43171 2944 44180 2972
rect 44174 2932 44180 2944
rect 44232 2972 44238 2984
rect 46952 2972 46980 3148
rect 48406 3136 48412 3148
rect 48464 3136 48470 3188
rect 48498 3136 48504 3188
rect 48556 3136 48562 3188
rect 48590 3136 48596 3188
rect 48648 3176 48654 3188
rect 48648 3148 52776 3176
rect 48648 3136 48654 3148
rect 47302 3068 47308 3120
rect 47360 3108 47366 3120
rect 50249 3111 50307 3117
rect 50249 3108 50261 3111
rect 47360 3080 50261 3108
rect 47360 3068 47366 3080
rect 50249 3077 50261 3080
rect 50295 3077 50307 3111
rect 52748 3108 52776 3148
rect 52822 3136 52828 3188
rect 52880 3176 52886 3188
rect 53101 3179 53159 3185
rect 53101 3176 53113 3179
rect 52880 3148 53113 3176
rect 52880 3136 52886 3148
rect 53101 3145 53113 3148
rect 53147 3145 53159 3179
rect 53101 3139 53159 3145
rect 54570 3136 54576 3188
rect 54628 3136 54634 3188
rect 55306 3136 55312 3188
rect 55364 3136 55370 3188
rect 56962 3136 56968 3188
rect 57020 3136 57026 3188
rect 58342 3108 58348 3120
rect 52748 3080 58348 3108
rect 50249 3071 50307 3077
rect 58342 3068 58348 3080
rect 58400 3068 58406 3120
rect 47854 3000 47860 3052
rect 47912 3000 47918 3052
rect 48038 3049 48044 3052
rect 48005 3043 48044 3049
rect 48005 3009 48017 3043
rect 48005 3003 48044 3009
rect 48038 3000 48044 3003
rect 48096 3000 48102 3052
rect 48133 3043 48191 3049
rect 48133 3009 48145 3043
rect 48179 3009 48191 3043
rect 48133 3003 48191 3009
rect 44232 2944 46980 2972
rect 44232 2932 44238 2944
rect 47210 2932 47216 2984
rect 47268 2972 47274 2984
rect 47762 2972 47768 2984
rect 47268 2944 47768 2972
rect 47268 2932 47274 2944
rect 47762 2932 47768 2944
rect 47820 2972 47826 2984
rect 48148 2972 48176 3003
rect 48222 3000 48228 3052
rect 48280 3000 48286 3052
rect 48406 3049 48412 3052
rect 48363 3043 48412 3049
rect 48363 3009 48375 3043
rect 48409 3009 48412 3043
rect 48363 3003 48412 3009
rect 48406 3000 48412 3003
rect 48464 3000 48470 3052
rect 48498 3000 48504 3052
rect 48556 3040 48562 3052
rect 49145 3043 49203 3049
rect 49145 3040 49157 3043
rect 48556 3012 49157 3040
rect 48556 3000 48562 3012
rect 49145 3009 49157 3012
rect 49191 3009 49203 3043
rect 49145 3003 49203 3009
rect 49418 3000 49424 3052
rect 49476 3040 49482 3052
rect 50065 3043 50123 3049
rect 50065 3040 50077 3043
rect 49476 3012 50077 3040
rect 49476 3000 49482 3012
rect 50065 3009 50077 3012
rect 50111 3009 50123 3043
rect 50065 3003 50123 3009
rect 50798 3000 50804 3052
rect 50856 3000 50862 3052
rect 51534 3000 51540 3052
rect 51592 3000 51598 3052
rect 52638 3000 52644 3052
rect 52696 3040 52702 3052
rect 52917 3043 52975 3049
rect 52917 3040 52929 3043
rect 52696 3012 52929 3040
rect 52696 3000 52702 3012
rect 52917 3009 52929 3012
rect 52963 3009 52975 3043
rect 52917 3003 52975 3009
rect 53006 3000 53012 3052
rect 53064 3040 53070 3052
rect 53745 3043 53803 3049
rect 53745 3040 53757 3043
rect 53064 3012 53757 3040
rect 53064 3000 53070 3012
rect 53745 3009 53757 3012
rect 53791 3009 53803 3043
rect 53745 3003 53803 3009
rect 54386 3000 54392 3052
rect 54444 3000 54450 3052
rect 55214 3000 55220 3052
rect 55272 3000 55278 3052
rect 55950 3000 55956 3052
rect 56008 3000 56014 3052
rect 56134 3000 56140 3052
rect 56192 3040 56198 3052
rect 56597 3043 56655 3049
rect 56597 3040 56609 3043
rect 56192 3012 56609 3040
rect 56192 3000 56198 3012
rect 56597 3009 56609 3012
rect 56643 3009 56655 3043
rect 56597 3003 56655 3009
rect 56778 3000 56784 3052
rect 56836 3000 56842 3052
rect 56962 3000 56968 3052
rect 57020 3040 57026 3052
rect 58161 3043 58219 3049
rect 58161 3040 58173 3043
rect 57020 3012 58173 3040
rect 57020 3000 57026 3012
rect 58161 3009 58173 3012
rect 58207 3009 58219 3043
rect 58161 3003 58219 3009
rect 48774 2972 48780 2984
rect 47820 2944 48780 2972
rect 47820 2932 47826 2944
rect 48774 2932 48780 2944
rect 48832 2932 48838 2984
rect 49050 2932 49056 2984
rect 49108 2972 49114 2984
rect 51721 2975 51779 2981
rect 51721 2972 51733 2975
rect 49108 2944 51733 2972
rect 49108 2932 49114 2944
rect 51721 2941 51733 2944
rect 51767 2941 51779 2975
rect 51721 2935 51779 2941
rect 33560 2876 35296 2904
rect 33560 2864 33566 2876
rect 38838 2864 38844 2916
rect 38896 2904 38902 2916
rect 38933 2907 38991 2913
rect 38933 2904 38945 2907
rect 38896 2876 38945 2904
rect 38896 2864 38902 2876
rect 38933 2873 38945 2876
rect 38979 2873 38991 2907
rect 38933 2867 38991 2873
rect 40586 2864 40592 2916
rect 40644 2904 40650 2916
rect 43165 2907 43223 2913
rect 43165 2904 43177 2907
rect 40644 2876 43177 2904
rect 40644 2864 40650 2876
rect 43165 2873 43177 2876
rect 43211 2873 43223 2907
rect 43165 2867 43223 2873
rect 43714 2864 43720 2916
rect 43772 2904 43778 2916
rect 53929 2907 53987 2913
rect 53929 2904 53941 2907
rect 43772 2876 53941 2904
rect 43772 2864 43778 2876
rect 53929 2873 53941 2876
rect 53975 2873 53987 2907
rect 58345 2907 58403 2913
rect 58345 2904 58357 2907
rect 53929 2867 53987 2873
rect 54036 2876 58357 2904
rect 22796 2808 25452 2836
rect 22796 2796 22802 2808
rect 25958 2796 25964 2848
rect 26016 2836 26022 2848
rect 28718 2836 28724 2848
rect 26016 2808 28724 2836
rect 26016 2796 26022 2808
rect 28718 2796 28724 2808
rect 28776 2796 28782 2848
rect 42886 2796 42892 2848
rect 42944 2836 42950 2848
rect 45278 2836 45284 2848
rect 42944 2808 45284 2836
rect 42944 2796 42950 2808
rect 45278 2796 45284 2808
rect 45336 2796 45342 2848
rect 49234 2796 49240 2848
rect 49292 2796 49298 2848
rect 49878 2796 49884 2848
rect 49936 2836 49942 2848
rect 50893 2839 50951 2845
rect 50893 2836 50905 2839
rect 49936 2808 50905 2836
rect 49936 2796 49942 2808
rect 50893 2805 50905 2808
rect 50939 2805 50951 2839
rect 50893 2799 50951 2805
rect 52454 2796 52460 2848
rect 52512 2836 52518 2848
rect 54036 2836 54064 2876
rect 58345 2873 58357 2876
rect 58391 2873 58403 2907
rect 58345 2867 58403 2873
rect 52512 2808 54064 2836
rect 52512 2796 52518 2808
rect 56042 2796 56048 2848
rect 56100 2796 56106 2848
rect 1104 2746 58880 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 58880 2746
rect 1104 2672 58880 2694
rect 7745 2635 7803 2641
rect 7745 2601 7757 2635
rect 7791 2632 7803 2635
rect 8386 2632 8392 2644
rect 7791 2604 8392 2632
rect 7791 2601 7803 2604
rect 7745 2595 7803 2601
rect 8386 2592 8392 2604
rect 8444 2592 8450 2644
rect 10321 2635 10379 2641
rect 10321 2601 10333 2635
rect 10367 2632 10379 2635
rect 12161 2635 12219 2641
rect 10367 2604 11376 2632
rect 10367 2601 10379 2604
rect 10321 2595 10379 2601
rect 7101 2567 7159 2573
rect 7101 2533 7113 2567
rect 7147 2564 7159 2567
rect 8294 2564 8300 2576
rect 7147 2536 8300 2564
rect 7147 2533 7159 2536
rect 7101 2527 7159 2533
rect 8294 2524 8300 2536
rect 8352 2524 8358 2576
rect 8573 2567 8631 2573
rect 8573 2533 8585 2567
rect 8619 2564 8631 2567
rect 8754 2564 8760 2576
rect 8619 2536 8760 2564
rect 8619 2533 8631 2536
rect 8573 2527 8631 2533
rect 8754 2524 8760 2536
rect 8812 2524 8818 2576
rect 9677 2567 9735 2573
rect 9677 2533 9689 2567
rect 9723 2564 9735 2567
rect 10594 2564 10600 2576
rect 9723 2536 10600 2564
rect 9723 2533 9735 2536
rect 9677 2527 9735 2533
rect 10594 2524 10600 2536
rect 10652 2524 10658 2576
rect 11348 2564 11376 2604
rect 12161 2601 12173 2635
rect 12207 2632 12219 2635
rect 13170 2632 13176 2644
rect 12207 2604 13176 2632
rect 12207 2601 12219 2604
rect 12161 2595 12219 2601
rect 13170 2592 13176 2604
rect 13228 2592 13234 2644
rect 13262 2592 13268 2644
rect 13320 2632 13326 2644
rect 13633 2635 13691 2641
rect 13633 2632 13645 2635
rect 13320 2604 13645 2632
rect 13320 2592 13326 2604
rect 13633 2601 13645 2604
rect 13679 2601 13691 2635
rect 13633 2595 13691 2601
rect 17880 2604 18460 2632
rect 12526 2564 12532 2576
rect 11348 2536 12532 2564
rect 12526 2524 12532 2536
rect 12584 2524 12590 2576
rect 12989 2567 13047 2573
rect 12989 2533 13001 2567
rect 13035 2564 13047 2567
rect 13446 2564 13452 2576
rect 13035 2536 13452 2564
rect 13035 2533 13047 2536
rect 12989 2527 13047 2533
rect 13446 2524 13452 2536
rect 13504 2524 13510 2576
rect 14461 2567 14519 2573
rect 14461 2533 14473 2567
rect 14507 2564 14519 2567
rect 17770 2564 17776 2576
rect 14507 2536 17776 2564
rect 14507 2533 14519 2536
rect 14461 2527 14519 2533
rect 17770 2524 17776 2536
rect 17828 2524 17834 2576
rect 5997 2499 6055 2505
rect 5997 2465 6009 2499
rect 6043 2496 6055 2499
rect 15197 2499 15255 2505
rect 6043 2468 13676 2496
rect 6043 2465 6055 2468
rect 5997 2459 6055 2465
rect 7653 2431 7711 2437
rect 7653 2397 7665 2431
rect 7699 2428 7711 2431
rect 9493 2431 9551 2437
rect 7699 2400 9444 2428
rect 7699 2397 7711 2400
rect 7653 2391 7711 2397
rect 5810 2320 5816 2372
rect 5868 2320 5874 2372
rect 6917 2363 6975 2369
rect 6917 2329 6929 2363
rect 6963 2360 6975 2363
rect 8018 2360 8024 2372
rect 6963 2332 8024 2360
rect 6963 2329 6975 2332
rect 6917 2323 6975 2329
rect 8018 2320 8024 2332
rect 8076 2320 8082 2372
rect 8386 2320 8392 2372
rect 8444 2320 8450 2372
rect 9416 2360 9444 2400
rect 9493 2397 9505 2431
rect 9539 2428 9551 2431
rect 10965 2431 11023 2437
rect 9539 2400 10916 2428
rect 9539 2397 9551 2400
rect 9493 2391 9551 2397
rect 10042 2360 10048 2372
rect 9416 2332 10048 2360
rect 10042 2320 10048 2332
rect 10100 2320 10106 2372
rect 10226 2320 10232 2372
rect 10284 2320 10290 2372
rect 10888 2360 10916 2400
rect 10965 2397 10977 2431
rect 11011 2428 11023 2431
rect 12526 2428 12532 2440
rect 11011 2400 12532 2428
rect 11011 2397 11023 2400
rect 10965 2391 11023 2397
rect 12526 2388 12532 2400
rect 12584 2388 12590 2440
rect 11698 2360 11704 2372
rect 10888 2332 11704 2360
rect 11698 2320 11704 2332
rect 11756 2320 11762 2372
rect 12066 2320 12072 2372
rect 12124 2320 12130 2372
rect 12805 2363 12863 2369
rect 12805 2329 12817 2363
rect 12851 2360 12863 2363
rect 13262 2360 13268 2372
rect 12851 2332 13268 2360
rect 12851 2329 12863 2332
rect 12805 2323 12863 2329
rect 13262 2320 13268 2332
rect 13320 2320 13326 2372
rect 13538 2320 13544 2372
rect 13596 2320 13602 2372
rect 13648 2360 13676 2468
rect 15197 2465 15209 2499
rect 15243 2496 15255 2499
rect 16390 2496 16396 2508
rect 15243 2468 16396 2496
rect 15243 2465 15255 2468
rect 15197 2459 15255 2465
rect 16390 2456 16396 2468
rect 16448 2456 16454 2508
rect 17880 2496 17908 2604
rect 17512 2468 17908 2496
rect 18432 2496 18460 2604
rect 19426 2592 19432 2644
rect 19484 2632 19490 2644
rect 22097 2635 22155 2641
rect 22097 2632 22109 2635
rect 19484 2604 22109 2632
rect 19484 2592 19490 2604
rect 22097 2601 22109 2604
rect 22143 2601 22155 2635
rect 22097 2595 22155 2601
rect 24581 2635 24639 2641
rect 24581 2601 24593 2635
rect 24627 2632 24639 2635
rect 27522 2632 27528 2644
rect 24627 2604 27528 2632
rect 24627 2601 24639 2604
rect 24581 2595 24639 2601
rect 27522 2592 27528 2604
rect 27580 2592 27586 2644
rect 39758 2632 39764 2644
rect 31726 2604 39764 2632
rect 31726 2564 31754 2604
rect 39758 2592 39764 2604
rect 39816 2592 39822 2644
rect 41414 2592 41420 2644
rect 41472 2592 41478 2644
rect 42981 2635 43039 2641
rect 42981 2601 42993 2635
rect 43027 2632 43039 2635
rect 43806 2632 43812 2644
rect 43027 2604 43812 2632
rect 43027 2601 43039 2604
rect 42981 2595 43039 2601
rect 43806 2592 43812 2604
rect 43864 2592 43870 2644
rect 44450 2592 44456 2644
rect 44508 2592 44514 2644
rect 45373 2635 45431 2641
rect 45373 2601 45385 2635
rect 45419 2632 45431 2635
rect 45419 2604 46060 2632
rect 45419 2601 45431 2604
rect 45373 2595 45431 2601
rect 21008 2536 31754 2564
rect 20806 2496 20812 2508
rect 18432 2468 20812 2496
rect 14918 2388 14924 2440
rect 14976 2388 14982 2440
rect 15838 2388 15844 2440
rect 15896 2388 15902 2440
rect 17037 2431 17095 2437
rect 15948 2400 16574 2428
rect 15948 2360 15976 2400
rect 13648 2332 15976 2360
rect 16117 2363 16175 2369
rect 16117 2329 16129 2363
rect 16163 2329 16175 2363
rect 16546 2360 16574 2400
rect 17037 2397 17049 2431
rect 17083 2428 17095 2431
rect 17402 2428 17408 2440
rect 17083 2400 17408 2428
rect 17083 2397 17095 2400
rect 17037 2391 17095 2397
rect 17402 2388 17408 2400
rect 17460 2388 17466 2440
rect 17512 2437 17540 2468
rect 20806 2456 20812 2468
rect 20864 2456 20870 2508
rect 17497 2431 17555 2437
rect 17497 2397 17509 2431
rect 17543 2397 17555 2431
rect 17497 2391 17555 2397
rect 17773 2431 17831 2437
rect 17773 2397 17785 2431
rect 17819 2428 17831 2431
rect 18230 2428 18236 2440
rect 17819 2400 18236 2428
rect 17819 2397 17831 2400
rect 17773 2391 17831 2397
rect 18230 2388 18236 2400
rect 18288 2388 18294 2440
rect 18414 2388 18420 2440
rect 18472 2388 18478 2440
rect 19334 2388 19340 2440
rect 19392 2428 19398 2440
rect 19613 2431 19671 2437
rect 19613 2428 19625 2431
rect 19392 2400 19625 2428
rect 19392 2388 19398 2400
rect 19613 2397 19625 2400
rect 19659 2397 19671 2431
rect 19613 2391 19671 2397
rect 20070 2388 20076 2440
rect 20128 2388 20134 2440
rect 21008 2437 21036 2536
rect 39206 2524 39212 2576
rect 39264 2564 39270 2576
rect 46032 2564 46060 2604
rect 46106 2592 46112 2644
rect 46164 2592 46170 2644
rect 47118 2632 47124 2644
rect 46216 2604 47124 2632
rect 46216 2564 46244 2604
rect 47118 2592 47124 2604
rect 47176 2592 47182 2644
rect 48593 2635 48651 2641
rect 48593 2601 48605 2635
rect 48639 2632 48651 2635
rect 49142 2632 49148 2644
rect 48639 2604 49148 2632
rect 48639 2601 48651 2604
rect 48593 2595 48651 2601
rect 49142 2592 49148 2604
rect 49200 2592 49206 2644
rect 49326 2592 49332 2644
rect 49384 2592 49390 2644
rect 49694 2592 49700 2644
rect 49752 2632 49758 2644
rect 50525 2635 50583 2641
rect 50525 2632 50537 2635
rect 49752 2604 50537 2632
rect 49752 2592 49758 2604
rect 50525 2601 50537 2604
rect 50571 2601 50583 2635
rect 50525 2595 50583 2601
rect 51626 2592 51632 2644
rect 51684 2592 51690 2644
rect 52730 2592 52736 2644
rect 52788 2632 52794 2644
rect 53101 2635 53159 2641
rect 53101 2632 53113 2635
rect 52788 2604 53113 2632
rect 52788 2592 52794 2604
rect 53101 2601 53113 2604
rect 53147 2601 53159 2635
rect 53101 2595 53159 2601
rect 39264 2536 44956 2564
rect 46032 2536 46244 2564
rect 46937 2567 46995 2573
rect 39264 2524 39270 2536
rect 21269 2499 21327 2505
rect 21269 2465 21281 2499
rect 21315 2496 21327 2499
rect 24118 2496 24124 2508
rect 21315 2468 24124 2496
rect 21315 2465 21327 2468
rect 21269 2459 21327 2465
rect 24118 2456 24124 2468
rect 24176 2456 24182 2508
rect 44818 2496 44824 2508
rect 26160 2468 44824 2496
rect 20993 2431 21051 2437
rect 20993 2397 21005 2431
rect 21039 2397 21051 2431
rect 20993 2391 21051 2397
rect 21818 2388 21824 2440
rect 21876 2428 21882 2440
rect 22005 2431 22063 2437
rect 22005 2428 22017 2431
rect 21876 2400 22017 2428
rect 21876 2388 21882 2400
rect 22005 2397 22017 2400
rect 22051 2397 22063 2431
rect 22005 2391 22063 2397
rect 22646 2388 22652 2440
rect 22704 2388 22710 2440
rect 23290 2428 23296 2440
rect 22848 2400 23296 2428
rect 18598 2360 18604 2372
rect 16546 2332 18604 2360
rect 16117 2323 16175 2329
rect 11057 2295 11115 2301
rect 11057 2261 11069 2295
rect 11103 2292 11115 2295
rect 15930 2292 15936 2304
rect 11103 2264 15936 2292
rect 11103 2261 11115 2264
rect 11057 2255 11115 2261
rect 15930 2252 15936 2264
rect 15988 2252 15994 2304
rect 16132 2292 16160 2323
rect 18598 2320 18604 2332
rect 18656 2320 18662 2372
rect 18693 2363 18751 2369
rect 18693 2329 18705 2363
rect 18739 2360 18751 2363
rect 20349 2363 20407 2369
rect 18739 2332 20300 2360
rect 18739 2329 18751 2332
rect 18693 2323 18751 2329
rect 19426 2292 19432 2304
rect 16132 2264 19432 2292
rect 19426 2252 19432 2264
rect 19484 2252 19490 2304
rect 20272 2292 20300 2332
rect 20349 2329 20361 2363
rect 20395 2360 20407 2363
rect 22848 2360 22876 2400
rect 23290 2388 23296 2400
rect 23348 2388 23354 2440
rect 23566 2388 23572 2440
rect 23624 2388 23630 2440
rect 24949 2431 25007 2437
rect 24949 2397 24961 2431
rect 24995 2428 25007 2431
rect 25222 2428 25228 2440
rect 24995 2400 25228 2428
rect 24995 2397 25007 2400
rect 24949 2391 25007 2397
rect 25222 2388 25228 2400
rect 25280 2388 25286 2440
rect 26160 2437 26188 2468
rect 44818 2456 44824 2468
rect 44876 2456 44882 2508
rect 44928 2496 44956 2536
rect 46937 2533 46949 2567
rect 46983 2564 46995 2567
rect 47026 2564 47032 2576
rect 46983 2536 47032 2564
rect 46983 2533 46995 2536
rect 46937 2527 46995 2533
rect 47026 2524 47032 2536
rect 47084 2524 47090 2576
rect 48038 2524 48044 2576
rect 48096 2564 48102 2576
rect 55769 2567 55827 2573
rect 55769 2564 55781 2567
rect 48096 2536 55781 2564
rect 48096 2524 48102 2536
rect 55769 2533 55781 2536
rect 55815 2533 55827 2567
rect 55769 2527 55827 2533
rect 56505 2567 56563 2573
rect 56505 2533 56517 2567
rect 56551 2564 56563 2567
rect 56870 2564 56876 2576
rect 56551 2536 56876 2564
rect 56551 2533 56563 2536
rect 56505 2527 56563 2533
rect 56870 2524 56876 2536
rect 56928 2524 56934 2576
rect 58250 2564 58256 2576
rect 57072 2536 58256 2564
rect 48866 2496 48872 2508
rect 44928 2468 48872 2496
rect 48866 2456 48872 2468
rect 48924 2456 48930 2508
rect 54294 2456 54300 2508
rect 54352 2456 54358 2508
rect 26145 2431 26203 2437
rect 26145 2397 26157 2431
rect 26191 2397 26203 2431
rect 26145 2391 26203 2397
rect 26970 2388 26976 2440
rect 27028 2428 27034 2440
rect 27157 2431 27215 2437
rect 27157 2428 27169 2431
rect 27028 2400 27169 2428
rect 27028 2388 27034 2400
rect 27157 2397 27169 2400
rect 27203 2397 27215 2431
rect 27157 2391 27215 2397
rect 28718 2388 28724 2440
rect 28776 2388 28782 2440
rect 30193 2431 30251 2437
rect 30193 2397 30205 2431
rect 30239 2428 30251 2431
rect 30282 2428 30288 2440
rect 30239 2400 30288 2428
rect 30239 2397 30251 2400
rect 30193 2391 30251 2397
rect 30282 2388 30288 2400
rect 30340 2388 30346 2440
rect 30834 2388 30840 2440
rect 30892 2428 30898 2440
rect 31113 2431 31171 2437
rect 31113 2428 31125 2431
rect 30892 2400 31125 2428
rect 30892 2388 30898 2400
rect 31113 2397 31125 2400
rect 31159 2397 31171 2431
rect 31113 2391 31171 2397
rect 31938 2388 31944 2440
rect 31996 2428 32002 2440
rect 32309 2431 32367 2437
rect 32309 2428 32321 2431
rect 31996 2400 32321 2428
rect 31996 2388 32002 2400
rect 32309 2397 32321 2400
rect 32355 2397 32367 2431
rect 33229 2431 33287 2437
rect 33229 2428 33241 2431
rect 32309 2391 32367 2397
rect 32416 2400 33241 2428
rect 20395 2332 22876 2360
rect 22925 2363 22983 2369
rect 20395 2329 20407 2332
rect 20349 2323 20407 2329
rect 22925 2329 22937 2363
rect 22971 2329 22983 2363
rect 22925 2323 22983 2329
rect 23845 2363 23903 2369
rect 23845 2329 23857 2363
rect 23891 2360 23903 2363
rect 24762 2360 24768 2372
rect 23891 2332 24768 2360
rect 23891 2329 23903 2332
rect 23845 2323 23903 2329
rect 22462 2292 22468 2304
rect 20272 2264 22468 2292
rect 22462 2252 22468 2264
rect 22520 2252 22526 2304
rect 22940 2292 22968 2323
rect 24762 2320 24768 2332
rect 24820 2320 24826 2372
rect 25501 2363 25559 2369
rect 25501 2329 25513 2363
rect 25547 2360 25559 2363
rect 26050 2360 26056 2372
rect 25547 2332 26056 2360
rect 25547 2329 25559 2332
rect 25501 2323 25559 2329
rect 26050 2320 26056 2332
rect 26108 2320 26114 2372
rect 26421 2363 26479 2369
rect 26421 2329 26433 2363
rect 26467 2360 26479 2363
rect 26602 2360 26608 2372
rect 26467 2332 26608 2360
rect 26467 2329 26479 2332
rect 26421 2323 26479 2329
rect 26602 2320 26608 2332
rect 26660 2320 26666 2372
rect 26878 2320 26884 2372
rect 26936 2360 26942 2372
rect 27433 2363 27491 2369
rect 27433 2360 27445 2363
rect 26936 2332 27445 2360
rect 26936 2320 26942 2332
rect 27433 2329 27445 2332
rect 27479 2329 27491 2363
rect 27433 2323 27491 2329
rect 28997 2363 29055 2369
rect 28997 2329 29009 2363
rect 29043 2360 29055 2363
rect 29914 2360 29920 2372
rect 29043 2332 29920 2360
rect 29043 2329 29055 2332
rect 28997 2323 29055 2329
rect 29914 2320 29920 2332
rect 29972 2320 29978 2372
rect 30466 2320 30472 2372
rect 30524 2320 30530 2372
rect 31018 2320 31024 2372
rect 31076 2360 31082 2372
rect 31389 2363 31447 2369
rect 31389 2360 31401 2363
rect 31076 2332 31401 2360
rect 31076 2320 31082 2332
rect 31389 2329 31401 2332
rect 31435 2329 31447 2363
rect 31389 2323 31447 2329
rect 31754 2320 31760 2372
rect 31812 2360 31818 2372
rect 32416 2360 32444 2400
rect 33229 2397 33241 2400
rect 33275 2397 33287 2431
rect 33229 2391 33287 2397
rect 33686 2388 33692 2440
rect 33744 2428 33750 2440
rect 34885 2431 34943 2437
rect 34885 2428 34897 2431
rect 33744 2400 34897 2428
rect 33744 2388 33750 2400
rect 34885 2397 34897 2400
rect 34931 2397 34943 2431
rect 34885 2391 34943 2397
rect 35805 2431 35863 2437
rect 35805 2397 35817 2431
rect 35851 2428 35863 2431
rect 36722 2428 36728 2440
rect 35851 2400 36728 2428
rect 35851 2397 35863 2400
rect 35805 2391 35863 2397
rect 36722 2388 36728 2400
rect 36780 2388 36786 2440
rect 37461 2431 37519 2437
rect 37461 2397 37473 2431
rect 37507 2397 37519 2431
rect 37461 2391 37519 2397
rect 31812 2332 32444 2360
rect 31812 2320 31818 2332
rect 32582 2320 32588 2372
rect 32640 2320 32646 2372
rect 33134 2320 33140 2372
rect 33192 2360 33198 2372
rect 33505 2363 33563 2369
rect 33505 2360 33517 2363
rect 33192 2332 33517 2360
rect 33192 2320 33198 2332
rect 33505 2329 33517 2332
rect 33551 2329 33563 2363
rect 33505 2323 33563 2329
rect 34514 2320 34520 2372
rect 34572 2360 34578 2372
rect 35161 2363 35219 2369
rect 35161 2360 35173 2363
rect 34572 2332 35173 2360
rect 34572 2320 34578 2332
rect 35161 2329 35173 2332
rect 35207 2329 35219 2363
rect 35161 2323 35219 2329
rect 36078 2320 36084 2372
rect 36136 2320 36142 2372
rect 24946 2292 24952 2304
rect 22940 2264 24952 2292
rect 24946 2252 24952 2264
rect 25004 2252 25010 2304
rect 28077 2295 28135 2301
rect 28077 2261 28089 2295
rect 28123 2292 28135 2295
rect 28902 2292 28908 2304
rect 28123 2264 28908 2292
rect 28123 2261 28135 2264
rect 28077 2255 28135 2261
rect 28902 2252 28908 2264
rect 28960 2252 28966 2304
rect 37476 2292 37504 2391
rect 37550 2388 37556 2440
rect 37608 2428 37614 2440
rect 38381 2431 38439 2437
rect 38381 2428 38393 2431
rect 37608 2400 38393 2428
rect 37608 2388 37614 2400
rect 38381 2397 38393 2400
rect 38427 2397 38439 2431
rect 38381 2391 38439 2397
rect 38488 2400 38792 2428
rect 37734 2320 37740 2372
rect 37792 2320 37798 2372
rect 37826 2320 37832 2372
rect 37884 2360 37890 2372
rect 38488 2360 38516 2400
rect 37884 2332 38516 2360
rect 37884 2320 37890 2332
rect 38654 2320 38660 2372
rect 38712 2320 38718 2372
rect 38764 2360 38792 2400
rect 39298 2388 39304 2440
rect 39356 2428 39362 2440
rect 40037 2431 40095 2437
rect 40037 2428 40049 2431
rect 39356 2400 40049 2428
rect 39356 2388 39362 2400
rect 40037 2397 40049 2400
rect 40083 2397 40095 2431
rect 40037 2391 40095 2397
rect 40144 2400 41276 2428
rect 40144 2360 40172 2400
rect 38764 2332 40172 2360
rect 40310 2320 40316 2372
rect 40368 2320 40374 2372
rect 40954 2320 40960 2372
rect 41012 2360 41018 2372
rect 41141 2363 41199 2369
rect 41141 2360 41153 2363
rect 41012 2332 41153 2360
rect 41012 2320 41018 2332
rect 41141 2329 41153 2332
rect 41187 2329 41199 2363
rect 41141 2323 41199 2329
rect 40862 2292 40868 2304
rect 37476 2264 40868 2292
rect 40862 2252 40868 2264
rect 40920 2252 40926 2304
rect 41248 2292 41276 2400
rect 41414 2388 41420 2440
rect 41472 2428 41478 2440
rect 43625 2431 43683 2437
rect 43625 2428 43637 2431
rect 41472 2400 43637 2428
rect 41472 2388 41478 2400
rect 43625 2397 43637 2400
rect 43671 2397 43683 2431
rect 43625 2391 43683 2397
rect 47946 2388 47952 2440
rect 48004 2388 48010 2440
rect 48130 2437 48136 2440
rect 48097 2431 48136 2437
rect 48097 2397 48109 2431
rect 48097 2391 48136 2397
rect 48130 2388 48136 2391
rect 48188 2388 48194 2440
rect 48314 2388 48320 2440
rect 48372 2388 48378 2440
rect 48414 2431 48472 2437
rect 48414 2397 48426 2431
rect 48460 2428 48472 2431
rect 48590 2428 48596 2440
rect 48460 2400 48596 2428
rect 48460 2397 48472 2400
rect 48414 2391 48472 2397
rect 48590 2388 48596 2400
rect 48648 2388 48654 2440
rect 51074 2388 51080 2440
rect 51132 2428 51138 2440
rect 51445 2431 51503 2437
rect 51445 2428 51457 2431
rect 51132 2400 51457 2428
rect 51132 2388 51138 2400
rect 51445 2397 51457 2400
rect 51491 2397 51503 2431
rect 51445 2391 51503 2397
rect 53926 2388 53932 2440
rect 53984 2428 53990 2440
rect 57072 2437 57100 2536
rect 58250 2524 58256 2536
rect 58308 2524 58314 2576
rect 58342 2524 58348 2576
rect 58400 2524 58406 2576
rect 57333 2499 57391 2505
rect 57333 2465 57345 2499
rect 57379 2496 57391 2499
rect 58894 2496 58900 2508
rect 57379 2468 58900 2496
rect 57379 2465 57391 2468
rect 57333 2459 57391 2465
rect 58894 2456 58900 2468
rect 58952 2456 58958 2508
rect 54021 2431 54079 2437
rect 54021 2428 54033 2431
rect 53984 2400 54033 2428
rect 53984 2388 53990 2400
rect 54021 2397 54033 2400
rect 54067 2397 54079 2431
rect 54021 2391 54079 2397
rect 57057 2431 57115 2437
rect 57057 2397 57069 2431
rect 57103 2397 57115 2431
rect 58986 2428 58992 2440
rect 57057 2391 57115 2397
rect 57256 2400 58992 2428
rect 41782 2320 41788 2372
rect 41840 2360 41846 2372
rect 42705 2363 42763 2369
rect 42705 2360 42717 2363
rect 41840 2332 42717 2360
rect 41840 2320 41846 2332
rect 42705 2329 42717 2332
rect 42751 2329 42763 2363
rect 42705 2323 42763 2329
rect 43806 2320 43812 2372
rect 43864 2360 43870 2372
rect 44361 2363 44419 2369
rect 44361 2360 44373 2363
rect 43864 2332 44373 2360
rect 43864 2320 43870 2332
rect 44361 2329 44373 2332
rect 44407 2329 44419 2363
rect 44361 2323 44419 2329
rect 44450 2320 44456 2372
rect 44508 2360 44514 2372
rect 45281 2363 45339 2369
rect 45281 2360 45293 2363
rect 44508 2332 45293 2360
rect 44508 2320 44514 2332
rect 45281 2329 45293 2332
rect 45327 2329 45339 2363
rect 45281 2323 45339 2329
rect 46014 2320 46020 2372
rect 46072 2320 46078 2372
rect 46106 2320 46112 2372
rect 46164 2360 46170 2372
rect 46753 2363 46811 2369
rect 46753 2360 46765 2363
rect 46164 2332 46765 2360
rect 46164 2320 46170 2332
rect 46753 2329 46765 2332
rect 46799 2329 46811 2363
rect 46753 2323 46811 2329
rect 47762 2320 47768 2372
rect 47820 2360 47826 2372
rect 48225 2363 48283 2369
rect 48225 2360 48237 2363
rect 47820 2332 48237 2360
rect 47820 2320 47826 2332
rect 48225 2329 48237 2332
rect 48271 2329 48283 2363
rect 48225 2323 48283 2329
rect 48498 2320 48504 2372
rect 48556 2360 48562 2372
rect 49237 2363 49295 2369
rect 49237 2360 49249 2363
rect 48556 2332 49249 2360
rect 48556 2320 48562 2332
rect 49237 2329 49249 2332
rect 49283 2329 49295 2363
rect 49237 2323 49295 2329
rect 49878 2320 49884 2372
rect 49936 2360 49942 2372
rect 50433 2363 50491 2369
rect 50433 2360 50445 2363
rect 49936 2332 50445 2360
rect 49936 2320 49942 2332
rect 50433 2329 50445 2332
rect 50479 2329 50491 2363
rect 50433 2323 50491 2329
rect 51258 2320 51264 2372
rect 51316 2360 51322 2372
rect 53009 2363 53067 2369
rect 53009 2360 53021 2363
rect 51316 2332 53021 2360
rect 51316 2320 51322 2332
rect 53009 2329 53021 2332
rect 53055 2329 53067 2363
rect 53009 2323 53067 2329
rect 55582 2320 55588 2372
rect 55640 2320 55646 2372
rect 56321 2363 56379 2369
rect 56321 2329 56333 2363
rect 56367 2360 56379 2363
rect 57256 2360 57284 2400
rect 58986 2388 58992 2400
rect 59044 2388 59050 2440
rect 56367 2332 57284 2360
rect 56367 2329 56379 2332
rect 56321 2323 56379 2329
rect 57330 2320 57336 2372
rect 57388 2360 57394 2372
rect 58161 2363 58219 2369
rect 58161 2360 58173 2363
rect 57388 2332 58173 2360
rect 57388 2320 57394 2332
rect 58161 2329 58173 2332
rect 58207 2329 58219 2363
rect 58161 2323 58219 2329
rect 43717 2295 43775 2301
rect 43717 2292 43729 2295
rect 41248 2264 43729 2292
rect 43717 2261 43729 2264
rect 43763 2261 43775 2295
rect 43717 2255 43775 2261
rect 1104 2202 58880 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 50294 2202
rect 50346 2150 50358 2202
rect 50410 2150 50422 2202
rect 50474 2150 50486 2202
rect 50538 2150 50550 2202
rect 50602 2150 58880 2202
rect 1104 2128 58880 2150
rect 18598 2048 18604 2100
rect 18656 2088 18662 2100
rect 22370 2088 22376 2100
rect 18656 2060 22376 2088
rect 18656 2048 18662 2060
rect 22370 2048 22376 2060
rect 22428 2048 22434 2100
rect 48130 2048 48136 2100
rect 48188 2088 48194 2100
rect 56042 2088 56048 2100
rect 48188 2060 56048 2088
rect 48188 2048 48194 2060
rect 56042 2048 56048 2060
rect 56100 2048 56106 2100
rect 18230 1980 18236 2032
rect 18288 2020 18294 2032
rect 20622 2020 20628 2032
rect 18288 1992 20628 2020
rect 18288 1980 18294 1992
rect 20622 1980 20628 1992
rect 20680 1980 20686 2032
rect 23566 1980 23572 2032
rect 23624 2020 23630 2032
rect 44634 2020 44640 2032
rect 23624 1992 44640 2020
rect 23624 1980 23630 1992
rect 44634 1980 44640 1992
rect 44692 1980 44698 2032
rect 15838 1912 15844 1964
rect 15896 1952 15902 1964
rect 30558 1952 30564 1964
rect 15896 1924 30564 1952
rect 15896 1912 15902 1924
rect 30558 1912 30564 1924
rect 30616 1912 30622 1964
rect 22646 1776 22652 1828
rect 22704 1816 22710 1828
rect 39482 1816 39488 1828
rect 22704 1788 39488 1816
rect 22704 1776 22710 1788
rect 39482 1776 39488 1788
rect 39540 1776 39546 1828
rect 22830 1504 22836 1556
rect 22888 1544 22894 1556
rect 24394 1544 24400 1556
rect 22888 1516 24400 1544
rect 22888 1504 22894 1516
rect 24394 1504 24400 1516
rect 24452 1504 24458 1556
rect 36262 1232 36268 1284
rect 36320 1272 36326 1284
rect 39666 1272 39672 1284
rect 36320 1244 39672 1272
rect 36320 1232 36326 1244
rect 39666 1232 39672 1244
rect 39724 1232 39730 1284
rect 50338 1232 50344 1284
rect 50396 1272 50402 1284
rect 54386 1272 54392 1284
rect 50396 1244 54392 1272
rect 50396 1232 50402 1244
rect 54386 1232 54392 1244
rect 54444 1232 54450 1284
rect 34330 1164 34336 1216
rect 34388 1204 34394 1216
rect 36170 1204 36176 1216
rect 34388 1176 36176 1204
rect 34388 1164 34394 1176
rect 36170 1164 36176 1176
rect 36228 1164 36234 1216
rect 36814 1164 36820 1216
rect 36872 1204 36878 1216
rect 38746 1204 38752 1216
rect 36872 1176 38752 1204
rect 36872 1164 36878 1176
rect 38746 1164 38752 1176
rect 38804 1164 38810 1216
rect 39022 1164 39028 1216
rect 39080 1204 39086 1216
rect 43346 1204 43352 1216
rect 39080 1176 43352 1204
rect 39080 1164 39086 1176
rect 43346 1164 43352 1176
rect 43404 1164 43410 1216
rect 47026 1164 47032 1216
rect 47084 1204 47090 1216
rect 51534 1204 51540 1216
rect 47084 1176 51540 1204
rect 47084 1164 47090 1176
rect 51534 1164 51540 1176
rect 51592 1164 51598 1216
rect 53650 1164 53656 1216
rect 53708 1204 53714 1216
rect 56962 1204 56968 1216
rect 53708 1176 56968 1204
rect 53708 1164 53714 1176
rect 56962 1164 56968 1176
rect 57020 1164 57026 1216
rect 7926 1096 7932 1148
rect 7984 1136 7990 1148
rect 9214 1136 9220 1148
rect 7984 1108 9220 1136
rect 7984 1096 7990 1108
rect 9214 1096 9220 1108
rect 9272 1096 9278 1148
rect 35710 1096 35716 1148
rect 35768 1136 35774 1148
rect 38654 1136 38660 1148
rect 35768 1108 38660 1136
rect 35768 1096 35774 1108
rect 38654 1096 38660 1108
rect 38712 1096 38718 1148
rect 39850 1096 39856 1148
rect 39908 1136 39914 1148
rect 44082 1136 44088 1148
rect 39908 1108 44088 1136
rect 39908 1096 39914 1108
rect 44082 1096 44088 1108
rect 44140 1096 44146 1148
rect 47578 1096 47584 1148
rect 47636 1136 47642 1148
rect 49970 1136 49976 1148
rect 47636 1108 49976 1136
rect 47636 1096 47642 1108
rect 49970 1096 49976 1108
rect 50028 1096 50034 1148
rect 52546 1096 52552 1148
rect 52604 1136 52610 1148
rect 55950 1136 55956 1148
rect 52604 1108 55956 1136
rect 52604 1096 52610 1108
rect 55950 1096 55956 1108
rect 56008 1096 56014 1148
rect 8386 1028 8392 1080
rect 8444 1068 8450 1080
rect 10870 1068 10876 1080
rect 8444 1040 10876 1068
rect 8444 1028 8450 1040
rect 10870 1028 10876 1040
rect 10928 1028 10934 1080
rect 13262 1028 13268 1080
rect 13320 1068 13326 1080
rect 13906 1068 13912 1080
rect 13320 1040 13912 1068
rect 13320 1028 13326 1040
rect 13906 1028 13912 1040
rect 13964 1028 13970 1080
rect 17862 1028 17868 1080
rect 17920 1068 17926 1080
rect 19978 1068 19984 1080
rect 17920 1040 19984 1068
rect 17920 1028 17926 1040
rect 19978 1028 19984 1040
rect 20036 1028 20042 1080
rect 20530 1028 20536 1080
rect 20588 1068 20594 1080
rect 22186 1068 22192 1080
rect 20588 1040 22192 1068
rect 20588 1028 20594 1040
rect 22186 1028 22192 1040
rect 22244 1028 22250 1080
rect 34882 1028 34888 1080
rect 34940 1068 34946 1080
rect 37734 1068 37740 1080
rect 34940 1040 37740 1068
rect 34940 1028 34946 1040
rect 37734 1028 37740 1040
rect 37792 1028 37798 1080
rect 39298 1028 39304 1080
rect 39356 1068 39362 1080
rect 43254 1068 43260 1080
rect 39356 1040 43260 1068
rect 39356 1028 39362 1040
rect 43254 1028 43260 1040
rect 43312 1028 43318 1080
rect 43714 1028 43720 1080
rect 43772 1068 43778 1080
rect 46290 1068 46296 1080
rect 43772 1040 46296 1068
rect 43772 1028 43778 1040
rect 46290 1028 46296 1040
rect 46348 1028 46354 1080
rect 47302 1028 47308 1080
rect 47360 1068 47366 1080
rect 51258 1068 51264 1080
rect 47360 1040 51264 1068
rect 47360 1028 47366 1040
rect 51258 1028 51264 1040
rect 51316 1028 51322 1080
rect 51718 1028 51724 1080
rect 51776 1068 51782 1080
rect 55214 1068 55220 1080
rect 51776 1040 55220 1068
rect 51776 1028 51782 1040
rect 55214 1028 55220 1040
rect 55272 1028 55278 1080
rect 6822 960 6828 1012
rect 6880 1000 6886 1012
rect 7834 1000 7840 1012
rect 6880 972 7840 1000
rect 6880 960 6886 972
rect 7834 960 7840 972
rect 7892 960 7898 1012
rect 9030 960 9036 1012
rect 9088 1000 9094 1012
rect 10594 1000 10600 1012
rect 9088 972 10600 1000
rect 9088 960 9094 972
rect 10594 960 10600 972
rect 10652 960 10658 1012
rect 10962 960 10968 1012
rect 11020 1000 11026 1012
rect 12250 1000 12256 1012
rect 11020 972 12256 1000
rect 11020 960 11026 972
rect 12250 960 12256 972
rect 12308 960 12314 1012
rect 13538 960 13544 1012
rect 13596 1000 13602 1012
rect 14734 1000 14740 1012
rect 13596 972 14740 1000
rect 13596 960 13602 972
rect 14734 960 14740 972
rect 14792 960 14798 1012
rect 17402 960 17408 1012
rect 17460 1000 17466 1012
rect 18874 1000 18880 1012
rect 17460 972 18880 1000
rect 17460 960 17466 972
rect 18874 960 18880 972
rect 18932 960 18938 1012
rect 20438 960 20444 1012
rect 20496 1000 20502 1012
rect 20806 1000 20812 1012
rect 20496 972 20812 1000
rect 20496 960 20502 972
rect 20806 960 20812 972
rect 20864 960 20870 1012
rect 21174 960 21180 1012
rect 21232 1000 21238 1012
rect 22738 1000 22744 1012
rect 21232 972 22744 1000
rect 21232 960 21238 972
rect 22738 960 22744 972
rect 22796 960 22802 1012
rect 23750 960 23756 1012
rect 23808 1000 23814 1012
rect 25222 1000 25228 1012
rect 23808 972 25228 1000
rect 23808 960 23814 972
rect 25222 960 25228 972
rect 25280 960 25286 1012
rect 31846 960 31852 1012
rect 31904 1000 31910 1012
rect 33134 1000 33140 1012
rect 31904 972 33140 1000
rect 31904 960 31910 972
rect 33134 960 33140 972
rect 33192 960 33198 1012
rect 33778 960 33784 1012
rect 33836 1000 33842 1012
rect 36078 1000 36084 1012
rect 33836 972 36084 1000
rect 33836 960 33842 972
rect 36078 960 36084 972
rect 36136 960 36142 1012
rect 36538 960 36544 1012
rect 36596 1000 36602 1012
rect 40310 1000 40316 1012
rect 36596 972 40316 1000
rect 36596 960 36602 972
rect 40310 960 40316 972
rect 40368 960 40374 1012
rect 42334 960 42340 1012
rect 42392 1000 42398 1012
rect 46014 1000 46020 1012
rect 42392 972 46020 1000
rect 42392 960 42398 972
rect 46014 960 46020 972
rect 46072 960 46078 1012
rect 48958 960 48964 1012
rect 49016 1000 49022 1012
rect 52638 1000 52644 1012
rect 49016 972 52644 1000
rect 49016 960 49022 972
rect 52638 960 52644 972
rect 52696 960 52702 1012
rect 52822 960 52828 1012
rect 52880 1000 52886 1012
rect 57330 1000 57336 1012
rect 52880 972 57336 1000
rect 52880 960 52886 972
rect 57330 960 57336 972
rect 57388 960 57394 1012
rect 5810 892 5816 944
rect 5868 932 5874 944
rect 7282 932 7288 944
rect 5868 904 7288 932
rect 5868 892 5874 904
rect 7282 892 7288 904
rect 7340 892 7346 944
rect 8018 892 8024 944
rect 8076 932 8082 944
rect 9490 932 9496 944
rect 8076 904 9496 932
rect 8076 892 8082 904
rect 9490 892 9496 904
rect 9548 892 9554 944
rect 10226 892 10232 944
rect 10284 932 10290 944
rect 11974 932 11980 944
rect 10284 904 11980 932
rect 10284 892 10290 904
rect 11974 892 11980 904
rect 12032 892 12038 944
rect 12066 892 12072 944
rect 12124 932 12130 944
rect 13078 932 13084 944
rect 12124 904 13084 932
rect 12124 892 12130 904
rect 13078 892 13084 904
rect 13136 892 13142 944
rect 13722 892 13728 944
rect 13780 932 13786 944
rect 14458 932 14464 944
rect 13780 904 14464 932
rect 13780 892 13786 904
rect 14458 892 14464 904
rect 14516 892 14522 944
rect 17034 892 17040 944
rect 17092 932 17098 944
rect 18598 932 18604 944
rect 17092 904 18604 932
rect 17092 892 17098 904
rect 18598 892 18604 904
rect 18656 892 18662 944
rect 18690 892 18696 944
rect 18748 932 18754 944
rect 20530 932 20536 944
rect 18748 904 20536 932
rect 18748 892 18754 904
rect 20530 892 20536 904
rect 20588 892 20594 944
rect 20622 892 20628 944
rect 20680 932 20686 944
rect 21634 932 21640 944
rect 20680 904 21640 932
rect 20680 892 20686 904
rect 21634 892 21640 904
rect 21692 892 21698 944
rect 24762 892 24768 944
rect 24820 932 24826 944
rect 25498 932 25504 944
rect 24820 904 25504 932
rect 24820 892 24826 904
rect 25498 892 25504 904
rect 25556 892 25562 944
rect 27522 892 27528 944
rect 27580 932 27586 944
rect 27982 932 27988 944
rect 27580 904 27988 932
rect 27580 892 27586 904
rect 27982 892 27988 904
rect 28040 892 28046 944
rect 31294 892 31300 944
rect 31352 932 31358 944
rect 32582 932 32588 944
rect 31352 904 32588 932
rect 31352 892 31358 904
rect 32582 892 32588 904
rect 32640 892 32646 944
rect 32950 892 32956 944
rect 33008 932 33014 944
rect 34514 932 34520 944
rect 33008 904 34520 932
rect 33008 892 33014 904
rect 34514 892 34520 904
rect 34572 892 34578 944
rect 35434 892 35440 944
rect 35492 932 35498 944
rect 37274 932 37280 944
rect 35492 904 37280 932
rect 35492 892 35498 904
rect 37274 892 37280 904
rect 37332 892 37338 944
rect 37642 892 37648 944
rect 37700 932 37706 944
rect 37700 904 37780 932
rect 37700 892 37706 904
rect 23198 824 23204 876
rect 23256 864 23262 876
rect 23750 864 23756 876
rect 23256 836 23756 864
rect 23256 824 23262 836
rect 23750 824 23756 836
rect 23808 824 23814 876
rect 37752 796 37780 904
rect 38746 892 38752 944
rect 38804 892 38810 944
rect 40678 892 40684 944
rect 40736 932 40742 944
rect 44450 932 44456 944
rect 40736 904 44456 932
rect 40736 892 40742 904
rect 44450 892 44456 904
rect 44508 892 44514 944
rect 44818 892 44824 944
rect 44876 932 44882 944
rect 46106 932 46112 944
rect 44876 904 46112 932
rect 44876 892 44882 904
rect 46106 892 46112 904
rect 46164 892 46170 944
rect 47854 892 47860 944
rect 47912 932 47918 944
rect 48498 932 48504 944
rect 47912 904 48504 932
rect 47912 892 47918 904
rect 48498 892 48504 904
rect 48556 892 48562 944
rect 49234 892 49240 944
rect 49292 932 49298 944
rect 49878 932 49884 944
rect 49292 904 49884 932
rect 49292 892 49298 904
rect 49878 892 49884 904
rect 49936 892 49942 944
rect 50890 892 50896 944
rect 50948 932 50954 944
rect 53006 932 53012 944
rect 50948 904 53012 932
rect 50948 892 50954 904
rect 53006 892 53012 904
rect 53064 892 53070 944
rect 53374 892 53380 944
rect 53432 932 53438 944
rect 55582 932 55588 944
rect 53432 904 55588 932
rect 53432 892 53438 904
rect 55582 892 55588 904
rect 55640 892 55646 944
rect 38764 864 38792 892
rect 43806 864 43812 876
rect 38764 836 43812 864
rect 43806 824 43812 836
rect 43864 824 43870 876
rect 48774 824 48780 876
rect 48832 864 48838 876
rect 51074 864 51080 876
rect 48832 836 51080 864
rect 48832 824 48838 836
rect 51074 824 51080 836
rect 51132 824 51138 876
rect 41414 796 41420 808
rect 37752 768 41420 796
rect 41414 756 41420 768
rect 41472 756 41478 808
rect 46658 756 46664 808
rect 46716 796 46722 808
rect 50798 796 50804 808
rect 46716 768 50804 796
rect 46716 756 46722 768
rect 50798 756 50804 768
rect 50856 756 50862 808
rect 44082 76 44088 128
rect 44140 116 44146 128
rect 49418 116 49424 128
rect 44140 88 49424 116
rect 44140 76 44146 88
rect 49418 76 49424 88
rect 49476 76 49482 128
<< via1 >>
rect 16396 59100 16448 59152
rect 16948 59100 17000 59152
rect 18972 59100 19024 59152
rect 19432 59100 19484 59152
rect 21548 59100 21600 59152
rect 22100 59100 22152 59152
rect 37004 59100 37056 59152
rect 37556 59100 37608 59152
rect 39580 59100 39632 59152
rect 40040 59100 40092 59152
rect 55036 59100 55088 59152
rect 55588 59100 55640 59152
rect 56784 57944 56836 57996
rect 58992 57944 59044 57996
rect 19574 57638 19626 57690
rect 19638 57638 19690 57690
rect 19702 57638 19754 57690
rect 19766 57638 19818 57690
rect 19830 57638 19882 57690
rect 50294 57638 50346 57690
rect 50358 57638 50410 57690
rect 50422 57638 50474 57690
rect 50486 57638 50538 57690
rect 50550 57638 50602 57690
rect 2228 57468 2280 57520
rect 3516 57468 3568 57520
rect 4804 57468 4856 57520
rect 7380 57468 7432 57520
rect 8668 57468 8720 57520
rect 9956 57468 10008 57520
rect 12532 57468 12584 57520
rect 16948 57511 17000 57520
rect 16948 57477 16957 57511
rect 16957 57477 16991 57511
rect 16991 57477 17000 57511
rect 16948 57468 17000 57477
rect 17684 57468 17736 57520
rect 20260 57468 20312 57520
rect 22100 57511 22152 57520
rect 22100 57477 22109 57511
rect 22109 57477 22143 57511
rect 22143 57477 22152 57511
rect 22100 57468 22152 57477
rect 22836 57468 22888 57520
rect 25412 57468 25464 57520
rect 26700 57468 26752 57520
rect 27988 57468 28040 57520
rect 29276 57468 29328 57520
rect 30564 57468 30616 57520
rect 31852 57468 31904 57520
rect 33140 57468 33192 57520
rect 34520 57468 34572 57520
rect 35900 57511 35952 57520
rect 35900 57477 35909 57511
rect 35909 57477 35943 57511
rect 35943 57477 35952 57511
rect 35900 57468 35952 57477
rect 37556 57511 37608 57520
rect 37556 57477 37565 57511
rect 37565 57477 37599 57511
rect 37599 57477 37608 57511
rect 37556 57468 37608 57477
rect 38292 57468 38344 57520
rect 40868 57468 40920 57520
rect 42156 57468 42208 57520
rect 43444 57468 43496 57520
rect 44732 57468 44784 57520
rect 47308 57468 47360 57520
rect 49884 57468 49936 57520
rect 53840 57468 53892 57520
rect 55588 57511 55640 57520
rect 55588 57477 55597 57511
rect 55597 57477 55631 57511
rect 55631 57477 55640 57511
rect 55588 57468 55640 57477
rect 56324 57468 56376 57520
rect 58992 57468 59044 57520
rect 6092 57400 6144 57452
rect 11244 57400 11296 57452
rect 13820 57400 13872 57452
rect 15200 57443 15252 57452
rect 15200 57409 15209 57443
rect 15209 57409 15243 57443
rect 15243 57409 15252 57443
rect 15200 57400 15252 57409
rect 19432 57443 19484 57452
rect 19432 57409 19441 57443
rect 19441 57409 19475 57443
rect 19475 57409 19484 57443
rect 19432 57400 19484 57409
rect 24124 57400 24176 57452
rect 40040 57443 40092 57452
rect 40040 57409 40049 57443
rect 40049 57409 40083 57443
rect 40083 57409 40092 57443
rect 40040 57400 40092 57409
rect 46020 57400 46072 57452
rect 48596 57400 48648 57452
rect 51172 57400 51224 57452
rect 52460 57400 52512 57452
rect 58900 57400 58952 57452
rect 26884 57332 26936 57384
rect 3424 57264 3476 57316
rect 17132 57307 17184 57316
rect 17132 57273 17141 57307
rect 17141 57273 17175 57307
rect 17175 57273 17184 57307
rect 17132 57264 17184 57273
rect 52644 57264 52696 57316
rect 56692 57264 56744 57316
rect 58808 57264 58860 57316
rect 3976 57196 4028 57248
rect 4712 57196 4764 57248
rect 6736 57239 6788 57248
rect 6736 57205 6745 57239
rect 6745 57205 6779 57239
rect 6779 57205 6788 57239
rect 6736 57196 6788 57205
rect 7380 57196 7432 57248
rect 9128 57196 9180 57248
rect 9956 57196 10008 57248
rect 11888 57239 11940 57248
rect 11888 57205 11897 57239
rect 11897 57205 11931 57239
rect 11931 57205 11940 57239
rect 11888 57196 11940 57205
rect 12808 57239 12860 57248
rect 12808 57205 12817 57239
rect 12817 57205 12851 57239
rect 12851 57205 12860 57239
rect 12808 57196 12860 57205
rect 15384 57239 15436 57248
rect 15384 57205 15393 57239
rect 15393 57205 15427 57239
rect 15427 57205 15436 57239
rect 15384 57196 15436 57205
rect 17960 57239 18012 57248
rect 17960 57205 17969 57239
rect 17969 57205 18003 57239
rect 18003 57205 18012 57239
rect 17960 57196 18012 57205
rect 19984 57196 20036 57248
rect 20168 57196 20220 57248
rect 22192 57239 22244 57248
rect 22192 57205 22201 57239
rect 22201 57205 22235 57239
rect 22235 57205 22244 57239
rect 22192 57196 22244 57205
rect 22652 57196 22704 57248
rect 24768 57239 24820 57248
rect 24768 57205 24777 57239
rect 24777 57205 24811 57239
rect 24811 57205 24820 57239
rect 24768 57196 24820 57205
rect 25688 57239 25740 57248
rect 25688 57205 25697 57239
rect 25697 57205 25731 57239
rect 25731 57205 25740 57239
rect 25688 57196 25740 57205
rect 26700 57196 26752 57248
rect 27988 57196 28040 57248
rect 29920 57239 29972 57248
rect 29920 57205 29929 57239
rect 29929 57205 29963 57239
rect 29963 57205 29972 57239
rect 29920 57196 29972 57205
rect 30840 57239 30892 57248
rect 30840 57205 30849 57239
rect 30849 57205 30883 57239
rect 30883 57205 30892 57239
rect 30840 57196 30892 57205
rect 31208 57196 31260 57248
rect 33416 57239 33468 57248
rect 33416 57205 33425 57239
rect 33425 57205 33459 57239
rect 33459 57205 33468 57239
rect 33416 57196 33468 57205
rect 34796 57196 34848 57248
rect 35624 57196 35676 57248
rect 37096 57196 37148 57248
rect 37924 57196 37976 57248
rect 39304 57196 39356 57248
rect 40316 57196 40368 57248
rect 41696 57196 41748 57248
rect 43628 57196 43680 57248
rect 45376 57239 45428 57248
rect 45376 57205 45385 57239
rect 45385 57205 45419 57239
rect 45419 57205 45428 57239
rect 45376 57196 45428 57205
rect 46296 57239 46348 57248
rect 46296 57205 46305 57239
rect 46305 57205 46339 57239
rect 46339 57205 46348 57239
rect 46296 57196 46348 57205
rect 46388 57196 46440 57248
rect 48872 57239 48924 57248
rect 48872 57205 48881 57239
rect 48881 57205 48915 57239
rect 48915 57205 48924 57239
rect 48872 57196 48924 57205
rect 49056 57196 49108 57248
rect 51448 57239 51500 57248
rect 51448 57205 51457 57239
rect 51457 57205 51491 57239
rect 51491 57205 51500 57239
rect 51448 57196 51500 57205
rect 51724 57196 51776 57248
rect 53932 57196 53984 57248
rect 54116 57196 54168 57248
rect 57244 57239 57296 57248
rect 57244 57205 57253 57239
rect 57253 57205 57287 57239
rect 57287 57205 57296 57239
rect 57244 57196 57296 57205
rect 58256 57239 58308 57248
rect 58256 57205 58265 57239
rect 58265 57205 58299 57239
rect 58299 57205 58308 57239
rect 58256 57196 58308 57205
rect 4214 57094 4266 57146
rect 4278 57094 4330 57146
rect 4342 57094 4394 57146
rect 4406 57094 4458 57146
rect 4470 57094 4522 57146
rect 34934 57094 34986 57146
rect 34998 57094 35050 57146
rect 35062 57094 35114 57146
rect 35126 57094 35178 57146
rect 35190 57094 35242 57146
rect 22192 56992 22244 57044
rect 31576 56992 31628 57044
rect 57428 56992 57480 57044
rect 58992 56992 59044 57044
rect 53564 56924 53616 56976
rect 58256 56924 58308 56976
rect 17960 56856 18012 56908
rect 30472 56856 30524 56908
rect 58992 56856 59044 56908
rect 56784 56831 56836 56840
rect 56784 56797 56793 56831
rect 56793 56797 56827 56831
rect 56827 56797 56836 56831
rect 56784 56788 56836 56797
rect 57612 56788 57664 56840
rect 52460 56720 52512 56772
rect 59452 56720 59504 56772
rect 56232 56695 56284 56704
rect 56232 56661 56241 56695
rect 56241 56661 56275 56695
rect 56275 56661 56284 56695
rect 56232 56652 56284 56661
rect 19574 56550 19626 56602
rect 19638 56550 19690 56602
rect 19702 56550 19754 56602
rect 19766 56550 19818 56602
rect 19830 56550 19882 56602
rect 50294 56550 50346 56602
rect 50358 56550 50410 56602
rect 50422 56550 50474 56602
rect 50486 56550 50538 56602
rect 50550 56550 50602 56602
rect 58716 56448 58768 56500
rect 56692 56380 56744 56432
rect 58992 56380 59044 56432
rect 940 56312 992 56364
rect 58164 56355 58216 56364
rect 58164 56321 58173 56355
rect 58173 56321 58207 56355
rect 58207 56321 58216 56355
rect 58164 56312 58216 56321
rect 18604 56244 18656 56296
rect 55220 56244 55272 56296
rect 53840 56176 53892 56228
rect 52552 56108 52604 56160
rect 56048 56108 56100 56160
rect 4214 56006 4266 56058
rect 4278 56006 4330 56058
rect 4342 56006 4394 56058
rect 4406 56006 4458 56058
rect 4470 56006 4522 56058
rect 34934 56006 34986 56058
rect 34998 56006 35050 56058
rect 35062 56006 35114 56058
rect 35126 56006 35178 56058
rect 35190 56006 35242 56058
rect 26792 55836 26844 55888
rect 52460 55836 52512 55888
rect 53196 55836 53248 55888
rect 940 55700 992 55752
rect 57428 55743 57480 55752
rect 57428 55709 57437 55743
rect 57437 55709 57471 55743
rect 57471 55709 57480 55743
rect 57428 55700 57480 55709
rect 58992 55700 59044 55752
rect 21364 55632 21416 55684
rect 57520 55607 57572 55616
rect 57520 55573 57529 55607
rect 57529 55573 57563 55607
rect 57563 55573 57572 55607
rect 57520 55564 57572 55573
rect 19574 55462 19626 55514
rect 19638 55462 19690 55514
rect 19702 55462 19754 55514
rect 19766 55462 19818 55514
rect 19830 55462 19882 55514
rect 50294 55462 50346 55514
rect 50358 55462 50410 55514
rect 50422 55462 50474 55514
rect 50486 55462 50538 55514
rect 50550 55462 50602 55514
rect 59084 55360 59136 55412
rect 1032 55224 1084 55276
rect 58808 55224 58860 55276
rect 1952 55063 2004 55072
rect 1952 55029 1961 55063
rect 1961 55029 1995 55063
rect 1995 55029 2004 55063
rect 1952 55020 2004 55029
rect 4214 54918 4266 54970
rect 4278 54918 4330 54970
rect 4342 54918 4394 54970
rect 4406 54918 4458 54970
rect 4470 54918 4522 54970
rect 34934 54918 34986 54970
rect 34998 54918 35050 54970
rect 35062 54918 35114 54970
rect 35126 54918 35178 54970
rect 35190 54918 35242 54970
rect 58992 54612 59044 54664
rect 940 54544 992 54596
rect 2688 54544 2740 54596
rect 58900 54544 58952 54596
rect 56600 54476 56652 54528
rect 58256 54519 58308 54528
rect 58256 54485 58265 54519
rect 58265 54485 58299 54519
rect 58299 54485 58308 54519
rect 58256 54476 58308 54485
rect 19574 54374 19626 54426
rect 19638 54374 19690 54426
rect 19702 54374 19754 54426
rect 19766 54374 19818 54426
rect 19830 54374 19882 54426
rect 50294 54374 50346 54426
rect 50358 54374 50410 54426
rect 50422 54374 50474 54426
rect 50486 54374 50538 54426
rect 50550 54374 50602 54426
rect 1032 54136 1084 54188
rect 58992 54136 59044 54188
rect 2596 53932 2648 53984
rect 58532 53932 58584 53984
rect 4214 53830 4266 53882
rect 4278 53830 4330 53882
rect 4342 53830 4394 53882
rect 4406 53830 4458 53882
rect 4470 53830 4522 53882
rect 34934 53830 34986 53882
rect 34998 53830 35050 53882
rect 35062 53830 35114 53882
rect 35126 53830 35178 53882
rect 35190 53830 35242 53882
rect 940 53456 992 53508
rect 58164 53499 58216 53508
rect 58164 53465 58173 53499
rect 58173 53465 58207 53499
rect 58207 53465 58216 53499
rect 58164 53456 58216 53465
rect 58440 53456 58492 53508
rect 47860 53388 47912 53440
rect 19574 53286 19626 53338
rect 19638 53286 19690 53338
rect 19702 53286 19754 53338
rect 19766 53286 19818 53338
rect 19830 53286 19882 53338
rect 50294 53286 50346 53338
rect 50358 53286 50410 53338
rect 50422 53286 50474 53338
rect 50486 53286 50538 53338
rect 50550 53286 50602 53338
rect 1952 53184 2004 53236
rect 1032 53048 1084 53100
rect 48136 52980 48188 53032
rect 52460 53048 52512 53100
rect 58900 53048 58952 53100
rect 48504 52980 48556 53032
rect 11704 52844 11756 52896
rect 48044 52887 48096 52896
rect 48044 52853 48053 52887
rect 48053 52853 48087 52887
rect 48087 52853 48096 52887
rect 48044 52844 48096 52853
rect 58072 52844 58124 52896
rect 4214 52742 4266 52794
rect 4278 52742 4330 52794
rect 4342 52742 4394 52794
rect 4406 52742 4458 52794
rect 4470 52742 4522 52794
rect 34934 52742 34986 52794
rect 34998 52742 35050 52794
rect 35062 52742 35114 52794
rect 35126 52742 35178 52794
rect 35190 52742 35242 52794
rect 47676 52683 47728 52692
rect 47676 52649 47685 52683
rect 47685 52649 47719 52683
rect 47719 52649 47728 52683
rect 47676 52640 47728 52649
rect 55956 52572 56008 52624
rect 58164 52572 58216 52624
rect 11888 52436 11940 52488
rect 42340 52479 42392 52488
rect 42340 52445 42349 52479
rect 42349 52445 42383 52479
rect 42383 52445 42392 52479
rect 42340 52436 42392 52445
rect 58256 52504 58308 52556
rect 42524 52479 42576 52488
rect 42524 52445 42533 52479
rect 42533 52445 42567 52479
rect 42567 52445 42576 52479
rect 42524 52436 42576 52445
rect 47860 52479 47912 52488
rect 47860 52445 47869 52479
rect 47869 52445 47903 52479
rect 47903 52445 47912 52479
rect 47860 52436 47912 52445
rect 48136 52436 48188 52488
rect 940 52368 992 52420
rect 2044 52411 2096 52420
rect 2044 52377 2053 52411
rect 2053 52377 2087 52411
rect 2087 52377 2096 52411
rect 2044 52368 2096 52377
rect 48504 52479 48556 52488
rect 48504 52445 48513 52479
rect 48513 52445 48547 52479
rect 48547 52445 48556 52479
rect 48504 52436 48556 52445
rect 57520 52436 57572 52488
rect 58992 52436 59044 52488
rect 58164 52411 58216 52420
rect 58164 52377 58173 52411
rect 58173 52377 58207 52411
rect 58207 52377 58216 52411
rect 58164 52368 58216 52377
rect 42708 52343 42760 52352
rect 42708 52309 42717 52343
rect 42717 52309 42751 52343
rect 42751 52309 42760 52343
rect 42708 52300 42760 52309
rect 19574 52198 19626 52250
rect 19638 52198 19690 52250
rect 19702 52198 19754 52250
rect 19766 52198 19818 52250
rect 19830 52198 19882 52250
rect 50294 52198 50346 52250
rect 50358 52198 50410 52250
rect 50422 52198 50474 52250
rect 50486 52198 50538 52250
rect 50550 52198 50602 52250
rect 58992 52028 59044 52080
rect 1032 51960 1084 52012
rect 2044 51892 2096 51944
rect 47768 51935 47820 51944
rect 47768 51901 47777 51935
rect 47777 51901 47811 51935
rect 47811 51901 47820 51935
rect 47768 51892 47820 51901
rect 48136 51892 48188 51944
rect 53564 51960 53616 52012
rect 58808 51960 58860 52012
rect 48504 51892 48556 51944
rect 37280 51824 37332 51876
rect 46848 51756 46900 51808
rect 57980 51756 58032 51808
rect 4214 51654 4266 51706
rect 4278 51654 4330 51706
rect 4342 51654 4394 51706
rect 4406 51654 4458 51706
rect 4470 51654 4522 51706
rect 34934 51654 34986 51706
rect 34998 51654 35050 51706
rect 35062 51654 35114 51706
rect 35126 51654 35178 51706
rect 35190 51654 35242 51706
rect 2688 51552 2740 51604
rect 47952 51484 48004 51536
rect 48136 51484 48188 51536
rect 36912 51391 36964 51400
rect 36912 51357 36921 51391
rect 36921 51357 36955 51391
rect 36955 51357 36964 51391
rect 36912 51348 36964 51357
rect 37096 51391 37148 51400
rect 37096 51357 37103 51391
rect 37103 51357 37148 51391
rect 37096 51348 37148 51357
rect 37280 51391 37332 51400
rect 37280 51357 37289 51391
rect 37289 51357 37323 51391
rect 37323 51357 37332 51391
rect 37280 51348 37332 51357
rect 42524 51348 42576 51400
rect 46848 51391 46900 51400
rect 46848 51357 46857 51391
rect 46857 51357 46891 51391
rect 46891 51357 46900 51391
rect 46848 51348 46900 51357
rect 48228 51348 48280 51400
rect 48596 51416 48648 51468
rect 940 51280 992 51332
rect 2044 51323 2096 51332
rect 2044 51289 2053 51323
rect 2053 51289 2087 51323
rect 2087 51289 2096 51323
rect 2044 51280 2096 51289
rect 37188 51323 37240 51332
rect 37188 51289 37197 51323
rect 37197 51289 37231 51323
rect 37231 51289 37240 51323
rect 37188 51280 37240 51289
rect 47032 51323 47084 51332
rect 47032 51289 47041 51323
rect 47041 51289 47075 51323
rect 47075 51289 47084 51323
rect 47032 51280 47084 51289
rect 37556 51255 37608 51264
rect 37556 51221 37565 51255
rect 37565 51221 37599 51255
rect 37599 51221 37608 51255
rect 37556 51212 37608 51221
rect 47492 51280 47544 51332
rect 48872 51348 48924 51400
rect 58992 51348 59044 51400
rect 52644 51280 52696 51332
rect 58900 51280 58952 51332
rect 53840 51212 53892 51264
rect 57520 51255 57572 51264
rect 57520 51221 57529 51255
rect 57529 51221 57563 51255
rect 57563 51221 57572 51255
rect 57520 51212 57572 51221
rect 58716 51212 58768 51264
rect 19574 51110 19626 51162
rect 19638 51110 19690 51162
rect 19702 51110 19754 51162
rect 19766 51110 19818 51162
rect 19830 51110 19882 51162
rect 50294 51110 50346 51162
rect 50358 51110 50410 51162
rect 50422 51110 50474 51162
rect 50486 51110 50538 51162
rect 50550 51110 50602 51162
rect 47032 50940 47084 50992
rect 48136 50940 48188 50992
rect 1032 50872 1084 50924
rect 55220 51008 55272 51060
rect 48688 50940 48740 50992
rect 54116 50940 54168 50992
rect 2044 50804 2096 50856
rect 48872 50872 48924 50924
rect 47308 50804 47360 50856
rect 48504 50847 48556 50856
rect 48504 50813 48513 50847
rect 48513 50813 48547 50847
rect 48547 50813 48556 50847
rect 48504 50804 48556 50813
rect 2412 50668 2464 50720
rect 2596 50668 2648 50720
rect 49240 50736 49292 50788
rect 58256 50872 58308 50924
rect 55864 50804 55916 50856
rect 58072 50804 58124 50856
rect 49148 50668 49200 50720
rect 58072 50668 58124 50720
rect 4214 50566 4266 50618
rect 4278 50566 4330 50618
rect 4342 50566 4394 50618
rect 4406 50566 4458 50618
rect 4470 50566 4522 50618
rect 34934 50566 34986 50618
rect 34998 50566 35050 50618
rect 35062 50566 35114 50618
rect 35126 50566 35178 50618
rect 35190 50566 35242 50618
rect 48504 50464 48556 50516
rect 49424 50464 49476 50516
rect 48596 50396 48648 50448
rect 49240 50396 49292 50448
rect 49148 50328 49200 50380
rect 56048 50396 56100 50448
rect 49424 50371 49476 50380
rect 49424 50337 49433 50371
rect 49433 50337 49467 50371
rect 49467 50337 49476 50371
rect 49424 50328 49476 50337
rect 58348 50328 58400 50380
rect 59084 50328 59136 50380
rect 940 50192 992 50244
rect 48780 50192 48832 50244
rect 49608 50192 49660 50244
rect 58164 50235 58216 50244
rect 58164 50201 58173 50235
rect 58173 50201 58207 50235
rect 58207 50201 58216 50235
rect 58164 50192 58216 50201
rect 43076 50124 43128 50176
rect 56140 50124 56192 50176
rect 19574 50022 19626 50074
rect 19638 50022 19690 50074
rect 19702 50022 19754 50074
rect 19766 50022 19818 50074
rect 19830 50022 19882 50074
rect 50294 50022 50346 50074
rect 50358 50022 50410 50074
rect 50422 50022 50474 50074
rect 50486 50022 50538 50074
rect 50550 50022 50602 50074
rect 47032 49852 47084 49904
rect 1032 49784 1084 49836
rect 42524 49784 42576 49836
rect 1860 49716 1912 49768
rect 42616 49759 42668 49768
rect 42616 49725 42625 49759
rect 42625 49725 42659 49759
rect 42659 49725 42668 49759
rect 42616 49716 42668 49725
rect 43076 49827 43128 49836
rect 43076 49793 43085 49827
rect 43085 49793 43119 49827
rect 43119 49793 43128 49827
rect 43076 49784 43128 49793
rect 43260 49827 43312 49836
rect 43260 49793 43269 49827
rect 43269 49793 43303 49827
rect 43303 49793 43312 49827
rect 43260 49784 43312 49793
rect 56600 49784 56652 49836
rect 58992 49784 59044 49836
rect 48504 49716 48556 49768
rect 58624 49716 58676 49768
rect 4214 49478 4266 49530
rect 4278 49478 4330 49530
rect 4342 49478 4394 49530
rect 4406 49478 4458 49530
rect 4470 49478 4522 49530
rect 34934 49478 34986 49530
rect 34998 49478 35050 49530
rect 35062 49478 35114 49530
rect 35126 49478 35178 49530
rect 35190 49478 35242 49530
rect 30840 49240 30892 49292
rect 30472 49215 30524 49224
rect 30472 49181 30481 49215
rect 30481 49181 30515 49215
rect 30515 49181 30524 49215
rect 30472 49172 30524 49181
rect 940 49104 992 49156
rect 30380 49147 30432 49156
rect 30380 49113 30389 49147
rect 30389 49113 30423 49147
rect 30423 49113 30432 49147
rect 30380 49104 30432 49113
rect 1952 49079 2004 49088
rect 1952 49045 1961 49079
rect 1961 49045 1995 49079
rect 1995 49045 2004 49079
rect 1952 49036 2004 49045
rect 28356 49036 28408 49088
rect 31392 49104 31444 49156
rect 57980 49147 58032 49156
rect 57980 49113 57989 49147
rect 57989 49113 58023 49147
rect 58023 49113 58032 49147
rect 57980 49104 58032 49113
rect 30932 49036 30984 49088
rect 58072 49079 58124 49088
rect 58072 49045 58081 49079
rect 58081 49045 58115 49079
rect 58115 49045 58124 49079
rect 58072 49036 58124 49045
rect 19574 48934 19626 48986
rect 19638 48934 19690 48986
rect 19702 48934 19754 48986
rect 19766 48934 19818 48986
rect 19830 48934 19882 48986
rect 50294 48934 50346 48986
rect 50358 48934 50410 48986
rect 50422 48934 50474 48986
rect 50486 48934 50538 48986
rect 50550 48934 50602 48986
rect 1032 48696 1084 48748
rect 9956 48739 10008 48748
rect 9956 48705 9965 48739
rect 9965 48705 9999 48739
rect 9999 48705 10008 48739
rect 9956 48696 10008 48705
rect 10140 48739 10192 48748
rect 10140 48705 10149 48739
rect 10149 48705 10183 48739
rect 10183 48705 10192 48739
rect 10140 48696 10192 48705
rect 2228 48628 2280 48680
rect 57888 48764 57940 48816
rect 31392 48739 31444 48748
rect 31392 48705 31401 48739
rect 31401 48705 31435 48739
rect 31435 48705 31444 48739
rect 31392 48696 31444 48705
rect 31576 48739 31628 48748
rect 31576 48705 31585 48739
rect 31585 48705 31619 48739
rect 31619 48705 31628 48739
rect 31576 48696 31628 48705
rect 58808 48696 58860 48748
rect 33048 48628 33100 48680
rect 31484 48560 31536 48612
rect 10508 48535 10560 48544
rect 10508 48501 10517 48535
rect 10517 48501 10551 48535
rect 10551 48501 10560 48535
rect 10508 48492 10560 48501
rect 30656 48492 30708 48544
rect 56048 48492 56100 48544
rect 4214 48390 4266 48442
rect 4278 48390 4330 48442
rect 4342 48390 4394 48442
rect 4406 48390 4458 48442
rect 4470 48390 4522 48442
rect 34934 48390 34986 48442
rect 34998 48390 35050 48442
rect 35062 48390 35114 48442
rect 35126 48390 35178 48442
rect 35190 48390 35242 48442
rect 35716 48288 35768 48340
rect 35900 48288 35952 48340
rect 57888 48288 57940 48340
rect 58992 48288 59044 48340
rect 31392 48220 31444 48272
rect 58164 48220 58216 48272
rect 10508 48152 10560 48204
rect 40960 48152 41012 48204
rect 30380 48084 30432 48136
rect 31208 48127 31260 48136
rect 31208 48093 31215 48127
rect 31215 48093 31260 48127
rect 31208 48084 31260 48093
rect 31392 48127 31444 48136
rect 31392 48093 31401 48127
rect 31401 48093 31435 48127
rect 31435 48093 31444 48127
rect 31392 48084 31444 48093
rect 31484 48127 31536 48136
rect 31484 48093 31498 48127
rect 31498 48093 31532 48127
rect 31532 48093 31536 48127
rect 31484 48084 31536 48093
rect 34888 48127 34940 48136
rect 34888 48093 34897 48127
rect 34897 48093 34931 48127
rect 34931 48093 34940 48127
rect 34888 48084 34940 48093
rect 940 48016 992 48068
rect 31300 48059 31352 48068
rect 31300 48025 31309 48059
rect 31309 48025 31343 48059
rect 31343 48025 31352 48059
rect 31300 48016 31352 48025
rect 34796 48016 34848 48068
rect 35900 48084 35952 48136
rect 37188 48084 37240 48136
rect 41788 48084 41840 48136
rect 30840 47948 30892 48000
rect 31668 47991 31720 48000
rect 31668 47957 31677 47991
rect 31677 47957 31711 47991
rect 31711 47957 31720 47991
rect 31668 47948 31720 47957
rect 41604 48016 41656 48068
rect 57888 48127 57940 48136
rect 57888 48093 57897 48127
rect 57897 48093 57931 48127
rect 57931 48093 57940 48127
rect 57888 48084 57940 48093
rect 58992 48084 59044 48136
rect 59084 48016 59136 48068
rect 35440 47991 35492 48000
rect 35440 47957 35449 47991
rect 35449 47957 35483 47991
rect 35483 47957 35492 47991
rect 35440 47948 35492 47957
rect 35900 47948 35952 48000
rect 57336 47991 57388 48000
rect 57336 47957 57345 47991
rect 57345 47957 57379 47991
rect 57379 47957 57388 47991
rect 57336 47948 57388 47957
rect 19574 47846 19626 47898
rect 19638 47846 19690 47898
rect 19702 47846 19754 47898
rect 19766 47846 19818 47898
rect 19830 47846 19882 47898
rect 50294 47846 50346 47898
rect 50358 47846 50410 47898
rect 50422 47846 50474 47898
rect 50486 47846 50538 47898
rect 50550 47846 50602 47898
rect 34888 47744 34940 47796
rect 35348 47744 35400 47796
rect 40960 47719 41012 47728
rect 40960 47685 40969 47719
rect 40969 47685 41003 47719
rect 41003 47685 41012 47719
rect 40960 47676 41012 47685
rect 41604 47719 41656 47728
rect 41604 47685 41613 47719
rect 41613 47685 41647 47719
rect 41647 47685 41656 47719
rect 41604 47676 41656 47685
rect 41696 47719 41748 47728
rect 41696 47685 41705 47719
rect 41705 47685 41739 47719
rect 41739 47685 41748 47719
rect 41696 47676 41748 47685
rect 58440 47676 58492 47728
rect 1032 47608 1084 47660
rect 30380 47608 30432 47660
rect 30840 47651 30892 47660
rect 30840 47617 30850 47651
rect 30850 47617 30884 47651
rect 30884 47617 30892 47651
rect 30840 47608 30892 47617
rect 31024 47651 31076 47660
rect 31024 47617 31033 47651
rect 31033 47617 31067 47651
rect 31067 47617 31076 47651
rect 31024 47608 31076 47617
rect 31484 47608 31536 47660
rect 32956 47608 33008 47660
rect 33048 47608 33100 47660
rect 35440 47608 35492 47660
rect 41788 47651 41840 47660
rect 41788 47617 41802 47651
rect 41802 47617 41836 47651
rect 41836 47617 41840 47651
rect 41788 47608 41840 47617
rect 43076 47540 43128 47592
rect 58900 47608 58952 47660
rect 58992 47540 59044 47592
rect 14464 47404 14516 47456
rect 31392 47447 31444 47456
rect 31392 47413 31401 47447
rect 31401 47413 31435 47447
rect 31435 47413 31444 47447
rect 31392 47404 31444 47413
rect 42156 47404 42208 47456
rect 57428 47447 57480 47456
rect 57428 47413 57437 47447
rect 57437 47413 57471 47447
rect 57471 47413 57480 47447
rect 57428 47404 57480 47413
rect 58440 47404 58492 47456
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 58808 47132 58860 47184
rect 30472 46996 30524 47048
rect 31300 46996 31352 47048
rect 32680 46996 32732 47048
rect 35716 46996 35768 47048
rect 58992 46996 59044 47048
rect 940 46928 992 46980
rect 32312 46928 32364 46980
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 50294 46758 50346 46810
rect 50358 46758 50410 46810
rect 50422 46758 50474 46810
rect 50486 46758 50538 46810
rect 50550 46758 50602 46810
rect 1032 46520 1084 46572
rect 32312 46563 32364 46572
rect 32312 46529 32321 46563
rect 32321 46529 32355 46563
rect 32355 46529 32364 46563
rect 32312 46520 32364 46529
rect 31024 46452 31076 46504
rect 32680 46563 32732 46572
rect 32680 46529 32689 46563
rect 32689 46529 32723 46563
rect 32723 46529 32732 46563
rect 32680 46520 32732 46529
rect 58164 46563 58216 46572
rect 58164 46529 58173 46563
rect 58173 46529 58207 46563
rect 58207 46529 58216 46563
rect 58164 46520 58216 46529
rect 37924 46452 37976 46504
rect 50712 46452 50764 46504
rect 58532 46452 58584 46504
rect 35532 46384 35584 46436
rect 26976 46316 27028 46368
rect 32312 46316 32364 46368
rect 58256 46359 58308 46368
rect 58256 46325 58265 46359
rect 58265 46325 58299 46359
rect 58299 46325 58308 46359
rect 58256 46316 58308 46325
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 36912 46112 36964 46164
rect 940 45908 992 45960
rect 26976 45908 27028 45960
rect 36820 45951 36872 45960
rect 36820 45917 36829 45951
rect 36829 45917 36863 45951
rect 36863 45917 36872 45951
rect 36820 45908 36872 45917
rect 58992 45908 59044 45960
rect 35532 45840 35584 45892
rect 1768 45815 1820 45824
rect 1768 45781 1777 45815
rect 1777 45781 1811 45815
rect 1811 45781 1820 45815
rect 1768 45772 1820 45781
rect 38292 45840 38344 45892
rect 58072 45840 58124 45892
rect 48688 45772 48740 45824
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 50294 45670 50346 45722
rect 50358 45670 50410 45722
rect 50422 45670 50474 45722
rect 50486 45670 50538 45722
rect 50550 45670 50602 45722
rect 35532 45568 35584 45620
rect 29736 45500 29788 45552
rect 1032 45432 1084 45484
rect 32312 45475 32364 45484
rect 32312 45441 32321 45475
rect 32321 45441 32355 45475
rect 32355 45441 32364 45475
rect 32312 45432 32364 45441
rect 32404 45475 32456 45484
rect 32404 45441 32414 45475
rect 32414 45441 32448 45475
rect 32448 45441 32456 45475
rect 32404 45432 32456 45441
rect 32588 45475 32640 45484
rect 32588 45441 32597 45475
rect 32597 45441 32631 45475
rect 32631 45441 32640 45475
rect 32588 45432 32640 45441
rect 32680 45475 32732 45484
rect 32680 45441 32689 45475
rect 32689 45441 32723 45475
rect 32723 45441 32732 45475
rect 32680 45432 32732 45441
rect 1768 45364 1820 45416
rect 35624 45543 35676 45552
rect 35624 45509 35633 45543
rect 35633 45509 35667 45543
rect 35667 45509 35676 45543
rect 35624 45500 35676 45509
rect 35900 45500 35952 45552
rect 36820 45500 36872 45552
rect 35716 45475 35768 45484
rect 35716 45441 35725 45475
rect 35725 45441 35759 45475
rect 35759 45441 35768 45475
rect 35716 45432 35768 45441
rect 58164 45475 58216 45484
rect 58164 45441 58173 45475
rect 58173 45441 58207 45475
rect 58207 45441 58216 45475
rect 58164 45432 58216 45441
rect 58348 45432 58400 45484
rect 58532 45432 58584 45484
rect 32588 45296 32640 45348
rect 42340 45296 42392 45348
rect 7196 45228 7248 45280
rect 32772 45228 32824 45280
rect 36452 45228 36504 45280
rect 58256 45271 58308 45280
rect 58256 45237 58265 45271
rect 58265 45237 58299 45271
rect 58299 45237 58308 45271
rect 58256 45228 58308 45237
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 6736 45024 6788 45076
rect 32404 45024 32456 45076
rect 39396 44956 39448 45008
rect 940 44752 992 44804
rect 2136 44752 2188 44804
rect 58348 45024 58400 45076
rect 47216 44820 47268 44872
rect 57336 44956 57388 45008
rect 49332 44931 49384 44940
rect 49332 44897 49341 44931
rect 49341 44897 49375 44931
rect 49375 44897 49384 44931
rect 49332 44888 49384 44897
rect 58900 44888 58952 44940
rect 58992 44820 59044 44872
rect 48688 44727 48740 44736
rect 48688 44693 48697 44727
rect 48697 44693 48731 44727
rect 48731 44693 48740 44727
rect 48688 44684 48740 44693
rect 57336 44727 57388 44736
rect 57336 44693 57345 44727
rect 57345 44693 57379 44727
rect 57379 44693 57388 44727
rect 57336 44684 57388 44693
rect 59268 44752 59320 44804
rect 58716 44684 58768 44736
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 50294 44582 50346 44634
rect 50358 44582 50410 44634
rect 50422 44582 50474 44634
rect 50486 44582 50538 44634
rect 50550 44582 50602 44634
rect 41696 44412 41748 44464
rect 42616 44412 42668 44464
rect 1032 44344 1084 44396
rect 41420 44387 41472 44396
rect 41420 44353 41429 44387
rect 41429 44353 41463 44387
rect 41463 44353 41472 44387
rect 41420 44344 41472 44353
rect 49332 44344 49384 44396
rect 58992 44344 59044 44396
rect 26976 44140 27028 44192
rect 58256 44183 58308 44192
rect 58256 44149 58265 44183
rect 58265 44149 58299 44183
rect 58299 44149 58308 44183
rect 58256 44140 58308 44149
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 41328 43775 41380 43784
rect 41328 43741 41337 43775
rect 41337 43741 41371 43775
rect 41371 43741 41380 43775
rect 41328 43732 41380 43741
rect 41696 43775 41748 43784
rect 41696 43741 41705 43775
rect 41705 43741 41739 43775
rect 41739 43741 41748 43775
rect 41696 43732 41748 43741
rect 940 43664 992 43716
rect 2320 43664 2372 43716
rect 37004 43664 37056 43716
rect 37924 43596 37976 43648
rect 56140 43732 56192 43784
rect 58072 43775 58124 43784
rect 58072 43741 58081 43775
rect 58081 43741 58115 43775
rect 58115 43741 58124 43775
rect 58072 43732 58124 43741
rect 42892 43707 42944 43716
rect 42892 43673 42901 43707
rect 42901 43673 42935 43707
rect 42935 43673 42944 43707
rect 42892 43664 42944 43673
rect 47216 43664 47268 43716
rect 57336 43596 57388 43648
rect 58716 43596 58768 43648
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 50294 43494 50346 43546
rect 50358 43494 50410 43546
rect 50422 43494 50474 43546
rect 50486 43494 50538 43546
rect 50550 43494 50602 43546
rect 11704 43392 11756 43444
rect 26148 43392 26200 43444
rect 33784 43392 33836 43444
rect 42892 43392 42944 43444
rect 57888 43392 57940 43444
rect 58072 43392 58124 43444
rect 1032 43256 1084 43308
rect 58992 43256 59044 43308
rect 11704 43052 11756 43104
rect 59176 43052 59228 43104
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 58900 42644 58952 42696
rect 940 42576 992 42628
rect 27896 42508 27948 42560
rect 58900 42508 58952 42560
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 50294 42406 50346 42458
rect 50358 42406 50410 42458
rect 50422 42406 50474 42458
rect 50486 42406 50538 42458
rect 50550 42406 50602 42458
rect 31024 42304 31076 42356
rect 28080 42279 28132 42288
rect 28080 42245 28089 42279
rect 28089 42245 28123 42279
rect 28123 42245 28132 42279
rect 28080 42236 28132 42245
rect 28172 42279 28224 42288
rect 28172 42245 28181 42279
rect 28181 42245 28215 42279
rect 28215 42245 28224 42279
rect 28172 42236 28224 42245
rect 50896 42236 50948 42288
rect 58532 42236 58584 42288
rect 1032 42168 1084 42220
rect 27896 42211 27948 42220
rect 27896 42177 27905 42211
rect 27905 42177 27939 42211
rect 27939 42177 27948 42211
rect 27896 42168 27948 42177
rect 28264 42211 28316 42220
rect 28264 42177 28273 42211
rect 28273 42177 28307 42211
rect 28307 42177 28316 42211
rect 28264 42168 28316 42177
rect 30472 42168 30524 42220
rect 58348 42211 58400 42220
rect 58348 42177 58357 42211
rect 58357 42177 58391 42211
rect 58391 42177 58400 42211
rect 58348 42168 58400 42177
rect 37740 42100 37792 42152
rect 56048 42100 56100 42152
rect 14464 42032 14516 42084
rect 22744 42032 22796 42084
rect 33508 42032 33560 42084
rect 55956 42032 56008 42084
rect 26424 41964 26476 42016
rect 28540 41964 28592 42016
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 31852 41692 31904 41744
rect 940 41556 992 41608
rect 26424 41599 26476 41608
rect 26424 41565 26433 41599
rect 26433 41565 26467 41599
rect 26467 41565 26476 41599
rect 26424 41556 26476 41565
rect 26700 41599 26752 41608
rect 26700 41565 26709 41599
rect 26709 41565 26743 41599
rect 26743 41565 26752 41599
rect 26700 41556 26752 41565
rect 28264 41556 28316 41608
rect 28724 41556 28776 41608
rect 58992 41556 59044 41608
rect 28080 41488 28132 41540
rect 21272 41420 21324 41472
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 50294 41318 50346 41370
rect 50358 41318 50410 41370
rect 50422 41318 50474 41370
rect 50486 41318 50538 41370
rect 50550 41318 50602 41370
rect 1032 41080 1084 41132
rect 9220 40876 9272 40928
rect 58532 40876 58584 40928
rect 58808 40876 58860 40928
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 58808 40672 58860 40724
rect 59084 40672 59136 40724
rect 9128 40511 9180 40520
rect 9128 40477 9137 40511
rect 9137 40477 9171 40511
rect 9171 40477 9180 40511
rect 9128 40468 9180 40477
rect 9588 40511 9640 40520
rect 9588 40477 9591 40511
rect 9591 40477 9640 40511
rect 9588 40468 9640 40477
rect 31392 40511 31444 40520
rect 31392 40477 31401 40511
rect 31401 40477 31435 40511
rect 31435 40477 31444 40511
rect 31392 40468 31444 40477
rect 940 40400 992 40452
rect 9312 40443 9364 40452
rect 9312 40409 9321 40443
rect 9321 40409 9355 40443
rect 9355 40409 9364 40443
rect 9312 40400 9364 40409
rect 10140 40400 10192 40452
rect 40316 40511 40368 40520
rect 40316 40477 40325 40511
rect 40325 40477 40359 40511
rect 40359 40477 40368 40511
rect 40316 40468 40368 40477
rect 40592 40511 40644 40520
rect 40592 40477 40601 40511
rect 40601 40477 40635 40511
rect 40635 40477 40644 40511
rect 40592 40468 40644 40477
rect 43720 40400 43772 40452
rect 49148 40400 49200 40452
rect 31484 40375 31536 40384
rect 31484 40341 31493 40375
rect 31493 40341 31527 40375
rect 31527 40341 31536 40375
rect 31484 40332 31536 40341
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 50294 40230 50346 40282
rect 50358 40230 50410 40282
rect 50422 40230 50474 40282
rect 50486 40230 50538 40282
rect 50550 40230 50602 40282
rect 1032 40060 1084 40112
rect 58348 39899 58400 39908
rect 58348 39865 58357 39899
rect 58357 39865 58391 39899
rect 58391 39865 58400 39899
rect 58348 39856 58400 39865
rect 7656 39788 7708 39840
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 7932 39559 7984 39568
rect 7932 39525 7941 39559
rect 7941 39525 7975 39559
rect 7975 39525 7984 39559
rect 7932 39516 7984 39525
rect 7380 39423 7432 39432
rect 7380 39389 7389 39423
rect 7389 39389 7423 39423
rect 7423 39389 7432 39423
rect 7380 39380 7432 39389
rect 7656 39423 7708 39432
rect 7656 39389 7665 39423
rect 7665 39389 7699 39423
rect 7699 39389 7708 39423
rect 7656 39380 7708 39389
rect 7840 39423 7892 39432
rect 7840 39389 7843 39423
rect 7843 39389 7892 39423
rect 7840 39380 7892 39389
rect 9220 39380 9272 39432
rect 29552 39380 29604 39432
rect 940 39312 992 39364
rect 4896 39312 4948 39364
rect 9312 39312 9364 39364
rect 11704 39312 11756 39364
rect 29368 39312 29420 39364
rect 32680 39244 32732 39296
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 50294 39142 50346 39194
rect 50358 39142 50410 39194
rect 50422 39142 50474 39194
rect 50486 39142 50538 39194
rect 50550 39142 50602 39194
rect 55864 38972 55916 39024
rect 1032 38904 1084 38956
rect 32680 38947 32732 38956
rect 32680 38913 32689 38947
rect 32689 38913 32723 38947
rect 32723 38913 32732 38947
rect 32680 38904 32732 38913
rect 32864 38947 32916 38956
rect 32864 38913 32873 38947
rect 32873 38913 32907 38947
rect 32907 38913 32916 38947
rect 32864 38904 32916 38913
rect 33048 38947 33100 38956
rect 33048 38913 33057 38947
rect 33057 38913 33091 38947
rect 33091 38913 33100 38947
rect 33048 38904 33100 38913
rect 4988 38768 5040 38820
rect 29460 38700 29512 38752
rect 31484 38700 31536 38752
rect 33692 38700 33744 38752
rect 58348 38743 58400 38752
rect 58348 38709 58357 38743
rect 58357 38709 58391 38743
rect 58391 38709 58400 38743
rect 58348 38700 58400 38709
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 7840 38496 7892 38548
rect 9588 38496 9640 38548
rect 11428 38496 11480 38548
rect 5264 38471 5316 38480
rect 5264 38437 5273 38471
rect 5273 38437 5307 38471
rect 5307 38437 5316 38471
rect 5264 38428 5316 38437
rect 58164 38428 58216 38480
rect 58440 38428 58492 38480
rect 33048 38360 33100 38412
rect 4712 38335 4764 38344
rect 4712 38301 4721 38335
rect 4721 38301 4755 38335
rect 4755 38301 4764 38335
rect 4712 38292 4764 38301
rect 4896 38335 4948 38344
rect 4896 38301 4905 38335
rect 4905 38301 4939 38335
rect 4939 38301 4948 38335
rect 4896 38292 4948 38301
rect 4988 38335 5040 38344
rect 4988 38301 4997 38335
rect 4997 38301 5031 38335
rect 5031 38301 5040 38335
rect 4988 38292 5040 38301
rect 940 38224 992 38276
rect 3608 38224 3660 38276
rect 7840 38292 7892 38344
rect 21272 38292 21324 38344
rect 27160 38292 27212 38344
rect 33232 38292 33284 38344
rect 41420 38224 41472 38276
rect 32680 38156 32732 38208
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 50294 38054 50346 38106
rect 50358 38054 50410 38106
rect 50422 38054 50474 38106
rect 50486 38054 50538 38106
rect 50550 38054 50602 38106
rect 7196 37884 7248 37936
rect 30564 37884 30616 37936
rect 1032 37816 1084 37868
rect 32680 37859 32732 37868
rect 32680 37825 32689 37859
rect 32689 37825 32723 37859
rect 32723 37825 32732 37859
rect 32680 37816 32732 37825
rect 32864 37859 32916 37868
rect 32864 37825 32873 37859
rect 32873 37825 32907 37859
rect 32907 37825 32916 37859
rect 32864 37816 32916 37825
rect 33048 37859 33100 37868
rect 33048 37825 33062 37859
rect 33062 37825 33096 37859
rect 33096 37825 33100 37859
rect 53288 37884 53340 37936
rect 58072 37884 58124 37936
rect 33048 37816 33100 37825
rect 57520 37816 57572 37868
rect 3700 37680 3752 37732
rect 33600 37612 33652 37664
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 19432 37272 19484 37324
rect 57520 37204 57572 37256
rect 58992 37204 59044 37256
rect 940 37136 992 37188
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 50294 36966 50346 37018
rect 50358 36966 50410 37018
rect 50422 36966 50474 37018
rect 50486 36966 50538 37018
rect 50550 36966 50602 37018
rect 3424 36864 3476 36916
rect 1032 36728 1084 36780
rect 3148 36728 3200 36780
rect 3608 36771 3660 36780
rect 3608 36737 3617 36771
rect 3617 36737 3651 36771
rect 3651 36737 3660 36771
rect 3608 36728 3660 36737
rect 3700 36771 3752 36780
rect 3700 36737 3709 36771
rect 3709 36737 3743 36771
rect 3743 36737 3752 36771
rect 3700 36728 3752 36737
rect 3884 36728 3936 36780
rect 19340 36728 19392 36780
rect 58072 36771 58124 36780
rect 58072 36737 58081 36771
rect 58081 36737 58115 36771
rect 58115 36737 58124 36771
rect 58072 36728 58124 36737
rect 4620 36660 4672 36712
rect 4896 36660 4948 36712
rect 11428 36660 11480 36712
rect 21456 36703 21508 36712
rect 21456 36669 21465 36703
rect 21465 36669 21499 36703
rect 21499 36669 21508 36703
rect 21456 36660 21508 36669
rect 2044 36592 2096 36644
rect 31024 36592 31076 36644
rect 59544 36524 59596 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 58164 36227 58216 36236
rect 58164 36193 58173 36227
rect 58173 36193 58207 36227
rect 58207 36193 58216 36227
rect 58164 36184 58216 36193
rect 940 36116 992 36168
rect 19432 36116 19484 36168
rect 20168 36159 20220 36168
rect 20168 36125 20177 36159
rect 20177 36125 20211 36159
rect 20211 36125 20220 36159
rect 20168 36116 20220 36125
rect 27804 36116 27856 36168
rect 28356 36116 28408 36168
rect 30380 36159 30432 36168
rect 30380 36125 30389 36159
rect 30389 36125 30423 36159
rect 30423 36125 30432 36159
rect 30380 36116 30432 36125
rect 30656 36159 30708 36168
rect 30656 36125 30665 36159
rect 30665 36125 30699 36159
rect 30699 36125 30708 36159
rect 30656 36116 30708 36125
rect 31024 36159 31076 36168
rect 31024 36125 31033 36159
rect 31033 36125 31067 36159
rect 31067 36125 31076 36159
rect 31024 36116 31076 36125
rect 31392 36159 31444 36168
rect 31392 36125 31401 36159
rect 31401 36125 31435 36159
rect 31435 36125 31444 36159
rect 31392 36116 31444 36125
rect 55956 36116 56008 36168
rect 21456 36048 21508 36100
rect 31300 36048 31352 36100
rect 32864 36048 32916 36100
rect 3424 35980 3476 36032
rect 28632 35980 28684 36032
rect 30472 36023 30524 36032
rect 30472 35989 30481 36023
rect 30481 35989 30515 36023
rect 30515 35989 30524 36023
rect 30472 35980 30524 35989
rect 45008 35980 45060 36032
rect 46296 35980 46348 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 50294 35878 50346 35930
rect 50358 35878 50410 35930
rect 50422 35878 50474 35930
rect 50486 35878 50538 35930
rect 50550 35878 50602 35930
rect 3884 35776 3936 35828
rect 28264 35776 28316 35828
rect 33416 35776 33468 35828
rect 1032 35640 1084 35692
rect 57980 35708 58032 35760
rect 58164 35751 58216 35760
rect 58164 35717 58173 35751
rect 58173 35717 58207 35751
rect 58207 35717 58216 35751
rect 58164 35708 58216 35717
rect 2872 35683 2924 35692
rect 2872 35649 2881 35683
rect 2881 35649 2915 35683
rect 2915 35649 2924 35683
rect 2872 35640 2924 35649
rect 2964 35683 3016 35692
rect 2964 35649 2973 35683
rect 2973 35649 3007 35683
rect 3007 35649 3016 35683
rect 2964 35640 3016 35649
rect 4068 35640 4120 35692
rect 1952 35572 2004 35624
rect 28264 35683 28316 35692
rect 28264 35649 28273 35683
rect 28273 35649 28307 35683
rect 28307 35649 28316 35683
rect 28264 35640 28316 35649
rect 28448 35683 28500 35692
rect 28448 35649 28457 35683
rect 28457 35649 28491 35683
rect 28491 35649 28500 35683
rect 28448 35640 28500 35649
rect 28632 35640 28684 35692
rect 29092 35683 29144 35692
rect 29092 35649 29101 35683
rect 29101 35649 29135 35683
rect 29135 35649 29144 35683
rect 29092 35640 29144 35649
rect 30840 35640 30892 35692
rect 28724 35572 28776 35624
rect 33324 35683 33376 35692
rect 33324 35649 33333 35683
rect 33333 35649 33367 35683
rect 33367 35649 33376 35683
rect 33324 35640 33376 35649
rect 33416 35640 33468 35692
rect 33692 35640 33744 35692
rect 34796 35640 34848 35692
rect 33876 35572 33928 35624
rect 43720 35572 43772 35624
rect 41144 35504 41196 35556
rect 59728 35504 59780 35556
rect 23204 35436 23256 35488
rect 27988 35479 28040 35488
rect 27988 35445 27997 35479
rect 27997 35445 28031 35479
rect 28031 35445 28040 35479
rect 27988 35436 28040 35445
rect 28448 35436 28500 35488
rect 30104 35436 30156 35488
rect 33140 35436 33192 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 1768 35232 1820 35284
rect 26700 35232 26752 35284
rect 31392 35232 31444 35284
rect 29092 35164 29144 35216
rect 33876 35232 33928 35284
rect 57428 35164 57480 35216
rect 30564 35028 30616 35080
rect 30840 35071 30892 35080
rect 30840 35037 30849 35071
rect 30849 35037 30883 35071
rect 30883 35037 30892 35071
rect 30840 35028 30892 35037
rect 33232 35096 33284 35148
rect 33416 35096 33468 35148
rect 33692 35096 33744 35148
rect 58348 35096 58400 35148
rect 940 34960 992 35012
rect 28080 34960 28132 35012
rect 30748 35003 30800 35012
rect 30748 34969 30757 35003
rect 30757 34969 30791 35003
rect 30791 34969 30800 35003
rect 30748 34960 30800 34969
rect 31576 34960 31628 35012
rect 32036 35003 32088 35012
rect 32036 34969 32045 35003
rect 32045 34969 32079 35003
rect 32079 34969 32088 35003
rect 32036 34960 32088 34969
rect 32772 35028 32824 35080
rect 33140 35071 33192 35080
rect 33140 35037 33149 35071
rect 33149 35037 33183 35071
rect 33183 35037 33192 35071
rect 33140 35028 33192 35037
rect 42248 35071 42300 35080
rect 42248 35037 42257 35071
rect 42257 35037 42291 35071
rect 42291 35037 42300 35071
rect 42248 35028 42300 35037
rect 42800 35028 42852 35080
rect 43260 35028 43312 35080
rect 57612 35028 57664 35080
rect 32956 34960 33008 35012
rect 58164 35003 58216 35012
rect 58164 34969 58173 35003
rect 58173 34969 58207 35003
rect 58207 34969 58216 35003
rect 58164 34960 58216 34969
rect 59084 34960 59136 35012
rect 59360 34960 59412 35012
rect 32220 34892 32272 34944
rect 32772 34892 32824 34944
rect 33416 34892 33468 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 50294 34790 50346 34842
rect 50358 34790 50410 34842
rect 50422 34790 50474 34842
rect 50486 34790 50538 34842
rect 50550 34790 50602 34842
rect 1768 34731 1820 34740
rect 1768 34697 1777 34731
rect 1777 34697 1811 34731
rect 1811 34697 1820 34731
rect 1768 34688 1820 34697
rect 10140 34688 10192 34740
rect 24400 34688 24452 34740
rect 5264 34620 5316 34672
rect 34060 34688 34112 34740
rect 41144 34731 41196 34740
rect 41144 34697 41153 34731
rect 41153 34697 41187 34731
rect 41187 34697 41196 34731
rect 41144 34688 41196 34697
rect 1032 34552 1084 34604
rect 24308 34595 24360 34604
rect 24308 34561 24317 34595
rect 24317 34561 24351 34595
rect 24351 34561 24360 34595
rect 24308 34552 24360 34561
rect 24584 34552 24636 34604
rect 32404 34552 32456 34604
rect 32496 34595 32548 34604
rect 32496 34561 32505 34595
rect 32505 34561 32539 34595
rect 32539 34561 32548 34595
rect 32496 34552 32548 34561
rect 33692 34620 33744 34672
rect 37556 34620 37608 34672
rect 32772 34595 32824 34604
rect 32772 34561 32781 34595
rect 32781 34561 32815 34595
rect 32815 34561 32824 34595
rect 32772 34552 32824 34561
rect 26700 34484 26752 34536
rect 32956 34595 33008 34604
rect 32956 34561 32970 34595
rect 32970 34561 33004 34595
rect 33004 34561 33008 34595
rect 32956 34552 33008 34561
rect 34704 34552 34756 34604
rect 42800 34688 42852 34740
rect 59084 34688 59136 34740
rect 42432 34620 42484 34672
rect 42800 34552 42852 34604
rect 43628 34595 43680 34604
rect 43628 34561 43637 34595
rect 43637 34561 43671 34595
rect 43671 34561 43680 34595
rect 43628 34552 43680 34561
rect 43720 34595 43772 34604
rect 43720 34561 43729 34595
rect 43729 34561 43763 34595
rect 43763 34561 43772 34595
rect 43720 34552 43772 34561
rect 58072 34595 58124 34604
rect 58072 34561 58081 34595
rect 58081 34561 58115 34595
rect 58115 34561 58124 34595
rect 58072 34552 58124 34561
rect 34336 34527 34388 34536
rect 34336 34493 34345 34527
rect 34345 34493 34379 34527
rect 34379 34493 34388 34527
rect 34336 34484 34388 34493
rect 41696 34484 41748 34536
rect 34060 34459 34112 34468
rect 34060 34425 34069 34459
rect 34069 34425 34103 34459
rect 34103 34425 34112 34459
rect 34060 34416 34112 34425
rect 42984 34348 43036 34400
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 34704 34144 34756 34196
rect 4068 34076 4120 34128
rect 3976 33983 4028 33992
rect 3976 33949 3985 33983
rect 3985 33949 4019 33983
rect 4019 33949 4028 33983
rect 3976 33940 4028 33949
rect 58532 34144 58584 34196
rect 42800 34119 42852 34128
rect 42800 34085 42809 34119
rect 42809 34085 42843 34119
rect 42843 34085 42852 34119
rect 42800 34076 42852 34085
rect 39948 34008 40000 34060
rect 42708 34008 42760 34060
rect 940 33872 992 33924
rect 4620 33872 4672 33924
rect 32772 33872 32824 33924
rect 33784 33872 33836 33924
rect 34796 33940 34848 33992
rect 43076 33983 43128 33992
rect 43076 33949 43085 33983
rect 43085 33949 43119 33983
rect 43119 33949 43128 33983
rect 43076 33940 43128 33949
rect 43168 33940 43220 33992
rect 47952 34051 48004 34060
rect 47952 34017 47961 34051
rect 47961 34017 47995 34051
rect 47995 34017 48004 34051
rect 47952 34008 48004 34017
rect 47676 33940 47728 33992
rect 49056 34008 49108 34060
rect 46020 33872 46072 33924
rect 56692 33940 56744 33992
rect 58164 33915 58216 33924
rect 58164 33881 58173 33915
rect 58173 33881 58207 33915
rect 58207 33881 58216 33915
rect 58164 33872 58216 33881
rect 33968 33847 34020 33856
rect 33968 33813 33983 33847
rect 33983 33813 34017 33847
rect 34017 33813 34020 33847
rect 33968 33804 34020 33813
rect 47860 33804 47912 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 50294 33702 50346 33754
rect 50358 33702 50410 33754
rect 50422 33702 50474 33754
rect 50486 33702 50538 33754
rect 50550 33702 50602 33754
rect 33232 33643 33284 33652
rect 33232 33609 33241 33643
rect 33241 33609 33275 33643
rect 33275 33609 33284 33643
rect 33232 33600 33284 33609
rect 2964 33532 3016 33584
rect 33968 33532 34020 33584
rect 1032 33464 1084 33516
rect 30104 33464 30156 33516
rect 33140 33464 33192 33516
rect 33600 33507 33652 33516
rect 33600 33473 33609 33507
rect 33609 33473 33643 33507
rect 33643 33473 33652 33507
rect 33600 33464 33652 33473
rect 58072 33507 58124 33516
rect 58072 33473 58081 33507
rect 58081 33473 58115 33507
rect 58115 33473 58124 33507
rect 58072 33464 58124 33473
rect 37096 33396 37148 33448
rect 50988 33260 51040 33312
rect 51448 33260 51500 33312
rect 59636 33260 59688 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 1952 33056 2004 33108
rect 2412 33056 2464 33108
rect 29736 33056 29788 33108
rect 30196 33056 30248 33108
rect 50804 33056 50856 33108
rect 57244 33056 57296 33108
rect 2228 32920 2280 32972
rect 2412 32920 2464 32972
rect 23020 32920 23072 32972
rect 29828 32920 29880 32972
rect 28264 32852 28316 32904
rect 42248 32852 42300 32904
rect 49884 32852 49936 32904
rect 940 32784 992 32836
rect 27712 32784 27764 32836
rect 28080 32784 28132 32836
rect 58164 32827 58216 32836
rect 58164 32793 58173 32827
rect 58173 32793 58207 32827
rect 58207 32793 58216 32827
rect 58164 32784 58216 32793
rect 2320 32716 2372 32768
rect 3424 32716 3476 32768
rect 59268 32716 59320 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 50294 32614 50346 32666
rect 50358 32614 50410 32666
rect 50422 32614 50474 32666
rect 50486 32614 50538 32666
rect 50550 32614 50602 32666
rect 2412 32512 2464 32564
rect 2872 32512 2924 32564
rect 3240 32512 3292 32564
rect 2320 32487 2372 32496
rect 2320 32453 2329 32487
rect 2329 32453 2363 32487
rect 2363 32453 2372 32487
rect 2320 32444 2372 32453
rect 28172 32512 28224 32564
rect 46480 32512 46532 32564
rect 19984 32444 20036 32496
rect 2136 32376 2188 32428
rect 2504 32376 2556 32428
rect 3332 32419 3384 32428
rect 3332 32385 3341 32419
rect 3341 32385 3375 32419
rect 3375 32385 3384 32419
rect 3332 32376 3384 32385
rect 3424 32419 3476 32428
rect 3424 32385 3434 32419
rect 3434 32385 3468 32419
rect 3468 32385 3476 32419
rect 3424 32376 3476 32385
rect 3700 32419 3752 32428
rect 3700 32385 3709 32419
rect 3709 32385 3743 32419
rect 3743 32385 3752 32419
rect 3700 32376 3752 32385
rect 4068 32376 4120 32428
rect 11796 32376 11848 32428
rect 27896 32419 27948 32428
rect 27896 32385 27905 32419
rect 27905 32385 27939 32419
rect 27939 32385 27948 32419
rect 27896 32376 27948 32385
rect 27620 32308 27672 32360
rect 28448 32376 28500 32428
rect 31484 32444 31536 32496
rect 2596 32215 2648 32224
rect 2596 32181 2605 32215
rect 2605 32181 2639 32215
rect 2639 32181 2648 32215
rect 2596 32172 2648 32181
rect 28080 32240 28132 32292
rect 29552 32351 29604 32360
rect 29552 32317 29561 32351
rect 29561 32317 29595 32351
rect 29595 32317 29604 32351
rect 29552 32308 29604 32317
rect 29828 32308 29880 32360
rect 43076 32444 43128 32496
rect 54576 32444 54628 32496
rect 39948 32376 40000 32428
rect 52828 32376 52880 32428
rect 58072 32419 58124 32428
rect 58072 32385 58081 32419
rect 58081 32385 58115 32419
rect 58115 32385 58124 32419
rect 58072 32376 58124 32385
rect 28632 32172 28684 32224
rect 30196 32172 30248 32224
rect 37832 32215 37884 32224
rect 37832 32181 37841 32215
rect 37841 32181 37875 32215
rect 37875 32181 37884 32215
rect 37832 32172 37884 32181
rect 57980 32172 58032 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 27620 31968 27672 32020
rect 27896 31968 27948 32020
rect 37096 32011 37148 32020
rect 37096 31977 37105 32011
rect 37105 31977 37139 32011
rect 37139 31977 37148 32011
rect 37096 31968 37148 31977
rect 37832 31968 37884 32020
rect 47768 31968 47820 32020
rect 3700 31900 3752 31952
rect 1032 31832 1084 31884
rect 940 31764 992 31816
rect 26976 31832 27028 31884
rect 27712 31764 27764 31816
rect 28172 31832 28224 31884
rect 54484 31900 54536 31952
rect 28080 31764 28132 31816
rect 30840 31764 30892 31816
rect 36452 31807 36504 31816
rect 36452 31773 36461 31807
rect 36461 31773 36495 31807
rect 36495 31773 36504 31807
rect 36452 31764 36504 31773
rect 36636 31807 36688 31816
rect 36636 31773 36643 31807
rect 36643 31773 36688 31807
rect 36636 31764 36688 31773
rect 36820 31807 36872 31816
rect 36820 31773 36829 31807
rect 36829 31773 36863 31807
rect 36863 31773 36872 31807
rect 36820 31764 36872 31773
rect 37004 31764 37056 31816
rect 57060 31764 57112 31816
rect 58900 31832 58952 31884
rect 58992 31764 59044 31816
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 50294 31526 50346 31578
rect 50358 31526 50410 31578
rect 50422 31526 50474 31578
rect 50486 31526 50538 31578
rect 50550 31526 50602 31578
rect 3332 31424 3384 31476
rect 58440 31356 58492 31408
rect 2044 31331 2096 31340
rect 2044 31297 2053 31331
rect 2053 31297 2087 31331
rect 2087 31297 2096 31331
rect 2044 31288 2096 31297
rect 2320 31331 2372 31340
rect 2320 31297 2329 31331
rect 2329 31297 2363 31331
rect 2363 31297 2372 31331
rect 2320 31288 2372 31297
rect 2688 31288 2740 31340
rect 48136 31288 48188 31340
rect 48320 31331 48372 31340
rect 48320 31297 48329 31331
rect 48329 31297 48363 31331
rect 48363 31297 48372 31331
rect 48320 31288 48372 31297
rect 58072 31331 58124 31340
rect 58072 31297 58081 31331
rect 58081 31297 58115 31331
rect 58115 31297 58124 31331
rect 58072 31288 58124 31297
rect 19432 31220 19484 31272
rect 45560 31084 45612 31136
rect 58256 31127 58308 31136
rect 58256 31093 58265 31127
rect 58265 31093 58299 31127
rect 58299 31093 58308 31127
rect 58256 31084 58308 31093
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 27620 30880 27672 30932
rect 30748 30880 30800 30932
rect 48136 30923 48188 30932
rect 48136 30889 48145 30923
rect 48145 30889 48179 30923
rect 48179 30889 48188 30923
rect 48136 30880 48188 30889
rect 940 30676 992 30728
rect 26240 30676 26292 30728
rect 29920 30812 29972 30864
rect 43904 30812 43956 30864
rect 58256 30880 58308 30932
rect 29368 30744 29420 30796
rect 28724 30719 28776 30728
rect 28724 30685 28738 30719
rect 28738 30685 28772 30719
rect 28772 30685 28776 30719
rect 28724 30676 28776 30685
rect 29644 30676 29696 30728
rect 41420 30744 41472 30796
rect 30288 30676 30340 30728
rect 46572 30676 46624 30728
rect 47584 30719 47636 30728
rect 47584 30685 47593 30719
rect 47593 30685 47627 30719
rect 47627 30685 47636 30719
rect 47584 30676 47636 30685
rect 47768 30719 47820 30728
rect 47768 30685 47777 30719
rect 47777 30685 47811 30719
rect 47811 30685 47820 30719
rect 47768 30676 47820 30685
rect 28172 30608 28224 30660
rect 28632 30651 28684 30660
rect 28632 30617 28641 30651
rect 28641 30617 28675 30651
rect 28675 30617 28684 30651
rect 28632 30608 28684 30617
rect 1768 30583 1820 30592
rect 1768 30549 1777 30583
rect 1777 30549 1811 30583
rect 1811 30549 1820 30583
rect 1768 30540 1820 30549
rect 27712 30540 27764 30592
rect 29736 30540 29788 30592
rect 30380 30583 30432 30592
rect 30380 30549 30389 30583
rect 30389 30549 30423 30583
rect 30423 30549 30432 30583
rect 30380 30540 30432 30549
rect 32128 30651 32180 30660
rect 32128 30617 32137 30651
rect 32137 30617 32171 30651
rect 32171 30617 32180 30651
rect 32128 30608 32180 30617
rect 36544 30540 36596 30592
rect 58624 30676 58676 30728
rect 58164 30651 58216 30660
rect 58164 30617 58173 30651
rect 58173 30617 58207 30651
rect 58207 30617 58216 30651
rect 58164 30608 58216 30617
rect 48688 30540 48740 30592
rect 56324 30540 56376 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 50294 30438 50346 30490
rect 50358 30438 50410 30490
rect 50422 30438 50474 30490
rect 50486 30438 50538 30490
rect 50550 30438 50602 30490
rect 1768 30336 1820 30388
rect 28632 30336 28684 30388
rect 29644 30336 29696 30388
rect 30104 30336 30156 30388
rect 30840 30336 30892 30388
rect 940 30268 992 30320
rect 2596 30243 2648 30252
rect 2596 30209 2605 30243
rect 2605 30209 2639 30243
rect 2639 30209 2648 30243
rect 2596 30200 2648 30209
rect 2688 30200 2740 30252
rect 13820 30200 13872 30252
rect 17132 30311 17184 30320
rect 17132 30277 17141 30311
rect 17141 30277 17175 30311
rect 17175 30277 17184 30311
rect 17132 30268 17184 30277
rect 22836 30311 22888 30320
rect 22836 30277 22845 30311
rect 22845 30277 22879 30311
rect 22879 30277 22888 30311
rect 22836 30268 22888 30277
rect 29736 30268 29788 30320
rect 17224 30243 17276 30252
rect 17224 30209 17233 30243
rect 17233 30209 17267 30243
rect 17267 30209 17276 30243
rect 17224 30200 17276 30209
rect 22468 30200 22520 30252
rect 22928 30243 22980 30252
rect 22928 30209 22937 30243
rect 22937 30209 22971 30243
rect 22971 30209 22980 30243
rect 22928 30200 22980 30209
rect 23112 30200 23164 30252
rect 23204 30243 23256 30252
rect 23204 30209 23213 30243
rect 23213 30209 23247 30243
rect 23247 30209 23256 30243
rect 23204 30200 23256 30209
rect 23296 30200 23348 30252
rect 24216 30200 24268 30252
rect 28724 30200 28776 30252
rect 22376 30132 22428 30184
rect 26240 30132 26292 30184
rect 30012 30132 30064 30184
rect 30380 30243 30432 30252
rect 30380 30209 30389 30243
rect 30389 30209 30423 30243
rect 30423 30209 30432 30243
rect 30380 30200 30432 30209
rect 48228 30268 48280 30320
rect 53196 30268 53248 30320
rect 31208 30243 31260 30252
rect 31208 30209 31217 30243
rect 31217 30209 31251 30243
rect 31251 30209 31260 30243
rect 31208 30200 31260 30209
rect 32128 30200 32180 30252
rect 36820 30200 36872 30252
rect 47584 30200 47636 30252
rect 52736 30200 52788 30252
rect 58072 30243 58124 30252
rect 58072 30209 58081 30243
rect 58081 30209 58115 30243
rect 58115 30209 58124 30243
rect 58072 30200 58124 30209
rect 22284 29996 22336 30048
rect 22836 29996 22888 30048
rect 23756 29996 23808 30048
rect 28172 29996 28224 30048
rect 28356 29996 28408 30048
rect 30564 29996 30616 30048
rect 45560 30064 45612 30116
rect 32588 29996 32640 30048
rect 41880 29996 41932 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 2320 29724 2372 29776
rect 7932 29724 7984 29776
rect 27988 29724 28040 29776
rect 30380 29724 30432 29776
rect 32588 29767 32640 29776
rect 32588 29733 32597 29767
rect 32597 29733 32631 29767
rect 32631 29733 32640 29767
rect 32588 29724 32640 29733
rect 33324 29724 33376 29776
rect 940 29588 992 29640
rect 1032 29520 1084 29572
rect 11796 29520 11848 29572
rect 23112 29656 23164 29708
rect 23296 29588 23348 29640
rect 31392 29656 31444 29708
rect 33968 29656 34020 29708
rect 36636 29724 36688 29776
rect 51540 29724 51592 29776
rect 49700 29656 49752 29708
rect 58164 29699 58216 29708
rect 58164 29665 58173 29699
rect 58173 29665 58207 29699
rect 58207 29665 58216 29699
rect 58164 29656 58216 29665
rect 28448 29631 28500 29640
rect 28448 29597 28457 29631
rect 28457 29597 28491 29631
rect 28491 29597 28500 29631
rect 28448 29588 28500 29597
rect 28724 29631 28776 29640
rect 28724 29597 28733 29631
rect 28733 29597 28767 29631
rect 28767 29597 28776 29631
rect 28724 29588 28776 29597
rect 29736 29631 29788 29640
rect 29736 29597 29745 29631
rect 29745 29597 29779 29631
rect 29779 29597 29788 29631
rect 29736 29588 29788 29597
rect 30012 29631 30064 29640
rect 30012 29597 30021 29631
rect 30021 29597 30055 29631
rect 30055 29597 30064 29631
rect 30012 29588 30064 29597
rect 32588 29588 32640 29640
rect 29184 29563 29236 29572
rect 29184 29529 29193 29563
rect 29193 29529 29227 29563
rect 29227 29529 29236 29563
rect 29184 29520 29236 29529
rect 2320 29452 2372 29504
rect 13912 29452 13964 29504
rect 15016 29452 15068 29504
rect 28632 29452 28684 29504
rect 30196 29495 30248 29504
rect 30196 29461 30205 29495
rect 30205 29461 30239 29495
rect 30239 29461 30248 29495
rect 30196 29452 30248 29461
rect 30564 29520 30616 29572
rect 57704 29588 57756 29640
rect 32036 29452 32088 29504
rect 39304 29452 39356 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 50294 29350 50346 29402
rect 50358 29350 50410 29402
rect 50422 29350 50474 29402
rect 50486 29350 50538 29402
rect 50550 29350 50602 29402
rect 2412 29248 2464 29300
rect 22284 29248 22336 29300
rect 22468 29291 22520 29300
rect 22468 29257 22477 29291
rect 22477 29257 22511 29291
rect 22511 29257 22520 29291
rect 22468 29248 22520 29257
rect 22744 29291 22796 29300
rect 22744 29257 22753 29291
rect 22753 29257 22787 29291
rect 22787 29257 22796 29291
rect 22744 29248 22796 29257
rect 22928 29248 22980 29300
rect 23388 29248 23440 29300
rect 2320 29223 2372 29232
rect 2320 29189 2329 29223
rect 2329 29189 2363 29223
rect 2363 29189 2372 29223
rect 2320 29180 2372 29189
rect 2136 29112 2188 29164
rect 2688 29112 2740 29164
rect 22744 29112 22796 29164
rect 23204 29155 23256 29164
rect 23204 29121 23213 29155
rect 23213 29121 23247 29155
rect 23247 29121 23256 29155
rect 23204 29112 23256 29121
rect 28908 29248 28960 29300
rect 23572 29180 23624 29232
rect 23756 29155 23808 29164
rect 23756 29121 23765 29155
rect 23765 29121 23799 29155
rect 23799 29121 23808 29155
rect 23756 29112 23808 29121
rect 3240 29044 3292 29096
rect 13912 29044 13964 29096
rect 2136 28976 2188 29028
rect 24952 29044 25004 29096
rect 28632 29155 28684 29164
rect 28632 29121 28641 29155
rect 28641 29121 28675 29155
rect 28675 29121 28684 29155
rect 28632 29112 28684 29121
rect 28724 29155 28776 29164
rect 28724 29121 28733 29155
rect 28733 29121 28767 29155
rect 28767 29121 28776 29155
rect 28724 29112 28776 29121
rect 28816 29155 28868 29164
rect 28816 29121 28825 29155
rect 28825 29121 28859 29155
rect 28859 29121 28868 29155
rect 28816 29112 28868 29121
rect 29644 29155 29696 29164
rect 29644 29121 29653 29155
rect 29653 29121 29687 29155
rect 29687 29121 29696 29155
rect 29644 29112 29696 29121
rect 31024 29112 31076 29164
rect 31668 29044 31720 29096
rect 58348 29180 58400 29232
rect 58072 29155 58124 29164
rect 58072 29121 58081 29155
rect 58081 29121 58115 29155
rect 58115 29121 58124 29155
rect 58072 29112 58124 29121
rect 58440 28976 58492 29028
rect 24492 28908 24544 28960
rect 29000 28951 29052 28960
rect 29000 28917 29009 28951
rect 29009 28917 29043 28951
rect 29043 28917 29052 28951
rect 29000 28908 29052 28917
rect 30932 28908 30984 28960
rect 31760 28951 31812 28960
rect 31760 28917 31769 28951
rect 31769 28917 31803 28951
rect 31803 28917 31812 28951
rect 31760 28908 31812 28917
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 28448 28704 28500 28756
rect 28816 28704 28868 28756
rect 29000 28704 29052 28756
rect 24308 28636 24360 28688
rect 30380 28636 30432 28688
rect 19432 28568 19484 28620
rect 23664 28568 23716 28620
rect 25504 28568 25556 28620
rect 940 28500 992 28552
rect 23296 28500 23348 28552
rect 23388 28432 23440 28484
rect 23756 28500 23808 28552
rect 24584 28500 24636 28552
rect 25872 28500 25924 28552
rect 28540 28500 28592 28552
rect 28816 28543 28868 28552
rect 28816 28509 28825 28543
rect 28825 28509 28859 28543
rect 28859 28509 28868 28543
rect 28816 28500 28868 28509
rect 30472 28568 30524 28620
rect 37004 28704 37056 28756
rect 31760 28636 31812 28688
rect 28724 28432 28776 28484
rect 30012 28432 30064 28484
rect 37924 28500 37976 28552
rect 42156 28500 42208 28552
rect 52184 28568 52236 28620
rect 58164 28611 58216 28620
rect 58164 28577 58173 28611
rect 58173 28577 58207 28611
rect 58207 28577 58216 28611
rect 58164 28568 58216 28577
rect 30288 28432 30340 28484
rect 41696 28432 41748 28484
rect 42064 28432 42116 28484
rect 13820 28364 13872 28416
rect 25412 28364 25464 28416
rect 27988 28364 28040 28416
rect 31576 28364 31628 28416
rect 31944 28364 31996 28416
rect 41236 28364 41288 28416
rect 49240 28500 49292 28552
rect 56600 28500 56652 28552
rect 48688 28475 48740 28484
rect 48688 28441 48697 28475
rect 48697 28441 48731 28475
rect 48731 28441 48740 28475
rect 48688 28432 48740 28441
rect 50712 28432 50764 28484
rect 48872 28364 48924 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 50294 28262 50346 28314
rect 50358 28262 50410 28314
rect 50422 28262 50474 28314
rect 50486 28262 50538 28314
rect 50550 28262 50602 28314
rect 18972 28160 19024 28212
rect 22284 28160 22336 28212
rect 22468 28160 22520 28212
rect 24308 28203 24360 28212
rect 24308 28169 24317 28203
rect 24317 28169 24351 28203
rect 24351 28169 24360 28203
rect 24308 28160 24360 28169
rect 28724 28160 28776 28212
rect 28816 28160 28868 28212
rect 30104 28160 30156 28212
rect 940 28092 992 28144
rect 15384 28092 15436 28144
rect 23296 28024 23348 28076
rect 23388 28067 23440 28076
rect 23388 28033 23397 28067
rect 23397 28033 23431 28067
rect 23431 28033 23440 28067
rect 23388 28024 23440 28033
rect 23756 28067 23808 28076
rect 23756 28033 23765 28067
rect 23765 28033 23799 28067
rect 23799 28033 23808 28067
rect 23756 28024 23808 28033
rect 24492 28067 24544 28076
rect 24492 28033 24501 28067
rect 24501 28033 24535 28067
rect 24535 28033 24544 28067
rect 24492 28024 24544 28033
rect 24952 28024 25004 28076
rect 25504 28067 25556 28076
rect 25504 28033 25513 28067
rect 25513 28033 25547 28067
rect 25547 28033 25556 28067
rect 25504 28024 25556 28033
rect 25596 28067 25648 28076
rect 25596 28033 25605 28067
rect 25605 28033 25639 28067
rect 25639 28033 25648 28067
rect 25596 28024 25648 28033
rect 25872 28024 25924 28076
rect 28540 28067 28592 28076
rect 28540 28033 28549 28067
rect 28549 28033 28583 28067
rect 28583 28033 28592 28067
rect 28540 28024 28592 28033
rect 22284 27956 22336 28008
rect 25044 27888 25096 27940
rect 26056 27931 26108 27940
rect 26056 27897 26065 27931
rect 26065 27897 26099 27931
rect 26099 27897 26108 27931
rect 26056 27888 26108 27897
rect 27344 27999 27396 28008
rect 27344 27965 27353 27999
rect 27353 27965 27387 27999
rect 27387 27965 27396 27999
rect 27344 27956 27396 27965
rect 27528 27956 27580 28008
rect 28908 28067 28960 28076
rect 28908 28033 28917 28067
rect 28917 28033 28951 28067
rect 28951 28033 28960 28067
rect 28908 28024 28960 28033
rect 29000 27956 29052 28008
rect 29368 28024 29420 28076
rect 30012 28024 30064 28076
rect 30472 28024 30524 28076
rect 31484 28160 31536 28212
rect 28632 27820 28684 27872
rect 29000 27820 29052 27872
rect 30288 27956 30340 28008
rect 31116 27956 31168 28008
rect 48320 28092 48372 28144
rect 58716 28092 58768 28144
rect 58072 28067 58124 28076
rect 58072 28033 58081 28067
rect 58081 28033 58115 28067
rect 58115 28033 58124 28067
rect 58072 28024 58124 28033
rect 42616 27820 42668 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 22376 27616 22428 27668
rect 23664 27548 23716 27600
rect 26332 27548 26384 27600
rect 23020 27480 23072 27532
rect 940 27412 992 27464
rect 22100 27412 22152 27464
rect 23296 27412 23348 27464
rect 23572 27455 23624 27464
rect 23572 27421 23581 27455
rect 23581 27421 23615 27455
rect 23615 27421 23624 27455
rect 23572 27412 23624 27421
rect 23664 27412 23716 27464
rect 24952 27412 25004 27464
rect 25228 27412 25280 27464
rect 25412 27455 25464 27464
rect 25412 27421 25421 27455
rect 25421 27421 25455 27455
rect 25455 27421 25464 27455
rect 25412 27412 25464 27421
rect 25504 27412 25556 27464
rect 27344 27548 27396 27600
rect 26976 27455 27028 27464
rect 26976 27421 26985 27455
rect 26985 27421 27019 27455
rect 27019 27421 27028 27455
rect 26976 27412 27028 27421
rect 27068 27455 27120 27464
rect 27068 27421 27077 27455
rect 27077 27421 27111 27455
rect 27111 27421 27120 27455
rect 27068 27412 27120 27421
rect 27712 27455 27764 27464
rect 27712 27421 27721 27455
rect 27721 27421 27755 27455
rect 27755 27421 27764 27455
rect 27712 27412 27764 27421
rect 28448 27616 28500 27668
rect 30104 27548 30156 27600
rect 30472 27616 30524 27668
rect 30380 27548 30432 27600
rect 33140 27616 33192 27668
rect 34152 27616 34204 27668
rect 31668 27548 31720 27600
rect 28632 27480 28684 27532
rect 33784 27480 33836 27532
rect 45468 27548 45520 27600
rect 48964 27480 49016 27532
rect 18972 27276 19024 27328
rect 25596 27344 25648 27396
rect 26240 27344 26292 27396
rect 23756 27276 23808 27328
rect 24860 27276 24912 27328
rect 26056 27276 26108 27328
rect 26332 27276 26384 27328
rect 26516 27276 26568 27328
rect 26608 27276 26660 27328
rect 28448 27412 28500 27464
rect 30656 27455 30708 27464
rect 30656 27421 30665 27455
rect 30665 27421 30699 27455
rect 30699 27421 30708 27455
rect 30656 27412 30708 27421
rect 30932 27412 30984 27464
rect 32220 27455 32272 27464
rect 32220 27421 32229 27455
rect 32229 27421 32263 27455
rect 32263 27421 32272 27455
rect 32220 27412 32272 27421
rect 32312 27455 32364 27464
rect 32312 27421 32321 27455
rect 32321 27421 32355 27455
rect 32355 27421 32364 27455
rect 32312 27412 32364 27421
rect 27896 27387 27948 27396
rect 27896 27353 27905 27387
rect 27905 27353 27939 27387
rect 27939 27353 27948 27387
rect 27896 27344 27948 27353
rect 33508 27455 33560 27464
rect 33508 27421 33517 27455
rect 33517 27421 33551 27455
rect 33551 27421 33560 27455
rect 33508 27412 33560 27421
rect 33968 27455 34020 27464
rect 33968 27421 33977 27455
rect 33977 27421 34011 27455
rect 34011 27421 34020 27455
rect 33968 27412 34020 27421
rect 51356 27480 51408 27532
rect 58992 27480 59044 27532
rect 49424 27455 49476 27464
rect 49424 27421 49438 27455
rect 49438 27421 49472 27455
rect 49472 27421 49476 27455
rect 49424 27412 49476 27421
rect 56876 27412 56928 27464
rect 35348 27344 35400 27396
rect 48688 27344 48740 27396
rect 50896 27344 50948 27396
rect 28172 27276 28224 27328
rect 28448 27276 28500 27328
rect 33600 27276 33652 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 50294 27174 50346 27226
rect 50358 27174 50410 27226
rect 50422 27174 50474 27226
rect 50486 27174 50538 27226
rect 50550 27174 50602 27226
rect 23572 27072 23624 27124
rect 25044 27072 25096 27124
rect 25320 27072 25372 27124
rect 26056 27115 26108 27124
rect 26056 27081 26065 27115
rect 26065 27081 26099 27115
rect 26099 27081 26108 27115
rect 26056 27072 26108 27081
rect 26240 27115 26292 27124
rect 26240 27081 26249 27115
rect 26249 27081 26283 27115
rect 26283 27081 26292 27115
rect 26240 27072 26292 27081
rect 26332 27115 26384 27124
rect 26332 27081 26341 27115
rect 26341 27081 26375 27115
rect 26375 27081 26384 27115
rect 26332 27072 26384 27081
rect 26424 27072 26476 27124
rect 30656 27072 30708 27124
rect 31024 27115 31076 27124
rect 31024 27081 31033 27115
rect 31033 27081 31067 27115
rect 31067 27081 31076 27115
rect 31024 27072 31076 27081
rect 940 27004 992 27056
rect 1860 27004 1912 27056
rect 25504 27004 25556 27056
rect 26148 27047 26200 27056
rect 26148 27013 26157 27047
rect 26157 27013 26191 27047
rect 26191 27013 26200 27047
rect 26148 27004 26200 27013
rect 1032 26936 1084 26988
rect 23020 26979 23072 26988
rect 23020 26945 23029 26979
rect 23029 26945 23063 26979
rect 23063 26945 23072 26979
rect 23020 26936 23072 26945
rect 23388 26979 23440 26988
rect 23388 26945 23397 26979
rect 23397 26945 23431 26979
rect 23431 26945 23440 26979
rect 23388 26936 23440 26945
rect 24584 26936 24636 26988
rect 24860 26979 24912 26988
rect 24860 26945 24869 26979
rect 24869 26945 24903 26979
rect 24903 26945 24912 26979
rect 24860 26936 24912 26945
rect 25044 26979 25096 26988
rect 25044 26945 25053 26979
rect 25053 26945 25087 26979
rect 25087 26945 25096 26979
rect 25044 26936 25096 26945
rect 25136 26979 25188 26988
rect 25136 26945 25145 26979
rect 25145 26945 25179 26979
rect 25179 26945 25188 26979
rect 25136 26936 25188 26945
rect 25228 26979 25280 26988
rect 25228 26945 25238 26979
rect 25238 26945 25272 26979
rect 25272 26945 25280 26979
rect 25228 26936 25280 26945
rect 22928 26911 22980 26920
rect 22928 26877 22937 26911
rect 22937 26877 22971 26911
rect 22971 26877 22980 26911
rect 22928 26868 22980 26877
rect 24492 26868 24544 26920
rect 24952 26868 25004 26920
rect 26608 26868 26660 26920
rect 25596 26800 25648 26852
rect 26976 27004 27028 27056
rect 27712 27004 27764 27056
rect 30564 27004 30616 27056
rect 32036 27004 32088 27056
rect 59176 27072 59228 27124
rect 58164 27047 58216 27056
rect 58164 27013 58173 27047
rect 58173 27013 58207 27047
rect 58207 27013 58216 27047
rect 58164 27004 58216 27013
rect 27988 26979 28040 26988
rect 27988 26945 27997 26979
rect 27997 26945 28031 26979
rect 28031 26945 28040 26979
rect 27988 26936 28040 26945
rect 29092 26936 29144 26988
rect 30656 26979 30708 26988
rect 30656 26945 30665 26979
rect 30665 26945 30699 26979
rect 30699 26945 30708 26979
rect 30656 26936 30708 26945
rect 30748 26979 30800 26988
rect 30748 26945 30757 26979
rect 30757 26945 30791 26979
rect 30791 26945 30800 26979
rect 30748 26936 30800 26945
rect 31392 26936 31444 26988
rect 32772 26979 32824 26988
rect 32772 26945 32781 26979
rect 32781 26945 32815 26979
rect 32815 26945 32824 26979
rect 32772 26936 32824 26945
rect 32956 26979 33008 26988
rect 32956 26945 32965 26979
rect 32965 26945 32999 26979
rect 32999 26945 33008 26979
rect 32956 26936 33008 26945
rect 33140 26979 33192 26988
rect 33140 26945 33149 26979
rect 33149 26945 33183 26979
rect 33183 26945 33192 26979
rect 33140 26936 33192 26945
rect 42800 26936 42852 26988
rect 43168 26936 43220 26988
rect 30932 26868 30984 26920
rect 31668 26868 31720 26920
rect 34152 26868 34204 26920
rect 47216 26868 47268 26920
rect 49424 26868 49476 26920
rect 27068 26800 27120 26852
rect 30012 26732 30064 26784
rect 32588 26843 32640 26852
rect 32588 26809 32597 26843
rect 32597 26809 32631 26843
rect 32631 26809 32640 26843
rect 32588 26800 32640 26809
rect 43720 26800 43772 26852
rect 45468 26732 45520 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 22928 26528 22980 26580
rect 25412 26528 25464 26580
rect 27896 26528 27948 26580
rect 29920 26528 29972 26580
rect 20168 26324 20220 26376
rect 940 26256 992 26308
rect 1952 26256 2004 26308
rect 25412 26367 25464 26376
rect 25412 26333 25461 26367
rect 25461 26333 25464 26367
rect 25412 26324 25464 26333
rect 25596 26367 25648 26376
rect 25596 26333 25605 26367
rect 25605 26333 25639 26367
rect 25639 26333 25648 26367
rect 25596 26324 25648 26333
rect 23204 26256 23256 26308
rect 24860 26256 24912 26308
rect 28172 26392 28224 26444
rect 28356 26435 28408 26444
rect 28356 26401 28365 26435
rect 28365 26401 28399 26435
rect 28399 26401 28408 26435
rect 28356 26392 28408 26401
rect 26516 26367 26568 26376
rect 26516 26333 26525 26367
rect 26525 26333 26559 26367
rect 26559 26333 26568 26367
rect 26516 26324 26568 26333
rect 29092 26324 29144 26376
rect 24768 26188 24820 26240
rect 26332 26299 26384 26308
rect 26332 26265 26341 26299
rect 26341 26265 26375 26299
rect 26375 26265 26384 26299
rect 26332 26256 26384 26265
rect 26700 26256 26752 26308
rect 59360 26528 59412 26580
rect 43260 26460 43312 26512
rect 47952 26460 48004 26512
rect 29920 26367 29972 26376
rect 29920 26333 29929 26367
rect 29929 26333 29963 26367
rect 29963 26333 29972 26367
rect 29920 26324 29972 26333
rect 30012 26367 30064 26376
rect 30012 26333 30021 26367
rect 30021 26333 30055 26367
rect 30055 26333 30064 26367
rect 30012 26324 30064 26333
rect 30104 26367 30156 26376
rect 30104 26333 30113 26367
rect 30113 26333 30147 26367
rect 30147 26333 30156 26367
rect 30104 26324 30156 26333
rect 31668 26392 31720 26444
rect 30656 26324 30708 26376
rect 32956 26392 33008 26444
rect 35348 26392 35400 26444
rect 37832 26392 37884 26444
rect 30748 26256 30800 26308
rect 42800 26324 42852 26376
rect 43076 26324 43128 26376
rect 43260 26324 43312 26376
rect 43168 26256 43220 26308
rect 43720 26256 43772 26308
rect 30288 26231 30340 26240
rect 30288 26197 30297 26231
rect 30297 26197 30331 26231
rect 30331 26197 30340 26231
rect 30288 26188 30340 26197
rect 48228 26367 48280 26376
rect 48228 26333 48237 26367
rect 48237 26333 48271 26367
rect 48271 26333 48280 26367
rect 48228 26324 48280 26333
rect 48780 26392 48832 26444
rect 49240 26392 49292 26444
rect 48964 26367 49016 26376
rect 48964 26333 48973 26367
rect 48973 26333 49007 26367
rect 49007 26333 49016 26367
rect 48964 26324 49016 26333
rect 52920 26392 52972 26444
rect 58164 26435 58216 26444
rect 58164 26401 58173 26435
rect 58173 26401 58207 26435
rect 58207 26401 58216 26435
rect 58164 26392 58216 26401
rect 49424 26367 49476 26376
rect 49424 26333 49438 26367
rect 49438 26333 49472 26367
rect 49472 26333 49476 26367
rect 49424 26324 49476 26333
rect 53104 26324 53156 26376
rect 48688 26256 48740 26308
rect 48228 26188 48280 26240
rect 48412 26188 48464 26240
rect 56232 26188 56284 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 50294 26086 50346 26138
rect 50358 26086 50410 26138
rect 50422 26086 50474 26138
rect 50486 26086 50538 26138
rect 50550 26086 50602 26138
rect 20168 25916 20220 25968
rect 1584 25891 1636 25900
rect 1584 25857 1593 25891
rect 1593 25857 1627 25891
rect 1627 25857 1636 25891
rect 1584 25848 1636 25857
rect 20996 25891 21048 25900
rect 20996 25857 21005 25891
rect 21005 25857 21039 25891
rect 21039 25857 21048 25891
rect 20996 25848 21048 25857
rect 23020 25984 23072 26036
rect 24584 26027 24636 26036
rect 24584 25993 24593 26027
rect 24593 25993 24627 26027
rect 24627 25993 24636 26027
rect 24584 25984 24636 25993
rect 32588 25984 32640 26036
rect 41788 25984 41840 26036
rect 22928 25959 22980 25968
rect 22928 25925 22937 25959
rect 22937 25925 22971 25959
rect 22971 25925 22980 25959
rect 22928 25916 22980 25925
rect 23664 25916 23716 25968
rect 23940 25916 23992 25968
rect 22376 25848 22428 25900
rect 23296 25848 23348 25900
rect 24032 25848 24084 25900
rect 29092 25916 29144 25968
rect 28172 25891 28224 25900
rect 28172 25857 28181 25891
rect 28181 25857 28215 25891
rect 28215 25857 28224 25891
rect 28172 25848 28224 25857
rect 30104 25891 30156 25900
rect 30104 25857 30113 25891
rect 30113 25857 30147 25891
rect 30147 25857 30156 25891
rect 30104 25848 30156 25857
rect 30288 25848 30340 25900
rect 30380 25891 30432 25900
rect 30380 25857 30389 25891
rect 30389 25857 30423 25891
rect 30423 25857 30432 25891
rect 30380 25848 30432 25857
rect 37004 25848 37056 25900
rect 42064 25916 42116 25968
rect 45376 25916 45428 25968
rect 58164 25959 58216 25968
rect 58164 25925 58173 25959
rect 58173 25925 58207 25959
rect 58207 25925 58216 25959
rect 58164 25916 58216 25925
rect 41788 25848 41840 25900
rect 43260 25891 43312 25900
rect 43260 25857 43269 25891
rect 43269 25857 43303 25891
rect 43303 25857 43312 25891
rect 43260 25848 43312 25857
rect 43444 25891 43496 25900
rect 43444 25857 43451 25891
rect 43451 25857 43496 25891
rect 43444 25848 43496 25857
rect 43812 25848 43864 25900
rect 940 25780 992 25832
rect 23572 25780 23624 25832
rect 24584 25780 24636 25832
rect 27712 25780 27764 25832
rect 28264 25780 28316 25832
rect 30564 25823 30616 25832
rect 30564 25789 30573 25823
rect 30573 25789 30607 25823
rect 30607 25789 30616 25823
rect 30564 25780 30616 25789
rect 37556 25780 37608 25832
rect 38476 25780 38528 25832
rect 38844 25823 38896 25832
rect 38844 25789 38853 25823
rect 38853 25789 38887 25823
rect 38887 25789 38896 25823
rect 38844 25780 38896 25789
rect 47124 25780 47176 25832
rect 48872 25780 48924 25832
rect 23112 25712 23164 25764
rect 27896 25712 27948 25764
rect 32220 25712 32272 25764
rect 50068 25712 50120 25764
rect 26332 25644 26384 25696
rect 46756 25644 46808 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 1584 25440 1636 25492
rect 28172 25440 28224 25492
rect 30104 25440 30156 25492
rect 23664 25372 23716 25424
rect 22928 25304 22980 25356
rect 23480 25304 23532 25356
rect 24584 25304 24636 25356
rect 940 25168 992 25220
rect 2504 25279 2556 25288
rect 2504 25245 2513 25279
rect 2513 25245 2547 25279
rect 2547 25245 2556 25279
rect 2504 25236 2556 25245
rect 3148 25236 3200 25288
rect 23572 25236 23624 25288
rect 24492 25236 24544 25288
rect 37648 25372 37700 25424
rect 43812 25372 43864 25424
rect 45100 25372 45152 25424
rect 47860 25440 47912 25492
rect 27160 25279 27212 25288
rect 27160 25245 27169 25279
rect 27169 25245 27203 25279
rect 27203 25245 27212 25279
rect 27160 25236 27212 25245
rect 27712 25304 27764 25356
rect 27896 25304 27948 25356
rect 27528 25279 27580 25288
rect 27528 25245 27537 25279
rect 27537 25245 27571 25279
rect 27571 25245 27580 25279
rect 27528 25236 27580 25245
rect 27620 25236 27672 25288
rect 28264 25279 28316 25288
rect 28264 25245 28273 25279
rect 28273 25245 28307 25279
rect 28307 25245 28316 25279
rect 28264 25236 28316 25245
rect 28448 25279 28500 25288
rect 28448 25245 28457 25279
rect 28457 25245 28491 25279
rect 28491 25245 28500 25279
rect 28448 25236 28500 25245
rect 30748 25236 30800 25288
rect 37280 25279 37332 25288
rect 37280 25245 37289 25279
rect 37289 25245 37323 25279
rect 37323 25245 37332 25279
rect 37280 25236 37332 25245
rect 39488 25304 39540 25356
rect 37648 25279 37700 25288
rect 37648 25245 37657 25279
rect 37657 25245 37691 25279
rect 37691 25245 37700 25279
rect 37648 25236 37700 25245
rect 38844 25236 38896 25288
rect 43260 25236 43312 25288
rect 45928 25236 45980 25288
rect 46204 25279 46256 25288
rect 46204 25245 46211 25279
rect 46211 25245 46256 25279
rect 46204 25236 46256 25245
rect 46388 25279 46440 25288
rect 46388 25245 46397 25279
rect 46397 25245 46431 25279
rect 46431 25245 46440 25279
rect 46388 25236 46440 25245
rect 23296 25168 23348 25220
rect 27436 25211 27488 25220
rect 27436 25177 27445 25211
rect 27445 25177 27479 25211
rect 27479 25177 27488 25211
rect 27436 25168 27488 25177
rect 28356 25168 28408 25220
rect 22284 25100 22336 25152
rect 28080 25100 28132 25152
rect 31024 25143 31076 25152
rect 31024 25109 31033 25143
rect 31033 25109 31067 25143
rect 31067 25109 31076 25143
rect 31024 25100 31076 25109
rect 37556 25211 37608 25220
rect 37556 25177 37565 25211
rect 37565 25177 37599 25211
rect 37599 25177 37608 25211
rect 37556 25168 37608 25177
rect 38476 25168 38528 25220
rect 46296 25211 46348 25220
rect 46296 25177 46305 25211
rect 46305 25177 46339 25211
rect 46339 25177 46348 25211
rect 46296 25168 46348 25177
rect 47124 25279 47176 25288
rect 47124 25245 47133 25279
rect 47133 25245 47167 25279
rect 47167 25245 47176 25279
rect 47124 25236 47176 25245
rect 47032 25168 47084 25220
rect 47400 25279 47452 25288
rect 47400 25245 47409 25279
rect 47409 25245 47443 25279
rect 47443 25245 47452 25279
rect 47400 25236 47452 25245
rect 51724 25304 51776 25356
rect 48412 25279 48464 25288
rect 48412 25245 48421 25279
rect 48421 25245 48455 25279
rect 48455 25245 48464 25279
rect 48412 25236 48464 25245
rect 57888 25279 57940 25288
rect 57888 25245 57897 25279
rect 57897 25245 57931 25279
rect 57931 25245 57940 25279
rect 57888 25236 57940 25245
rect 49056 25168 49108 25220
rect 58164 25211 58216 25220
rect 58164 25177 58173 25211
rect 58173 25177 58207 25211
rect 58207 25177 58216 25211
rect 58164 25168 58216 25177
rect 47768 25143 47820 25152
rect 47768 25109 47777 25143
rect 47777 25109 47811 25143
rect 47811 25109 47820 25143
rect 47768 25100 47820 25109
rect 47860 25100 47912 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 50294 24998 50346 25050
rect 50358 24998 50410 25050
rect 50422 24998 50474 25050
rect 50486 24998 50538 25050
rect 50550 24998 50602 25050
rect 2504 24896 2556 24948
rect 1584 24803 1636 24812
rect 1584 24769 1593 24803
rect 1593 24769 1627 24803
rect 1627 24769 1636 24803
rect 1584 24760 1636 24769
rect 2412 24760 2464 24812
rect 23296 24896 23348 24948
rect 22284 24871 22336 24880
rect 22284 24837 22293 24871
rect 22293 24837 22327 24871
rect 22327 24837 22336 24871
rect 22284 24828 22336 24837
rect 940 24692 992 24744
rect 2136 24692 2188 24744
rect 15752 24760 15804 24812
rect 20996 24760 21048 24812
rect 22192 24760 22244 24812
rect 23664 24828 23716 24880
rect 24216 24939 24268 24948
rect 24216 24905 24225 24939
rect 24225 24905 24259 24939
rect 24259 24905 24268 24939
rect 24216 24896 24268 24905
rect 37280 24896 37332 24948
rect 46296 24896 46348 24948
rect 47400 24896 47452 24948
rect 47584 24896 47636 24948
rect 24032 24803 24084 24812
rect 24032 24769 24041 24803
rect 24041 24769 24075 24803
rect 24075 24769 24084 24803
rect 24032 24760 24084 24769
rect 2964 24624 3016 24676
rect 23480 24624 23532 24676
rect 23204 24556 23256 24608
rect 24860 24760 24912 24812
rect 25136 24760 25188 24812
rect 25688 24760 25740 24812
rect 27620 24760 27672 24812
rect 28356 24828 28408 24880
rect 24308 24624 24360 24676
rect 28080 24803 28132 24812
rect 28080 24769 28089 24803
rect 28089 24769 28123 24803
rect 28123 24769 28132 24803
rect 28080 24760 28132 24769
rect 28908 24760 28960 24812
rect 28632 24692 28684 24744
rect 30748 24828 30800 24880
rect 32772 24828 32824 24880
rect 29736 24692 29788 24744
rect 31024 24692 31076 24744
rect 28080 24624 28132 24676
rect 37372 24692 37424 24744
rect 37740 24803 37792 24812
rect 37740 24769 37749 24803
rect 37749 24769 37783 24803
rect 37783 24769 37792 24803
rect 37740 24760 37792 24769
rect 37832 24803 37884 24812
rect 37832 24769 37841 24803
rect 37841 24769 37875 24803
rect 37875 24769 37884 24803
rect 37832 24760 37884 24769
rect 47768 24871 47820 24880
rect 47768 24837 47777 24871
rect 47777 24837 47811 24871
rect 47811 24837 47820 24871
rect 47768 24828 47820 24837
rect 48228 24828 48280 24880
rect 51448 24828 51500 24880
rect 40684 24760 40736 24812
rect 47952 24803 48004 24812
rect 47952 24769 47961 24803
rect 47961 24769 47995 24803
rect 47995 24769 48004 24803
rect 47952 24760 48004 24769
rect 58072 24803 58124 24812
rect 58072 24769 58081 24803
rect 58081 24769 58115 24803
rect 58115 24769 58124 24803
rect 58072 24760 58124 24769
rect 39304 24692 39356 24744
rect 29736 24556 29788 24608
rect 31024 24556 31076 24608
rect 42984 24624 43036 24676
rect 36544 24556 36596 24608
rect 40776 24556 40828 24608
rect 48044 24599 48096 24608
rect 48044 24565 48053 24599
rect 48053 24565 48087 24599
rect 48087 24565 48096 24599
rect 48044 24556 48096 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 1584 24352 1636 24404
rect 12808 24284 12860 24336
rect 16120 24216 16172 24268
rect 17224 24284 17276 24336
rect 17776 24284 17828 24336
rect 27804 24352 27856 24404
rect 28264 24352 28316 24404
rect 30380 24395 30432 24404
rect 30380 24361 30389 24395
rect 30389 24361 30423 24395
rect 30423 24361 30432 24395
rect 30380 24352 30432 24361
rect 28172 24284 28224 24336
rect 28448 24284 28500 24336
rect 28540 24284 28592 24336
rect 36544 24352 36596 24404
rect 37096 24352 37148 24404
rect 41328 24352 41380 24404
rect 47676 24395 47728 24404
rect 47676 24361 47685 24395
rect 47685 24361 47719 24395
rect 47719 24361 47728 24395
rect 47676 24352 47728 24361
rect 33140 24284 33192 24336
rect 2412 24148 2464 24200
rect 2688 24191 2740 24200
rect 2688 24157 2701 24191
rect 2701 24157 2740 24191
rect 2688 24148 2740 24157
rect 23112 24191 23164 24200
rect 23112 24157 23121 24191
rect 23121 24157 23155 24191
rect 23155 24157 23164 24191
rect 23112 24148 23164 24157
rect 23296 24148 23348 24200
rect 23664 24148 23716 24200
rect 28172 24191 28224 24200
rect 28172 24157 28181 24191
rect 28181 24157 28215 24191
rect 28215 24157 28224 24191
rect 28172 24148 28224 24157
rect 940 24080 992 24132
rect 23204 24080 23256 24132
rect 27988 24080 28040 24132
rect 28448 24191 28500 24200
rect 28448 24157 28457 24191
rect 28457 24157 28491 24191
rect 28491 24157 28500 24191
rect 28448 24148 28500 24157
rect 28632 24191 28684 24200
rect 28632 24157 28646 24191
rect 28646 24157 28680 24191
rect 28680 24157 28684 24191
rect 28632 24148 28684 24157
rect 29736 24191 29788 24200
rect 29736 24157 29745 24191
rect 29745 24157 29779 24191
rect 29779 24157 29788 24191
rect 29736 24148 29788 24157
rect 29828 24191 29880 24200
rect 29828 24157 29838 24191
rect 29838 24157 29872 24191
rect 29872 24157 29880 24191
rect 29828 24148 29880 24157
rect 30288 24148 30340 24200
rect 29092 24080 29144 24132
rect 45192 24216 45244 24268
rect 37280 24191 37332 24200
rect 37280 24157 37289 24191
rect 37289 24157 37323 24191
rect 37323 24157 37332 24191
rect 37280 24148 37332 24157
rect 37372 24148 37424 24200
rect 37648 24191 37700 24200
rect 37648 24157 37657 24191
rect 37657 24157 37691 24191
rect 37691 24157 37700 24191
rect 37648 24148 37700 24157
rect 24032 24012 24084 24064
rect 27712 24012 27764 24064
rect 36636 24080 36688 24132
rect 32036 24012 32088 24064
rect 42800 24148 42852 24200
rect 46940 24148 46992 24200
rect 47584 24148 47636 24200
rect 39396 24080 39448 24132
rect 37924 24012 37976 24064
rect 47400 24123 47452 24132
rect 47400 24089 47409 24123
rect 47409 24089 47443 24123
rect 47443 24089 47452 24123
rect 47400 24080 47452 24089
rect 40224 24012 40276 24064
rect 54300 24216 54352 24268
rect 55220 24148 55272 24200
rect 58164 24123 58216 24132
rect 58164 24089 58173 24123
rect 58173 24089 58207 24123
rect 58207 24089 58216 24123
rect 58164 24080 58216 24089
rect 53380 24012 53432 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 50294 23910 50346 23962
rect 50358 23910 50410 23962
rect 50422 23910 50474 23962
rect 50486 23910 50538 23962
rect 50550 23910 50602 23962
rect 16120 23851 16172 23860
rect 16120 23817 16129 23851
rect 16129 23817 16163 23851
rect 16163 23817 16172 23851
rect 16120 23808 16172 23817
rect 23204 23808 23256 23860
rect 24400 23851 24452 23860
rect 24400 23817 24409 23851
rect 24409 23817 24443 23851
rect 24443 23817 24452 23851
rect 24400 23808 24452 23817
rect 28172 23808 28224 23860
rect 36636 23808 36688 23860
rect 20996 23740 21048 23792
rect 2872 23672 2924 23724
rect 15752 23715 15804 23724
rect 15752 23681 15761 23715
rect 15761 23681 15795 23715
rect 15795 23681 15804 23715
rect 15752 23672 15804 23681
rect 17776 23672 17828 23724
rect 23664 23672 23716 23724
rect 940 23604 992 23656
rect 23296 23604 23348 23656
rect 24032 23715 24084 23724
rect 24032 23681 24041 23715
rect 24041 23681 24075 23715
rect 24075 23681 24084 23715
rect 24032 23672 24084 23681
rect 27804 23740 27856 23792
rect 28632 23740 28684 23792
rect 37372 23740 37424 23792
rect 34428 23672 34480 23724
rect 36912 23672 36964 23724
rect 42156 23808 42208 23860
rect 42708 23740 42760 23792
rect 40868 23672 40920 23724
rect 35900 23604 35952 23656
rect 41696 23715 41748 23724
rect 41696 23681 41705 23715
rect 41705 23681 41739 23715
rect 41739 23681 41748 23715
rect 41696 23672 41748 23681
rect 42156 23672 42208 23724
rect 58072 23715 58124 23724
rect 58072 23681 58081 23715
rect 58081 23681 58115 23715
rect 58115 23681 58124 23715
rect 58072 23672 58124 23681
rect 36728 23536 36780 23588
rect 34152 23511 34204 23520
rect 34152 23477 34161 23511
rect 34161 23477 34195 23511
rect 34195 23477 34204 23511
rect 34152 23468 34204 23477
rect 36360 23468 36412 23520
rect 40132 23536 40184 23588
rect 42892 23604 42944 23656
rect 37464 23468 37516 23520
rect 40040 23468 40092 23520
rect 41328 23536 41380 23588
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 21364 23264 21416 23316
rect 24676 23264 24728 23316
rect 2872 23239 2924 23248
rect 2872 23205 2881 23239
rect 2881 23205 2915 23239
rect 2915 23205 2924 23239
rect 2872 23196 2924 23205
rect 23848 23196 23900 23248
rect 26700 23196 26752 23248
rect 36452 23264 36504 23316
rect 39120 23264 39172 23316
rect 2412 23128 2464 23180
rect 940 22992 992 23044
rect 3424 23060 3476 23112
rect 29736 23103 29788 23112
rect 29736 23069 29745 23103
rect 29745 23069 29779 23103
rect 29779 23069 29788 23103
rect 29736 23060 29788 23069
rect 31392 23128 31444 23180
rect 30656 23103 30708 23112
rect 30656 23069 30665 23103
rect 30665 23069 30699 23103
rect 30699 23069 30708 23103
rect 30656 23060 30708 23069
rect 33784 23060 33836 23112
rect 36452 23128 36504 23180
rect 34888 23103 34940 23112
rect 34888 23069 34897 23103
rect 34897 23069 34931 23103
rect 34931 23069 34940 23103
rect 34888 23060 34940 23069
rect 35900 23103 35952 23112
rect 35900 23069 35909 23103
rect 35909 23069 35943 23103
rect 35943 23069 35952 23103
rect 35900 23060 35952 23069
rect 36820 23060 36872 23112
rect 39948 23128 40000 23180
rect 2780 22992 2832 23044
rect 29828 22992 29880 23044
rect 32772 22992 32824 23044
rect 29552 22924 29604 22976
rect 33508 22924 33560 22976
rect 33692 22924 33744 22976
rect 35256 22992 35308 23044
rect 36176 22992 36228 23044
rect 36912 22992 36964 23044
rect 35164 22924 35216 22976
rect 38844 22967 38896 22976
rect 38844 22933 38853 22967
rect 38853 22933 38887 22967
rect 38887 22933 38896 22967
rect 38844 22924 38896 22933
rect 39212 23103 39264 23112
rect 39212 23069 39221 23103
rect 39221 23069 39255 23103
rect 39255 23069 39264 23103
rect 39212 23060 39264 23069
rect 39580 23060 39632 23112
rect 40040 23103 40092 23112
rect 40040 23069 40049 23103
rect 40049 23069 40083 23103
rect 40083 23069 40092 23103
rect 40040 23060 40092 23069
rect 42892 23307 42944 23316
rect 42892 23273 42901 23307
rect 42901 23273 42935 23307
rect 42935 23273 42944 23307
rect 42892 23264 42944 23273
rect 45744 23264 45796 23316
rect 41420 23128 41472 23180
rect 43444 23128 43496 23180
rect 56968 23196 57020 23248
rect 51908 23128 51960 23180
rect 41880 23103 41932 23112
rect 41880 23069 41889 23103
rect 41889 23069 41923 23103
rect 41923 23069 41932 23103
rect 41880 23060 41932 23069
rect 41972 23103 42024 23112
rect 41972 23069 41981 23103
rect 41981 23069 42015 23103
rect 42015 23069 42024 23103
rect 41972 23060 42024 23069
rect 42064 23103 42116 23112
rect 42064 23069 42073 23103
rect 42073 23069 42107 23103
rect 42107 23069 42116 23103
rect 42064 23060 42116 23069
rect 42248 23103 42300 23112
rect 42248 23069 42257 23103
rect 42257 23069 42291 23103
rect 42291 23069 42300 23103
rect 42248 23060 42300 23069
rect 42524 23060 42576 23112
rect 48228 23103 48280 23112
rect 48228 23069 48237 23103
rect 48237 23069 48271 23103
rect 48271 23069 48280 23103
rect 48228 23060 48280 23069
rect 49240 23060 49292 23112
rect 51632 23060 51684 23112
rect 55404 23060 55456 23112
rect 58256 23128 58308 23180
rect 40132 22992 40184 23044
rect 41144 22992 41196 23044
rect 41328 22992 41380 23044
rect 48320 22992 48372 23044
rect 48504 23035 48556 23044
rect 48504 23001 48513 23035
rect 48513 23001 48547 23035
rect 48547 23001 48556 23035
rect 48504 22992 48556 23001
rect 41512 22924 41564 22976
rect 42340 22924 42392 22976
rect 43812 22924 43864 22976
rect 53748 22992 53800 23044
rect 53840 22992 53892 23044
rect 48688 22924 48740 22976
rect 52000 22924 52052 22976
rect 56416 22924 56468 22976
rect 58164 23035 58216 23044
rect 58164 23001 58173 23035
rect 58173 23001 58207 23035
rect 58207 23001 58216 23035
rect 58164 22992 58216 23001
rect 58992 22924 59044 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 50294 22822 50346 22874
rect 50358 22822 50410 22874
rect 50422 22822 50474 22874
rect 50486 22822 50538 22874
rect 50550 22822 50602 22874
rect 2412 22720 2464 22772
rect 18512 22720 18564 22772
rect 30196 22720 30248 22772
rect 22468 22652 22520 22704
rect 24124 22695 24176 22704
rect 24124 22661 24133 22695
rect 24133 22661 24167 22695
rect 24167 22661 24176 22695
rect 24124 22652 24176 22661
rect 24768 22652 24820 22704
rect 10508 22584 10560 22636
rect 24400 22584 24452 22636
rect 29552 22627 29604 22636
rect 29552 22593 29561 22627
rect 29561 22593 29595 22627
rect 29595 22593 29604 22627
rect 29552 22584 29604 22593
rect 30288 22627 30340 22636
rect 30288 22593 30297 22627
rect 30297 22593 30331 22627
rect 30331 22593 30340 22627
rect 30288 22584 30340 22593
rect 32772 22627 32824 22636
rect 32772 22593 32781 22627
rect 32781 22593 32815 22627
rect 32815 22593 32824 22627
rect 32772 22584 32824 22593
rect 31576 22516 31628 22568
rect 33784 22763 33836 22772
rect 33784 22729 33793 22763
rect 33793 22729 33827 22763
rect 33827 22729 33836 22763
rect 33784 22720 33836 22729
rect 34888 22720 34940 22772
rect 37740 22720 37792 22772
rect 39948 22720 40000 22772
rect 40040 22720 40092 22772
rect 41604 22720 41656 22772
rect 42616 22720 42668 22772
rect 42708 22720 42760 22772
rect 35440 22652 35492 22704
rect 35256 22584 35308 22636
rect 38200 22652 38252 22704
rect 35348 22516 35400 22568
rect 35440 22516 35492 22568
rect 36084 22584 36136 22636
rect 37464 22627 37516 22636
rect 37464 22593 37473 22627
rect 37473 22593 37507 22627
rect 37507 22593 37516 22627
rect 37464 22584 37516 22593
rect 38844 22652 38896 22704
rect 40960 22652 41012 22704
rect 44272 22720 44324 22772
rect 44364 22720 44416 22772
rect 46664 22763 46716 22772
rect 46664 22729 46673 22763
rect 46673 22729 46707 22763
rect 46707 22729 46716 22763
rect 46664 22720 46716 22729
rect 48044 22720 48096 22772
rect 48504 22720 48556 22772
rect 49792 22720 49844 22772
rect 32220 22448 32272 22500
rect 36912 22491 36964 22500
rect 36912 22457 36921 22491
rect 36921 22457 36955 22491
rect 36955 22457 36964 22491
rect 36912 22448 36964 22457
rect 30012 22380 30064 22432
rect 30380 22380 30432 22432
rect 32772 22380 32824 22432
rect 35900 22380 35952 22432
rect 38844 22380 38896 22432
rect 41604 22627 41656 22636
rect 41604 22593 41613 22627
rect 41613 22593 41647 22627
rect 41647 22593 41656 22627
rect 41604 22584 41656 22593
rect 41328 22516 41380 22568
rect 43444 22652 43496 22704
rect 51632 22763 51684 22772
rect 51632 22729 51641 22763
rect 51641 22729 51675 22763
rect 51675 22729 51684 22763
rect 51632 22720 51684 22729
rect 53748 22720 53800 22772
rect 42248 22584 42300 22636
rect 42708 22584 42760 22636
rect 43352 22627 43404 22636
rect 43352 22593 43361 22627
rect 43361 22593 43395 22627
rect 43395 22593 43404 22627
rect 43352 22584 43404 22593
rect 44180 22584 44232 22636
rect 48780 22627 48832 22636
rect 48780 22593 48814 22627
rect 48814 22593 48832 22627
rect 48780 22584 48832 22593
rect 49240 22584 49292 22636
rect 51080 22627 51132 22636
rect 51080 22593 51089 22627
rect 51089 22593 51123 22627
rect 51123 22593 51132 22627
rect 51080 22584 51132 22593
rect 57980 22652 58032 22704
rect 41420 22448 41472 22500
rect 42524 22448 42576 22500
rect 42708 22380 42760 22432
rect 43536 22423 43588 22432
rect 43536 22389 43545 22423
rect 43545 22389 43579 22423
rect 43579 22389 43588 22423
rect 43536 22380 43588 22389
rect 44088 22559 44140 22568
rect 44088 22525 44097 22559
rect 44097 22525 44131 22559
rect 44131 22525 44140 22559
rect 44088 22516 44140 22525
rect 46572 22516 46624 22568
rect 46848 22516 46900 22568
rect 48412 22516 48464 22568
rect 51724 22584 51776 22636
rect 53012 22584 53064 22636
rect 54116 22584 54168 22636
rect 56324 22584 56376 22636
rect 58072 22627 58124 22636
rect 58072 22593 58081 22627
rect 58081 22593 58115 22627
rect 58115 22593 58124 22627
rect 58072 22584 58124 22593
rect 51908 22516 51960 22568
rect 55404 22516 55456 22568
rect 56416 22516 56468 22568
rect 53012 22448 53064 22500
rect 45560 22380 45612 22432
rect 49148 22380 49200 22432
rect 49792 22380 49844 22432
rect 55220 22448 55272 22500
rect 53288 22423 53340 22432
rect 53288 22389 53297 22423
rect 53297 22389 53331 22423
rect 53331 22389 53340 22423
rect 53288 22380 53340 22389
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 2780 22176 2832 22228
rect 29736 22176 29788 22228
rect 30840 22176 30892 22228
rect 940 22040 992 22092
rect 31116 22108 31168 22160
rect 31392 22108 31444 22160
rect 23480 22040 23532 22092
rect 28080 22040 28132 22092
rect 31576 22219 31628 22228
rect 31576 22185 31585 22219
rect 31585 22185 31619 22219
rect 31619 22185 31628 22219
rect 31576 22176 31628 22185
rect 32220 22219 32272 22228
rect 32220 22185 32229 22219
rect 32229 22185 32263 22219
rect 32263 22185 32272 22219
rect 32220 22176 32272 22185
rect 35440 22219 35492 22228
rect 35440 22185 35449 22219
rect 35449 22185 35483 22219
rect 35483 22185 35492 22219
rect 35440 22176 35492 22185
rect 32956 22108 33008 22160
rect 37740 22176 37792 22228
rect 38108 22176 38160 22228
rect 39856 22176 39908 22228
rect 48780 22176 48832 22228
rect 49148 22176 49200 22228
rect 35808 22108 35860 22160
rect 38752 22151 38804 22160
rect 38752 22117 38761 22151
rect 38761 22117 38795 22151
rect 38795 22117 38804 22151
rect 38752 22108 38804 22117
rect 38936 22108 38988 22160
rect 39120 22108 39172 22160
rect 2504 22015 2556 22024
rect 2504 21981 2513 22015
rect 2513 21981 2547 22015
rect 2547 21981 2556 22015
rect 2504 21972 2556 21981
rect 2596 22015 2648 22024
rect 2596 21981 2606 22015
rect 2606 21981 2640 22015
rect 2640 21981 2648 22015
rect 2596 21972 2648 21981
rect 10140 21972 10192 22024
rect 10508 21972 10560 22024
rect 22008 22015 22060 22024
rect 22008 21981 22017 22015
rect 22017 21981 22051 22015
rect 22051 21981 22060 22015
rect 22008 21972 22060 21981
rect 24124 21972 24176 22024
rect 26608 21972 26660 22024
rect 28264 21972 28316 22024
rect 29276 21972 29328 22024
rect 30932 21972 30984 22024
rect 33692 22040 33744 22092
rect 31392 22015 31444 22024
rect 31392 21981 31401 22015
rect 31401 21981 31435 22015
rect 31435 21981 31444 22015
rect 31392 21972 31444 21981
rect 31024 21947 31076 21956
rect 31024 21913 31033 21947
rect 31033 21913 31067 21947
rect 31067 21913 31076 21947
rect 31024 21904 31076 21913
rect 32772 22015 32824 22024
rect 32772 21981 32781 22015
rect 32781 21981 32815 22015
rect 32815 21981 32824 22015
rect 32772 21972 32824 21981
rect 33048 21972 33100 22024
rect 34796 21972 34848 22024
rect 23940 21836 23992 21888
rect 25228 21836 25280 21888
rect 28172 21879 28224 21888
rect 28172 21845 28181 21879
rect 28181 21845 28215 21879
rect 28215 21845 28224 21879
rect 28172 21836 28224 21845
rect 31392 21836 31444 21888
rect 32864 21836 32916 21888
rect 35900 22012 35952 22024
rect 35900 21978 35930 22012
rect 35930 21978 35952 22012
rect 35900 21972 35952 21978
rect 36268 21972 36320 22024
rect 36912 21972 36964 22024
rect 37096 21904 37148 21956
rect 38752 21972 38804 22024
rect 39028 22015 39080 22024
rect 39028 21981 39037 22015
rect 39037 21981 39071 22015
rect 39071 21981 39080 22015
rect 39028 21972 39080 21981
rect 39672 22040 39724 22092
rect 42800 22040 42852 22092
rect 51724 22108 51776 22160
rect 53104 22219 53156 22228
rect 53104 22185 53113 22219
rect 53113 22185 53147 22219
rect 53147 22185 53156 22219
rect 53104 22176 53156 22185
rect 54116 22219 54168 22228
rect 54116 22185 54125 22219
rect 54125 22185 54159 22219
rect 54159 22185 54168 22219
rect 54116 22176 54168 22185
rect 57152 22176 57204 22228
rect 58256 22219 58308 22228
rect 58256 22185 58265 22219
rect 58265 22185 58299 22219
rect 58299 22185 58308 22219
rect 58256 22176 58308 22185
rect 39580 21972 39632 22024
rect 39856 21972 39908 22024
rect 40500 21972 40552 22024
rect 41328 22015 41380 22024
rect 41328 21981 41337 22015
rect 41337 21981 41371 22015
rect 41371 21981 41380 22015
rect 41328 21972 41380 21981
rect 42340 22015 42392 22024
rect 42340 21981 42349 22015
rect 42349 21981 42383 22015
rect 42383 21981 42392 22015
rect 42340 21972 42392 21981
rect 42616 21972 42668 22024
rect 44088 21972 44140 22024
rect 44640 21972 44692 22024
rect 47676 22083 47728 22092
rect 47676 22049 47685 22083
rect 47685 22049 47719 22083
rect 47719 22049 47728 22083
rect 47676 22040 47728 22049
rect 51080 22040 51132 22092
rect 48596 22015 48648 22024
rect 48596 21981 48605 22015
rect 48605 21981 48639 22015
rect 48639 21981 48648 22015
rect 48596 21972 48648 21981
rect 48688 22015 48740 22024
rect 48688 21981 48697 22015
rect 48697 21981 48731 22015
rect 48731 21981 48740 22015
rect 48688 21972 48740 21981
rect 36636 21836 36688 21888
rect 37648 21836 37700 21888
rect 38108 21947 38160 21956
rect 38108 21913 38117 21947
rect 38117 21913 38151 21947
rect 38151 21913 38160 21947
rect 38108 21904 38160 21913
rect 38568 21836 38620 21888
rect 40408 21904 40460 21956
rect 41420 21904 41472 21956
rect 43444 21904 43496 21956
rect 44364 21947 44416 21956
rect 44364 21913 44373 21947
rect 44373 21913 44407 21947
rect 44407 21913 44416 21947
rect 44364 21904 44416 21913
rect 45284 21904 45336 21956
rect 47860 21904 47912 21956
rect 39120 21836 39172 21888
rect 40224 21879 40276 21888
rect 40224 21845 40233 21879
rect 40233 21845 40267 21879
rect 40267 21845 40276 21879
rect 40224 21836 40276 21845
rect 41604 21836 41656 21888
rect 43352 21836 43404 21888
rect 44548 21879 44600 21888
rect 44548 21845 44557 21879
rect 44557 21845 44591 21879
rect 44591 21845 44600 21879
rect 44548 21836 44600 21845
rect 46572 21879 46624 21888
rect 46572 21845 46581 21879
rect 46581 21845 46615 21879
rect 46615 21845 46624 21879
rect 46572 21836 46624 21845
rect 53012 22040 53064 22092
rect 53748 22040 53800 22092
rect 54024 22040 54076 22092
rect 57060 22040 57112 22092
rect 57796 22040 57848 22092
rect 52368 21972 52420 22024
rect 53564 22015 53616 22024
rect 53564 21981 53573 22015
rect 53573 21981 53607 22015
rect 53607 21981 53616 22015
rect 53564 21972 53616 21981
rect 53932 22015 53984 22024
rect 52000 21947 52052 21956
rect 52000 21913 52034 21947
rect 52034 21913 52052 21947
rect 52000 21904 52052 21913
rect 53932 21981 53941 22015
rect 53941 21981 53975 22015
rect 53975 21981 53984 22015
rect 53932 21972 53984 21981
rect 54208 21972 54260 22024
rect 55772 21972 55824 22024
rect 57152 21972 57204 22024
rect 53748 21947 53800 21956
rect 53748 21913 53757 21947
rect 53757 21913 53791 21947
rect 53791 21913 53800 21947
rect 53748 21904 53800 21913
rect 54024 21904 54076 21956
rect 55680 21904 55732 21956
rect 56324 21904 56376 21956
rect 55864 21836 55916 21888
rect 56784 21836 56836 21888
rect 57428 21904 57480 21956
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 50294 21734 50346 21786
rect 50358 21734 50410 21786
rect 50422 21734 50474 21786
rect 50486 21734 50538 21786
rect 50550 21734 50602 21786
rect 23204 21564 23256 21616
rect 23480 21564 23532 21616
rect 24032 21632 24084 21684
rect 28264 21675 28316 21684
rect 28264 21641 28273 21675
rect 28273 21641 28307 21675
rect 28307 21641 28316 21675
rect 28264 21632 28316 21641
rect 30288 21675 30340 21684
rect 30288 21641 30297 21675
rect 30297 21641 30331 21675
rect 30331 21641 30340 21675
rect 30288 21632 30340 21641
rect 30932 21675 30984 21684
rect 30932 21641 30941 21675
rect 30941 21641 30975 21675
rect 30975 21641 30984 21675
rect 30932 21632 30984 21641
rect 31024 21632 31076 21684
rect 11704 21496 11756 21548
rect 22100 21539 22152 21548
rect 22100 21505 22109 21539
rect 22109 21505 22143 21539
rect 22143 21505 22152 21539
rect 22100 21496 22152 21505
rect 22284 21496 22336 21548
rect 24860 21564 24912 21616
rect 27712 21564 27764 21616
rect 28080 21564 28132 21616
rect 940 21428 992 21480
rect 24584 21496 24636 21548
rect 25412 21496 25464 21548
rect 22468 21360 22520 21412
rect 24492 21428 24544 21480
rect 28448 21428 28500 21480
rect 29736 21496 29788 21548
rect 30840 21564 30892 21616
rect 31116 21539 31168 21548
rect 28356 21360 28408 21412
rect 29276 21471 29328 21480
rect 29276 21437 29285 21471
rect 29285 21437 29319 21471
rect 29319 21437 29328 21471
rect 29276 21428 29328 21437
rect 29828 21471 29880 21480
rect 29828 21437 29837 21471
rect 29837 21437 29871 21471
rect 29871 21437 29880 21471
rect 29828 21428 29880 21437
rect 29092 21360 29144 21412
rect 31116 21505 31125 21539
rect 31125 21505 31159 21539
rect 31159 21505 31168 21539
rect 31116 21496 31168 21505
rect 30656 21428 30708 21480
rect 36728 21675 36780 21684
rect 36728 21641 36737 21675
rect 36737 21641 36771 21675
rect 36771 21641 36780 21675
rect 36728 21632 36780 21641
rect 37004 21632 37056 21684
rect 41604 21632 41656 21684
rect 42064 21632 42116 21684
rect 31576 21564 31628 21616
rect 33048 21564 33100 21616
rect 32312 21539 32364 21548
rect 32312 21505 32321 21539
rect 32321 21505 32355 21539
rect 32355 21505 32364 21539
rect 32312 21496 32364 21505
rect 33692 21496 33744 21548
rect 36360 21564 36412 21616
rect 33048 21471 33100 21480
rect 33048 21437 33057 21471
rect 33057 21437 33091 21471
rect 33091 21437 33100 21471
rect 33048 21428 33100 21437
rect 34152 21428 34204 21480
rect 37188 21496 37240 21548
rect 31576 21360 31628 21412
rect 38844 21564 38896 21616
rect 37372 21496 37424 21548
rect 39672 21564 39724 21616
rect 40868 21564 40920 21616
rect 41236 21564 41288 21616
rect 42616 21632 42668 21684
rect 42800 21632 42852 21684
rect 43352 21632 43404 21684
rect 39396 21539 39448 21548
rect 39396 21505 39419 21539
rect 39419 21505 39448 21539
rect 39396 21496 39448 21505
rect 40408 21496 40460 21548
rect 42524 21496 42576 21548
rect 44088 21564 44140 21616
rect 53564 21632 53616 21684
rect 54024 21632 54076 21684
rect 46572 21564 46624 21616
rect 53288 21564 53340 21616
rect 55680 21675 55732 21684
rect 55680 21641 55689 21675
rect 55689 21641 55723 21675
rect 55723 21641 55732 21675
rect 55680 21632 55732 21641
rect 55864 21632 55916 21684
rect 57428 21632 57480 21684
rect 56600 21564 56652 21616
rect 42708 21496 42760 21548
rect 43444 21496 43496 21548
rect 48780 21539 48832 21548
rect 48780 21505 48789 21539
rect 48789 21505 48823 21539
rect 48823 21505 48832 21539
rect 48780 21496 48832 21505
rect 49792 21496 49844 21548
rect 55404 21539 55456 21548
rect 55404 21505 55413 21539
rect 55413 21505 55447 21539
rect 55447 21505 55456 21539
rect 55404 21496 55456 21505
rect 55496 21539 55548 21548
rect 55496 21505 55505 21539
rect 55505 21505 55539 21539
rect 55539 21505 55548 21539
rect 55496 21496 55548 21505
rect 56232 21496 56284 21548
rect 57428 21496 57480 21548
rect 57704 21496 57756 21548
rect 58072 21539 58124 21548
rect 58072 21505 58081 21539
rect 58081 21505 58115 21539
rect 58115 21505 58124 21539
rect 58072 21496 58124 21505
rect 26240 21292 26292 21344
rect 27344 21292 27396 21344
rect 30288 21292 30340 21344
rect 30840 21292 30892 21344
rect 37740 21360 37792 21412
rect 36728 21292 36780 21344
rect 37556 21292 37608 21344
rect 41420 21360 41472 21412
rect 40500 21335 40552 21344
rect 40500 21301 40509 21335
rect 40509 21301 40543 21335
rect 40543 21301 40552 21335
rect 40500 21292 40552 21301
rect 46020 21471 46072 21480
rect 46020 21437 46029 21471
rect 46029 21437 46063 21471
rect 46063 21437 46072 21471
rect 46020 21428 46072 21437
rect 46940 21428 46992 21480
rect 47676 21428 47728 21480
rect 52368 21428 52420 21480
rect 56140 21471 56192 21480
rect 56140 21437 56149 21471
rect 56149 21437 56183 21471
rect 56183 21437 56192 21471
rect 56140 21428 56192 21437
rect 45652 21360 45704 21412
rect 48688 21292 48740 21344
rect 57520 21335 57572 21344
rect 57520 21301 57529 21335
rect 57529 21301 57563 21335
rect 57563 21301 57572 21335
rect 57520 21292 57572 21301
rect 57612 21292 57664 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 23204 21131 23256 21140
rect 23204 21097 23213 21131
rect 23213 21097 23247 21131
rect 23247 21097 23256 21131
rect 23204 21088 23256 21097
rect 24860 21088 24912 21140
rect 25412 21131 25464 21140
rect 25412 21097 25421 21131
rect 25421 21097 25455 21131
rect 25455 21097 25464 21131
rect 25412 21088 25464 21097
rect 27344 21131 27396 21140
rect 27344 21097 27353 21131
rect 27353 21097 27387 21131
rect 27387 21097 27396 21131
rect 27344 21088 27396 21097
rect 30656 21088 30708 21140
rect 29092 21063 29144 21072
rect 29092 21029 29101 21063
rect 29101 21029 29135 21063
rect 29135 21029 29144 21063
rect 29092 21020 29144 21029
rect 31208 21020 31260 21072
rect 31392 21020 31444 21072
rect 32956 21088 33008 21140
rect 33692 21131 33744 21140
rect 33692 21097 33701 21131
rect 33701 21097 33735 21131
rect 33735 21097 33744 21131
rect 33692 21088 33744 21097
rect 36084 21088 36136 21140
rect 36912 21131 36964 21140
rect 36912 21097 36921 21131
rect 36921 21097 36955 21131
rect 36955 21097 36964 21131
rect 36912 21088 36964 21097
rect 37188 21088 37240 21140
rect 38384 21088 38436 21140
rect 43536 21088 43588 21140
rect 44180 21088 44232 21140
rect 45284 21088 45336 21140
rect 49884 21088 49936 21140
rect 55496 21088 55548 21140
rect 57796 21088 57848 21140
rect 37740 21020 37792 21072
rect 940 20952 992 21004
rect 22008 20927 22060 20936
rect 22008 20893 22017 20927
rect 22017 20893 22051 20927
rect 22051 20893 22060 20927
rect 22008 20884 22060 20893
rect 22468 20927 22520 20936
rect 22468 20893 22477 20927
rect 22477 20893 22511 20927
rect 22511 20893 22520 20927
rect 22468 20884 22520 20893
rect 23756 20927 23808 20936
rect 23756 20893 23765 20927
rect 23765 20893 23799 20927
rect 23799 20893 23808 20927
rect 23756 20884 23808 20893
rect 25228 20927 25280 20936
rect 25228 20893 25237 20927
rect 25237 20893 25271 20927
rect 25271 20893 25280 20927
rect 25228 20884 25280 20893
rect 28632 20952 28684 21004
rect 28540 20884 28592 20936
rect 33048 20952 33100 21004
rect 40316 21020 40368 21072
rect 40500 21020 40552 21072
rect 43260 21020 43312 21072
rect 29736 20927 29788 20936
rect 29736 20893 29745 20927
rect 29745 20893 29779 20927
rect 29779 20893 29788 20927
rect 29736 20884 29788 20893
rect 33508 20927 33560 20936
rect 33508 20893 33517 20927
rect 33517 20893 33551 20927
rect 33551 20893 33560 20927
rect 33508 20884 33560 20893
rect 36636 20884 36688 20936
rect 36728 20927 36780 20936
rect 36728 20893 36737 20927
rect 36737 20893 36771 20927
rect 36771 20893 36780 20927
rect 36728 20884 36780 20893
rect 24124 20816 24176 20868
rect 26240 20859 26292 20868
rect 26240 20825 26274 20859
rect 26274 20825 26292 20859
rect 26240 20816 26292 20825
rect 26332 20816 26384 20868
rect 27620 20748 27672 20800
rect 30012 20859 30064 20868
rect 30012 20825 30046 20859
rect 30046 20825 30064 20859
rect 30012 20816 30064 20825
rect 32864 20816 32916 20868
rect 32956 20816 33008 20868
rect 37464 20927 37516 20936
rect 37464 20893 37473 20927
rect 37473 20893 37507 20927
rect 37507 20893 37516 20927
rect 37464 20884 37516 20893
rect 38384 20884 38436 20936
rect 38568 20884 38620 20936
rect 38844 20884 38896 20936
rect 37832 20816 37884 20868
rect 32312 20748 32364 20800
rect 38660 20816 38712 20868
rect 39028 20816 39080 20868
rect 40224 20884 40276 20936
rect 40316 20884 40368 20936
rect 41236 20816 41288 20868
rect 41512 20927 41564 20936
rect 41512 20893 41521 20927
rect 41521 20893 41555 20927
rect 41555 20893 41564 20927
rect 41512 20884 41564 20893
rect 42524 20884 42576 20936
rect 43352 20884 43404 20936
rect 42156 20816 42208 20868
rect 42800 20859 42852 20868
rect 42800 20825 42809 20859
rect 42809 20825 42843 20859
rect 42843 20825 42852 20859
rect 42800 20816 42852 20825
rect 40224 20791 40276 20800
rect 40224 20757 40233 20791
rect 40233 20757 40267 20791
rect 40267 20757 40276 20791
rect 40224 20748 40276 20757
rect 40316 20748 40368 20800
rect 43352 20748 43404 20800
rect 43628 20884 43680 20936
rect 43904 20927 43956 20936
rect 43904 20893 43913 20927
rect 43913 20893 43947 20927
rect 43947 20893 43956 20927
rect 43904 20884 43956 20893
rect 43996 20927 44048 20936
rect 43996 20893 44005 20927
rect 44005 20893 44039 20927
rect 44039 20893 44048 20927
rect 43996 20884 44048 20893
rect 44548 20952 44600 21004
rect 44272 20927 44324 20936
rect 44272 20893 44281 20927
rect 44281 20893 44315 20927
rect 44315 20893 44324 20927
rect 44272 20884 44324 20893
rect 45836 21020 45888 21072
rect 46756 21020 46808 21072
rect 55772 20952 55824 21004
rect 56140 20952 56192 21004
rect 45560 20927 45612 20936
rect 45560 20893 45569 20927
rect 45569 20893 45603 20927
rect 45603 20893 45612 20927
rect 45560 20884 45612 20893
rect 45652 20927 45704 20936
rect 45652 20893 45661 20927
rect 45661 20893 45695 20927
rect 45695 20893 45704 20927
rect 45652 20884 45704 20893
rect 48412 20927 48464 20936
rect 48412 20893 48421 20927
rect 48421 20893 48455 20927
rect 48455 20893 48464 20927
rect 48412 20884 48464 20893
rect 48688 20927 48740 20936
rect 48688 20893 48722 20927
rect 48722 20893 48740 20927
rect 48688 20884 48740 20893
rect 55864 20884 55916 20936
rect 56784 20884 56836 20936
rect 56968 20884 57020 20936
rect 56048 20859 56100 20868
rect 56048 20825 56057 20859
rect 56057 20825 56091 20859
rect 56091 20825 56100 20859
rect 56048 20816 56100 20825
rect 48136 20748 48188 20800
rect 56324 20816 56376 20868
rect 56416 20748 56468 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 50294 20646 50346 20698
rect 50358 20646 50410 20698
rect 50422 20646 50474 20698
rect 50486 20646 50538 20698
rect 50550 20646 50602 20698
rect 24308 20544 24360 20596
rect 26608 20587 26660 20596
rect 26608 20553 26617 20587
rect 26617 20553 26651 20587
rect 26651 20553 26660 20587
rect 26608 20544 26660 20553
rect 23664 20519 23716 20528
rect 23664 20485 23673 20519
rect 23673 20485 23707 20519
rect 23707 20485 23716 20519
rect 23664 20476 23716 20485
rect 23940 20476 23992 20528
rect 28816 20544 28868 20596
rect 34428 20544 34480 20596
rect 37464 20544 37516 20596
rect 38844 20544 38896 20596
rect 40408 20544 40460 20596
rect 40868 20544 40920 20596
rect 47768 20544 47820 20596
rect 48780 20544 48832 20596
rect 49148 20587 49200 20596
rect 49148 20553 49157 20587
rect 49157 20553 49191 20587
rect 49191 20553 49200 20587
rect 49148 20544 49200 20553
rect 50528 20544 50580 20596
rect 28172 20519 28224 20528
rect 2964 20408 3016 20460
rect 940 20340 992 20392
rect 24400 20451 24452 20460
rect 24400 20417 24409 20451
rect 24409 20417 24443 20451
rect 24443 20417 24452 20451
rect 24400 20408 24452 20417
rect 24676 20451 24728 20460
rect 24676 20417 24685 20451
rect 24685 20417 24719 20451
rect 24719 20417 24728 20451
rect 24676 20408 24728 20417
rect 28172 20485 28206 20519
rect 28206 20485 28224 20519
rect 28172 20476 28224 20485
rect 28448 20408 28500 20460
rect 28724 20408 28776 20460
rect 29736 20408 29788 20460
rect 30656 20408 30708 20460
rect 33048 20408 33100 20460
rect 34796 20408 34848 20460
rect 35256 20451 35308 20460
rect 35256 20417 35265 20451
rect 35265 20417 35299 20451
rect 35299 20417 35308 20451
rect 35256 20408 35308 20417
rect 35532 20408 35584 20460
rect 27620 20340 27672 20392
rect 27896 20383 27948 20392
rect 27896 20349 27905 20383
rect 27905 20349 27939 20383
rect 27939 20349 27948 20383
rect 27896 20340 27948 20349
rect 31208 20340 31260 20392
rect 32956 20340 33008 20392
rect 35992 20340 36044 20392
rect 36728 20451 36780 20460
rect 36728 20417 36737 20451
rect 36737 20417 36771 20451
rect 36771 20417 36780 20451
rect 36728 20408 36780 20417
rect 37188 20408 37240 20460
rect 37464 20451 37516 20460
rect 37464 20417 37473 20451
rect 37473 20417 37507 20451
rect 37507 20417 37516 20451
rect 37464 20408 37516 20417
rect 41972 20476 42024 20528
rect 38844 20408 38896 20460
rect 38936 20451 38988 20460
rect 38936 20417 38945 20451
rect 38945 20417 38979 20451
rect 38979 20417 38988 20451
rect 38936 20408 38988 20417
rect 38568 20340 38620 20392
rect 38752 20340 38804 20392
rect 39120 20451 39172 20460
rect 39120 20417 39129 20451
rect 39129 20417 39163 20451
rect 39163 20417 39172 20451
rect 39120 20408 39172 20417
rect 39580 20408 39632 20460
rect 39672 20408 39724 20460
rect 40500 20408 40552 20460
rect 41052 20408 41104 20460
rect 41696 20451 41748 20460
rect 41696 20417 41705 20451
rect 41705 20417 41739 20451
rect 41739 20417 41748 20451
rect 41696 20408 41748 20417
rect 42616 20451 42668 20460
rect 42616 20417 42625 20451
rect 42625 20417 42659 20451
rect 42659 20417 42668 20451
rect 42616 20408 42668 20417
rect 44640 20476 44692 20528
rect 48412 20476 48464 20528
rect 43536 20451 43588 20460
rect 43536 20417 43570 20451
rect 43570 20417 43588 20451
rect 41972 20340 42024 20392
rect 43536 20408 43588 20417
rect 24676 20272 24728 20324
rect 17408 20204 17460 20256
rect 23664 20204 23716 20256
rect 28264 20204 28316 20256
rect 28908 20204 28960 20256
rect 34060 20204 34112 20256
rect 36268 20272 36320 20324
rect 36636 20272 36688 20324
rect 37832 20272 37884 20324
rect 41512 20272 41564 20324
rect 34704 20247 34756 20256
rect 34704 20213 34713 20247
rect 34713 20213 34747 20247
rect 34747 20213 34756 20247
rect 34704 20204 34756 20213
rect 35440 20247 35492 20256
rect 35440 20213 35449 20247
rect 35449 20213 35483 20247
rect 35483 20213 35492 20247
rect 35440 20204 35492 20213
rect 37004 20204 37056 20256
rect 41144 20247 41196 20256
rect 41144 20213 41153 20247
rect 41153 20213 41187 20247
rect 41187 20213 41196 20247
rect 41144 20204 41196 20213
rect 41880 20247 41932 20256
rect 41880 20213 41889 20247
rect 41889 20213 41923 20247
rect 41923 20213 41932 20247
rect 41880 20204 41932 20213
rect 42064 20204 42116 20256
rect 45928 20451 45980 20460
rect 45928 20417 45937 20451
rect 45937 20417 45971 20451
rect 45971 20417 45980 20451
rect 45928 20408 45980 20417
rect 47952 20451 48004 20460
rect 47952 20417 47958 20451
rect 47958 20417 47992 20451
rect 47992 20417 48004 20451
rect 47952 20408 48004 20417
rect 48688 20408 48740 20460
rect 49884 20408 49936 20460
rect 51080 20476 51132 20528
rect 53104 20587 53156 20596
rect 53104 20553 53113 20587
rect 53113 20553 53147 20587
rect 53147 20553 53156 20587
rect 53104 20544 53156 20553
rect 57428 20544 57480 20596
rect 55220 20476 55272 20528
rect 50160 20408 50212 20460
rect 44548 20340 44600 20392
rect 45376 20340 45428 20392
rect 44364 20272 44416 20324
rect 52276 20408 52328 20460
rect 53840 20408 53892 20460
rect 55680 20408 55732 20460
rect 55864 20408 55916 20460
rect 44548 20204 44600 20256
rect 44732 20204 44784 20256
rect 53472 20340 53524 20392
rect 53564 20383 53616 20392
rect 53564 20349 53573 20383
rect 53573 20349 53607 20383
rect 53607 20349 53616 20383
rect 53564 20340 53616 20349
rect 53012 20272 53064 20324
rect 53104 20272 53156 20324
rect 56324 20451 56376 20460
rect 56324 20417 56359 20451
rect 56359 20417 56376 20451
rect 56324 20408 56376 20417
rect 57520 20408 57572 20460
rect 58164 20451 58216 20460
rect 58164 20417 58173 20451
rect 58173 20417 58207 20451
rect 58207 20417 58216 20451
rect 58164 20408 58216 20417
rect 51264 20204 51316 20256
rect 52000 20204 52052 20256
rect 53472 20247 53524 20256
rect 53472 20213 53481 20247
rect 53481 20213 53515 20247
rect 53515 20213 53524 20247
rect 53472 20204 53524 20213
rect 56048 20204 56100 20256
rect 56416 20272 56468 20324
rect 56324 20204 56376 20256
rect 57980 20204 58032 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 28448 20043 28500 20052
rect 28448 20009 28457 20043
rect 28457 20009 28491 20043
rect 28491 20009 28500 20043
rect 28448 20000 28500 20009
rect 940 19864 992 19916
rect 22192 19864 22244 19916
rect 23112 19864 23164 19916
rect 28632 20000 28684 20052
rect 28816 20000 28868 20052
rect 30840 20000 30892 20052
rect 31208 20043 31260 20052
rect 31208 20009 31217 20043
rect 31217 20009 31251 20043
rect 31251 20009 31260 20043
rect 31208 20000 31260 20009
rect 28816 19907 28868 19916
rect 28816 19873 28825 19907
rect 28825 19873 28859 19907
rect 28859 19873 28868 19907
rect 28816 19864 28868 19873
rect 28908 19907 28960 19916
rect 28908 19873 28917 19907
rect 28917 19873 28951 19907
rect 28951 19873 28960 19907
rect 28908 19864 28960 19873
rect 22376 19796 22428 19848
rect 24492 19796 24544 19848
rect 24768 19796 24820 19848
rect 17224 19728 17276 19780
rect 24124 19728 24176 19780
rect 25320 19796 25372 19848
rect 26332 19839 26384 19848
rect 26332 19805 26341 19839
rect 26341 19805 26375 19839
rect 26375 19805 26384 19839
rect 26332 19796 26384 19805
rect 27896 19796 27948 19848
rect 25504 19728 25556 19780
rect 27068 19728 27120 19780
rect 940 19660 992 19712
rect 24676 19703 24728 19712
rect 24676 19669 24685 19703
rect 24685 19669 24719 19703
rect 24719 19669 24728 19703
rect 24676 19660 24728 19669
rect 27804 19660 27856 19712
rect 30288 19839 30340 19848
rect 30288 19805 30297 19839
rect 30297 19805 30331 19839
rect 30331 19805 30340 19839
rect 30288 19796 30340 19805
rect 30656 19932 30708 19984
rect 35440 20000 35492 20052
rect 36820 19932 36872 19984
rect 37372 20000 37424 20052
rect 37556 20000 37608 20052
rect 37740 20000 37792 20052
rect 38476 20000 38528 20052
rect 39120 20000 39172 20052
rect 43536 20000 43588 20052
rect 44180 20000 44232 20052
rect 44548 20000 44600 20052
rect 48320 20000 48372 20052
rect 49148 20000 49200 20052
rect 50436 20000 50488 20052
rect 51172 20000 51224 20052
rect 41880 19932 41932 19984
rect 42156 19932 42208 19984
rect 44364 19932 44416 19984
rect 53472 20000 53524 20052
rect 53656 20000 53708 20052
rect 56232 20043 56284 20052
rect 56232 20009 56241 20043
rect 56241 20009 56275 20043
rect 56275 20009 56284 20043
rect 56232 20000 56284 20009
rect 37372 19864 37424 19916
rect 28540 19728 28592 19780
rect 28816 19728 28868 19780
rect 30472 19728 30524 19780
rect 28724 19660 28776 19712
rect 29000 19660 29052 19712
rect 33048 19796 33100 19848
rect 34336 19728 34388 19780
rect 36176 19796 36228 19848
rect 36636 19796 36688 19848
rect 37004 19839 37056 19848
rect 37004 19805 37007 19839
rect 37007 19805 37041 19839
rect 37041 19805 37056 19839
rect 37004 19796 37056 19805
rect 37188 19796 37240 19848
rect 40040 19864 40092 19916
rect 41144 19864 41196 19916
rect 42064 19864 42116 19916
rect 42616 19864 42668 19916
rect 38476 19839 38528 19848
rect 38476 19805 38485 19839
rect 38485 19805 38519 19839
rect 38519 19805 38528 19839
rect 38476 19796 38528 19805
rect 38660 19796 38712 19848
rect 40132 19796 40184 19848
rect 40224 19839 40276 19848
rect 40224 19805 40233 19839
rect 40233 19805 40267 19839
rect 40267 19805 40276 19839
rect 40224 19796 40276 19805
rect 40868 19839 40920 19848
rect 40868 19805 40877 19839
rect 40877 19805 40911 19839
rect 40911 19805 40920 19839
rect 40868 19796 40920 19805
rect 41420 19796 41472 19848
rect 42984 19796 43036 19848
rect 43168 19839 43220 19848
rect 43168 19805 43177 19839
rect 43177 19805 43211 19839
rect 43211 19805 43220 19839
rect 43168 19796 43220 19805
rect 43996 19864 44048 19916
rect 43352 19839 43404 19848
rect 43352 19805 43361 19839
rect 43361 19805 43395 19839
rect 43395 19805 43404 19839
rect 43352 19796 43404 19805
rect 44180 19796 44232 19848
rect 44272 19839 44324 19848
rect 44272 19805 44281 19839
rect 44281 19805 44315 19839
rect 44315 19805 44324 19839
rect 44272 19796 44324 19805
rect 44456 19839 44508 19848
rect 44456 19805 44465 19839
rect 44465 19805 44499 19839
rect 44499 19805 44508 19839
rect 44456 19796 44508 19805
rect 44548 19796 44600 19848
rect 45560 19796 45612 19848
rect 47768 19839 47820 19848
rect 47768 19805 47777 19839
rect 47777 19805 47811 19839
rect 47811 19805 47820 19839
rect 47768 19796 47820 19805
rect 47860 19839 47912 19848
rect 47860 19805 47869 19839
rect 47869 19805 47903 19839
rect 47903 19805 47912 19839
rect 47860 19796 47912 19805
rect 35440 19703 35492 19712
rect 35440 19669 35449 19703
rect 35449 19669 35483 19703
rect 35483 19669 35492 19703
rect 35440 19660 35492 19669
rect 35532 19703 35584 19712
rect 35532 19669 35541 19703
rect 35541 19669 35575 19703
rect 35575 19669 35584 19703
rect 35532 19660 35584 19669
rect 35900 19660 35952 19712
rect 36452 19660 36504 19712
rect 36544 19703 36596 19712
rect 36544 19669 36553 19703
rect 36553 19669 36587 19703
rect 36587 19669 36596 19703
rect 36544 19660 36596 19669
rect 37372 19660 37424 19712
rect 38844 19660 38896 19712
rect 40500 19728 40552 19780
rect 40960 19728 41012 19780
rect 41328 19660 41380 19712
rect 41696 19660 41748 19712
rect 42156 19660 42208 19712
rect 43720 19660 43772 19712
rect 44916 19660 44968 19712
rect 53932 19932 53984 19984
rect 53564 19864 53616 19916
rect 55404 19864 55456 19916
rect 58256 19864 58308 19916
rect 48136 19839 48188 19848
rect 48136 19805 48145 19839
rect 48145 19805 48179 19839
rect 48179 19805 48188 19839
rect 48136 19796 48188 19805
rect 48596 19796 48648 19848
rect 48964 19728 49016 19780
rect 49148 19839 49200 19848
rect 49148 19805 49157 19839
rect 49157 19805 49191 19839
rect 49191 19805 49200 19839
rect 49148 19796 49200 19805
rect 50528 19839 50580 19848
rect 50528 19805 50534 19839
rect 50534 19805 50568 19839
rect 50568 19805 50580 19839
rect 50528 19796 50580 19805
rect 51264 19796 51316 19848
rect 51908 19796 51960 19848
rect 49240 19728 49292 19780
rect 49516 19728 49568 19780
rect 49332 19703 49384 19712
rect 49332 19669 49341 19703
rect 49341 19669 49375 19703
rect 49375 19669 49384 19703
rect 49332 19660 49384 19669
rect 50160 19660 50212 19712
rect 50436 19660 50488 19712
rect 51080 19728 51132 19780
rect 54116 19796 54168 19848
rect 54392 19839 54444 19848
rect 54392 19805 54401 19839
rect 54401 19805 54435 19839
rect 54435 19805 54444 19839
rect 54392 19796 54444 19805
rect 56048 19839 56100 19848
rect 56048 19805 56057 19839
rect 56057 19805 56091 19839
rect 56091 19805 56100 19839
rect 56048 19796 56100 19805
rect 52092 19728 52144 19780
rect 52368 19728 52420 19780
rect 54024 19703 54076 19712
rect 54024 19669 54033 19703
rect 54033 19669 54067 19703
rect 54067 19669 54076 19703
rect 54024 19660 54076 19669
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 50294 19558 50346 19610
rect 50358 19558 50410 19610
rect 50422 19558 50474 19610
rect 50486 19558 50538 19610
rect 50550 19558 50602 19610
rect 1032 19388 1084 19440
rect 18788 19320 18840 19372
rect 20536 19320 20588 19372
rect 22376 19456 22428 19508
rect 24400 19431 24452 19440
rect 24400 19397 24409 19431
rect 24409 19397 24443 19431
rect 24443 19397 24452 19431
rect 24400 19388 24452 19397
rect 27620 19456 27672 19508
rect 28356 19456 28408 19508
rect 28632 19456 28684 19508
rect 34336 19456 34388 19508
rect 29368 19388 29420 19440
rect 34796 19456 34848 19508
rect 36084 19499 36136 19508
rect 36084 19465 36093 19499
rect 36093 19465 36127 19499
rect 36127 19465 36136 19499
rect 36084 19456 36136 19465
rect 37188 19456 37240 19508
rect 37464 19456 37516 19508
rect 37832 19456 37884 19508
rect 23112 19363 23164 19372
rect 23112 19329 23121 19363
rect 23121 19329 23155 19363
rect 23155 19329 23164 19363
rect 23112 19320 23164 19329
rect 11704 19252 11756 19304
rect 24124 19363 24176 19372
rect 24124 19329 24134 19363
rect 24134 19329 24168 19363
rect 24168 19329 24176 19363
rect 24124 19320 24176 19329
rect 24584 19320 24636 19372
rect 25320 19320 25372 19372
rect 22928 19227 22980 19236
rect 22928 19193 22937 19227
rect 22937 19193 22971 19227
rect 22971 19193 22980 19227
rect 22928 19184 22980 19193
rect 22100 19116 22152 19168
rect 28264 19363 28316 19372
rect 28264 19329 28273 19363
rect 28273 19329 28307 19363
rect 28307 19329 28316 19363
rect 28264 19320 28316 19329
rect 30656 19320 30708 19372
rect 33048 19320 33100 19372
rect 34612 19320 34664 19372
rect 35348 19320 35400 19372
rect 35900 19388 35952 19440
rect 36544 19388 36596 19440
rect 35992 19363 36044 19372
rect 35992 19329 36001 19363
rect 36001 19329 36035 19363
rect 36035 19329 36044 19363
rect 35992 19320 36044 19329
rect 37556 19320 37608 19372
rect 38476 19431 38528 19440
rect 38476 19397 38510 19431
rect 38510 19397 38528 19431
rect 38476 19388 38528 19397
rect 40040 19456 40092 19508
rect 40960 19499 41012 19508
rect 40960 19465 40969 19499
rect 40969 19465 41003 19499
rect 41003 19465 41012 19499
rect 40960 19456 41012 19465
rect 41144 19499 41196 19508
rect 41144 19465 41153 19499
rect 41153 19465 41187 19499
rect 41187 19465 41196 19499
rect 41144 19456 41196 19465
rect 44456 19456 44508 19508
rect 38200 19363 38252 19372
rect 38200 19329 38209 19363
rect 38209 19329 38243 19363
rect 38243 19329 38252 19363
rect 38200 19320 38252 19329
rect 28632 19184 28684 19236
rect 36360 19184 36412 19236
rect 36912 19184 36964 19236
rect 40040 19363 40092 19372
rect 40040 19329 40049 19363
rect 40049 19329 40083 19363
rect 40083 19329 40092 19363
rect 40040 19320 40092 19329
rect 40224 19320 40276 19372
rect 41236 19320 41288 19372
rect 42708 19388 42760 19440
rect 43444 19388 43496 19440
rect 39672 19252 39724 19304
rect 41972 19252 42024 19304
rect 43996 19431 44048 19440
rect 43996 19397 44005 19431
rect 44005 19397 44039 19431
rect 44039 19397 44048 19431
rect 46020 19456 46072 19508
rect 49148 19456 49200 19508
rect 49516 19456 49568 19508
rect 50068 19456 50120 19508
rect 44916 19431 44968 19440
rect 43996 19388 44048 19397
rect 44916 19397 44950 19431
rect 44950 19397 44968 19431
rect 44916 19388 44968 19397
rect 46848 19431 46900 19440
rect 46848 19397 46857 19431
rect 46857 19397 46891 19431
rect 46891 19397 46900 19431
rect 46848 19388 46900 19397
rect 48044 19388 48096 19440
rect 44456 19320 44508 19372
rect 44640 19363 44692 19372
rect 44640 19329 44649 19363
rect 44649 19329 44683 19363
rect 44683 19329 44692 19363
rect 44640 19320 44692 19329
rect 44364 19252 44416 19304
rect 48136 19320 48188 19372
rect 48412 19320 48464 19372
rect 49332 19388 49384 19440
rect 49792 19388 49844 19440
rect 50160 19363 50212 19372
rect 50160 19329 50169 19363
rect 50169 19329 50203 19363
rect 50203 19329 50212 19363
rect 50160 19320 50212 19329
rect 52092 19499 52144 19508
rect 52092 19465 52101 19499
rect 52101 19465 52135 19499
rect 52135 19465 52144 19499
rect 52092 19456 52144 19465
rect 51908 19388 51960 19440
rect 53564 19456 53616 19508
rect 54116 19456 54168 19508
rect 56508 19456 56560 19508
rect 56600 19456 56652 19508
rect 57888 19456 57940 19508
rect 52368 19388 52420 19440
rect 52000 19363 52052 19372
rect 52000 19329 52009 19363
rect 52009 19329 52043 19363
rect 52043 19329 52052 19363
rect 52000 19320 52052 19329
rect 52092 19320 52144 19372
rect 53012 19320 53064 19372
rect 55772 19363 55824 19372
rect 55772 19329 55781 19363
rect 55781 19329 55815 19363
rect 55815 19329 55824 19363
rect 55772 19320 55824 19329
rect 55864 19320 55916 19372
rect 58992 19320 59044 19372
rect 52276 19252 52328 19304
rect 41328 19116 41380 19168
rect 41604 19116 41656 19168
rect 44272 19116 44324 19168
rect 46020 19159 46072 19168
rect 46020 19125 46029 19159
rect 46029 19125 46063 19159
rect 46063 19125 46072 19159
rect 46020 19116 46072 19125
rect 47124 19184 47176 19236
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 20720 18912 20772 18964
rect 26424 18912 26476 18964
rect 27068 18955 27120 18964
rect 27068 18921 27077 18955
rect 27077 18921 27111 18955
rect 27111 18921 27120 18955
rect 27068 18912 27120 18921
rect 34428 18912 34480 18964
rect 35348 18912 35400 18964
rect 36544 18955 36596 18964
rect 36544 18921 36553 18955
rect 36553 18921 36587 18955
rect 36587 18921 36596 18955
rect 36544 18912 36596 18921
rect 24768 18844 24820 18896
rect 22100 18776 22152 18828
rect 24400 18776 24452 18828
rect 12256 18708 12308 18760
rect 20812 18751 20864 18760
rect 20812 18717 20821 18751
rect 20821 18717 20855 18751
rect 20855 18717 20864 18751
rect 20812 18708 20864 18717
rect 21548 18708 21600 18760
rect 21732 18708 21784 18760
rect 24584 18708 24636 18760
rect 940 18640 992 18692
rect 24860 18640 24912 18692
rect 27620 18751 27672 18760
rect 27620 18717 27629 18751
rect 27629 18717 27663 18751
rect 27663 18717 27672 18751
rect 27620 18708 27672 18717
rect 33416 18844 33468 18896
rect 34796 18844 34848 18896
rect 35992 18844 36044 18896
rect 38476 18912 38528 18964
rect 40408 18912 40460 18964
rect 45928 18912 45980 18964
rect 47124 18912 47176 18964
rect 55680 18912 55732 18964
rect 33876 18776 33928 18828
rect 26332 18572 26384 18624
rect 29552 18640 29604 18692
rect 32496 18751 32548 18760
rect 32496 18717 32505 18751
rect 32505 18717 32539 18751
rect 32539 18717 32548 18751
rect 32496 18708 32548 18717
rect 34888 18708 34940 18760
rect 35716 18751 35768 18760
rect 35716 18717 35725 18751
rect 35725 18717 35759 18751
rect 35759 18717 35768 18751
rect 35716 18708 35768 18717
rect 36176 18708 36228 18760
rect 36452 18708 36504 18760
rect 27896 18572 27948 18624
rect 32220 18572 32272 18624
rect 34704 18572 34756 18624
rect 38752 18751 38804 18760
rect 38752 18717 38761 18751
rect 38761 18717 38795 18751
rect 38795 18717 38804 18751
rect 38752 18708 38804 18717
rect 39672 18708 39724 18760
rect 36728 18615 36780 18624
rect 36728 18581 36737 18615
rect 36737 18581 36771 18615
rect 36771 18581 36780 18615
rect 36728 18572 36780 18581
rect 39580 18640 39632 18692
rect 40868 18844 40920 18896
rect 40132 18708 40184 18760
rect 41512 18776 41564 18828
rect 41696 18819 41748 18828
rect 41696 18785 41705 18819
rect 41705 18785 41739 18819
rect 41739 18785 41748 18819
rect 41696 18776 41748 18785
rect 45008 18844 45060 18896
rect 52460 18844 52512 18896
rect 56140 18844 56192 18896
rect 46756 18776 46808 18828
rect 48504 18819 48556 18828
rect 48504 18785 48513 18819
rect 48513 18785 48547 18819
rect 48547 18785 48556 18819
rect 48504 18776 48556 18785
rect 49056 18819 49108 18828
rect 49056 18785 49065 18819
rect 49065 18785 49099 18819
rect 49099 18785 49108 18819
rect 49056 18776 49108 18785
rect 55680 18819 55732 18828
rect 55680 18785 55689 18819
rect 55689 18785 55723 18819
rect 55723 18785 55732 18819
rect 55680 18776 55732 18785
rect 40408 18708 40460 18760
rect 41144 18708 41196 18760
rect 42064 18751 42116 18760
rect 42064 18717 42073 18751
rect 42073 18717 42107 18751
rect 42107 18717 42116 18751
rect 42064 18708 42116 18717
rect 42708 18751 42760 18760
rect 42708 18717 42717 18751
rect 42717 18717 42751 18751
rect 42751 18717 42760 18751
rect 42708 18708 42760 18717
rect 43444 18708 43496 18760
rect 46020 18708 46072 18760
rect 38660 18572 38712 18624
rect 38844 18572 38896 18624
rect 39120 18572 39172 18624
rect 41972 18572 42024 18624
rect 42064 18572 42116 18624
rect 46940 18683 46992 18692
rect 46940 18649 46949 18683
rect 46949 18649 46983 18683
rect 46983 18649 46992 18683
rect 46940 18640 46992 18649
rect 43260 18572 43312 18624
rect 46020 18572 46072 18624
rect 47952 18683 48004 18692
rect 47952 18649 47961 18683
rect 47961 18649 47995 18683
rect 47995 18649 48004 18683
rect 47952 18640 48004 18649
rect 48780 18708 48832 18760
rect 54208 18708 54260 18760
rect 58164 18819 58216 18828
rect 58164 18785 58173 18819
rect 58173 18785 58207 18819
rect 58207 18785 58216 18819
rect 58164 18776 58216 18785
rect 56048 18751 56100 18760
rect 56048 18717 56062 18751
rect 56062 18717 56096 18751
rect 56096 18717 56100 18751
rect 56048 18708 56100 18717
rect 56324 18708 56376 18760
rect 56784 18708 56836 18760
rect 56600 18640 56652 18692
rect 49516 18572 49568 18624
rect 58992 18572 59044 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 50294 18470 50346 18522
rect 50358 18470 50410 18522
rect 50422 18470 50474 18522
rect 50486 18470 50538 18522
rect 50550 18470 50602 18522
rect 20904 18368 20956 18420
rect 29552 18368 29604 18420
rect 29644 18411 29696 18420
rect 29644 18377 29653 18411
rect 29653 18377 29687 18411
rect 29687 18377 29696 18411
rect 29644 18368 29696 18377
rect 20536 18300 20588 18352
rect 34612 18368 34664 18420
rect 34980 18368 35032 18420
rect 940 18164 992 18216
rect 22284 18232 22336 18284
rect 24308 18232 24360 18284
rect 26332 18275 26384 18284
rect 26332 18241 26341 18275
rect 26341 18241 26375 18275
rect 26375 18241 26384 18275
rect 26332 18232 26384 18241
rect 27896 18232 27948 18284
rect 29000 18232 29052 18284
rect 29092 18232 29144 18284
rect 29644 18232 29696 18284
rect 30380 18275 30432 18284
rect 30380 18241 30389 18275
rect 30389 18241 30423 18275
rect 30423 18241 30432 18275
rect 30380 18232 30432 18241
rect 32404 18275 32456 18284
rect 32404 18241 32413 18275
rect 32413 18241 32447 18275
rect 32447 18241 32456 18275
rect 32404 18232 32456 18241
rect 24400 18207 24452 18216
rect 24400 18173 24409 18207
rect 24409 18173 24443 18207
rect 24443 18173 24452 18207
rect 24400 18164 24452 18173
rect 24768 18164 24820 18216
rect 26700 18164 26752 18216
rect 34612 18232 34664 18284
rect 34704 18275 34756 18284
rect 34704 18241 34713 18275
rect 34713 18241 34747 18275
rect 34747 18241 34756 18275
rect 34704 18232 34756 18241
rect 35532 18232 35584 18284
rect 36176 18300 36228 18352
rect 37648 18300 37700 18352
rect 39948 18368 40000 18420
rect 40224 18368 40276 18420
rect 41420 18368 41472 18420
rect 42708 18368 42760 18420
rect 37372 18232 37424 18284
rect 36820 18164 36872 18216
rect 37924 18232 37976 18284
rect 39120 18232 39172 18284
rect 44732 18300 44784 18352
rect 45008 18411 45060 18420
rect 45008 18377 45017 18411
rect 45017 18377 45051 18411
rect 45051 18377 45060 18411
rect 45008 18368 45060 18377
rect 45376 18411 45428 18420
rect 45376 18377 45385 18411
rect 45385 18377 45419 18411
rect 45419 18377 45428 18411
rect 45376 18368 45428 18377
rect 46940 18368 46992 18420
rect 47676 18368 47728 18420
rect 48964 18368 49016 18420
rect 51080 18368 51132 18420
rect 55864 18411 55916 18420
rect 55864 18377 55873 18411
rect 55873 18377 55907 18411
rect 55907 18377 55916 18411
rect 55864 18368 55916 18377
rect 56048 18368 56100 18420
rect 41604 18232 41656 18284
rect 40316 18164 40368 18216
rect 41880 18275 41932 18284
rect 41880 18241 41889 18275
rect 41889 18241 41923 18275
rect 41923 18241 41932 18275
rect 41880 18232 41932 18241
rect 43996 18275 44048 18284
rect 43996 18241 44005 18275
rect 44005 18241 44039 18275
rect 44039 18241 44048 18275
rect 43996 18232 44048 18241
rect 44916 18232 44968 18284
rect 48688 18232 48740 18284
rect 50988 18300 51040 18352
rect 52276 18300 52328 18352
rect 48872 18232 48924 18284
rect 49056 18232 49108 18284
rect 49424 18275 49476 18284
rect 49424 18241 49433 18275
rect 49433 18241 49467 18275
rect 49467 18241 49476 18275
rect 49424 18232 49476 18241
rect 55680 18232 55732 18284
rect 56416 18300 56468 18352
rect 56692 18343 56744 18352
rect 56692 18309 56701 18343
rect 56701 18309 56735 18343
rect 56735 18309 56744 18343
rect 56692 18300 56744 18309
rect 56968 18343 57020 18352
rect 56968 18309 56977 18343
rect 56977 18309 57011 18343
rect 57011 18309 57020 18343
rect 56968 18300 57020 18309
rect 41972 18164 42024 18216
rect 42616 18164 42668 18216
rect 43076 18164 43128 18216
rect 43904 18207 43956 18216
rect 43904 18173 43913 18207
rect 43913 18173 43947 18207
rect 43947 18173 43956 18207
rect 43904 18164 43956 18173
rect 45100 18164 45152 18216
rect 45468 18207 45520 18216
rect 45468 18173 45477 18207
rect 45477 18173 45511 18207
rect 45511 18173 45520 18207
rect 45468 18164 45520 18173
rect 46940 18164 46992 18216
rect 48504 18207 48556 18216
rect 48504 18173 48513 18207
rect 48513 18173 48547 18207
rect 48547 18173 48556 18207
rect 48504 18164 48556 18173
rect 18604 18028 18656 18080
rect 24124 18028 24176 18080
rect 24768 18028 24820 18080
rect 26884 18028 26936 18080
rect 30104 18028 30156 18080
rect 30656 18028 30708 18080
rect 32588 18071 32640 18080
rect 32588 18037 32597 18071
rect 32597 18037 32631 18071
rect 32631 18037 32640 18071
rect 32588 18028 32640 18037
rect 32680 18028 32732 18080
rect 37464 18096 37516 18148
rect 40132 18096 40184 18148
rect 41696 18096 41748 18148
rect 54392 18096 54444 18148
rect 36636 18028 36688 18080
rect 37556 18028 37608 18080
rect 37832 18028 37884 18080
rect 40868 18028 40920 18080
rect 43076 18028 43128 18080
rect 43444 18071 43496 18080
rect 43444 18037 43453 18071
rect 43453 18037 43487 18071
rect 43487 18037 43496 18071
rect 43444 18028 43496 18037
rect 46480 18028 46532 18080
rect 47860 18071 47912 18080
rect 47860 18037 47869 18071
rect 47869 18037 47903 18071
rect 47903 18037 47912 18071
rect 47860 18028 47912 18037
rect 48320 18028 48372 18080
rect 54944 18028 54996 18080
rect 55404 18096 55456 18148
rect 56416 18096 56468 18148
rect 56692 18071 56744 18080
rect 56692 18037 56701 18071
rect 56701 18037 56735 18071
rect 56735 18037 56744 18071
rect 56692 18028 56744 18037
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 35624 17824 35676 17876
rect 36820 17824 36872 17876
rect 39028 17824 39080 17876
rect 41880 17824 41932 17876
rect 43720 17824 43772 17876
rect 44180 17824 44232 17876
rect 44364 17824 44416 17876
rect 45560 17824 45612 17876
rect 47768 17824 47820 17876
rect 56876 17824 56928 17876
rect 24676 17799 24728 17808
rect 24676 17765 24685 17799
rect 24685 17765 24719 17799
rect 24719 17765 24728 17799
rect 24676 17756 24728 17765
rect 22744 17688 22796 17740
rect 27528 17756 27580 17808
rect 29000 17756 29052 17808
rect 36176 17756 36228 17808
rect 17960 17620 18012 17672
rect 18420 17620 18472 17672
rect 21180 17620 21232 17672
rect 940 17552 992 17604
rect 22652 17620 22704 17672
rect 24584 17663 24636 17672
rect 24584 17629 24593 17663
rect 24593 17629 24627 17663
rect 24627 17629 24636 17663
rect 24584 17620 24636 17629
rect 24768 17620 24820 17672
rect 28264 17688 28316 17740
rect 28356 17688 28408 17740
rect 26148 17663 26200 17672
rect 26148 17629 26157 17663
rect 26157 17629 26191 17663
rect 26191 17629 26200 17663
rect 26148 17620 26200 17629
rect 26240 17620 26292 17672
rect 28540 17663 28592 17672
rect 28540 17629 28549 17663
rect 28549 17629 28583 17663
rect 28583 17629 28592 17663
rect 28540 17620 28592 17629
rect 30104 17620 30156 17672
rect 32680 17688 32732 17740
rect 36084 17688 36136 17740
rect 36268 17731 36320 17740
rect 36268 17697 36277 17731
rect 36277 17697 36311 17731
rect 36311 17697 36320 17731
rect 36268 17688 36320 17697
rect 36912 17799 36964 17808
rect 36912 17765 36921 17799
rect 36921 17765 36955 17799
rect 36955 17765 36964 17799
rect 36912 17756 36964 17765
rect 37188 17688 37240 17740
rect 38568 17756 38620 17808
rect 41972 17756 42024 17808
rect 43904 17756 43956 17808
rect 31760 17620 31812 17672
rect 32128 17663 32180 17672
rect 32128 17629 32137 17663
rect 32137 17629 32171 17663
rect 32171 17629 32180 17663
rect 32128 17620 32180 17629
rect 32956 17620 33008 17672
rect 34796 17620 34848 17672
rect 36544 17620 36596 17672
rect 21640 17552 21692 17604
rect 23756 17552 23808 17604
rect 24216 17552 24268 17604
rect 18328 17484 18380 17536
rect 20352 17484 20404 17536
rect 21364 17527 21416 17536
rect 21364 17493 21373 17527
rect 21373 17493 21407 17527
rect 21407 17493 21416 17527
rect 21364 17484 21416 17493
rect 24032 17484 24084 17536
rect 24768 17484 24820 17536
rect 25872 17484 25924 17536
rect 26608 17552 26660 17604
rect 26240 17484 26292 17536
rect 26516 17484 26568 17536
rect 30012 17484 30064 17536
rect 31576 17527 31628 17536
rect 31576 17493 31585 17527
rect 31585 17493 31619 17527
rect 31619 17493 31628 17527
rect 31576 17484 31628 17493
rect 32312 17527 32364 17536
rect 32312 17493 32321 17527
rect 32321 17493 32355 17527
rect 32355 17493 32364 17527
rect 32312 17484 32364 17493
rect 37372 17620 37424 17672
rect 38476 17663 38528 17672
rect 38476 17629 38485 17663
rect 38485 17629 38519 17663
rect 38519 17629 38528 17663
rect 38476 17620 38528 17629
rect 39672 17552 39724 17604
rect 40224 17663 40276 17672
rect 40224 17629 40233 17663
rect 40233 17629 40267 17663
rect 40267 17629 40276 17663
rect 40224 17620 40276 17629
rect 40408 17731 40460 17740
rect 40408 17697 40417 17731
rect 40417 17697 40451 17731
rect 40451 17697 40460 17731
rect 40408 17688 40460 17697
rect 40500 17688 40552 17740
rect 41328 17688 41380 17740
rect 41880 17620 41932 17672
rect 42248 17663 42300 17672
rect 42248 17629 42257 17663
rect 42257 17629 42291 17663
rect 42291 17629 42300 17663
rect 42248 17620 42300 17629
rect 44180 17688 44232 17740
rect 45468 17688 45520 17740
rect 55772 17756 55824 17808
rect 48964 17688 49016 17740
rect 51080 17688 51132 17740
rect 44088 17620 44140 17672
rect 44456 17620 44508 17672
rect 45652 17663 45704 17672
rect 45652 17629 45661 17663
rect 45661 17629 45695 17663
rect 45695 17629 45704 17663
rect 45652 17620 45704 17629
rect 47584 17620 47636 17672
rect 48412 17663 48464 17672
rect 48412 17629 48421 17663
rect 48421 17629 48455 17663
rect 48455 17629 48464 17663
rect 48412 17620 48464 17629
rect 48872 17620 48924 17672
rect 49056 17663 49108 17672
rect 49056 17629 49065 17663
rect 49065 17629 49099 17663
rect 49099 17629 49108 17663
rect 49056 17620 49108 17629
rect 49240 17663 49292 17672
rect 49240 17629 49249 17663
rect 49249 17629 49283 17663
rect 49283 17629 49292 17663
rect 49240 17620 49292 17629
rect 51724 17620 51776 17672
rect 52000 17620 52052 17672
rect 38108 17484 38160 17536
rect 40868 17484 40920 17536
rect 41236 17527 41288 17536
rect 41236 17493 41245 17527
rect 41245 17493 41279 17527
rect 41279 17493 41288 17527
rect 41236 17484 41288 17493
rect 42616 17552 42668 17604
rect 45284 17595 45336 17604
rect 45284 17561 45293 17595
rect 45293 17561 45327 17595
rect 45327 17561 45336 17595
rect 45284 17552 45336 17561
rect 42708 17484 42760 17536
rect 52092 17484 52144 17536
rect 56416 17663 56468 17672
rect 56416 17629 56425 17663
rect 56425 17629 56459 17663
rect 56459 17629 56468 17663
rect 56416 17620 56468 17629
rect 59452 17620 59504 17672
rect 56692 17484 56744 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 50294 17382 50346 17434
rect 50358 17382 50410 17434
rect 50422 17382 50474 17434
rect 50486 17382 50538 17434
rect 50550 17382 50602 17434
rect 3516 17212 3568 17264
rect 11704 17212 11756 17264
rect 12348 17144 12400 17196
rect 17592 17187 17644 17196
rect 17592 17153 17601 17187
rect 17601 17153 17635 17187
rect 17635 17153 17644 17187
rect 17592 17144 17644 17153
rect 18328 17187 18380 17196
rect 18328 17153 18337 17187
rect 18337 17153 18371 17187
rect 18371 17153 18380 17187
rect 18328 17144 18380 17153
rect 21180 17280 21232 17332
rect 24124 17323 24176 17332
rect 24124 17289 24133 17323
rect 24133 17289 24167 17323
rect 24167 17289 24176 17323
rect 24124 17280 24176 17289
rect 24768 17280 24820 17332
rect 28632 17280 28684 17332
rect 32128 17280 32180 17332
rect 32404 17280 32456 17332
rect 940 17076 992 17128
rect 23572 17144 23624 17196
rect 24124 17144 24176 17196
rect 24308 17144 24360 17196
rect 24584 17144 24636 17196
rect 21364 17076 21416 17128
rect 23020 17076 23072 17128
rect 23664 17008 23716 17060
rect 23940 17119 23949 17128
rect 23949 17119 23983 17128
rect 23983 17119 23992 17128
rect 23940 17076 23992 17119
rect 25688 17144 25740 17196
rect 26608 17187 26660 17196
rect 26608 17153 26617 17187
rect 26617 17153 26651 17187
rect 26651 17153 26660 17187
rect 26608 17144 26660 17153
rect 25780 17076 25832 17128
rect 26148 17076 26200 17128
rect 26792 17076 26844 17128
rect 27528 17144 27580 17196
rect 27620 17187 27672 17196
rect 27620 17153 27629 17187
rect 27629 17153 27663 17187
rect 27663 17153 27672 17187
rect 27620 17144 27672 17153
rect 30012 17212 30064 17264
rect 28264 17076 28316 17128
rect 28724 17119 28776 17128
rect 28724 17085 28733 17119
rect 28733 17085 28767 17119
rect 28767 17085 28776 17119
rect 28724 17076 28776 17085
rect 30656 17187 30708 17196
rect 30656 17153 30665 17187
rect 30665 17153 30699 17187
rect 30699 17153 30708 17187
rect 30656 17144 30708 17153
rect 32220 17212 32272 17264
rect 31576 17144 31628 17196
rect 32956 17144 33008 17196
rect 36084 17280 36136 17332
rect 36544 17280 36596 17332
rect 39028 17280 39080 17332
rect 36912 17212 36964 17264
rect 39672 17280 39724 17332
rect 42616 17323 42668 17332
rect 42616 17289 42625 17323
rect 42625 17289 42659 17323
rect 42659 17289 42668 17323
rect 42616 17280 42668 17289
rect 42708 17280 42760 17332
rect 46112 17280 46164 17332
rect 48504 17280 48556 17332
rect 34796 17144 34848 17196
rect 36176 17144 36228 17196
rect 40316 17212 40368 17264
rect 40776 17212 40828 17264
rect 40868 17212 40920 17264
rect 45652 17212 45704 17264
rect 45744 17212 45796 17264
rect 45928 17212 45980 17264
rect 14924 16940 14976 16992
rect 17408 16940 17460 16992
rect 17500 16940 17552 16992
rect 17868 16940 17920 16992
rect 22468 16940 22520 16992
rect 23480 16940 23532 16992
rect 26332 16940 26384 16992
rect 27160 16983 27212 16992
rect 27160 16949 27169 16983
rect 27169 16949 27203 16983
rect 27203 16949 27212 16983
rect 27160 16940 27212 16949
rect 27252 16940 27304 16992
rect 29736 16940 29788 16992
rect 30840 16983 30892 16992
rect 30840 16949 30849 16983
rect 30849 16949 30883 16983
rect 30883 16949 30892 16983
rect 30840 16940 30892 16949
rect 33324 16940 33376 16992
rect 35900 17119 35952 17128
rect 35900 17085 35909 17119
rect 35909 17085 35943 17119
rect 35943 17085 35952 17119
rect 35900 17076 35952 17085
rect 38568 17187 38620 17196
rect 38568 17153 38577 17187
rect 38577 17153 38611 17187
rect 38611 17153 38620 17187
rect 38568 17144 38620 17153
rect 38752 17187 38804 17196
rect 38752 17153 38761 17187
rect 38761 17153 38795 17187
rect 38795 17153 38804 17187
rect 38752 17144 38804 17153
rect 41236 17144 41288 17196
rect 42800 17144 42852 17196
rect 36544 17008 36596 17060
rect 35900 16940 35952 16992
rect 37832 17076 37884 17128
rect 41880 17076 41932 17128
rect 38476 17008 38528 17060
rect 37648 16983 37700 16992
rect 37648 16949 37657 16983
rect 37657 16949 37691 16983
rect 37691 16949 37700 16983
rect 37648 16940 37700 16949
rect 38660 16940 38712 16992
rect 43076 17187 43128 17196
rect 43076 17153 43085 17187
rect 43085 17153 43119 17187
rect 43119 17153 43128 17187
rect 43076 17144 43128 17153
rect 43260 17187 43312 17196
rect 43260 17153 43269 17187
rect 43269 17153 43303 17187
rect 43303 17153 43312 17187
rect 43260 17144 43312 17153
rect 43720 17144 43772 17196
rect 43076 17008 43128 17060
rect 44088 17187 44140 17196
rect 44088 17153 44097 17187
rect 44097 17153 44131 17187
rect 44131 17153 44140 17187
rect 44088 17144 44140 17153
rect 48320 17144 48372 17196
rect 48504 17144 48556 17196
rect 51724 17323 51776 17332
rect 51724 17289 51733 17323
rect 51733 17289 51767 17323
rect 51767 17289 51776 17323
rect 51724 17280 51776 17289
rect 51080 17212 51132 17264
rect 51172 17212 51224 17264
rect 53012 17280 53064 17332
rect 44180 17076 44232 17128
rect 45284 17076 45336 17128
rect 45652 17076 45704 17128
rect 48228 17076 48280 17128
rect 48412 17076 48464 17128
rect 45560 17008 45612 17060
rect 48964 17076 49016 17128
rect 53472 17144 53524 17196
rect 56140 17187 56192 17196
rect 56140 17153 56149 17187
rect 56149 17153 56183 17187
rect 56183 17153 56192 17187
rect 56140 17144 56192 17153
rect 58164 17255 58216 17264
rect 58164 17221 58173 17255
rect 58173 17221 58207 17255
rect 58207 17221 58216 17255
rect 58164 17212 58216 17221
rect 52276 17051 52328 17060
rect 52276 17017 52285 17051
rect 52285 17017 52319 17051
rect 52319 17017 52328 17051
rect 52276 17008 52328 17017
rect 48412 16940 48464 16992
rect 51540 16940 51592 16992
rect 51908 16940 51960 16992
rect 54668 17076 54720 17128
rect 56048 17076 56100 17128
rect 58256 17144 58308 17196
rect 58992 17076 59044 17128
rect 56232 16940 56284 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 17592 16736 17644 16788
rect 17224 16643 17276 16652
rect 17224 16609 17233 16643
rect 17233 16609 17267 16643
rect 17267 16609 17276 16643
rect 17224 16600 17276 16609
rect 19432 16600 19484 16652
rect 21548 16600 21600 16652
rect 25044 16736 25096 16788
rect 27252 16736 27304 16788
rect 1584 16575 1636 16584
rect 1584 16541 1593 16575
rect 1593 16541 1627 16575
rect 1627 16541 1636 16575
rect 1584 16532 1636 16541
rect 16212 16532 16264 16584
rect 17500 16575 17552 16584
rect 17500 16541 17509 16575
rect 17509 16541 17543 16575
rect 17543 16541 17552 16575
rect 17500 16532 17552 16541
rect 20352 16575 20404 16584
rect 20352 16541 20361 16575
rect 20361 16541 20395 16575
rect 20395 16541 20404 16575
rect 20352 16532 20404 16541
rect 22468 16575 22520 16584
rect 22468 16541 22502 16575
rect 22502 16541 22520 16575
rect 22468 16532 22520 16541
rect 22836 16532 22888 16584
rect 35716 16736 35768 16788
rect 37740 16736 37792 16788
rect 38752 16736 38804 16788
rect 39580 16736 39632 16788
rect 44180 16736 44232 16788
rect 44548 16736 44600 16788
rect 49056 16736 49108 16788
rect 51172 16736 51224 16788
rect 36084 16668 36136 16720
rect 25504 16643 25556 16652
rect 25504 16609 25513 16643
rect 25513 16609 25547 16643
rect 25547 16609 25556 16643
rect 25504 16600 25556 16609
rect 26516 16643 26568 16652
rect 26516 16609 26522 16643
rect 26522 16609 26568 16643
rect 26516 16600 26568 16609
rect 26700 16643 26752 16652
rect 26700 16609 26709 16643
rect 26709 16609 26743 16643
rect 26743 16609 26752 16643
rect 26700 16600 26752 16609
rect 24860 16532 24912 16584
rect 25320 16575 25372 16584
rect 25320 16541 25329 16575
rect 25329 16541 25363 16575
rect 25363 16541 25372 16575
rect 25320 16532 25372 16541
rect 25688 16575 25740 16584
rect 25688 16541 25697 16575
rect 25697 16541 25731 16575
rect 25731 16541 25740 16575
rect 25688 16532 25740 16541
rect 26332 16575 26384 16584
rect 26332 16541 26341 16575
rect 26341 16541 26375 16575
rect 26375 16541 26384 16575
rect 26332 16532 26384 16541
rect 27160 16600 27212 16652
rect 28724 16600 28776 16652
rect 33416 16600 33468 16652
rect 940 16464 992 16516
rect 25596 16464 25648 16516
rect 27252 16464 27304 16516
rect 28356 16532 28408 16584
rect 18696 16396 18748 16448
rect 24768 16396 24820 16448
rect 25872 16396 25924 16448
rect 30104 16464 30156 16516
rect 28172 16396 28224 16448
rect 28540 16396 28592 16448
rect 29092 16439 29144 16448
rect 29092 16405 29101 16439
rect 29101 16405 29135 16439
rect 29135 16405 29144 16439
rect 29092 16396 29144 16405
rect 31116 16439 31168 16448
rect 31116 16405 31125 16439
rect 31125 16405 31159 16439
rect 31159 16405 31168 16439
rect 31116 16396 31168 16405
rect 32680 16532 32732 16584
rect 32956 16532 33008 16584
rect 33692 16575 33744 16584
rect 33692 16541 33701 16575
rect 33701 16541 33735 16575
rect 33735 16541 33744 16575
rect 33692 16532 33744 16541
rect 34796 16532 34848 16584
rect 35900 16532 35952 16584
rect 36268 16532 36320 16584
rect 36728 16668 36780 16720
rect 32312 16464 32364 16516
rect 32772 16396 32824 16448
rect 34520 16464 34572 16516
rect 33876 16439 33928 16448
rect 33876 16405 33885 16439
rect 33885 16405 33919 16439
rect 33919 16405 33928 16439
rect 33876 16396 33928 16405
rect 34244 16396 34296 16448
rect 35164 16507 35216 16516
rect 35164 16473 35173 16507
rect 35173 16473 35207 16507
rect 35207 16473 35216 16507
rect 35164 16464 35216 16473
rect 36912 16532 36964 16584
rect 37556 16600 37608 16652
rect 44456 16668 44508 16720
rect 44640 16668 44692 16720
rect 38108 16643 38160 16652
rect 38108 16609 38117 16643
rect 38117 16609 38151 16643
rect 38151 16609 38160 16643
rect 38108 16600 38160 16609
rect 41144 16600 41196 16652
rect 45192 16643 45244 16652
rect 41052 16532 41104 16584
rect 42248 16532 42300 16584
rect 45192 16609 45201 16643
rect 45201 16609 45235 16643
rect 45235 16609 45244 16643
rect 45192 16600 45244 16609
rect 51540 16668 51592 16720
rect 44272 16575 44324 16584
rect 44272 16541 44281 16575
rect 44281 16541 44315 16575
rect 44315 16541 44324 16575
rect 44272 16532 44324 16541
rect 44364 16575 44416 16584
rect 44364 16541 44373 16575
rect 44373 16541 44407 16575
rect 44407 16541 44416 16575
rect 44364 16532 44416 16541
rect 44456 16575 44508 16584
rect 44456 16541 44465 16575
rect 44465 16541 44499 16575
rect 44499 16541 44508 16575
rect 44456 16532 44508 16541
rect 44732 16532 44784 16584
rect 37372 16464 37424 16516
rect 37740 16464 37792 16516
rect 38568 16464 38620 16516
rect 38752 16464 38804 16516
rect 40040 16439 40092 16448
rect 40040 16405 40049 16439
rect 40049 16405 40083 16439
rect 40083 16405 40092 16439
rect 40040 16396 40092 16405
rect 40132 16396 40184 16448
rect 41972 16464 42024 16516
rect 43352 16507 43404 16516
rect 43352 16473 43361 16507
rect 43361 16473 43395 16507
rect 43395 16473 43404 16507
rect 43352 16464 43404 16473
rect 47124 16507 47176 16516
rect 47124 16473 47133 16507
rect 47133 16473 47167 16507
rect 47167 16473 47176 16507
rect 47124 16464 47176 16473
rect 46572 16439 46624 16448
rect 46572 16405 46581 16439
rect 46581 16405 46615 16439
rect 46615 16405 46624 16439
rect 48412 16507 48464 16516
rect 48412 16473 48421 16507
rect 48421 16473 48455 16507
rect 48455 16473 48464 16507
rect 48412 16464 48464 16473
rect 49240 16532 49292 16584
rect 53472 16736 53524 16788
rect 56784 16736 56836 16788
rect 58256 16779 58308 16788
rect 58256 16745 58265 16779
rect 58265 16745 58299 16779
rect 58299 16745 58308 16779
rect 58256 16736 58308 16745
rect 53012 16668 53064 16720
rect 51816 16575 51868 16584
rect 51816 16541 51825 16575
rect 51825 16541 51859 16575
rect 51859 16541 51868 16575
rect 51816 16532 51868 16541
rect 52092 16575 52144 16584
rect 52092 16541 52126 16575
rect 52126 16541 52144 16575
rect 52092 16532 52144 16541
rect 54668 16575 54720 16584
rect 54668 16541 54677 16575
rect 54677 16541 54711 16575
rect 54711 16541 54720 16575
rect 54668 16532 54720 16541
rect 55956 16600 56008 16652
rect 56048 16643 56100 16652
rect 56048 16609 56057 16643
rect 56057 16609 56091 16643
rect 56091 16609 56100 16643
rect 56048 16600 56100 16609
rect 56232 16575 56284 16584
rect 56232 16541 56241 16575
rect 56241 16541 56275 16575
rect 56275 16541 56284 16575
rect 56232 16532 56284 16541
rect 56876 16643 56928 16652
rect 56876 16609 56885 16643
rect 56885 16609 56919 16643
rect 56919 16609 56928 16643
rect 56876 16600 56928 16609
rect 50988 16464 51040 16516
rect 46572 16396 46624 16405
rect 47676 16396 47728 16448
rect 51080 16396 51132 16448
rect 53656 16396 53708 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 50294 16294 50346 16346
rect 50358 16294 50410 16346
rect 50422 16294 50474 16346
rect 50486 16294 50538 16346
rect 50550 16294 50602 16346
rect 16212 16235 16264 16244
rect 16212 16201 16221 16235
rect 16221 16201 16255 16235
rect 16255 16201 16264 16235
rect 16212 16192 16264 16201
rect 11336 16124 11388 16176
rect 23572 16235 23624 16244
rect 23572 16201 23581 16235
rect 23581 16201 23615 16235
rect 23615 16201 23624 16235
rect 23572 16192 23624 16201
rect 28356 16192 28408 16244
rect 25872 16124 25924 16176
rect 27804 16124 27856 16176
rect 14556 16056 14608 16108
rect 17776 16056 17828 16108
rect 19432 16056 19484 16108
rect 20720 16056 20772 16108
rect 940 15988 992 16040
rect 17224 15988 17276 16040
rect 17684 15988 17736 16040
rect 18420 15988 18472 16040
rect 20352 15988 20404 16040
rect 20628 15988 20680 16040
rect 22284 16031 22336 16040
rect 22284 15997 22293 16031
rect 22293 15997 22327 16031
rect 22327 15997 22336 16031
rect 22284 15988 22336 15997
rect 18236 15852 18288 15904
rect 21364 15920 21416 15972
rect 23112 16031 23164 16040
rect 23112 15997 23121 16031
rect 23121 15997 23155 16031
rect 23155 15997 23164 16031
rect 23112 15988 23164 15997
rect 23388 15963 23440 15972
rect 23388 15929 23397 15963
rect 23397 15929 23431 15963
rect 23431 15929 23440 15963
rect 23388 15920 23440 15929
rect 21180 15895 21232 15904
rect 21180 15861 21189 15895
rect 21189 15861 21223 15895
rect 21223 15861 21232 15895
rect 21180 15852 21232 15861
rect 23480 15852 23532 15904
rect 24124 16056 24176 16108
rect 23848 15988 23900 16040
rect 24400 16056 24452 16108
rect 30840 16124 30892 16176
rect 31392 16167 31444 16176
rect 24308 15988 24360 16040
rect 25504 16031 25556 16040
rect 25504 15997 25529 16031
rect 25529 15997 25556 16031
rect 25504 15988 25556 15997
rect 25964 16031 26016 16040
rect 25964 15997 25973 16031
rect 25973 15997 26007 16031
rect 26007 15997 26016 16031
rect 25964 15988 26016 15997
rect 27896 15988 27948 16040
rect 28172 16099 28224 16108
rect 28172 16065 28181 16099
rect 28181 16065 28215 16099
rect 28215 16065 28224 16099
rect 28172 16056 28224 16065
rect 28264 16099 28316 16108
rect 28264 16065 28273 16099
rect 28273 16065 28307 16099
rect 28307 16065 28316 16099
rect 28264 16056 28316 16065
rect 28356 15988 28408 16040
rect 28724 16031 28776 16040
rect 28724 15997 28733 16031
rect 28733 15997 28767 16031
rect 28767 15997 28776 16031
rect 28724 15988 28776 15997
rect 24952 15920 25004 15972
rect 25044 15920 25096 15972
rect 31024 15988 31076 16040
rect 31392 16133 31401 16167
rect 31401 16133 31435 16167
rect 31435 16133 31444 16167
rect 31392 16124 31444 16133
rect 32496 16192 32548 16244
rect 32128 16124 32180 16176
rect 32588 16124 32640 16176
rect 32680 16099 32732 16108
rect 32680 16065 32689 16099
rect 32689 16065 32723 16099
rect 32723 16065 32732 16099
rect 32680 16056 32732 16065
rect 33508 16056 33560 16108
rect 34612 16235 34664 16244
rect 34612 16201 34621 16235
rect 34621 16201 34655 16235
rect 34655 16201 34664 16235
rect 34612 16192 34664 16201
rect 36912 16192 36964 16244
rect 37464 16192 37516 16244
rect 37740 16192 37792 16244
rect 34704 16099 34756 16108
rect 34704 16065 34713 16099
rect 34713 16065 34747 16099
rect 34747 16065 34756 16099
rect 34704 16056 34756 16065
rect 37648 16124 37700 16176
rect 35532 16056 35584 16108
rect 36820 16056 36872 16108
rect 37832 16099 37884 16108
rect 37832 16065 37841 16099
rect 37841 16065 37875 16099
rect 37875 16065 37884 16099
rect 37832 16056 37884 16065
rect 38660 16124 38712 16176
rect 40040 16124 40092 16176
rect 41788 16192 41840 16244
rect 42800 16192 42852 16244
rect 43076 16124 43128 16176
rect 44364 16124 44416 16176
rect 45192 16124 45244 16176
rect 47124 16192 47176 16244
rect 47768 16192 47820 16244
rect 48136 16192 48188 16244
rect 49516 16192 49568 16244
rect 53656 16235 53708 16244
rect 53656 16201 53665 16235
rect 53665 16201 53699 16235
rect 53699 16201 53708 16235
rect 53656 16192 53708 16201
rect 55956 16192 56008 16244
rect 39764 16056 39816 16108
rect 38568 15988 38620 16040
rect 38660 16031 38712 16040
rect 38660 15997 38669 16031
rect 38669 15997 38703 16031
rect 38703 15997 38712 16031
rect 38660 15988 38712 15997
rect 35164 15920 35216 15972
rect 37924 15920 37976 15972
rect 28264 15852 28316 15904
rect 30288 15852 30340 15904
rect 30380 15852 30432 15904
rect 30656 15852 30708 15904
rect 31024 15852 31076 15904
rect 34704 15852 34756 15904
rect 36084 15852 36136 15904
rect 37740 15852 37792 15904
rect 38200 15852 38252 15904
rect 43352 16056 43404 16108
rect 39948 15988 40000 16040
rect 41696 16031 41748 16040
rect 41696 15997 41705 16031
rect 41705 15997 41739 16031
rect 41739 15997 41748 16031
rect 41696 15988 41748 15997
rect 44180 16099 44232 16108
rect 44180 16065 44189 16099
rect 44189 16065 44223 16099
rect 44223 16065 44232 16099
rect 44180 16056 44232 16065
rect 46756 16099 46808 16108
rect 46756 16065 46765 16099
rect 46765 16065 46799 16099
rect 46799 16065 46808 16099
rect 46756 16056 46808 16065
rect 48320 16124 48372 16176
rect 52460 16124 52512 16176
rect 53564 16124 53616 16176
rect 58164 16167 58216 16176
rect 58164 16133 58173 16167
rect 58173 16133 58207 16167
rect 58207 16133 58216 16167
rect 58164 16124 58216 16133
rect 59084 16124 59136 16176
rect 59728 16124 59780 16176
rect 48044 16099 48096 16108
rect 48044 16065 48078 16099
rect 48078 16065 48096 16099
rect 48044 16056 48096 16065
rect 50160 16056 50212 16108
rect 50620 16056 50672 16108
rect 51080 16056 51132 16108
rect 46572 15988 46624 16040
rect 46848 16031 46900 16040
rect 46848 15997 46857 16031
rect 46857 15997 46891 16031
rect 46891 15997 46900 16031
rect 46848 15988 46900 15997
rect 44088 15920 44140 15972
rect 51816 15988 51868 16040
rect 56876 16056 56928 16108
rect 40040 15895 40092 15904
rect 40040 15861 40049 15895
rect 40049 15861 40083 15895
rect 40083 15861 40092 15895
rect 40040 15852 40092 15861
rect 41236 15895 41288 15904
rect 41236 15861 41245 15895
rect 41245 15861 41279 15895
rect 41279 15861 41288 15895
rect 41236 15852 41288 15861
rect 43076 15852 43128 15904
rect 43260 15852 43312 15904
rect 44732 15852 44784 15904
rect 46388 15895 46440 15904
rect 46388 15861 46397 15895
rect 46397 15861 46431 15895
rect 46431 15861 46440 15895
rect 46388 15852 46440 15861
rect 46572 15852 46624 15904
rect 51540 15852 51592 15904
rect 53472 15895 53524 15904
rect 53472 15861 53481 15895
rect 53481 15861 53515 15895
rect 53515 15861 53524 15895
rect 53472 15852 53524 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 14556 15691 14608 15700
rect 14556 15657 14565 15691
rect 14565 15657 14599 15691
rect 14599 15657 14608 15691
rect 14556 15648 14608 15657
rect 11428 15555 11480 15564
rect 11428 15521 11437 15555
rect 11437 15521 11471 15555
rect 11471 15521 11480 15555
rect 11428 15512 11480 15521
rect 11796 15555 11848 15564
rect 11796 15521 11805 15555
rect 11805 15521 11839 15555
rect 11839 15521 11848 15555
rect 11796 15512 11848 15521
rect 23204 15648 23256 15700
rect 23388 15648 23440 15700
rect 25044 15691 25096 15700
rect 25044 15657 25053 15691
rect 25053 15657 25087 15691
rect 25087 15657 25096 15691
rect 25044 15648 25096 15657
rect 25596 15648 25648 15700
rect 29000 15648 29052 15700
rect 29184 15648 29236 15700
rect 30012 15648 30064 15700
rect 31024 15648 31076 15700
rect 32220 15691 32272 15700
rect 32220 15657 32229 15691
rect 32229 15657 32263 15691
rect 32263 15657 32272 15691
rect 32220 15648 32272 15657
rect 33692 15648 33744 15700
rect 15476 15580 15528 15632
rect 15844 15555 15896 15564
rect 15844 15521 15853 15555
rect 15853 15521 15887 15555
rect 15887 15521 15896 15555
rect 15844 15512 15896 15521
rect 17776 15623 17828 15632
rect 17776 15589 17785 15623
rect 17785 15589 17819 15623
rect 17819 15589 17828 15623
rect 17776 15580 17828 15589
rect 17868 15512 17920 15564
rect 28724 15580 28776 15632
rect 39948 15648 40000 15700
rect 38660 15580 38712 15632
rect 42248 15648 42300 15700
rect 21272 15512 21324 15564
rect 2688 15444 2740 15496
rect 11336 15487 11388 15496
rect 11336 15453 11345 15487
rect 11345 15453 11379 15487
rect 11379 15453 11388 15487
rect 11336 15444 11388 15453
rect 11704 15487 11756 15496
rect 11704 15453 11713 15487
rect 11713 15453 11747 15487
rect 11747 15453 11756 15487
rect 11704 15444 11756 15453
rect 940 15376 992 15428
rect 10508 15376 10560 15428
rect 15660 15444 15712 15496
rect 15752 15487 15804 15496
rect 15752 15453 15761 15487
rect 15761 15453 15795 15487
rect 15795 15453 15804 15487
rect 15752 15444 15804 15453
rect 16212 15444 16264 15496
rect 20720 15444 20772 15496
rect 17960 15376 18012 15428
rect 12256 15308 12308 15360
rect 18420 15419 18472 15428
rect 18420 15385 18429 15419
rect 18429 15385 18463 15419
rect 18463 15385 18472 15419
rect 18420 15376 18472 15385
rect 20628 15376 20680 15428
rect 21456 15487 21508 15496
rect 21456 15453 21465 15487
rect 21465 15453 21499 15487
rect 21499 15453 21508 15487
rect 21456 15444 21508 15453
rect 25044 15512 25096 15564
rect 21640 15376 21692 15428
rect 22192 15376 22244 15428
rect 22376 15376 22428 15428
rect 22744 15376 22796 15428
rect 23112 15376 23164 15428
rect 18604 15351 18656 15360
rect 18604 15317 18613 15351
rect 18613 15317 18647 15351
rect 18647 15317 18656 15351
rect 18604 15308 18656 15317
rect 20260 15308 20312 15360
rect 20996 15308 21048 15360
rect 22468 15351 22520 15360
rect 22468 15317 22477 15351
rect 22477 15317 22511 15351
rect 22511 15317 22520 15351
rect 22468 15308 22520 15317
rect 22560 15351 22612 15360
rect 22560 15317 22569 15351
rect 22569 15317 22603 15351
rect 22603 15317 22612 15351
rect 22560 15308 22612 15317
rect 23480 15487 23532 15496
rect 23480 15453 23489 15487
rect 23489 15453 23523 15487
rect 23523 15453 23532 15487
rect 23480 15444 23532 15453
rect 23756 15376 23808 15428
rect 25504 15419 25556 15428
rect 25504 15385 25513 15419
rect 25513 15385 25547 15419
rect 25547 15385 25556 15419
rect 25504 15376 25556 15385
rect 26700 15376 26752 15428
rect 29276 15512 29328 15564
rect 30656 15512 30708 15564
rect 34704 15512 34756 15564
rect 41696 15580 41748 15632
rect 46848 15580 46900 15632
rect 47492 15580 47544 15632
rect 47768 15580 47820 15632
rect 28908 15487 28960 15496
rect 28908 15453 28917 15487
rect 28917 15453 28951 15487
rect 28951 15453 28960 15487
rect 28908 15444 28960 15453
rect 30196 15444 30248 15496
rect 30932 15487 30984 15496
rect 30932 15453 30941 15487
rect 30941 15453 30975 15487
rect 30975 15453 30984 15487
rect 30932 15444 30984 15453
rect 31024 15444 31076 15496
rect 32956 15444 33008 15496
rect 26148 15308 26200 15360
rect 27896 15308 27948 15360
rect 28264 15308 28316 15360
rect 28356 15351 28408 15360
rect 28356 15317 28365 15351
rect 28365 15317 28399 15351
rect 28399 15317 28408 15351
rect 33508 15376 33560 15428
rect 34796 15444 34848 15496
rect 38476 15444 38528 15496
rect 45192 15512 45244 15564
rect 40776 15444 40828 15496
rect 41236 15444 41288 15496
rect 46388 15444 46440 15496
rect 47492 15487 47544 15496
rect 47492 15453 47501 15487
rect 47501 15453 47535 15487
rect 47535 15453 47544 15487
rect 47492 15444 47544 15453
rect 47676 15487 47728 15496
rect 47676 15453 47685 15487
rect 47685 15453 47719 15487
rect 47719 15453 47728 15487
rect 47676 15444 47728 15453
rect 51908 15648 51960 15700
rect 48136 15487 48188 15496
rect 48136 15453 48145 15487
rect 48145 15453 48179 15487
rect 48179 15453 48188 15487
rect 48136 15444 48188 15453
rect 55864 15580 55916 15632
rect 56140 15580 56192 15632
rect 51540 15512 51592 15564
rect 37832 15376 37884 15428
rect 28356 15308 28408 15317
rect 29828 15308 29880 15360
rect 29920 15308 29972 15360
rect 31024 15308 31076 15360
rect 31392 15308 31444 15360
rect 32128 15308 32180 15360
rect 38200 15351 38252 15360
rect 38200 15317 38209 15351
rect 38209 15317 38243 15351
rect 38243 15317 38252 15351
rect 38200 15308 38252 15317
rect 38384 15308 38436 15360
rect 39764 15376 39816 15428
rect 43076 15376 43128 15428
rect 43536 15376 43588 15428
rect 46572 15376 46624 15428
rect 44364 15351 44416 15360
rect 44364 15317 44373 15351
rect 44373 15317 44407 15351
rect 44407 15317 44416 15351
rect 44364 15308 44416 15317
rect 44456 15308 44508 15360
rect 47952 15419 48004 15428
rect 47952 15385 47987 15419
rect 47987 15385 48004 15419
rect 51080 15487 51132 15496
rect 51080 15453 51089 15487
rect 51089 15453 51123 15487
rect 51123 15453 51132 15487
rect 51080 15444 51132 15453
rect 47952 15376 48004 15385
rect 46848 15308 46900 15360
rect 51172 15376 51224 15428
rect 52092 15444 52144 15496
rect 54484 15444 54536 15496
rect 51908 15376 51960 15428
rect 58164 15419 58216 15428
rect 58164 15385 58173 15419
rect 58173 15385 58207 15419
rect 58207 15385 58216 15419
rect 58164 15376 58216 15385
rect 48872 15308 48924 15360
rect 49240 15308 49292 15360
rect 50068 15308 50120 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 50294 15206 50346 15258
rect 50358 15206 50410 15258
rect 50422 15206 50474 15258
rect 50486 15206 50538 15258
rect 50550 15206 50602 15258
rect 12348 15104 12400 15156
rect 15752 15104 15804 15156
rect 17408 15104 17460 15156
rect 5448 15036 5500 15088
rect 12440 14968 12492 15020
rect 15752 14968 15804 15020
rect 17868 15036 17920 15088
rect 20352 15104 20404 15156
rect 20812 15104 20864 15156
rect 21456 15104 21508 15156
rect 23940 15104 23992 15156
rect 24124 15104 24176 15156
rect 940 14900 992 14952
rect 15476 14943 15528 14952
rect 15476 14909 15485 14943
rect 15485 14909 15519 14943
rect 15519 14909 15528 14943
rect 15476 14900 15528 14909
rect 15568 14943 15620 14952
rect 15568 14909 15577 14943
rect 15577 14909 15611 14943
rect 15611 14909 15620 14943
rect 15568 14900 15620 14909
rect 18604 14968 18656 15020
rect 20260 15011 20312 15020
rect 20260 14977 20269 15011
rect 20269 14977 20303 15011
rect 20303 14977 20312 15011
rect 20260 14968 20312 14977
rect 20996 15011 21048 15020
rect 20996 14977 21005 15011
rect 21005 14977 21039 15011
rect 21039 14977 21048 15011
rect 20996 14968 21048 14977
rect 22652 15036 22704 15088
rect 22744 15079 22796 15088
rect 22744 15045 22753 15079
rect 22753 15045 22787 15079
rect 22787 15045 22796 15079
rect 22744 15036 22796 15045
rect 27896 15104 27948 15156
rect 28540 15104 28592 15156
rect 30104 15147 30156 15156
rect 30104 15113 30113 15147
rect 30113 15113 30147 15147
rect 30147 15113 30156 15147
rect 30104 15104 30156 15113
rect 24584 15036 24636 15088
rect 32404 15104 32456 15156
rect 23204 15011 23256 15020
rect 23204 14977 23213 15011
rect 23213 14977 23247 15011
rect 23247 14977 23256 15011
rect 23204 14968 23256 14977
rect 23940 14968 23992 15020
rect 25412 14968 25464 15020
rect 25872 15011 25924 15020
rect 25872 14977 25881 15011
rect 25881 14977 25915 15011
rect 25915 14977 25924 15011
rect 25872 14968 25924 14977
rect 21732 14900 21784 14952
rect 22008 14943 22060 14952
rect 22008 14909 22017 14943
rect 22017 14909 22051 14943
rect 22051 14909 22060 14943
rect 22008 14900 22060 14909
rect 22376 14943 22428 14952
rect 22376 14909 22385 14943
rect 22385 14909 22419 14943
rect 22419 14909 22428 14943
rect 22376 14900 22428 14909
rect 25136 14900 25188 14952
rect 17500 14764 17552 14816
rect 24676 14832 24728 14884
rect 25320 14943 25372 14952
rect 25320 14909 25329 14943
rect 25329 14909 25363 14943
rect 25363 14909 25372 14943
rect 25320 14900 25372 14909
rect 25688 14900 25740 14952
rect 28448 15011 28500 15020
rect 28448 14977 28457 15011
rect 28457 14977 28491 15011
rect 28491 14977 28500 15011
rect 28448 14968 28500 14977
rect 26516 14943 26568 14952
rect 26516 14909 26525 14943
rect 26525 14909 26559 14943
rect 26559 14909 26568 14943
rect 26516 14900 26568 14909
rect 28908 14900 28960 14952
rect 25872 14832 25924 14884
rect 21088 14764 21140 14816
rect 22652 14764 22704 14816
rect 23204 14764 23256 14816
rect 24124 14764 24176 14816
rect 24492 14764 24544 14816
rect 27068 14832 27120 14884
rect 29920 15011 29972 15020
rect 29920 14977 29929 15011
rect 29929 14977 29963 15011
rect 29963 14977 29972 15011
rect 29920 14968 29972 14977
rect 31760 14968 31812 15020
rect 32404 14968 32456 15020
rect 33600 15011 33652 15020
rect 33600 14977 33609 15011
rect 33609 14977 33643 15011
rect 33643 14977 33652 15011
rect 33600 14968 33652 14977
rect 33692 14968 33744 15020
rect 36360 15036 36412 15088
rect 38108 15036 38160 15088
rect 34428 15011 34480 15020
rect 34428 14977 34437 15011
rect 34437 14977 34471 15011
rect 34471 14977 34480 15011
rect 34428 14968 34480 14977
rect 37648 15011 37700 15020
rect 37648 14977 37657 15011
rect 37657 14977 37691 15011
rect 37691 14977 37700 15011
rect 37648 14968 37700 14977
rect 38200 14968 38252 15020
rect 42800 15036 42852 15088
rect 43536 15147 43588 15156
rect 43536 15113 43545 15147
rect 43545 15113 43579 15147
rect 43579 15113 43588 15147
rect 43536 15104 43588 15113
rect 44824 15104 44876 15156
rect 44916 15104 44968 15156
rect 44456 15036 44508 15088
rect 44732 15036 44784 15088
rect 40500 14968 40552 15020
rect 29552 14764 29604 14816
rect 29644 14764 29696 14816
rect 30840 14764 30892 14816
rect 31392 14832 31444 14884
rect 43536 14900 43588 14952
rect 44364 14968 44416 15020
rect 44088 14943 44140 14952
rect 44088 14909 44097 14943
rect 44097 14909 44131 14943
rect 44131 14909 44140 14943
rect 44088 14900 44140 14909
rect 48044 15104 48096 15156
rect 50620 15104 50672 15156
rect 49884 15036 49936 15088
rect 50988 15036 51040 15088
rect 54668 15036 54720 15088
rect 45928 14968 45980 15020
rect 47492 14968 47544 15020
rect 50068 14968 50120 15020
rect 31668 14764 31720 14816
rect 33968 14832 34020 14884
rect 49792 14832 49844 14884
rect 50896 14968 50948 15020
rect 54484 15011 54536 15020
rect 54484 14977 54493 15011
rect 54493 14977 54527 15011
rect 54527 14977 54536 15011
rect 54484 14968 54536 14977
rect 54944 15079 54996 15088
rect 54944 15045 54953 15079
rect 54953 15045 54987 15079
rect 54987 15045 54996 15079
rect 54944 15036 54996 15045
rect 58072 15011 58124 15020
rect 58072 14977 58081 15011
rect 58081 14977 58115 15011
rect 58115 14977 58124 15011
rect 58072 14968 58124 14977
rect 52000 14832 52052 14884
rect 56048 14832 56100 14884
rect 34704 14764 34756 14816
rect 38384 14764 38436 14816
rect 39948 14764 40000 14816
rect 40960 14764 41012 14816
rect 58256 14807 58308 14816
rect 58256 14773 58265 14807
rect 58265 14773 58299 14807
rect 58299 14773 58308 14807
rect 58256 14764 58308 14773
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 15660 14560 15712 14612
rect 13360 14492 13412 14544
rect 15108 14424 15160 14476
rect 24584 14560 24636 14612
rect 24952 14560 25004 14612
rect 28448 14560 28500 14612
rect 30932 14560 30984 14612
rect 31116 14603 31168 14612
rect 31116 14569 31125 14603
rect 31125 14569 31159 14603
rect 31159 14569 31168 14603
rect 31116 14560 31168 14569
rect 31760 14603 31812 14612
rect 31760 14569 31769 14603
rect 31769 14569 31803 14603
rect 31803 14569 31812 14603
rect 31760 14560 31812 14569
rect 32128 14560 32180 14612
rect 32680 14560 32732 14612
rect 33692 14560 33744 14612
rect 33784 14560 33836 14612
rect 40500 14603 40552 14612
rect 40500 14569 40509 14603
rect 40509 14569 40543 14603
rect 40543 14569 40552 14603
rect 40500 14560 40552 14569
rect 17684 14535 17736 14544
rect 17684 14501 17693 14535
rect 17693 14501 17727 14535
rect 17727 14501 17736 14535
rect 17684 14492 17736 14501
rect 18788 14492 18840 14544
rect 21272 14535 21324 14544
rect 21272 14501 21281 14535
rect 21281 14501 21315 14535
rect 21315 14501 21324 14535
rect 21272 14492 21324 14501
rect 21640 14492 21692 14544
rect 29644 14492 29696 14544
rect 30840 14492 30892 14544
rect 5448 14356 5500 14408
rect 15016 14399 15068 14408
rect 15016 14365 15025 14399
rect 15025 14365 15059 14399
rect 15059 14365 15068 14399
rect 15016 14356 15068 14365
rect 17316 14424 17368 14476
rect 17408 14424 17460 14476
rect 22284 14424 22336 14476
rect 22376 14424 22428 14476
rect 940 14288 992 14340
rect 12532 14288 12584 14340
rect 17500 14399 17552 14408
rect 17500 14365 17509 14399
rect 17509 14365 17543 14399
rect 17543 14365 17552 14399
rect 17500 14356 17552 14365
rect 15844 14331 15896 14340
rect 15844 14297 15853 14331
rect 15853 14297 15887 14331
rect 15887 14297 15896 14331
rect 15844 14288 15896 14297
rect 20444 14331 20496 14340
rect 20444 14297 20493 14331
rect 20493 14297 20496 14331
rect 20444 14288 20496 14297
rect 20628 14331 20680 14340
rect 20628 14297 20637 14331
rect 20637 14297 20671 14331
rect 20671 14297 20680 14331
rect 20628 14288 20680 14297
rect 21088 14399 21140 14408
rect 21088 14365 21097 14399
rect 21097 14365 21131 14399
rect 21131 14365 21140 14399
rect 21088 14356 21140 14365
rect 25412 14424 25464 14476
rect 26884 14467 26936 14476
rect 26884 14433 26893 14467
rect 26893 14433 26927 14467
rect 26927 14433 26936 14467
rect 26884 14424 26936 14433
rect 25044 14399 25096 14408
rect 25044 14365 25053 14399
rect 25053 14365 25087 14399
rect 25087 14365 25096 14399
rect 25044 14356 25096 14365
rect 26516 14356 26568 14408
rect 26608 14356 26660 14408
rect 28816 14356 28868 14408
rect 29460 14356 29512 14408
rect 25228 14288 25280 14340
rect 27712 14288 27764 14340
rect 29552 14288 29604 14340
rect 31116 14356 31168 14408
rect 29828 14288 29880 14340
rect 14464 14220 14516 14272
rect 15108 14263 15160 14272
rect 15108 14229 15117 14263
rect 15117 14229 15151 14263
rect 15151 14229 15160 14263
rect 15108 14220 15160 14229
rect 23388 14220 23440 14272
rect 23664 14220 23716 14272
rect 26240 14263 26292 14272
rect 26240 14229 26249 14263
rect 26249 14229 26283 14263
rect 26283 14229 26292 14263
rect 26240 14220 26292 14229
rect 29092 14220 29144 14272
rect 29184 14220 29236 14272
rect 30104 14288 30156 14340
rect 30196 14288 30248 14340
rect 31116 14220 31168 14272
rect 31300 14220 31352 14272
rect 34428 14492 34480 14544
rect 33232 14399 33284 14408
rect 33232 14365 33241 14399
rect 33241 14365 33275 14399
rect 33275 14365 33284 14399
rect 33232 14356 33284 14365
rect 32588 14288 32640 14340
rect 33784 14356 33836 14408
rect 34520 14356 34572 14408
rect 35348 14356 35400 14408
rect 34060 14220 34112 14272
rect 35808 14492 35860 14544
rect 44916 14560 44968 14612
rect 59544 14560 59596 14612
rect 40960 14467 41012 14476
rect 40960 14433 40969 14467
rect 40969 14433 41003 14467
rect 41003 14433 41012 14467
rect 40960 14424 41012 14433
rect 41144 14467 41196 14476
rect 41144 14433 41153 14467
rect 41153 14433 41187 14467
rect 41187 14433 41196 14467
rect 41144 14424 41196 14433
rect 45284 14424 45336 14476
rect 48412 14424 48464 14476
rect 46848 14288 46900 14340
rect 49792 14399 49844 14408
rect 49792 14365 49801 14399
rect 49801 14365 49835 14399
rect 49835 14365 49844 14399
rect 49792 14356 49844 14365
rect 50160 14356 50212 14408
rect 50068 14220 50120 14272
rect 51724 14263 51776 14272
rect 51724 14229 51733 14263
rect 51733 14229 51767 14263
rect 51767 14229 51776 14263
rect 58164 14331 58216 14340
rect 58164 14297 58173 14331
rect 58173 14297 58207 14331
rect 58207 14297 58216 14331
rect 58164 14288 58216 14297
rect 51724 14220 51776 14229
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 50294 14118 50346 14170
rect 50358 14118 50410 14170
rect 50422 14118 50474 14170
rect 50486 14118 50538 14170
rect 50550 14118 50602 14170
rect 15568 14059 15620 14068
rect 15568 14025 15577 14059
rect 15577 14025 15611 14059
rect 15611 14025 15620 14059
rect 15568 14016 15620 14025
rect 20720 14016 20772 14068
rect 22284 14016 22336 14068
rect 26332 14016 26384 14068
rect 26608 14059 26660 14068
rect 26608 14025 26617 14059
rect 26617 14025 26651 14059
rect 26651 14025 26660 14059
rect 26608 14016 26660 14025
rect 27712 14059 27764 14068
rect 27712 14025 27721 14059
rect 27721 14025 27755 14059
rect 27755 14025 27764 14059
rect 27712 14016 27764 14025
rect 29184 14016 29236 14068
rect 30196 14016 30248 14068
rect 31024 14016 31076 14068
rect 31668 14016 31720 14068
rect 15476 13948 15528 14000
rect 17316 13948 17368 14000
rect 940 13812 992 13864
rect 22192 13880 22244 13932
rect 22468 13880 22520 13932
rect 22100 13812 22152 13864
rect 24124 13948 24176 14000
rect 24860 13948 24912 14000
rect 25964 13948 26016 14000
rect 23940 13923 23992 13932
rect 23940 13889 23949 13923
rect 23949 13889 23983 13923
rect 23983 13889 23992 13923
rect 23940 13880 23992 13889
rect 24492 13880 24544 13932
rect 25228 13923 25280 13932
rect 25228 13889 25237 13923
rect 25237 13889 25271 13923
rect 25271 13889 25280 13923
rect 25228 13880 25280 13889
rect 26240 13880 26292 13932
rect 29828 13948 29880 14000
rect 28908 13880 28960 13932
rect 24308 13812 24360 13864
rect 26332 13812 26384 13864
rect 28724 13812 28776 13864
rect 15292 13744 15344 13796
rect 22744 13744 22796 13796
rect 23572 13676 23624 13728
rect 24216 13676 24268 13728
rect 28816 13744 28868 13796
rect 29552 13923 29604 13932
rect 29552 13889 29561 13923
rect 29561 13889 29595 13923
rect 29595 13889 29604 13923
rect 29552 13880 29604 13889
rect 29644 13880 29696 13932
rect 29920 13880 29972 13932
rect 31392 13923 31444 13932
rect 31392 13889 31401 13923
rect 31401 13889 31435 13923
rect 31435 13889 31444 13923
rect 31392 13880 31444 13889
rect 30104 13812 30156 13864
rect 30656 13812 30708 13864
rect 32588 13923 32640 13932
rect 32588 13889 32597 13923
rect 32597 13889 32631 13923
rect 32631 13889 32640 13923
rect 32588 13880 32640 13889
rect 32864 13923 32916 13932
rect 32864 13889 32873 13923
rect 32873 13889 32907 13923
rect 32907 13889 32916 13923
rect 32864 13880 32916 13889
rect 33324 13923 33376 13932
rect 33324 13889 33333 13923
rect 33333 13889 33367 13923
rect 33367 13889 33376 13923
rect 33324 13880 33376 13889
rect 33784 13880 33836 13932
rect 34060 13880 34112 13932
rect 35348 14059 35400 14068
rect 35348 14025 35357 14059
rect 35357 14025 35391 14059
rect 35391 14025 35400 14059
rect 35348 14016 35400 14025
rect 38936 14016 38988 14068
rect 34428 13948 34480 14000
rect 44916 13948 44968 14000
rect 46664 13948 46716 14000
rect 49884 13991 49936 14000
rect 49884 13957 49893 13991
rect 49893 13957 49927 13991
rect 49927 13957 49936 13991
rect 49884 13948 49936 13957
rect 50896 14016 50948 14068
rect 58256 13948 58308 14000
rect 35808 13880 35860 13932
rect 42708 13880 42760 13932
rect 43168 13880 43220 13932
rect 30380 13744 30432 13796
rect 37924 13855 37976 13864
rect 37924 13821 37933 13855
rect 37933 13821 37967 13855
rect 37967 13821 37976 13855
rect 37924 13812 37976 13821
rect 38108 13855 38160 13864
rect 38108 13821 38117 13855
rect 38117 13821 38151 13855
rect 38151 13821 38160 13855
rect 38108 13812 38160 13821
rect 38476 13812 38528 13864
rect 50068 13812 50120 13864
rect 32680 13744 32732 13796
rect 51724 13880 51776 13932
rect 56416 13923 56468 13932
rect 56416 13889 56425 13923
rect 56425 13889 56459 13923
rect 56459 13889 56468 13923
rect 56416 13880 56468 13889
rect 57060 13923 57112 13932
rect 57060 13889 57069 13923
rect 57069 13889 57103 13923
rect 57103 13889 57112 13923
rect 57060 13880 57112 13889
rect 58072 13923 58124 13932
rect 58072 13889 58081 13923
rect 58081 13889 58115 13923
rect 58115 13889 58124 13923
rect 58072 13880 58124 13889
rect 50620 13812 50672 13864
rect 51080 13812 51132 13864
rect 56232 13855 56284 13864
rect 56232 13821 56241 13855
rect 56241 13821 56275 13855
rect 56275 13821 56284 13855
rect 56232 13812 56284 13821
rect 58992 13812 59044 13864
rect 58164 13744 58216 13796
rect 30012 13676 30064 13728
rect 31760 13676 31812 13728
rect 34152 13676 34204 13728
rect 37464 13719 37516 13728
rect 37464 13685 37473 13719
rect 37473 13685 37507 13719
rect 37507 13685 37516 13719
rect 37464 13676 37516 13685
rect 43904 13676 43956 13728
rect 56600 13719 56652 13728
rect 56600 13685 56609 13719
rect 56609 13685 56643 13719
rect 56643 13685 56652 13719
rect 56600 13676 56652 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 16212 13515 16264 13524
rect 16212 13481 16221 13515
rect 16221 13481 16255 13515
rect 16255 13481 16264 13515
rect 16212 13472 16264 13481
rect 21364 13472 21416 13524
rect 21456 13472 21508 13524
rect 28172 13472 28224 13524
rect 29276 13472 29328 13524
rect 32588 13472 32640 13524
rect 34060 13472 34112 13524
rect 16028 13447 16080 13456
rect 16028 13413 16037 13447
rect 16037 13413 16071 13447
rect 16071 13413 16080 13447
rect 16028 13404 16080 13413
rect 23112 13404 23164 13456
rect 24124 13404 24176 13456
rect 15476 13336 15528 13388
rect 4252 13268 4304 13320
rect 8484 13268 8536 13320
rect 23756 13336 23808 13388
rect 24584 13336 24636 13388
rect 25228 13379 25280 13388
rect 25228 13345 25237 13379
rect 25237 13345 25271 13379
rect 25271 13345 25280 13379
rect 25228 13336 25280 13345
rect 22560 13268 22612 13320
rect 23664 13311 23716 13320
rect 23664 13277 23673 13311
rect 23673 13277 23707 13311
rect 23707 13277 23716 13311
rect 23664 13268 23716 13277
rect 940 13200 992 13252
rect 20536 13200 20588 13252
rect 23296 13132 23348 13184
rect 25320 13132 25372 13184
rect 27160 13404 27212 13456
rect 37924 13472 37976 13524
rect 48320 13472 48372 13524
rect 49884 13404 49936 13456
rect 56416 13472 56468 13524
rect 57704 13472 57756 13524
rect 26884 13336 26936 13388
rect 27896 13336 27948 13388
rect 28816 13200 28868 13252
rect 30288 13268 30340 13320
rect 30656 13268 30708 13320
rect 28172 13132 28224 13184
rect 30380 13132 30432 13184
rect 33416 13268 33468 13320
rect 34428 13336 34480 13388
rect 37188 13336 37240 13388
rect 49792 13336 49844 13388
rect 34060 13311 34112 13320
rect 34060 13277 34069 13311
rect 34069 13277 34103 13311
rect 34103 13277 34112 13311
rect 34060 13268 34112 13277
rect 34152 13311 34204 13320
rect 34152 13277 34161 13311
rect 34161 13277 34195 13311
rect 34195 13277 34204 13311
rect 34152 13268 34204 13277
rect 34244 13268 34296 13320
rect 36268 13268 36320 13320
rect 37464 13268 37516 13320
rect 51540 13336 51592 13388
rect 32312 13200 32364 13252
rect 41144 13200 41196 13252
rect 43352 13200 43404 13252
rect 36912 13132 36964 13184
rect 43076 13175 43128 13184
rect 43076 13141 43085 13175
rect 43085 13141 43119 13175
rect 43119 13141 43128 13175
rect 43076 13132 43128 13141
rect 44180 13132 44232 13184
rect 49424 13200 49476 13252
rect 49792 13200 49844 13252
rect 50620 13311 50672 13320
rect 50620 13277 50629 13311
rect 50629 13277 50663 13311
rect 50663 13277 50672 13311
rect 50620 13268 50672 13277
rect 55864 13311 55916 13320
rect 55864 13277 55873 13311
rect 55873 13277 55907 13311
rect 55907 13277 55916 13311
rect 55864 13268 55916 13277
rect 47492 13132 47544 13184
rect 50160 13132 50212 13184
rect 50896 13243 50948 13252
rect 50896 13209 50905 13243
rect 50905 13209 50939 13243
rect 50939 13209 50948 13243
rect 50896 13200 50948 13209
rect 51724 13200 51776 13252
rect 55956 13243 56008 13252
rect 55956 13209 55965 13243
rect 55965 13209 55999 13243
rect 55999 13209 56008 13243
rect 55956 13200 56008 13209
rect 56784 13379 56836 13388
rect 56784 13345 56793 13379
rect 56793 13345 56827 13379
rect 56827 13345 56836 13379
rect 56784 13336 56836 13345
rect 56140 13243 56192 13252
rect 56140 13209 56175 13243
rect 56175 13209 56192 13243
rect 56600 13268 56652 13320
rect 56140 13200 56192 13209
rect 57704 13200 57756 13252
rect 57152 13132 57204 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 50294 13030 50346 13082
rect 50358 13030 50410 13082
rect 50422 13030 50474 13082
rect 50486 13030 50538 13082
rect 50550 13030 50602 13082
rect 4252 12860 4304 12912
rect 12348 12792 12400 12844
rect 940 12724 992 12776
rect 20812 12588 20864 12640
rect 22744 12588 22796 12640
rect 23296 12971 23348 12980
rect 23296 12937 23305 12971
rect 23305 12937 23339 12971
rect 23339 12937 23348 12971
rect 23296 12928 23348 12937
rect 23664 12928 23716 12980
rect 26148 12971 26200 12980
rect 26148 12937 26157 12971
rect 26157 12937 26191 12971
rect 26191 12937 26200 12971
rect 26148 12928 26200 12937
rect 26516 12928 26568 12980
rect 26884 12928 26936 12980
rect 29460 12928 29512 12980
rect 30012 12928 30064 12980
rect 35624 12928 35676 12980
rect 23020 12860 23072 12912
rect 24584 12860 24636 12912
rect 30656 12903 30708 12912
rect 30656 12869 30665 12903
rect 30665 12869 30699 12903
rect 30699 12869 30708 12903
rect 30656 12860 30708 12869
rect 31024 12860 31076 12912
rect 23388 12767 23440 12776
rect 23388 12733 23397 12767
rect 23397 12733 23431 12767
rect 23431 12733 23440 12767
rect 23388 12724 23440 12733
rect 25136 12792 25188 12844
rect 25964 12835 26016 12844
rect 25964 12801 25973 12835
rect 25973 12801 26007 12835
rect 26007 12801 26016 12835
rect 25964 12792 26016 12801
rect 29736 12792 29788 12844
rect 30288 12792 30340 12844
rect 30380 12835 30432 12844
rect 30380 12801 30389 12835
rect 30389 12801 30423 12835
rect 30423 12801 30432 12835
rect 30380 12792 30432 12801
rect 31668 12792 31720 12844
rect 33784 12903 33836 12912
rect 33784 12869 33793 12903
rect 33793 12869 33827 12903
rect 33827 12869 33836 12903
rect 33784 12860 33836 12869
rect 43076 12860 43128 12912
rect 49424 12903 49476 12912
rect 49424 12869 49433 12903
rect 49433 12869 49467 12903
rect 49467 12869 49476 12903
rect 49424 12860 49476 12869
rect 51816 12860 51868 12912
rect 55772 12903 55824 12912
rect 55772 12869 55781 12903
rect 55781 12869 55815 12903
rect 55815 12869 55824 12903
rect 55772 12860 55824 12869
rect 57060 12860 57112 12912
rect 57152 12903 57204 12912
rect 57152 12869 57161 12903
rect 57161 12869 57195 12903
rect 57195 12869 57204 12903
rect 57152 12860 57204 12869
rect 37188 12792 37240 12844
rect 39304 12792 39356 12844
rect 42984 12835 43036 12844
rect 42984 12801 42993 12835
rect 42993 12801 43027 12835
rect 43027 12801 43036 12835
rect 42984 12792 43036 12801
rect 46940 12792 46992 12844
rect 47952 12792 48004 12844
rect 55588 12835 55640 12844
rect 55588 12801 55597 12835
rect 55597 12801 55631 12835
rect 55631 12801 55640 12835
rect 55588 12792 55640 12801
rect 25872 12724 25924 12776
rect 34612 12724 34664 12776
rect 36268 12724 36320 12776
rect 37556 12724 37608 12776
rect 38108 12767 38160 12776
rect 38108 12733 38117 12767
rect 38117 12733 38151 12767
rect 38151 12733 38160 12767
rect 38108 12724 38160 12733
rect 29276 12656 29328 12708
rect 40040 12656 40092 12708
rect 43352 12724 43404 12776
rect 45836 12724 45888 12776
rect 50896 12724 50948 12776
rect 56140 12792 56192 12844
rect 56416 12792 56468 12844
rect 56508 12792 56560 12844
rect 58072 12835 58124 12844
rect 58072 12801 58081 12835
rect 58081 12801 58115 12835
rect 58115 12801 58124 12835
rect 58072 12792 58124 12801
rect 43904 12656 43956 12708
rect 51540 12656 51592 12708
rect 55864 12656 55916 12708
rect 25872 12588 25924 12640
rect 26056 12588 26108 12640
rect 32312 12588 32364 12640
rect 36636 12588 36688 12640
rect 38568 12588 38620 12640
rect 41696 12588 41748 12640
rect 43168 12588 43220 12640
rect 56508 12588 56560 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 12348 12384 12400 12436
rect 22560 12384 22612 12436
rect 23664 12384 23716 12436
rect 23940 12384 23992 12436
rect 24768 12384 24820 12436
rect 23020 12316 23072 12368
rect 13544 12291 13596 12300
rect 13544 12257 13553 12291
rect 13553 12257 13587 12291
rect 13587 12257 13596 12291
rect 13544 12248 13596 12257
rect 15476 12248 15528 12300
rect 13084 12180 13136 12232
rect 940 12112 992 12164
rect 13176 12112 13228 12164
rect 13452 12223 13504 12232
rect 13452 12189 13461 12223
rect 13461 12189 13495 12223
rect 13495 12189 13504 12223
rect 13452 12180 13504 12189
rect 13636 12223 13688 12232
rect 13636 12189 13645 12223
rect 13645 12189 13679 12223
rect 13679 12189 13688 12223
rect 13636 12180 13688 12189
rect 23480 12180 23532 12232
rect 23664 12223 23716 12232
rect 23664 12189 23673 12223
rect 23673 12189 23707 12223
rect 23707 12189 23716 12223
rect 23664 12180 23716 12189
rect 24584 12291 24636 12300
rect 24584 12257 24593 12291
rect 24593 12257 24627 12291
rect 24627 12257 24636 12291
rect 24584 12248 24636 12257
rect 26148 12180 26200 12232
rect 28908 12384 28960 12436
rect 29184 12384 29236 12436
rect 35716 12384 35768 12436
rect 38108 12384 38160 12436
rect 56600 12384 56652 12436
rect 57060 12384 57112 12436
rect 32404 12316 32456 12368
rect 37372 12316 37424 12368
rect 39764 12316 39816 12368
rect 31024 12248 31076 12300
rect 42984 12248 43036 12300
rect 44088 12248 44140 12300
rect 50160 12248 50212 12300
rect 55772 12248 55824 12300
rect 56784 12291 56836 12300
rect 56784 12257 56793 12291
rect 56793 12257 56827 12291
rect 56827 12257 56836 12291
rect 56784 12248 56836 12257
rect 30380 12180 30432 12232
rect 30932 12223 30984 12232
rect 30932 12189 30941 12223
rect 30941 12189 30975 12223
rect 30975 12189 30984 12223
rect 30932 12180 30984 12189
rect 31024 12112 31076 12164
rect 23756 12087 23808 12096
rect 23756 12053 23765 12087
rect 23765 12053 23799 12087
rect 23799 12053 23808 12087
rect 23756 12044 23808 12053
rect 23940 12044 23992 12096
rect 30288 12044 30340 12096
rect 31760 12180 31812 12232
rect 32680 12180 32732 12232
rect 32956 12180 33008 12232
rect 36268 12180 36320 12232
rect 37648 12180 37700 12232
rect 41880 12223 41932 12232
rect 41880 12189 41889 12223
rect 41889 12189 41923 12223
rect 41923 12189 41932 12223
rect 41880 12180 41932 12189
rect 44272 12180 44324 12232
rect 47124 12180 47176 12232
rect 49332 12180 49384 12232
rect 37464 12112 37516 12164
rect 32496 12044 32548 12096
rect 41328 12112 41380 12164
rect 37740 12087 37792 12096
rect 37740 12053 37749 12087
rect 37749 12053 37783 12087
rect 37783 12053 37792 12087
rect 37740 12044 37792 12053
rect 41512 12087 41564 12096
rect 41512 12053 41521 12087
rect 41521 12053 41555 12087
rect 41555 12053 41564 12087
rect 41512 12044 41564 12053
rect 41972 12087 42024 12096
rect 41972 12053 41981 12087
rect 41981 12053 42015 12087
rect 42015 12053 42024 12087
rect 41972 12044 42024 12053
rect 42708 12087 42760 12096
rect 42708 12053 42717 12087
rect 42717 12053 42751 12087
rect 42751 12053 42760 12087
rect 42708 12044 42760 12053
rect 43076 12044 43128 12096
rect 49884 12180 49936 12232
rect 54944 12180 54996 12232
rect 56140 12112 56192 12164
rect 56692 12112 56744 12164
rect 51724 12087 51776 12096
rect 51724 12053 51733 12087
rect 51733 12053 51767 12087
rect 51767 12053 51776 12087
rect 51724 12044 51776 12053
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 50294 11942 50346 11994
rect 50358 11942 50410 11994
rect 50422 11942 50474 11994
rect 50486 11942 50538 11994
rect 50550 11942 50602 11994
rect 1584 11840 1636 11892
rect 11704 11840 11756 11892
rect 13084 11883 13136 11892
rect 13084 11849 13093 11883
rect 13093 11849 13127 11883
rect 13127 11849 13136 11883
rect 13084 11840 13136 11849
rect 13452 11840 13504 11892
rect 23296 11840 23348 11892
rect 23664 11840 23716 11892
rect 24952 11840 25004 11892
rect 25412 11840 25464 11892
rect 30656 11840 30708 11892
rect 22744 11772 22796 11824
rect 23940 11815 23992 11824
rect 23940 11781 23949 11815
rect 23949 11781 23983 11815
rect 23983 11781 23992 11815
rect 23940 11772 23992 11781
rect 940 11636 992 11688
rect 13176 11636 13228 11688
rect 13452 11679 13504 11688
rect 13452 11645 13461 11679
rect 13461 11645 13495 11679
rect 13495 11645 13504 11679
rect 13452 11636 13504 11645
rect 13544 11679 13596 11688
rect 13544 11645 13553 11679
rect 13553 11645 13587 11679
rect 13587 11645 13596 11679
rect 13544 11636 13596 11645
rect 18052 11679 18104 11688
rect 18052 11645 18061 11679
rect 18061 11645 18095 11679
rect 18095 11645 18104 11679
rect 18052 11636 18104 11645
rect 18144 11679 18196 11688
rect 18144 11645 18153 11679
rect 18153 11645 18187 11679
rect 18187 11645 18196 11679
rect 18144 11636 18196 11645
rect 20720 11568 20772 11620
rect 25136 11747 25188 11756
rect 25136 11713 25145 11747
rect 25145 11713 25179 11747
rect 25179 11713 25188 11747
rect 25136 11704 25188 11713
rect 29644 11772 29696 11824
rect 29828 11747 29880 11756
rect 29828 11713 29862 11747
rect 29862 11713 29880 11747
rect 29828 11704 29880 11713
rect 31024 11840 31076 11892
rect 32128 11840 32180 11892
rect 37464 11883 37516 11892
rect 37464 11849 37473 11883
rect 37473 11849 37507 11883
rect 37507 11849 37516 11883
rect 37464 11840 37516 11849
rect 38844 11840 38896 11892
rect 42984 11883 43036 11892
rect 42984 11849 42993 11883
rect 42993 11849 43027 11883
rect 43027 11849 43036 11883
rect 42984 11840 43036 11849
rect 47768 11840 47820 11892
rect 49056 11840 49108 11892
rect 56692 11883 56744 11892
rect 56692 11849 56701 11883
rect 56701 11849 56735 11883
rect 56735 11849 56744 11883
rect 56692 11840 56744 11849
rect 32496 11704 32548 11756
rect 32680 11704 32732 11756
rect 32772 11747 32824 11756
rect 32772 11713 32781 11747
rect 32781 11713 32815 11747
rect 32815 11713 32824 11747
rect 32772 11704 32824 11713
rect 34796 11704 34848 11756
rect 35348 11704 35400 11756
rect 36268 11772 36320 11824
rect 37740 11772 37792 11824
rect 41512 11772 41564 11824
rect 46480 11772 46532 11824
rect 36636 11704 36688 11756
rect 37648 11704 37700 11756
rect 29552 11679 29604 11688
rect 29552 11645 29561 11679
rect 29561 11645 29595 11679
rect 29595 11645 29604 11679
rect 29552 11636 29604 11645
rect 30932 11636 30984 11688
rect 31852 11636 31904 11688
rect 32220 11636 32272 11688
rect 42800 11747 42852 11756
rect 42800 11713 42809 11747
rect 42809 11713 42843 11747
rect 42843 11713 42852 11747
rect 42800 11704 42852 11713
rect 45192 11704 45244 11756
rect 46664 11704 46716 11756
rect 34520 11636 34572 11688
rect 29092 11568 29144 11620
rect 38016 11679 38068 11688
rect 38016 11645 38025 11679
rect 38025 11645 38059 11679
rect 38059 11645 38068 11679
rect 38016 11636 38068 11645
rect 38200 11636 38252 11688
rect 40592 11679 40644 11688
rect 40592 11645 40601 11679
rect 40601 11645 40635 11679
rect 40635 11645 40644 11679
rect 40592 11636 40644 11645
rect 42892 11636 42944 11688
rect 44088 11679 44140 11688
rect 44088 11645 44097 11679
rect 44097 11645 44131 11679
rect 44131 11645 44140 11679
rect 44088 11636 44140 11645
rect 23020 11500 23072 11552
rect 28540 11500 28592 11552
rect 28816 11500 28868 11552
rect 31852 11500 31904 11552
rect 35440 11500 35492 11552
rect 39120 11568 39172 11620
rect 55956 11772 56008 11824
rect 48780 11704 48832 11756
rect 54208 11704 54260 11756
rect 56508 11747 56560 11756
rect 56508 11713 56517 11747
rect 56517 11713 56551 11747
rect 56551 11713 56560 11747
rect 56508 11704 56560 11713
rect 58072 11747 58124 11756
rect 58072 11713 58081 11747
rect 58081 11713 58115 11747
rect 58115 11713 58124 11747
rect 58072 11704 58124 11713
rect 49056 11679 49108 11688
rect 49056 11645 49065 11679
rect 49065 11645 49099 11679
rect 49099 11645 49108 11679
rect 49056 11636 49108 11645
rect 37556 11500 37608 11552
rect 37740 11500 37792 11552
rect 41972 11543 42024 11552
rect 41972 11509 41981 11543
rect 41981 11509 42015 11543
rect 42015 11509 42024 11543
rect 41972 11500 42024 11509
rect 48872 11568 48924 11620
rect 56140 11636 56192 11688
rect 45468 11543 45520 11552
rect 45468 11509 45477 11543
rect 45477 11509 45511 11543
rect 45511 11509 45520 11543
rect 45468 11500 45520 11509
rect 48320 11500 48372 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 13636 11296 13688 11348
rect 15476 11339 15528 11348
rect 15476 11305 15485 11339
rect 15485 11305 15519 11339
rect 15519 11305 15528 11339
rect 15476 11296 15528 11305
rect 18144 11296 18196 11348
rect 20628 11296 20680 11348
rect 23388 11296 23440 11348
rect 29828 11296 29880 11348
rect 13176 11228 13228 11280
rect 14464 11203 14516 11212
rect 14464 11169 14473 11203
rect 14473 11169 14507 11203
rect 14507 11169 14516 11203
rect 14464 11160 14516 11169
rect 14556 11203 14608 11212
rect 14556 11169 14565 11203
rect 14565 11169 14599 11203
rect 14599 11169 14608 11203
rect 14556 11160 14608 11169
rect 15936 11228 15988 11280
rect 16120 11160 16172 11212
rect 22192 11228 22244 11280
rect 28540 11228 28592 11280
rect 30472 11296 30524 11348
rect 30104 11228 30156 11280
rect 23848 11203 23900 11212
rect 23848 11169 23857 11203
rect 23857 11169 23891 11203
rect 23891 11169 23900 11203
rect 23848 11160 23900 11169
rect 13452 11092 13504 11144
rect 14740 11135 14792 11144
rect 14740 11101 14749 11135
rect 14749 11101 14783 11135
rect 14783 11101 14792 11135
rect 14740 11092 14792 11101
rect 940 11024 992 11076
rect 12440 11024 12492 11076
rect 15844 11092 15896 11144
rect 29184 11160 29236 11212
rect 29828 11160 29880 11212
rect 27528 11092 27580 11144
rect 28816 11135 28868 11144
rect 28816 11101 28825 11135
rect 28825 11101 28859 11135
rect 28859 11101 28868 11135
rect 28816 11092 28868 11101
rect 28908 11092 28960 11144
rect 30012 11135 30064 11144
rect 30012 11101 30021 11135
rect 30021 11101 30055 11135
rect 30055 11101 30064 11135
rect 30012 11092 30064 11101
rect 30932 11160 30984 11212
rect 30472 11092 30524 11144
rect 32128 11203 32180 11212
rect 32128 11169 32137 11203
rect 32137 11169 32171 11203
rect 32171 11169 32180 11203
rect 32128 11160 32180 11169
rect 31944 11135 31996 11144
rect 31944 11101 31953 11135
rect 31953 11101 31987 11135
rect 31987 11101 31996 11135
rect 31944 11092 31996 11101
rect 32404 11135 32456 11144
rect 32404 11101 32413 11135
rect 32413 11101 32447 11135
rect 32447 11101 32456 11135
rect 32404 11092 32456 11101
rect 15108 10956 15160 11008
rect 18052 11024 18104 11076
rect 20444 11024 20496 11076
rect 23848 11024 23900 11076
rect 29920 11024 29972 11076
rect 33232 11160 33284 11212
rect 32772 11135 32824 11144
rect 32772 11101 32781 11135
rect 32781 11101 32815 11135
rect 32815 11101 32824 11135
rect 32772 11092 32824 11101
rect 33692 11135 33744 11144
rect 33692 11101 33701 11135
rect 33701 11101 33735 11135
rect 33735 11101 33744 11135
rect 33692 11092 33744 11101
rect 32956 11024 33008 11076
rect 23664 10956 23716 11008
rect 27620 10956 27672 11008
rect 27988 10956 28040 11008
rect 29092 10956 29144 11008
rect 33416 10999 33468 11008
rect 33416 10965 33425 10999
rect 33425 10965 33459 10999
rect 33459 10965 33468 10999
rect 33416 10956 33468 10965
rect 34152 11024 34204 11076
rect 35256 11092 35308 11144
rect 35440 11135 35492 11144
rect 35440 11101 35474 11135
rect 35474 11101 35492 11135
rect 35440 11092 35492 11101
rect 35716 11092 35768 11144
rect 38108 11271 38160 11280
rect 38108 11237 38117 11271
rect 38117 11237 38151 11271
rect 38151 11237 38160 11271
rect 38108 11228 38160 11237
rect 38292 11135 38344 11144
rect 38292 11101 38301 11135
rect 38301 11101 38335 11135
rect 38335 11101 38344 11135
rect 38292 11092 38344 11101
rect 45192 11339 45244 11348
rect 45192 11305 45201 11339
rect 45201 11305 45235 11339
rect 45235 11305 45244 11339
rect 45192 11296 45244 11305
rect 48780 11339 48832 11348
rect 48780 11305 48789 11339
rect 48789 11305 48823 11339
rect 48823 11305 48832 11339
rect 48780 11296 48832 11305
rect 43076 11271 43128 11280
rect 43076 11237 43085 11271
rect 43085 11237 43119 11271
rect 43119 11237 43128 11271
rect 43076 11228 43128 11237
rect 46296 11228 46348 11280
rect 49332 11228 49384 11280
rect 40592 11160 40644 11212
rect 43996 11160 44048 11212
rect 39120 11135 39172 11144
rect 39120 11101 39129 11135
rect 39129 11101 39163 11135
rect 39163 11101 39172 11135
rect 39120 11092 39172 11101
rect 39304 11135 39356 11144
rect 39304 11101 39313 11135
rect 39313 11101 39347 11135
rect 39347 11101 39356 11135
rect 39304 11092 39356 11101
rect 42708 11092 42760 11144
rect 39212 11024 39264 11076
rect 39396 11024 39448 11076
rect 45468 11092 45520 11144
rect 45836 11203 45888 11212
rect 45836 11169 45845 11203
rect 45845 11169 45879 11203
rect 45879 11169 45888 11203
rect 46756 11203 46808 11212
rect 45836 11160 45888 11169
rect 46756 11169 46765 11203
rect 46765 11169 46799 11203
rect 46799 11169 46808 11203
rect 46756 11160 46808 11169
rect 45744 11024 45796 11076
rect 46480 11135 46532 11144
rect 46480 11101 46489 11135
rect 46489 11101 46523 11135
rect 46523 11101 46532 11135
rect 46480 11092 46532 11101
rect 46848 11092 46900 11144
rect 58164 11203 58216 11212
rect 58164 11169 58173 11203
rect 58173 11169 58207 11203
rect 58207 11169 58216 11203
rect 58164 11160 58216 11169
rect 48596 11135 48648 11144
rect 48596 11101 48605 11135
rect 48605 11101 48639 11135
rect 48639 11101 48648 11135
rect 48596 11092 48648 11101
rect 51724 11092 51776 11144
rect 37372 10956 37424 11008
rect 39488 10999 39540 11008
rect 39488 10965 39497 10999
rect 39497 10965 39531 10999
rect 39531 10965 39540 10999
rect 39488 10956 39540 10965
rect 39580 10956 39632 11008
rect 44456 10956 44508 11008
rect 50804 11024 50856 11076
rect 58900 11024 58952 11076
rect 49240 10956 49292 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 50294 10854 50346 10906
rect 50358 10854 50410 10906
rect 50422 10854 50474 10906
rect 50486 10854 50538 10906
rect 50550 10854 50602 10906
rect 13544 10752 13596 10804
rect 14740 10752 14792 10804
rect 2688 10684 2740 10736
rect 23388 10752 23440 10804
rect 23756 10752 23808 10804
rect 30012 10752 30064 10804
rect 30288 10752 30340 10804
rect 30472 10752 30524 10804
rect 12348 10616 12400 10668
rect 12440 10659 12492 10668
rect 12440 10625 12449 10659
rect 12449 10625 12483 10659
rect 12483 10625 12492 10659
rect 12440 10616 12492 10625
rect 13452 10616 13504 10668
rect 18696 10616 18748 10668
rect 28080 10684 28132 10736
rect 940 10548 992 10600
rect 13084 10480 13136 10532
rect 13544 10412 13596 10464
rect 17040 10412 17092 10464
rect 25412 10616 25464 10668
rect 29092 10684 29144 10736
rect 23940 10591 23992 10600
rect 23940 10557 23949 10591
rect 23949 10557 23983 10591
rect 23983 10557 23992 10591
rect 23940 10548 23992 10557
rect 23664 10480 23716 10532
rect 25780 10591 25832 10600
rect 25780 10557 25789 10591
rect 25789 10557 25823 10591
rect 25823 10557 25832 10591
rect 25780 10548 25832 10557
rect 25964 10591 26016 10600
rect 25964 10557 25973 10591
rect 25973 10557 26007 10591
rect 26007 10557 26016 10591
rect 25964 10548 26016 10557
rect 23388 10412 23440 10464
rect 27620 10480 27672 10532
rect 27712 10480 27764 10532
rect 25320 10455 25372 10464
rect 25320 10421 25329 10455
rect 25329 10421 25363 10455
rect 25363 10421 25372 10455
rect 25320 10412 25372 10421
rect 28540 10659 28592 10668
rect 28540 10625 28549 10659
rect 28549 10625 28583 10659
rect 28583 10625 28592 10659
rect 28540 10616 28592 10625
rect 28632 10616 28684 10668
rect 29552 10616 29604 10668
rect 33416 10684 33468 10736
rect 34796 10752 34848 10804
rect 35716 10752 35768 10804
rect 29000 10591 29052 10600
rect 29000 10557 29009 10591
rect 29009 10557 29043 10591
rect 29043 10557 29052 10591
rect 29000 10548 29052 10557
rect 35624 10616 35676 10668
rect 38200 10659 38252 10668
rect 38200 10625 38209 10659
rect 38209 10625 38243 10659
rect 38243 10625 38252 10659
rect 38200 10616 38252 10625
rect 39488 10684 39540 10736
rect 59636 10752 59688 10804
rect 39028 10616 39080 10668
rect 32680 10591 32732 10600
rect 32680 10557 32689 10591
rect 32689 10557 32723 10591
rect 32723 10557 32732 10591
rect 32680 10548 32732 10557
rect 33692 10548 33744 10600
rect 28816 10480 28868 10532
rect 30472 10412 30524 10464
rect 32404 10412 32456 10464
rect 46756 10616 46808 10668
rect 44088 10548 44140 10600
rect 44548 10591 44600 10600
rect 44548 10557 44557 10591
rect 44557 10557 44591 10591
rect 44591 10557 44600 10591
rect 44548 10548 44600 10557
rect 56048 10616 56100 10668
rect 56508 10659 56560 10668
rect 56508 10625 56517 10659
rect 56517 10625 56551 10659
rect 56551 10625 56560 10659
rect 56508 10616 56560 10625
rect 56600 10659 56652 10668
rect 56600 10625 56609 10659
rect 56609 10625 56643 10659
rect 56643 10625 56652 10659
rect 56600 10616 56652 10625
rect 57060 10659 57112 10668
rect 57060 10625 57069 10659
rect 57069 10625 57103 10659
rect 57103 10625 57112 10659
rect 57060 10616 57112 10625
rect 38384 10412 38436 10464
rect 39580 10455 39632 10464
rect 39580 10421 39589 10455
rect 39589 10421 39623 10455
rect 39623 10421 39632 10455
rect 39580 10412 39632 10421
rect 40224 10455 40276 10464
rect 40224 10421 40233 10455
rect 40233 10421 40267 10455
rect 40267 10421 40276 10455
rect 40224 10412 40276 10421
rect 44824 10412 44876 10464
rect 56416 10548 56468 10600
rect 58256 10659 58308 10668
rect 58256 10625 58265 10659
rect 58265 10625 58299 10659
rect 58299 10625 58308 10659
rect 58256 10616 58308 10625
rect 57888 10548 57940 10600
rect 56508 10480 56560 10532
rect 56876 10412 56928 10464
rect 57980 10412 58032 10464
rect 58992 10412 59044 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 12348 10251 12400 10260
rect 12348 10217 12357 10251
rect 12357 10217 12391 10251
rect 12391 10217 12400 10251
rect 12348 10208 12400 10217
rect 23940 10208 23992 10260
rect 23572 10183 23624 10192
rect 23572 10149 23581 10183
rect 23581 10149 23615 10183
rect 23615 10149 23624 10183
rect 23572 10140 23624 10149
rect 26056 10140 26108 10192
rect 27528 10140 27580 10192
rect 32680 10251 32732 10260
rect 32680 10217 32689 10251
rect 32689 10217 32723 10251
rect 32723 10217 32732 10251
rect 32680 10208 32732 10217
rect 39304 10208 39356 10260
rect 45836 10208 45888 10260
rect 57060 10208 57112 10260
rect 58256 10208 58308 10260
rect 12532 10115 12584 10124
rect 12532 10081 12541 10115
rect 12541 10081 12575 10115
rect 12575 10081 12584 10115
rect 12532 10072 12584 10081
rect 12624 10115 12676 10124
rect 12624 10081 12633 10115
rect 12633 10081 12667 10115
rect 12667 10081 12676 10115
rect 12624 10072 12676 10081
rect 25964 10072 26016 10124
rect 12348 10004 12400 10056
rect 12440 10004 12492 10056
rect 940 9936 992 9988
rect 13820 10004 13872 10056
rect 24584 10047 24636 10056
rect 24584 10013 24593 10047
rect 24593 10013 24627 10047
rect 24627 10013 24636 10047
rect 24584 10004 24636 10013
rect 25320 10004 25372 10056
rect 13360 9936 13412 9988
rect 25228 9936 25280 9988
rect 28080 10047 28132 10056
rect 28080 10013 28089 10047
rect 28089 10013 28123 10047
rect 28123 10013 28132 10047
rect 28080 10004 28132 10013
rect 30380 10004 30432 10056
rect 33232 10072 33284 10124
rect 38568 10004 38620 10056
rect 39580 10140 39632 10192
rect 56692 10140 56744 10192
rect 39028 10115 39080 10124
rect 39028 10081 39037 10115
rect 39037 10081 39071 10115
rect 39071 10081 39080 10115
rect 39028 10072 39080 10081
rect 28908 9936 28960 9988
rect 31208 9979 31260 9988
rect 31208 9945 31217 9979
rect 31217 9945 31251 9979
rect 31251 9945 31260 9979
rect 31208 9936 31260 9945
rect 32864 9936 32916 9988
rect 34152 9936 34204 9988
rect 34336 9936 34388 9988
rect 23296 9868 23348 9920
rect 25780 9868 25832 9920
rect 29276 9868 29328 9920
rect 36268 9868 36320 9920
rect 36452 9936 36504 9988
rect 38384 9936 38436 9988
rect 56784 10115 56836 10124
rect 56784 10081 56793 10115
rect 56793 10081 56827 10115
rect 56827 10081 56836 10115
rect 56784 10072 56836 10081
rect 44548 10004 44600 10056
rect 47492 10004 47544 10056
rect 56324 10047 56376 10056
rect 56324 10013 56333 10047
rect 56333 10013 56367 10047
rect 56367 10013 56376 10047
rect 56324 10004 56376 10013
rect 56876 10004 56928 10056
rect 45468 9979 45520 9988
rect 45468 9945 45502 9979
rect 45502 9945 45520 9979
rect 45468 9936 45520 9945
rect 38016 9868 38068 9920
rect 39028 9868 39080 9920
rect 48320 9936 48372 9988
rect 56048 9979 56100 9988
rect 56048 9945 56057 9979
rect 56057 9945 56091 9979
rect 56091 9945 56100 9979
rect 56048 9936 56100 9945
rect 56232 9911 56284 9920
rect 56232 9877 56241 9911
rect 56241 9877 56275 9911
rect 56275 9877 56284 9911
rect 56232 9868 56284 9877
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 50294 9766 50346 9818
rect 50358 9766 50410 9818
rect 50422 9766 50474 9818
rect 50486 9766 50538 9818
rect 50550 9766 50602 9818
rect 17960 9664 18012 9716
rect 18696 9664 18748 9716
rect 25228 9664 25280 9716
rect 28540 9664 28592 9716
rect 23572 9596 23624 9648
rect 12256 9528 12308 9580
rect 12532 9571 12584 9580
rect 12532 9537 12541 9571
rect 12541 9537 12575 9571
rect 12575 9537 12584 9571
rect 12532 9528 12584 9537
rect 17316 9528 17368 9580
rect 22744 9528 22796 9580
rect 23020 9528 23072 9580
rect 24584 9596 24636 9648
rect 29000 9596 29052 9648
rect 29460 9596 29512 9648
rect 30196 9596 30248 9648
rect 31024 9664 31076 9716
rect 940 9460 992 9512
rect 12348 9503 12400 9512
rect 12348 9469 12357 9503
rect 12357 9469 12391 9503
rect 12391 9469 12400 9503
rect 12348 9460 12400 9469
rect 12808 9503 12860 9512
rect 12808 9469 12817 9503
rect 12817 9469 12851 9503
rect 12851 9469 12860 9503
rect 12808 9460 12860 9469
rect 12624 9392 12676 9444
rect 13820 9503 13872 9512
rect 13820 9469 13829 9503
rect 13829 9469 13863 9503
rect 13863 9469 13872 9503
rect 13820 9460 13872 9469
rect 23204 9503 23256 9512
rect 23204 9469 23213 9503
rect 23213 9469 23247 9503
rect 23247 9469 23256 9503
rect 23204 9460 23256 9469
rect 26332 9571 26384 9580
rect 26332 9537 26341 9571
rect 26341 9537 26375 9571
rect 26375 9537 26384 9571
rect 26332 9528 26384 9537
rect 27160 9571 27212 9580
rect 27160 9537 27169 9571
rect 27169 9537 27203 9571
rect 27203 9537 27212 9571
rect 27160 9528 27212 9537
rect 27712 9528 27764 9580
rect 27988 9528 28040 9580
rect 29184 9528 29236 9580
rect 30288 9571 30340 9580
rect 30288 9537 30297 9571
rect 30297 9537 30331 9571
rect 30331 9537 30340 9571
rect 30288 9528 30340 9537
rect 30012 9460 30064 9512
rect 30932 9528 30984 9580
rect 30840 9460 30892 9512
rect 12900 9324 12952 9376
rect 26148 9392 26200 9444
rect 28540 9435 28592 9444
rect 28540 9401 28549 9435
rect 28549 9401 28583 9435
rect 28583 9401 28592 9435
rect 28540 9392 28592 9401
rect 28632 9392 28684 9444
rect 29920 9392 29972 9444
rect 31116 9392 31168 9444
rect 31576 9634 31628 9686
rect 32404 9664 32456 9716
rect 45468 9664 45520 9716
rect 56232 9664 56284 9716
rect 32128 9596 32180 9648
rect 32864 9596 32916 9648
rect 31576 9571 31628 9580
rect 31576 9537 31585 9571
rect 31585 9537 31619 9571
rect 31619 9537 31628 9571
rect 31576 9528 31628 9537
rect 32496 9528 32548 9580
rect 33232 9571 33284 9580
rect 33232 9537 33241 9571
rect 33241 9537 33275 9571
rect 33275 9537 33284 9571
rect 33232 9528 33284 9537
rect 33692 9528 33744 9580
rect 35624 9596 35676 9648
rect 35716 9596 35768 9648
rect 37096 9596 37148 9648
rect 31852 9392 31904 9444
rect 32404 9392 32456 9444
rect 24308 9324 24360 9376
rect 26608 9324 26660 9376
rect 36452 9503 36504 9512
rect 36452 9469 36461 9503
rect 36461 9469 36495 9503
rect 36495 9469 36504 9503
rect 36452 9460 36504 9469
rect 35440 9367 35492 9376
rect 35440 9333 35449 9367
rect 35449 9333 35483 9367
rect 35483 9333 35492 9367
rect 35440 9324 35492 9333
rect 35716 9324 35768 9376
rect 38844 9596 38896 9648
rect 38292 9528 38344 9580
rect 40224 9596 40276 9648
rect 40868 9596 40920 9648
rect 44640 9596 44692 9648
rect 58808 9596 58860 9648
rect 39304 9571 39356 9580
rect 39304 9537 39313 9571
rect 39313 9537 39347 9571
rect 39347 9537 39356 9571
rect 39304 9528 39356 9537
rect 38936 9460 38988 9512
rect 43904 9460 43956 9512
rect 45836 9503 45888 9512
rect 45836 9469 45845 9503
rect 45845 9469 45879 9503
rect 45879 9469 45888 9503
rect 45836 9460 45888 9469
rect 46756 9460 46808 9512
rect 41880 9392 41932 9444
rect 56416 9571 56468 9580
rect 56416 9537 56425 9571
rect 56425 9537 56459 9571
rect 56459 9537 56468 9571
rect 56416 9528 56468 9537
rect 57060 9571 57112 9580
rect 57060 9537 57069 9571
rect 57069 9537 57103 9571
rect 57103 9537 57112 9571
rect 57060 9528 57112 9537
rect 58992 9460 59044 9512
rect 52092 9392 52144 9444
rect 56324 9324 56376 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 12256 9163 12308 9172
rect 12256 9129 12265 9163
rect 12265 9129 12299 9163
rect 12299 9129 12308 9163
rect 12256 9120 12308 9129
rect 24308 9120 24360 9172
rect 25136 9120 25188 9172
rect 27344 9120 27396 9172
rect 25872 9052 25924 9104
rect 12164 8916 12216 8968
rect 940 8848 992 8900
rect 12348 8848 12400 8900
rect 12624 8959 12676 8968
rect 12624 8925 12633 8959
rect 12633 8925 12667 8959
rect 12667 8925 12676 8959
rect 12624 8916 12676 8925
rect 12716 8959 12768 8968
rect 12716 8925 12725 8959
rect 12725 8925 12759 8959
rect 12759 8925 12768 8959
rect 12716 8916 12768 8925
rect 18420 8916 18472 8968
rect 22836 8916 22888 8968
rect 23572 8984 23624 9036
rect 25688 9027 25740 9036
rect 25688 8993 25697 9027
rect 25697 8993 25731 9027
rect 25731 8993 25740 9027
rect 25688 8984 25740 8993
rect 26976 8984 27028 9036
rect 27160 9027 27212 9036
rect 27160 8993 27169 9027
rect 27169 8993 27203 9027
rect 27203 8993 27212 9027
rect 27160 8984 27212 8993
rect 23020 8959 23072 8968
rect 23020 8925 23029 8959
rect 23029 8925 23063 8959
rect 23063 8925 23072 8959
rect 23020 8916 23072 8925
rect 23112 8916 23164 8968
rect 25412 8959 25464 8968
rect 25412 8925 25421 8959
rect 25421 8925 25455 8959
rect 25455 8925 25464 8959
rect 25412 8916 25464 8925
rect 26424 8959 26476 8968
rect 26424 8925 26433 8959
rect 26433 8925 26467 8959
rect 26467 8925 26476 8959
rect 26424 8916 26476 8925
rect 17316 8848 17368 8900
rect 28356 8916 28408 8968
rect 29644 9052 29696 9104
rect 31484 9120 31536 9172
rect 36452 9120 36504 9172
rect 36636 9120 36688 9172
rect 39028 9120 39080 9172
rect 45192 9120 45244 9172
rect 57060 9120 57112 9172
rect 29552 8984 29604 9036
rect 29736 8984 29788 9036
rect 29644 8916 29696 8968
rect 29828 8916 29880 8968
rect 30288 8984 30340 9036
rect 30196 8959 30248 8968
rect 30196 8925 30205 8959
rect 30205 8925 30239 8959
rect 30239 8925 30248 8959
rect 30196 8916 30248 8925
rect 34428 8984 34480 9036
rect 30472 8916 30524 8968
rect 31116 8916 31168 8968
rect 27804 8848 27856 8900
rect 27988 8848 28040 8900
rect 31484 8848 31536 8900
rect 31668 8959 31720 8968
rect 31668 8925 31677 8959
rect 31677 8925 31711 8959
rect 31711 8925 31720 8959
rect 31668 8916 31720 8925
rect 35348 8916 35400 8968
rect 35808 8959 35860 8968
rect 35808 8925 35817 8959
rect 35817 8925 35851 8959
rect 35851 8925 35860 8959
rect 35808 8916 35860 8925
rect 44824 9052 44876 9104
rect 35992 8984 36044 9036
rect 38568 8984 38620 9036
rect 42800 8984 42852 9036
rect 43260 8984 43312 9036
rect 48596 8984 48648 9036
rect 48964 8984 49016 9036
rect 56784 9027 56836 9036
rect 56784 8993 56793 9027
rect 56793 8993 56827 9027
rect 56827 8993 56836 9027
rect 56784 8984 56836 8993
rect 37648 8916 37700 8968
rect 42340 8916 42392 8968
rect 43904 8916 43956 8968
rect 44364 8916 44416 8968
rect 56692 8916 56744 8968
rect 36268 8891 36320 8900
rect 36268 8857 36277 8891
rect 36277 8857 36311 8891
rect 36311 8857 36320 8891
rect 36268 8848 36320 8857
rect 37924 8848 37976 8900
rect 46204 8848 46256 8900
rect 48412 8848 48464 8900
rect 48964 8848 49016 8900
rect 12440 8780 12492 8832
rect 20536 8780 20588 8832
rect 25044 8823 25096 8832
rect 25044 8789 25053 8823
rect 25053 8789 25087 8823
rect 25087 8789 25096 8823
rect 25044 8780 25096 8789
rect 25596 8780 25648 8832
rect 28264 8780 28316 8832
rect 29092 8823 29144 8832
rect 29092 8789 29101 8823
rect 29101 8789 29135 8823
rect 29135 8789 29144 8823
rect 29092 8780 29144 8789
rect 30288 8780 30340 8832
rect 30380 8780 30432 8832
rect 31576 8780 31628 8832
rect 33140 8780 33192 8832
rect 33784 8780 33836 8832
rect 40684 8823 40736 8832
rect 40684 8789 40693 8823
rect 40693 8789 40727 8823
rect 40727 8789 40736 8823
rect 40684 8780 40736 8789
rect 41144 8823 41196 8832
rect 41144 8789 41153 8823
rect 41153 8789 41187 8823
rect 41187 8789 41196 8823
rect 41144 8780 41196 8789
rect 46112 8780 46164 8832
rect 48780 8780 48832 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 50294 8678 50346 8730
rect 50358 8678 50410 8730
rect 50422 8678 50474 8730
rect 50486 8678 50538 8730
rect 50550 8678 50602 8730
rect 11152 8576 11204 8628
rect 11336 8576 11388 8628
rect 12164 8619 12216 8628
rect 12164 8585 12173 8619
rect 12173 8585 12207 8619
rect 12207 8585 12216 8619
rect 12164 8576 12216 8585
rect 23296 8576 23348 8628
rect 27712 8576 27764 8628
rect 28448 8576 28500 8628
rect 28908 8576 28960 8628
rect 29644 8576 29696 8628
rect 30656 8576 30708 8628
rect 31576 8619 31628 8628
rect 31576 8585 31585 8619
rect 31585 8585 31619 8619
rect 31619 8585 31628 8619
rect 31576 8576 31628 8585
rect 33048 8576 33100 8628
rect 12532 8508 12584 8560
rect 940 8372 992 8424
rect 12348 8483 12400 8492
rect 12348 8449 12357 8483
rect 12357 8449 12391 8483
rect 12391 8449 12400 8483
rect 12348 8440 12400 8449
rect 12440 8483 12492 8492
rect 12440 8449 12449 8483
rect 12449 8449 12483 8483
rect 12483 8449 12492 8483
rect 12440 8440 12492 8449
rect 10968 8415 11020 8424
rect 10968 8381 10977 8415
rect 10977 8381 11011 8415
rect 11011 8381 11020 8415
rect 10968 8372 11020 8381
rect 11060 8415 11112 8424
rect 11060 8381 11069 8415
rect 11069 8381 11103 8415
rect 11103 8381 11112 8415
rect 11060 8372 11112 8381
rect 12532 8415 12584 8424
rect 12532 8381 12541 8415
rect 12541 8381 12575 8415
rect 12575 8381 12584 8415
rect 12532 8372 12584 8381
rect 12624 8415 12676 8424
rect 12624 8381 12633 8415
rect 12633 8381 12667 8415
rect 12667 8381 12676 8415
rect 12624 8372 12676 8381
rect 10876 8304 10928 8356
rect 24124 8440 24176 8492
rect 24584 8508 24636 8560
rect 24768 8508 24820 8560
rect 27988 8508 28040 8560
rect 25044 8440 25096 8492
rect 27068 8440 27120 8492
rect 29276 8483 29328 8492
rect 29276 8449 29285 8483
rect 29285 8449 29319 8483
rect 29319 8449 29328 8483
rect 29276 8440 29328 8449
rect 21180 8372 21232 8424
rect 21548 8372 21600 8424
rect 28356 8415 28408 8424
rect 28356 8381 28365 8415
rect 28365 8381 28399 8415
rect 28399 8381 28408 8415
rect 28356 8372 28408 8381
rect 28632 8372 28684 8424
rect 29000 8372 29052 8424
rect 29920 8372 29972 8424
rect 31852 8508 31904 8560
rect 33692 8551 33744 8560
rect 33692 8517 33701 8551
rect 33701 8517 33735 8551
rect 33735 8517 33744 8551
rect 33692 8508 33744 8517
rect 30288 8483 30340 8492
rect 30288 8449 30297 8483
rect 30297 8449 30331 8483
rect 30331 8449 30340 8483
rect 30288 8440 30340 8449
rect 30380 8440 30432 8492
rect 31208 8440 31260 8492
rect 33140 8440 33192 8492
rect 33324 8483 33376 8492
rect 33324 8449 33333 8483
rect 33333 8449 33367 8483
rect 33367 8449 33376 8483
rect 33324 8440 33376 8449
rect 33416 8483 33468 8492
rect 33416 8449 33426 8483
rect 33426 8449 33460 8483
rect 33460 8449 33468 8483
rect 33416 8440 33468 8449
rect 33876 8440 33928 8492
rect 34612 8440 34664 8492
rect 35532 8508 35584 8560
rect 41144 8576 41196 8628
rect 46204 8576 46256 8628
rect 36176 8508 36228 8560
rect 35808 8483 35860 8492
rect 35808 8449 35817 8483
rect 35817 8449 35851 8483
rect 35851 8449 35860 8483
rect 35808 8440 35860 8449
rect 35348 8372 35400 8424
rect 39120 8440 39172 8492
rect 40684 8440 40736 8492
rect 47676 8508 47728 8560
rect 53196 8508 53248 8560
rect 42708 8440 42760 8492
rect 42892 8483 42944 8492
rect 42892 8449 42926 8483
rect 42926 8449 42944 8483
rect 42892 8440 42944 8449
rect 47860 8440 47912 8492
rect 17316 8236 17368 8288
rect 18236 8236 18288 8288
rect 22100 8304 22152 8356
rect 25596 8347 25648 8356
rect 25596 8313 25605 8347
rect 25605 8313 25639 8347
rect 25639 8313 25648 8347
rect 25596 8304 25648 8313
rect 28448 8304 28500 8356
rect 29736 8304 29788 8356
rect 33140 8304 33192 8356
rect 20996 8236 21048 8288
rect 26608 8236 26660 8288
rect 26792 8236 26844 8288
rect 31944 8236 31996 8288
rect 34520 8347 34572 8356
rect 34520 8313 34529 8347
rect 34529 8313 34563 8347
rect 34563 8313 34572 8347
rect 37648 8415 37700 8424
rect 37648 8381 37657 8415
rect 37657 8381 37691 8415
rect 37691 8381 37700 8415
rect 37648 8372 37700 8381
rect 45100 8372 45152 8424
rect 46480 8372 46532 8424
rect 47216 8372 47268 8424
rect 48320 8440 48372 8492
rect 48964 8483 49016 8492
rect 48964 8449 48973 8483
rect 48973 8449 49007 8483
rect 49007 8449 49016 8483
rect 48964 8440 49016 8449
rect 58072 8483 58124 8492
rect 58072 8449 58081 8483
rect 58081 8449 58115 8483
rect 58115 8449 58124 8483
rect 58072 8440 58124 8449
rect 49056 8372 49108 8424
rect 34520 8304 34572 8313
rect 36452 8347 36504 8356
rect 36452 8313 36461 8347
rect 36461 8313 36495 8347
rect 36495 8313 36504 8347
rect 36452 8304 36504 8313
rect 37372 8304 37424 8356
rect 48136 8304 48188 8356
rect 48780 8347 48832 8356
rect 48780 8313 48789 8347
rect 48789 8313 48823 8347
rect 48823 8313 48832 8347
rect 48780 8304 48832 8313
rect 53380 8304 53432 8356
rect 55312 8304 55364 8356
rect 35440 8236 35492 8288
rect 42616 8236 42668 8288
rect 43536 8236 43588 8288
rect 48964 8236 49016 8288
rect 56600 8236 56652 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 11060 8032 11112 8084
rect 12624 8032 12676 8084
rect 23204 8032 23256 8084
rect 8760 7964 8812 8016
rect 10600 7964 10652 8016
rect 12808 7964 12860 8016
rect 11152 7939 11204 7948
rect 11152 7905 11161 7939
rect 11161 7905 11195 7939
rect 11195 7905 11204 7939
rect 11152 7896 11204 7905
rect 11244 7939 11296 7948
rect 11244 7905 11253 7939
rect 11253 7905 11287 7939
rect 11287 7905 11296 7939
rect 11244 7896 11296 7905
rect 12440 7896 12492 7948
rect 940 7760 992 7812
rect 10968 7760 11020 7812
rect 11428 7871 11480 7880
rect 11428 7837 11437 7871
rect 11437 7837 11471 7871
rect 11471 7837 11480 7871
rect 11428 7828 11480 7837
rect 11520 7828 11572 7880
rect 13360 7896 13412 7948
rect 19156 7896 19208 7948
rect 26792 8032 26844 8084
rect 27804 8032 27856 8084
rect 30472 8032 30524 8084
rect 32404 8032 32456 8084
rect 35440 8032 35492 8084
rect 35900 8032 35952 8084
rect 39396 8032 39448 8084
rect 42892 8032 42944 8084
rect 26608 7964 26660 8016
rect 36636 7964 36688 8016
rect 36912 7964 36964 8016
rect 38108 8007 38160 8016
rect 38108 7973 38117 8007
rect 38117 7973 38151 8007
rect 38151 7973 38160 8007
rect 38108 7964 38160 7973
rect 23572 7896 23624 7948
rect 11244 7692 11296 7744
rect 25596 7760 25648 7812
rect 27712 7896 27764 7948
rect 28632 7896 28684 7948
rect 29092 7896 29144 7948
rect 28816 7828 28868 7880
rect 30104 7828 30156 7880
rect 27252 7803 27304 7812
rect 27252 7769 27261 7803
rect 27261 7769 27295 7803
rect 27295 7769 27304 7803
rect 27252 7760 27304 7769
rect 28264 7803 28316 7812
rect 28264 7769 28273 7803
rect 28273 7769 28307 7803
rect 28307 7769 28316 7803
rect 28264 7760 28316 7769
rect 29184 7760 29236 7812
rect 30656 7871 30708 7880
rect 30656 7837 30670 7871
rect 30670 7837 30704 7871
rect 30704 7837 30708 7871
rect 30656 7828 30708 7837
rect 31576 7828 31628 7880
rect 31852 7896 31904 7948
rect 35992 7896 36044 7948
rect 42984 7896 43036 7948
rect 43260 7896 43312 7948
rect 31760 7871 31812 7880
rect 31760 7837 31769 7871
rect 31769 7837 31803 7871
rect 31803 7837 31812 7871
rect 31760 7828 31812 7837
rect 31944 7871 31996 7880
rect 31944 7837 31953 7871
rect 31953 7837 31987 7871
rect 31987 7837 31996 7871
rect 31944 7828 31996 7837
rect 32128 7828 32180 7880
rect 34520 7828 34572 7880
rect 35440 7828 35492 7880
rect 35808 7871 35860 7880
rect 35808 7837 35817 7871
rect 35817 7837 35851 7871
rect 35851 7837 35860 7871
rect 35808 7828 35860 7837
rect 37372 7828 37424 7880
rect 37464 7871 37516 7880
rect 37464 7837 37473 7871
rect 37473 7837 37507 7871
rect 37507 7837 37516 7871
rect 37464 7828 37516 7837
rect 37556 7871 37608 7880
rect 37556 7837 37565 7871
rect 37565 7837 37599 7871
rect 37599 7837 37608 7871
rect 37556 7828 37608 7837
rect 37832 7828 37884 7880
rect 38844 7828 38896 7880
rect 43628 7828 43680 7880
rect 44824 7828 44876 7880
rect 47492 7939 47544 7948
rect 47492 7905 47501 7939
rect 47501 7905 47535 7939
rect 47535 7905 47544 7939
rect 47492 7896 47544 7905
rect 46940 7828 46992 7880
rect 30472 7803 30524 7812
rect 30472 7769 30481 7803
rect 30481 7769 30515 7803
rect 30515 7769 30524 7803
rect 30472 7760 30524 7769
rect 22468 7692 22520 7744
rect 27528 7692 27580 7744
rect 28448 7692 28500 7744
rect 29000 7692 29052 7744
rect 34152 7803 34204 7812
rect 34152 7769 34161 7803
rect 34161 7769 34195 7803
rect 34195 7769 34204 7803
rect 34152 7760 34204 7769
rect 35900 7803 35952 7812
rect 35900 7769 35909 7803
rect 35909 7769 35943 7803
rect 35943 7769 35952 7803
rect 35900 7760 35952 7769
rect 36268 7803 36320 7812
rect 36268 7769 36277 7803
rect 36277 7769 36311 7803
rect 36311 7769 36320 7803
rect 36268 7760 36320 7769
rect 36636 7760 36688 7812
rect 48136 7760 48188 7812
rect 56416 7828 56468 7880
rect 57980 7896 58032 7948
rect 58164 7939 58216 7948
rect 58164 7905 58173 7939
rect 58173 7905 58207 7939
rect 58207 7905 58216 7939
rect 58164 7896 58216 7905
rect 43444 7735 43496 7744
rect 43444 7701 43453 7735
rect 43453 7701 43487 7735
rect 43487 7701 43496 7735
rect 43444 7692 43496 7701
rect 47952 7692 48004 7744
rect 56508 7692 56560 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 50294 7590 50346 7642
rect 50358 7590 50410 7642
rect 50422 7590 50474 7642
rect 50486 7590 50538 7642
rect 50550 7590 50602 7642
rect 11428 7488 11480 7540
rect 12716 7488 12768 7540
rect 10968 7420 11020 7472
rect 12348 7352 12400 7404
rect 24124 7395 24176 7404
rect 24124 7361 24133 7395
rect 24133 7361 24167 7395
rect 24167 7361 24176 7395
rect 24124 7352 24176 7361
rect 24952 7352 25004 7404
rect 29920 7531 29972 7540
rect 29920 7497 29929 7531
rect 29929 7497 29963 7531
rect 29963 7497 29972 7531
rect 29920 7488 29972 7497
rect 30748 7488 30800 7540
rect 31484 7488 31536 7540
rect 35348 7488 35400 7540
rect 35808 7488 35860 7540
rect 37464 7488 37516 7540
rect 30380 7420 30432 7472
rect 30656 7420 30708 7472
rect 30932 7352 30984 7404
rect 33784 7463 33836 7472
rect 33784 7429 33793 7463
rect 33793 7429 33827 7463
rect 33827 7429 33836 7463
rect 33784 7420 33836 7429
rect 940 7284 992 7336
rect 20444 7284 20496 7336
rect 27528 7284 27580 7336
rect 30748 7284 30800 7336
rect 31116 7327 31168 7336
rect 31116 7293 31125 7327
rect 31125 7293 31159 7327
rect 31159 7293 31168 7327
rect 31116 7284 31168 7293
rect 32404 7395 32456 7404
rect 32404 7361 32413 7395
rect 32413 7361 32447 7395
rect 32447 7361 32456 7395
rect 32404 7352 32456 7361
rect 32772 7395 32824 7404
rect 32772 7361 32781 7395
rect 32781 7361 32815 7395
rect 32815 7361 32824 7395
rect 32772 7352 32824 7361
rect 37372 7352 37424 7404
rect 43444 7420 43496 7472
rect 44824 7531 44876 7540
rect 44824 7497 44833 7531
rect 44833 7497 44867 7531
rect 44867 7497 44876 7531
rect 44824 7488 44876 7497
rect 46940 7488 46992 7540
rect 48136 7531 48188 7540
rect 48136 7497 48145 7531
rect 48145 7497 48179 7531
rect 48179 7497 48188 7531
rect 48136 7488 48188 7497
rect 56508 7531 56560 7540
rect 56508 7497 56517 7531
rect 56517 7497 56551 7531
rect 56551 7497 56560 7531
rect 56508 7488 56560 7497
rect 48964 7420 49016 7472
rect 38200 7395 38252 7404
rect 38200 7361 38209 7395
rect 38209 7361 38243 7395
rect 38243 7361 38252 7395
rect 38200 7352 38252 7361
rect 44272 7352 44324 7404
rect 45192 7395 45244 7404
rect 45192 7361 45201 7395
rect 45201 7361 45235 7395
rect 45235 7361 45244 7395
rect 45192 7352 45244 7361
rect 9128 7216 9180 7268
rect 12072 7259 12124 7268
rect 12072 7225 12081 7259
rect 12081 7225 12115 7259
rect 12115 7225 12124 7259
rect 12072 7216 12124 7225
rect 13452 7216 13504 7268
rect 30472 7216 30524 7268
rect 30932 7259 30984 7268
rect 30932 7225 30941 7259
rect 30941 7225 30975 7259
rect 30975 7225 30984 7259
rect 30932 7216 30984 7225
rect 31024 7216 31076 7268
rect 25044 7148 25096 7200
rect 25136 7148 25188 7200
rect 27252 7148 27304 7200
rect 29000 7148 29052 7200
rect 30012 7148 30064 7200
rect 35624 7284 35676 7336
rect 34796 7216 34848 7268
rect 39488 7327 39540 7336
rect 39488 7293 39497 7327
rect 39497 7293 39531 7327
rect 39531 7293 39540 7327
rect 39488 7284 39540 7293
rect 44456 7284 44508 7336
rect 44824 7284 44876 7336
rect 45008 7284 45060 7336
rect 46020 7352 46072 7404
rect 46572 7395 46624 7404
rect 46572 7361 46581 7395
rect 46581 7361 46615 7395
rect 46615 7361 46624 7395
rect 46572 7352 46624 7361
rect 47952 7395 48004 7404
rect 47952 7361 47961 7395
rect 47961 7361 47995 7395
rect 47995 7361 48004 7395
rect 47952 7352 48004 7361
rect 55496 7352 55548 7404
rect 56048 7420 56100 7472
rect 56324 7463 56376 7472
rect 56324 7429 56333 7463
rect 56333 7429 56367 7463
rect 56367 7429 56376 7463
rect 56324 7420 56376 7429
rect 55772 7395 55824 7404
rect 55772 7361 55781 7395
rect 55781 7361 55815 7395
rect 55815 7361 55824 7395
rect 55772 7352 55824 7361
rect 47124 7284 47176 7336
rect 47492 7284 47544 7336
rect 38384 7259 38436 7268
rect 38384 7225 38393 7259
rect 38393 7225 38427 7259
rect 38427 7225 38436 7259
rect 38384 7216 38436 7225
rect 31760 7148 31812 7200
rect 39672 7191 39724 7200
rect 39672 7157 39681 7191
rect 39681 7157 39715 7191
rect 39715 7157 39724 7191
rect 39672 7148 39724 7157
rect 42708 7216 42760 7268
rect 56600 7395 56652 7404
rect 56600 7361 56609 7395
rect 56609 7361 56643 7395
rect 56643 7361 56652 7395
rect 56600 7352 56652 7361
rect 57980 7352 58032 7404
rect 58072 7395 58124 7404
rect 58072 7361 58081 7395
rect 58081 7361 58115 7395
rect 58115 7361 58124 7395
rect 58072 7352 58124 7361
rect 58992 7284 59044 7336
rect 58256 7259 58308 7268
rect 58256 7225 58265 7259
rect 58265 7225 58299 7259
rect 58299 7225 58308 7259
rect 58256 7216 58308 7225
rect 42984 7148 43036 7200
rect 47676 7148 47728 7200
rect 48136 7148 48188 7200
rect 56048 7148 56100 7200
rect 56968 7148 57020 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 20996 6944 21048 6996
rect 24952 6987 25004 6996
rect 24952 6953 24961 6987
rect 24961 6953 24995 6987
rect 24995 6953 25004 6987
rect 24952 6944 25004 6953
rect 14464 6808 14516 6860
rect 10416 6740 10468 6792
rect 13912 6740 13964 6792
rect 21180 6876 21232 6928
rect 31392 6987 31444 6996
rect 31392 6953 31401 6987
rect 31401 6953 31435 6987
rect 31435 6953 31444 6987
rect 31392 6944 31444 6953
rect 38200 6944 38252 6996
rect 39672 6944 39724 6996
rect 41420 6944 41472 6996
rect 46940 6944 46992 6996
rect 47216 6944 47268 6996
rect 31576 6876 31628 6928
rect 31944 6876 31996 6928
rect 32772 6876 32824 6928
rect 25688 6808 25740 6860
rect 27160 6808 27212 6860
rect 27528 6851 27580 6860
rect 27528 6817 27537 6851
rect 27537 6817 27571 6851
rect 27571 6817 27580 6851
rect 27528 6808 27580 6817
rect 940 6672 992 6724
rect 20444 6715 20496 6724
rect 20444 6681 20453 6715
rect 20453 6681 20487 6715
rect 20487 6681 20496 6715
rect 20444 6672 20496 6681
rect 27620 6740 27672 6792
rect 28172 6808 28224 6860
rect 29000 6851 29052 6860
rect 29000 6817 29009 6851
rect 29009 6817 29043 6851
rect 29043 6817 29052 6851
rect 29000 6808 29052 6817
rect 29276 6808 29328 6860
rect 30472 6808 30524 6860
rect 30656 6851 30708 6860
rect 30656 6817 30665 6851
rect 30665 6817 30699 6851
rect 30699 6817 30708 6851
rect 30656 6808 30708 6817
rect 27896 6740 27948 6792
rect 30748 6783 30800 6792
rect 30748 6749 30757 6783
rect 30757 6749 30791 6783
rect 30791 6749 30800 6783
rect 30748 6740 30800 6749
rect 31024 6740 31076 6792
rect 25136 6672 25188 6724
rect 29828 6672 29880 6724
rect 31576 6783 31628 6792
rect 31576 6749 31585 6783
rect 31585 6749 31619 6783
rect 31619 6749 31628 6783
rect 31576 6740 31628 6749
rect 32036 6740 32088 6792
rect 32496 6783 32548 6792
rect 32496 6749 32505 6783
rect 32505 6749 32539 6783
rect 32539 6749 32548 6783
rect 32496 6740 32548 6749
rect 32772 6783 32824 6792
rect 32772 6749 32781 6783
rect 32781 6749 32815 6783
rect 32815 6749 32824 6783
rect 32772 6740 32824 6749
rect 37280 6808 37332 6860
rect 37924 6851 37976 6860
rect 37924 6817 37933 6851
rect 37933 6817 37967 6851
rect 37967 6817 37976 6851
rect 37924 6808 37976 6817
rect 38292 6876 38344 6928
rect 40684 6876 40736 6928
rect 38108 6808 38160 6860
rect 46020 6876 46072 6928
rect 57980 6944 58032 6996
rect 35624 6783 35676 6792
rect 35624 6749 35633 6783
rect 35633 6749 35667 6783
rect 35667 6749 35676 6783
rect 35624 6740 35676 6749
rect 35716 6740 35768 6792
rect 39856 6740 39908 6792
rect 39948 6740 40000 6792
rect 40500 6740 40552 6792
rect 43904 6808 43956 6860
rect 44272 6740 44324 6792
rect 44456 6783 44508 6792
rect 44456 6749 44465 6783
rect 44465 6749 44499 6783
rect 44499 6749 44508 6783
rect 44456 6740 44508 6749
rect 44916 6740 44968 6792
rect 33140 6672 33192 6724
rect 34152 6672 34204 6724
rect 34704 6672 34756 6724
rect 31024 6604 31076 6656
rect 31760 6647 31812 6656
rect 31760 6613 31769 6647
rect 31769 6613 31803 6647
rect 31803 6613 31812 6647
rect 31760 6604 31812 6613
rect 32772 6604 32824 6656
rect 34060 6647 34112 6656
rect 34060 6613 34069 6647
rect 34069 6613 34103 6647
rect 34103 6613 34112 6647
rect 34060 6604 34112 6613
rect 34612 6604 34664 6656
rect 39304 6672 39356 6724
rect 43996 6672 44048 6724
rect 45008 6672 45060 6724
rect 37096 6604 37148 6656
rect 40224 6604 40276 6656
rect 42708 6604 42760 6656
rect 43260 6647 43312 6656
rect 43260 6613 43269 6647
rect 43269 6613 43303 6647
rect 43303 6613 43312 6647
rect 43260 6604 43312 6613
rect 44548 6647 44600 6656
rect 44548 6613 44557 6647
rect 44557 6613 44591 6647
rect 44591 6613 44600 6647
rect 44548 6604 44600 6613
rect 45376 6604 45428 6656
rect 45744 6783 45796 6792
rect 45744 6749 45753 6783
rect 45753 6749 45787 6783
rect 45787 6749 45796 6783
rect 45744 6740 45796 6749
rect 46112 6783 46164 6792
rect 46112 6749 46121 6783
rect 46121 6749 46155 6783
rect 46155 6749 46164 6783
rect 46112 6740 46164 6749
rect 46664 6740 46716 6792
rect 45836 6604 45888 6656
rect 46388 6604 46440 6656
rect 46664 6604 46716 6656
rect 47216 6604 47268 6656
rect 47676 6715 47728 6724
rect 47676 6681 47685 6715
rect 47685 6681 47719 6715
rect 47719 6681 47728 6715
rect 47676 6672 47728 6681
rect 47860 6783 47912 6792
rect 47860 6749 47869 6783
rect 47869 6749 47903 6783
rect 47903 6749 47912 6783
rect 47860 6740 47912 6749
rect 48596 6740 48648 6792
rect 55404 6672 55456 6724
rect 56784 6740 56836 6792
rect 56968 6783 57020 6792
rect 56968 6749 57002 6783
rect 57002 6749 57020 6783
rect 56968 6740 57020 6749
rect 58992 6672 59044 6724
rect 48228 6604 48280 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 50294 6502 50346 6554
rect 50358 6502 50410 6554
rect 50422 6502 50474 6554
rect 50486 6502 50538 6554
rect 50550 6502 50602 6554
rect 10416 6443 10468 6452
rect 10416 6409 10425 6443
rect 10425 6409 10459 6443
rect 10459 6409 10468 6443
rect 10416 6400 10468 6409
rect 18328 6400 18380 6452
rect 10692 6332 10744 6384
rect 25136 6332 25188 6384
rect 25228 6375 25280 6384
rect 25228 6341 25237 6375
rect 25237 6341 25271 6375
rect 25271 6341 25280 6375
rect 25228 6332 25280 6341
rect 28172 6400 28224 6452
rect 29184 6400 29236 6452
rect 29644 6400 29696 6452
rect 26056 6264 26108 6316
rect 940 6196 992 6248
rect 10508 6196 10560 6248
rect 10692 6239 10744 6248
rect 10692 6205 10701 6239
rect 10701 6205 10735 6239
rect 10735 6205 10744 6239
rect 10692 6196 10744 6205
rect 10784 6239 10836 6248
rect 10784 6205 10793 6239
rect 10793 6205 10827 6239
rect 10827 6205 10836 6239
rect 10784 6196 10836 6205
rect 11060 6196 11112 6248
rect 20444 6196 20496 6248
rect 25320 6239 25372 6248
rect 25320 6205 25329 6239
rect 25329 6205 25363 6239
rect 25363 6205 25372 6239
rect 25320 6196 25372 6205
rect 25688 6196 25740 6248
rect 26332 6196 26384 6248
rect 26792 6196 26844 6248
rect 30840 6400 30892 6452
rect 34612 6400 34664 6452
rect 34704 6443 34756 6452
rect 34704 6409 34713 6443
rect 34713 6409 34747 6443
rect 34747 6409 34756 6443
rect 34704 6400 34756 6409
rect 39488 6400 39540 6452
rect 39856 6443 39908 6452
rect 39856 6409 39865 6443
rect 39865 6409 39899 6443
rect 39899 6409 39908 6443
rect 39856 6400 39908 6409
rect 40500 6443 40552 6452
rect 40500 6409 40509 6443
rect 40509 6409 40543 6443
rect 40543 6409 40552 6443
rect 40500 6400 40552 6409
rect 44272 6443 44324 6452
rect 44272 6409 44281 6443
rect 44281 6409 44315 6443
rect 44315 6409 44324 6443
rect 44272 6400 44324 6409
rect 45192 6400 45244 6452
rect 45468 6400 45520 6452
rect 45652 6400 45704 6452
rect 46388 6400 46440 6452
rect 48412 6400 48464 6452
rect 31116 6332 31168 6384
rect 31760 6332 31812 6384
rect 28356 6264 28408 6316
rect 27804 6239 27856 6248
rect 27804 6205 27813 6239
rect 27813 6205 27847 6239
rect 27847 6205 27856 6239
rect 27804 6196 27856 6205
rect 28080 6196 28132 6248
rect 28540 6196 28592 6248
rect 28816 6307 28868 6316
rect 28816 6273 28825 6307
rect 28825 6273 28859 6307
rect 28859 6273 28868 6307
rect 28816 6264 28868 6273
rect 29460 6264 29512 6316
rect 29644 6307 29696 6316
rect 29644 6273 29653 6307
rect 29653 6273 29687 6307
rect 29687 6273 29696 6307
rect 29644 6264 29696 6273
rect 29828 6307 29880 6316
rect 29828 6273 29837 6307
rect 29837 6273 29871 6307
rect 29871 6273 29880 6307
rect 29828 6264 29880 6273
rect 30656 6307 30708 6316
rect 30656 6273 30665 6307
rect 30665 6273 30699 6307
rect 30699 6273 30708 6307
rect 30656 6264 30708 6273
rect 30748 6307 30800 6316
rect 30748 6273 30757 6307
rect 30757 6273 30791 6307
rect 30791 6273 30800 6307
rect 30748 6264 30800 6273
rect 32588 6307 32640 6316
rect 32588 6273 32597 6307
rect 32597 6273 32631 6307
rect 32631 6273 32640 6307
rect 32588 6264 32640 6273
rect 32772 6307 32824 6316
rect 32772 6273 32781 6307
rect 32781 6273 32815 6307
rect 32815 6273 32824 6307
rect 32772 6264 32824 6273
rect 37096 6332 37148 6384
rect 35348 6264 35400 6316
rect 35532 6307 35584 6316
rect 35532 6273 35541 6307
rect 35541 6273 35575 6307
rect 35575 6273 35584 6307
rect 35532 6264 35584 6273
rect 35900 6307 35952 6316
rect 35900 6273 35909 6307
rect 35909 6273 35943 6307
rect 35943 6273 35952 6307
rect 35900 6264 35952 6273
rect 36360 6264 36412 6316
rect 43352 6332 43404 6384
rect 37464 6307 37516 6316
rect 37464 6273 37473 6307
rect 37473 6273 37507 6307
rect 37507 6273 37516 6307
rect 37464 6264 37516 6273
rect 30564 6239 30616 6248
rect 30564 6205 30573 6239
rect 30573 6205 30607 6239
rect 30607 6205 30616 6239
rect 30564 6196 30616 6205
rect 30932 6196 30984 6248
rect 33140 6196 33192 6248
rect 16580 6128 16632 6180
rect 29000 6128 29052 6180
rect 30288 6128 30340 6180
rect 24584 6060 24636 6112
rect 24676 6060 24728 6112
rect 25688 6060 25740 6112
rect 28724 6060 28776 6112
rect 34060 6128 34112 6180
rect 34612 6196 34664 6248
rect 34428 6128 34480 6180
rect 35716 6128 35768 6180
rect 36268 6171 36320 6180
rect 36268 6137 36277 6171
rect 36277 6137 36311 6171
rect 36311 6137 36320 6171
rect 36268 6128 36320 6137
rect 37556 6196 37608 6248
rect 38200 6128 38252 6180
rect 39028 6264 39080 6316
rect 39304 6307 39356 6316
rect 39304 6273 39313 6307
rect 39313 6273 39347 6307
rect 39347 6273 39356 6307
rect 39304 6264 39356 6273
rect 40040 6264 40092 6316
rect 39304 6128 39356 6180
rect 40500 6264 40552 6316
rect 42800 6264 42852 6316
rect 43444 6264 43496 6316
rect 44364 6264 44416 6316
rect 45744 6332 45796 6384
rect 45100 6307 45152 6316
rect 45100 6273 45109 6307
rect 45109 6273 45143 6307
rect 45143 6273 45152 6307
rect 45100 6264 45152 6273
rect 45192 6264 45244 6316
rect 45468 6196 45520 6248
rect 47676 6264 47728 6316
rect 54668 6332 54720 6384
rect 43904 6128 43956 6180
rect 46664 6128 46716 6180
rect 48596 6128 48648 6180
rect 32956 6103 33008 6112
rect 32956 6069 32965 6103
rect 32965 6069 32999 6103
rect 32999 6069 33008 6103
rect 32956 6060 33008 6069
rect 35808 6060 35860 6112
rect 37556 6060 37608 6112
rect 37832 6060 37884 6112
rect 40040 6060 40092 6112
rect 44088 6060 44140 6112
rect 46388 6060 46440 6112
rect 47860 6060 47912 6112
rect 54760 6060 54812 6112
rect 55680 6264 55732 6316
rect 56784 6332 56836 6384
rect 56048 6307 56100 6316
rect 56048 6273 56082 6307
rect 56082 6273 56100 6307
rect 56048 6264 56100 6273
rect 56324 6264 56376 6316
rect 57152 6196 57204 6248
rect 56416 6060 56468 6112
rect 57060 6060 57112 6112
rect 58072 6103 58124 6112
rect 58072 6069 58081 6103
rect 58081 6069 58115 6103
rect 58115 6069 58124 6103
rect 58072 6060 58124 6069
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 11060 5899 11112 5908
rect 11060 5865 11069 5899
rect 11069 5865 11103 5899
rect 11103 5865 11112 5899
rect 11060 5856 11112 5865
rect 12348 5856 12400 5908
rect 23112 5899 23164 5908
rect 23112 5865 23121 5899
rect 23121 5865 23155 5899
rect 23155 5865 23164 5899
rect 23112 5856 23164 5865
rect 24584 5856 24636 5908
rect 8392 5788 8444 5840
rect 13820 5788 13872 5840
rect 24768 5788 24820 5840
rect 26792 5899 26844 5908
rect 26792 5865 26801 5899
rect 26801 5865 26835 5899
rect 26835 5865 26844 5899
rect 26792 5856 26844 5865
rect 29920 5856 29972 5908
rect 30840 5856 30892 5908
rect 30932 5899 30984 5908
rect 30932 5865 30941 5899
rect 30941 5865 30975 5899
rect 30975 5865 30984 5899
rect 30932 5856 30984 5865
rect 31024 5856 31076 5908
rect 39948 5856 40000 5908
rect 40316 5856 40368 5908
rect 45100 5856 45152 5908
rect 27712 5788 27764 5840
rect 31392 5788 31444 5840
rect 32588 5788 32640 5840
rect 10140 5763 10192 5772
rect 10140 5729 10149 5763
rect 10149 5729 10183 5763
rect 10183 5729 10192 5763
rect 10140 5720 10192 5729
rect 4620 5652 4672 5704
rect 9404 5695 9456 5704
rect 9404 5661 9413 5695
rect 9413 5661 9447 5695
rect 9447 5661 9456 5695
rect 9404 5652 9456 5661
rect 9496 5695 9548 5704
rect 9496 5661 9505 5695
rect 9505 5661 9539 5695
rect 9539 5661 9548 5695
rect 9496 5652 9548 5661
rect 10784 5720 10836 5772
rect 25320 5720 25372 5772
rect 30012 5763 30064 5772
rect 30012 5729 30021 5763
rect 30021 5729 30055 5763
rect 30055 5729 30064 5763
rect 30012 5720 30064 5729
rect 30104 5720 30156 5772
rect 940 5584 992 5636
rect 10140 5584 10192 5636
rect 18144 5695 18196 5704
rect 18144 5661 18153 5695
rect 18153 5661 18187 5695
rect 18187 5661 18196 5695
rect 18144 5652 18196 5661
rect 18236 5695 18288 5704
rect 18236 5661 18245 5695
rect 18245 5661 18279 5695
rect 18279 5661 18288 5695
rect 18236 5652 18288 5661
rect 20444 5652 20496 5704
rect 27528 5652 27580 5704
rect 27712 5695 27764 5704
rect 27712 5661 27721 5695
rect 27721 5661 27755 5695
rect 27755 5661 27764 5695
rect 27712 5652 27764 5661
rect 24768 5584 24820 5636
rect 25688 5627 25740 5636
rect 25688 5593 25722 5627
rect 25722 5593 25740 5627
rect 25688 5584 25740 5593
rect 25872 5584 25924 5636
rect 26424 5584 26476 5636
rect 29184 5652 29236 5704
rect 32496 5720 32548 5772
rect 30104 5584 30156 5636
rect 31944 5652 31996 5704
rect 32036 5652 32088 5704
rect 32680 5652 32732 5704
rect 33048 5720 33100 5772
rect 28172 5516 28224 5568
rect 29184 5516 29236 5568
rect 30380 5559 30432 5568
rect 30380 5525 30389 5559
rect 30389 5525 30423 5559
rect 30423 5525 30432 5559
rect 30380 5516 30432 5525
rect 32128 5584 32180 5636
rect 32956 5695 33008 5704
rect 32956 5661 32965 5695
rect 32965 5661 32999 5695
rect 32999 5661 33008 5695
rect 32956 5652 33008 5661
rect 33140 5695 33192 5704
rect 33140 5661 33149 5695
rect 33149 5661 33183 5695
rect 33183 5661 33192 5695
rect 33140 5652 33192 5661
rect 34152 5695 34204 5704
rect 34152 5661 34161 5695
rect 34161 5661 34195 5695
rect 34195 5661 34204 5695
rect 34152 5652 34204 5661
rect 34612 5652 34664 5704
rect 35532 5695 35584 5704
rect 35532 5661 35541 5695
rect 35541 5661 35575 5695
rect 35575 5661 35584 5695
rect 35532 5652 35584 5661
rect 35808 5695 35860 5704
rect 35808 5661 35817 5695
rect 35817 5661 35851 5695
rect 35851 5661 35860 5695
rect 35808 5652 35860 5661
rect 43812 5788 43864 5840
rect 45560 5899 45612 5908
rect 45560 5865 45569 5899
rect 45569 5865 45603 5899
rect 45603 5865 45612 5899
rect 45560 5856 45612 5865
rect 46572 5856 46624 5908
rect 46756 5899 46808 5908
rect 46756 5865 46765 5899
rect 46765 5865 46799 5899
rect 46799 5865 46808 5899
rect 46756 5856 46808 5865
rect 55772 5856 55824 5908
rect 36084 5720 36136 5772
rect 35440 5584 35492 5636
rect 36268 5627 36320 5636
rect 36268 5593 36277 5627
rect 36277 5593 36311 5627
rect 36311 5593 36320 5627
rect 36268 5584 36320 5593
rect 32588 5516 32640 5568
rect 33416 5516 33468 5568
rect 39580 5652 39632 5704
rect 40224 5720 40276 5772
rect 46388 5788 46440 5840
rect 47492 5788 47544 5840
rect 54668 5788 54720 5840
rect 58440 5856 58492 5908
rect 43168 5652 43220 5704
rect 44548 5652 44600 5704
rect 38200 5627 38252 5636
rect 38200 5593 38209 5627
rect 38209 5593 38243 5627
rect 38243 5593 38252 5627
rect 38200 5584 38252 5593
rect 38292 5584 38344 5636
rect 38936 5627 38988 5636
rect 38936 5593 38945 5627
rect 38945 5593 38979 5627
rect 38979 5593 38988 5627
rect 38936 5584 38988 5593
rect 42892 5584 42944 5636
rect 44088 5584 44140 5636
rect 45192 5627 45244 5636
rect 45192 5593 45201 5627
rect 45201 5593 45235 5627
rect 45235 5593 45244 5627
rect 45192 5584 45244 5593
rect 46020 5695 46072 5704
rect 46020 5661 46029 5695
rect 46029 5661 46063 5695
rect 46063 5661 46072 5695
rect 46020 5652 46072 5661
rect 53656 5720 53708 5772
rect 46664 5695 46716 5704
rect 46664 5661 46673 5695
rect 46673 5661 46707 5695
rect 46707 5661 46716 5695
rect 46664 5652 46716 5661
rect 56416 5720 56468 5772
rect 56784 5763 56836 5772
rect 56784 5729 56793 5763
rect 56793 5729 56827 5763
rect 56827 5729 56836 5763
rect 56784 5720 56836 5729
rect 56876 5652 56928 5704
rect 58072 5652 58124 5704
rect 57152 5584 57204 5636
rect 57336 5584 57388 5636
rect 58992 5584 59044 5636
rect 38016 5516 38068 5568
rect 40040 5516 40092 5568
rect 43352 5516 43404 5568
rect 47216 5516 47268 5568
rect 55680 5516 55732 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 50294 5414 50346 5466
rect 50358 5414 50410 5466
rect 50422 5414 50474 5466
rect 50486 5414 50538 5466
rect 50550 5414 50602 5466
rect 23112 5312 23164 5364
rect 24308 5312 24360 5364
rect 25044 5312 25096 5364
rect 25320 5312 25372 5364
rect 26332 5355 26384 5364
rect 26332 5321 26341 5355
rect 26341 5321 26375 5355
rect 26375 5321 26384 5355
rect 26332 5312 26384 5321
rect 26424 5355 26476 5364
rect 26424 5321 26433 5355
rect 26433 5321 26467 5355
rect 26467 5321 26476 5355
rect 26424 5312 26476 5321
rect 24676 5244 24728 5296
rect 26056 5287 26108 5296
rect 26056 5253 26065 5287
rect 26065 5253 26099 5287
rect 26099 5253 26108 5287
rect 26056 5244 26108 5253
rect 29184 5355 29236 5364
rect 29184 5321 29193 5355
rect 29193 5321 29227 5355
rect 29227 5321 29236 5355
rect 29184 5312 29236 5321
rect 29828 5244 29880 5296
rect 9588 5176 9640 5228
rect 19800 5219 19852 5228
rect 19800 5185 19809 5219
rect 19809 5185 19843 5219
rect 19843 5185 19852 5219
rect 19800 5176 19852 5185
rect 20812 5176 20864 5228
rect 24124 5219 24176 5228
rect 24124 5185 24133 5219
rect 24133 5185 24167 5219
rect 24167 5185 24176 5219
rect 24124 5176 24176 5185
rect 26608 5219 26660 5228
rect 26608 5185 26617 5219
rect 26617 5185 26651 5219
rect 26651 5185 26660 5219
rect 26608 5176 26660 5185
rect 27620 5176 27672 5228
rect 29184 5176 29236 5228
rect 30656 5176 30708 5228
rect 31300 5219 31352 5228
rect 31300 5185 31309 5219
rect 31309 5185 31343 5219
rect 31343 5185 31352 5219
rect 31300 5176 31352 5185
rect 34612 5287 34664 5296
rect 34612 5253 34621 5287
rect 34621 5253 34655 5287
rect 34655 5253 34664 5287
rect 34612 5244 34664 5253
rect 31760 5176 31812 5228
rect 32220 5176 32272 5228
rect 32588 5219 32640 5228
rect 32588 5185 32597 5219
rect 32597 5185 32631 5219
rect 32631 5185 32640 5219
rect 32588 5176 32640 5185
rect 32680 5176 32732 5228
rect 40224 5312 40276 5364
rect 40500 5355 40552 5364
rect 40500 5321 40509 5355
rect 40509 5321 40543 5355
rect 40543 5321 40552 5355
rect 40500 5312 40552 5321
rect 41236 5355 41288 5364
rect 41236 5321 41245 5355
rect 41245 5321 41279 5355
rect 41279 5321 41288 5355
rect 41236 5312 41288 5321
rect 35624 5244 35676 5296
rect 36176 5244 36228 5296
rect 43444 5287 43496 5296
rect 43444 5253 43453 5287
rect 43453 5253 43487 5287
rect 43487 5253 43496 5287
rect 43444 5244 43496 5253
rect 44456 5244 44508 5296
rect 47952 5244 48004 5296
rect 49608 5244 49660 5296
rect 57336 5287 57388 5296
rect 57336 5253 57345 5287
rect 57345 5253 57379 5287
rect 57379 5253 57388 5287
rect 57336 5244 57388 5253
rect 35532 5219 35584 5228
rect 35532 5185 35541 5219
rect 35541 5185 35575 5219
rect 35575 5185 35584 5219
rect 35532 5176 35584 5185
rect 35808 5219 35860 5228
rect 35808 5185 35817 5219
rect 35817 5185 35851 5219
rect 35851 5185 35860 5219
rect 35808 5176 35860 5185
rect 940 5108 992 5160
rect 19984 5151 20036 5160
rect 19984 5117 19993 5151
rect 19993 5117 20027 5151
rect 20027 5117 20036 5151
rect 19984 5108 20036 5117
rect 21272 5151 21324 5160
rect 21272 5117 21281 5151
rect 21281 5117 21315 5151
rect 21315 5117 21324 5151
rect 21272 5108 21324 5117
rect 21732 5108 21784 5160
rect 22836 5151 22888 5160
rect 22836 5117 22845 5151
rect 22845 5117 22879 5151
rect 22879 5117 22888 5151
rect 22836 5108 22888 5117
rect 27712 5108 27764 5160
rect 30104 5108 30156 5160
rect 31944 5108 31996 5160
rect 32312 5151 32364 5160
rect 32312 5117 32321 5151
rect 32321 5117 32355 5151
rect 32355 5117 32364 5151
rect 32312 5108 32364 5117
rect 36268 5219 36320 5228
rect 36268 5185 36277 5219
rect 36277 5185 36311 5219
rect 36311 5185 36320 5219
rect 36268 5176 36320 5185
rect 36728 5219 36780 5228
rect 36728 5185 36737 5219
rect 36737 5185 36771 5219
rect 36771 5185 36780 5219
rect 36728 5176 36780 5185
rect 37556 5219 37608 5228
rect 37556 5185 37565 5219
rect 37565 5185 37599 5219
rect 37599 5185 37608 5219
rect 37556 5176 37608 5185
rect 39120 5219 39172 5228
rect 39120 5185 39129 5219
rect 39129 5185 39163 5219
rect 39163 5185 39172 5219
rect 39120 5176 39172 5185
rect 39396 5219 39448 5228
rect 39396 5185 39430 5219
rect 39430 5185 39448 5219
rect 39396 5176 39448 5185
rect 41052 5219 41104 5228
rect 41052 5185 41061 5219
rect 41061 5185 41095 5219
rect 41095 5185 41104 5219
rect 41052 5176 41104 5185
rect 41236 5176 41288 5228
rect 43260 5219 43312 5228
rect 43260 5185 43269 5219
rect 43269 5185 43303 5219
rect 43303 5185 43312 5219
rect 43260 5176 43312 5185
rect 44548 5176 44600 5228
rect 44824 5176 44876 5228
rect 1584 5040 1636 5092
rect 20352 5040 20404 5092
rect 23480 5040 23532 5092
rect 22100 4972 22152 5024
rect 24860 4972 24912 5024
rect 25044 4972 25096 5024
rect 26608 4972 26660 5024
rect 26700 4972 26752 5024
rect 30196 4972 30248 5024
rect 33692 5083 33744 5092
rect 33692 5049 33701 5083
rect 33701 5049 33735 5083
rect 33735 5049 33744 5083
rect 33692 5040 33744 5049
rect 35348 5040 35400 5092
rect 34704 5015 34756 5024
rect 34704 4981 34713 5015
rect 34713 4981 34747 5015
rect 34747 4981 34756 5015
rect 34704 4972 34756 4981
rect 37832 5151 37884 5160
rect 37832 5117 37841 5151
rect 37841 5117 37875 5151
rect 37875 5117 37884 5151
rect 37832 5108 37884 5117
rect 42892 5108 42944 5160
rect 45376 5176 45428 5228
rect 46204 5176 46256 5228
rect 45468 5108 45520 5160
rect 46664 5108 46716 5160
rect 41880 5040 41932 5092
rect 41972 5083 42024 5092
rect 41972 5049 41981 5083
rect 41981 5049 42015 5083
rect 42015 5049 42024 5083
rect 41972 5040 42024 5049
rect 42432 5040 42484 5092
rect 45376 5040 45428 5092
rect 46480 5083 46532 5092
rect 46480 5049 46489 5083
rect 46489 5049 46523 5083
rect 46523 5049 46532 5083
rect 46480 5040 46532 5049
rect 55680 5176 55732 5228
rect 57060 5219 57112 5228
rect 57060 5185 57069 5219
rect 57069 5185 57103 5219
rect 57103 5185 57112 5219
rect 57060 5176 57112 5185
rect 58072 5219 58124 5228
rect 58072 5185 58081 5219
rect 58081 5185 58115 5219
rect 58115 5185 58124 5219
rect 58072 5176 58124 5185
rect 58992 5108 59044 5160
rect 57336 5040 57388 5092
rect 58900 4972 58952 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 15844 4768 15896 4820
rect 12072 4700 12124 4752
rect 18236 4768 18288 4820
rect 21732 4768 21784 4820
rect 27712 4811 27764 4820
rect 27712 4777 27721 4811
rect 27721 4777 27755 4811
rect 27755 4777 27764 4811
rect 27712 4768 27764 4777
rect 27804 4768 27856 4820
rect 38108 4768 38160 4820
rect 39396 4768 39448 4820
rect 22008 4700 22060 4752
rect 18144 4632 18196 4684
rect 24308 4700 24360 4752
rect 25596 4700 25648 4752
rect 31208 4700 31260 4752
rect 32772 4700 32824 4752
rect 33692 4700 33744 4752
rect 35348 4700 35400 4752
rect 1584 4607 1636 4616
rect 1584 4573 1593 4607
rect 1593 4573 1627 4607
rect 1627 4573 1636 4607
rect 1584 4564 1636 4573
rect 18052 4564 18104 4616
rect 22284 4632 22336 4684
rect 23296 4632 23348 4684
rect 24124 4632 24176 4684
rect 27896 4632 27948 4684
rect 28448 4632 28500 4684
rect 20352 4607 20404 4616
rect 20352 4573 20361 4607
rect 20361 4573 20395 4607
rect 20395 4573 20404 4607
rect 20352 4564 20404 4573
rect 20904 4564 20956 4616
rect 940 4496 992 4548
rect 10324 4496 10376 4548
rect 11428 4496 11480 4548
rect 20260 4496 20312 4548
rect 20812 4496 20864 4548
rect 21364 4539 21416 4548
rect 21364 4505 21373 4539
rect 21373 4505 21407 4539
rect 21407 4505 21416 4539
rect 21364 4496 21416 4505
rect 23572 4496 23624 4548
rect 24584 4607 24636 4616
rect 24584 4573 24593 4607
rect 24593 4573 24627 4607
rect 24627 4573 24636 4607
rect 24584 4564 24636 4573
rect 24860 4607 24912 4616
rect 24860 4573 24894 4607
rect 24894 4573 24912 4607
rect 24860 4564 24912 4573
rect 27068 4564 27120 4616
rect 27712 4564 27764 4616
rect 27988 4607 28040 4616
rect 27988 4573 27997 4607
rect 27997 4573 28031 4607
rect 28031 4573 28040 4607
rect 27988 4564 28040 4573
rect 28080 4607 28132 4616
rect 28080 4573 28089 4607
rect 28089 4573 28123 4607
rect 28123 4573 28132 4607
rect 28080 4564 28132 4573
rect 28172 4607 28224 4616
rect 28172 4573 28181 4607
rect 28181 4573 28215 4607
rect 28215 4573 28224 4607
rect 28172 4564 28224 4573
rect 29460 4564 29512 4616
rect 31760 4564 31812 4616
rect 36360 4632 36412 4684
rect 27804 4496 27856 4548
rect 17132 4428 17184 4480
rect 20904 4428 20956 4480
rect 22560 4471 22612 4480
rect 22560 4437 22569 4471
rect 22569 4437 22603 4471
rect 22603 4437 22612 4471
rect 22560 4428 22612 4437
rect 23296 4428 23348 4480
rect 24768 4428 24820 4480
rect 27988 4428 28040 4480
rect 29552 4496 29604 4548
rect 31852 4496 31904 4548
rect 32128 4607 32180 4616
rect 32128 4573 32137 4607
rect 32137 4573 32171 4607
rect 32171 4573 32180 4607
rect 32128 4564 32180 4573
rect 32220 4496 32272 4548
rect 32404 4564 32456 4616
rect 32956 4564 33008 4616
rect 33508 4564 33560 4616
rect 33692 4564 33744 4616
rect 34060 4564 34112 4616
rect 35164 4607 35216 4616
rect 35164 4573 35173 4607
rect 35173 4573 35207 4607
rect 35207 4573 35216 4607
rect 35164 4564 35216 4573
rect 35716 4564 35768 4616
rect 35900 4607 35952 4616
rect 35900 4573 35909 4607
rect 35909 4573 35943 4607
rect 35943 4573 35952 4607
rect 35900 4564 35952 4573
rect 35992 4607 36044 4616
rect 35992 4573 36001 4607
rect 36001 4573 36035 4607
rect 36035 4573 36044 4607
rect 35992 4564 36044 4573
rect 37832 4700 37884 4752
rect 37188 4675 37240 4684
rect 37188 4641 37197 4675
rect 37197 4641 37231 4675
rect 37231 4641 37240 4675
rect 37188 4632 37240 4641
rect 37096 4564 37148 4616
rect 37740 4564 37792 4616
rect 40132 4700 40184 4752
rect 40868 4700 40920 4752
rect 42156 4811 42208 4820
rect 42156 4777 42165 4811
rect 42165 4777 42199 4811
rect 42199 4777 42208 4811
rect 42156 4768 42208 4777
rect 43168 4768 43220 4820
rect 46848 4768 46900 4820
rect 48688 4811 48740 4820
rect 48688 4777 48697 4811
rect 48697 4777 48731 4811
rect 48731 4777 48740 4811
rect 48688 4768 48740 4777
rect 42892 4700 42944 4752
rect 48228 4700 48280 4752
rect 48412 4700 48464 4752
rect 40224 4632 40276 4684
rect 40684 4675 40736 4684
rect 40684 4641 40693 4675
rect 40693 4641 40727 4675
rect 40727 4641 40736 4675
rect 40684 4632 40736 4641
rect 46388 4632 46440 4684
rect 28264 4428 28316 4480
rect 32588 4428 32640 4480
rect 33048 4539 33100 4548
rect 33048 4505 33057 4539
rect 33057 4505 33091 4539
rect 33091 4505 33100 4539
rect 33048 4496 33100 4505
rect 34152 4496 34204 4548
rect 37556 4496 37608 4548
rect 33140 4428 33192 4480
rect 36360 4428 36412 4480
rect 36636 4471 36688 4480
rect 36636 4437 36645 4471
rect 36645 4437 36679 4471
rect 36679 4437 36688 4471
rect 36636 4428 36688 4437
rect 37188 4428 37240 4480
rect 40408 4564 40460 4616
rect 43352 4564 43404 4616
rect 46480 4564 46532 4616
rect 48044 4607 48096 4616
rect 48044 4573 48053 4607
rect 48053 4573 48087 4607
rect 48087 4573 48096 4607
rect 48044 4564 48096 4573
rect 38660 4496 38712 4548
rect 40132 4428 40184 4480
rect 40316 4428 40368 4480
rect 41328 4539 41380 4548
rect 41328 4505 41337 4539
rect 41337 4505 41371 4539
rect 41371 4505 41380 4539
rect 41328 4496 41380 4505
rect 42064 4496 42116 4548
rect 45652 4496 45704 4548
rect 46020 4496 46072 4548
rect 42892 4471 42944 4480
rect 42892 4437 42901 4471
rect 42901 4437 42935 4471
rect 42935 4437 42944 4471
rect 42892 4428 42944 4437
rect 47400 4471 47452 4480
rect 47400 4437 47409 4471
rect 47409 4437 47443 4471
rect 47443 4437 47452 4471
rect 47400 4428 47452 4437
rect 48320 4607 48372 4616
rect 48320 4573 48329 4607
rect 48329 4573 48363 4607
rect 48363 4573 48372 4607
rect 48320 4564 48372 4573
rect 56416 4632 56468 4684
rect 56784 4632 56836 4684
rect 49240 4564 49292 4616
rect 55404 4564 55456 4616
rect 56324 4564 56376 4616
rect 48780 4496 48832 4548
rect 55496 4496 55548 4548
rect 56968 4496 57020 4548
rect 53472 4428 53524 4480
rect 58256 4471 58308 4480
rect 58256 4437 58265 4471
rect 58265 4437 58299 4471
rect 58299 4437 58308 4471
rect 58256 4428 58308 4437
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 50294 4326 50346 4378
rect 50358 4326 50410 4378
rect 50422 4326 50474 4378
rect 50486 4326 50538 4378
rect 50550 4326 50602 4378
rect 8944 4156 8996 4208
rect 8116 4088 8168 4140
rect 11060 4156 11112 4208
rect 10140 4131 10192 4140
rect 10140 4097 10149 4131
rect 10149 4097 10183 4131
rect 10183 4097 10192 4131
rect 10140 4088 10192 4097
rect 9680 4020 9732 4072
rect 4620 3952 4672 4004
rect 10048 4063 10100 4072
rect 10048 4029 10057 4063
rect 10057 4029 10091 4063
rect 10091 4029 10100 4063
rect 10048 4020 10100 4029
rect 10232 4063 10284 4072
rect 10232 4029 10241 4063
rect 10241 4029 10275 4063
rect 10275 4029 10284 4063
rect 10232 4020 10284 4029
rect 11520 4088 11572 4140
rect 25044 4224 25096 4276
rect 25228 4267 25280 4276
rect 25228 4233 25237 4267
rect 25237 4233 25271 4267
rect 25271 4233 25280 4267
rect 25228 4224 25280 4233
rect 27988 4224 28040 4276
rect 15568 4156 15620 4208
rect 21364 4156 21416 4208
rect 22928 4156 22980 4208
rect 11980 3995 12032 4004
rect 11980 3961 11989 3995
rect 11989 3961 12023 3995
rect 12023 3961 12032 3995
rect 11980 3952 12032 3961
rect 11888 3884 11940 3936
rect 15108 4088 15160 4140
rect 15660 4088 15712 4140
rect 17040 4088 17092 4140
rect 17316 4131 17368 4140
rect 17316 4097 17325 4131
rect 17325 4097 17359 4131
rect 17359 4097 17368 4131
rect 17316 4088 17368 4097
rect 19156 4131 19208 4140
rect 19156 4097 19165 4131
rect 19165 4097 19199 4131
rect 19199 4097 19208 4131
rect 19156 4088 19208 4097
rect 19432 4131 19484 4140
rect 19432 4097 19441 4131
rect 19441 4097 19475 4131
rect 19475 4097 19484 4131
rect 19432 4088 19484 4097
rect 20444 4088 20496 4140
rect 22284 4088 22336 4140
rect 12716 4020 12768 4072
rect 16120 4020 16172 4072
rect 17224 4020 17276 4072
rect 19892 3952 19944 4004
rect 12716 3884 12768 3936
rect 12992 3884 13044 3936
rect 13360 3884 13412 3936
rect 18144 3884 18196 3936
rect 18328 3884 18380 3936
rect 18696 3884 18748 3936
rect 20444 3952 20496 4004
rect 21548 3952 21600 4004
rect 22560 4088 22612 4140
rect 24492 4088 24544 4140
rect 24676 4088 24728 4140
rect 25780 4156 25832 4208
rect 27896 4156 27948 4208
rect 28540 4199 28592 4208
rect 28540 4165 28549 4199
rect 28549 4165 28583 4199
rect 28583 4165 28592 4199
rect 28540 4156 28592 4165
rect 23204 4020 23256 4072
rect 23572 4063 23624 4072
rect 23572 4029 23581 4063
rect 23581 4029 23615 4063
rect 23615 4029 23624 4063
rect 23572 4020 23624 4029
rect 25688 4063 25740 4072
rect 25688 4029 25697 4063
rect 25697 4029 25731 4063
rect 25731 4029 25740 4063
rect 25688 4020 25740 4029
rect 25780 4063 25832 4072
rect 25780 4029 25789 4063
rect 25789 4029 25823 4063
rect 25823 4029 25832 4063
rect 25780 4020 25832 4029
rect 24032 3952 24084 4004
rect 24584 3952 24636 4004
rect 25872 3952 25924 4004
rect 27436 3952 27488 4004
rect 27620 4063 27672 4072
rect 27620 4029 27629 4063
rect 27629 4029 27663 4063
rect 27663 4029 27672 4063
rect 27620 4020 27672 4029
rect 29184 4131 29236 4140
rect 29184 4097 29193 4131
rect 29193 4097 29227 4131
rect 29227 4097 29236 4131
rect 29184 4088 29236 4097
rect 30472 4224 30524 4276
rect 32128 4224 32180 4276
rect 29552 4156 29604 4208
rect 37188 4224 37240 4276
rect 37280 4224 37332 4276
rect 30012 4088 30064 4140
rect 31392 4131 31444 4140
rect 31392 4097 31401 4131
rect 31401 4097 31435 4131
rect 31435 4097 31444 4131
rect 31392 4088 31444 4097
rect 30380 4020 30432 4072
rect 32312 4131 32364 4140
rect 32312 4097 32321 4131
rect 32321 4097 32355 4131
rect 32355 4097 32364 4131
rect 36176 4156 36228 4208
rect 36544 4156 36596 4208
rect 39212 4224 39264 4276
rect 32312 4088 32364 4097
rect 34704 4131 34756 4140
rect 34704 4097 34713 4131
rect 34713 4097 34747 4131
rect 34747 4097 34756 4131
rect 34704 4088 34756 4097
rect 35440 4088 35492 4140
rect 22836 3884 22888 3936
rect 23756 3884 23808 3936
rect 26976 3884 27028 3936
rect 27160 3927 27212 3936
rect 27160 3893 27169 3927
rect 27169 3893 27203 3927
rect 27203 3893 27212 3927
rect 27160 3884 27212 3893
rect 32220 3952 32272 4004
rect 30288 3884 30340 3936
rect 32588 4063 32640 4072
rect 32588 4029 32597 4063
rect 32597 4029 32631 4063
rect 32631 4029 32640 4063
rect 32588 4020 32640 4029
rect 34612 4020 34664 4072
rect 35348 4020 35400 4072
rect 36084 4020 36136 4072
rect 39120 4156 39172 4208
rect 38200 4088 38252 4140
rect 38568 4088 38620 4140
rect 39028 4088 39080 4140
rect 40132 4224 40184 4276
rect 41052 4224 41104 4276
rect 44640 4224 44692 4276
rect 45192 4224 45244 4276
rect 44364 4156 44416 4208
rect 48044 4224 48096 4276
rect 40040 4088 40092 4140
rect 41052 4131 41104 4140
rect 41052 4097 41061 4131
rect 41061 4097 41095 4131
rect 41095 4097 41104 4131
rect 41052 4088 41104 4097
rect 41788 4131 41840 4140
rect 41788 4097 41797 4131
rect 41797 4097 41831 4131
rect 41831 4097 41840 4131
rect 41788 4088 41840 4097
rect 42708 4131 42760 4140
rect 42708 4097 42717 4131
rect 42717 4097 42751 4131
rect 42751 4097 42760 4131
rect 42708 4088 42760 4097
rect 42984 4088 43036 4140
rect 43352 4131 43404 4140
rect 43352 4097 43361 4131
rect 43361 4097 43395 4131
rect 43395 4097 43404 4131
rect 43352 4088 43404 4097
rect 38752 4020 38804 4072
rect 39120 4020 39172 4072
rect 40776 4020 40828 4072
rect 42616 4020 42668 4072
rect 43536 3995 43588 4004
rect 43536 3961 43545 3995
rect 43545 3961 43579 3995
rect 43579 3961 43588 3995
rect 43536 3952 43588 3961
rect 44272 3995 44324 4004
rect 44272 3961 44281 3995
rect 44281 3961 44315 3995
rect 44315 3961 44324 3995
rect 44272 3952 44324 3961
rect 36728 3927 36780 3936
rect 36728 3893 36737 3927
rect 36737 3893 36771 3927
rect 36771 3893 36780 3927
rect 36728 3884 36780 3893
rect 38200 3884 38252 3936
rect 40040 3884 40092 3936
rect 40224 3884 40276 3936
rect 43168 3884 43220 3936
rect 47492 4088 47544 4140
rect 47768 4131 47820 4140
rect 47768 4097 47777 4131
rect 47777 4097 47811 4131
rect 47811 4097 47820 4131
rect 47768 4088 47820 4097
rect 48320 4088 48372 4140
rect 47124 4020 47176 4072
rect 48596 4131 48648 4140
rect 48596 4097 48605 4131
rect 48605 4097 48639 4131
rect 48639 4097 48648 4131
rect 48596 4088 48648 4097
rect 48872 4131 48924 4140
rect 48872 4097 48881 4131
rect 48881 4097 48915 4131
rect 48915 4097 48924 4131
rect 48872 4088 48924 4097
rect 51172 4224 51224 4276
rect 50528 4199 50580 4208
rect 50528 4165 50537 4199
rect 50537 4165 50571 4199
rect 50571 4165 50580 4199
rect 50528 4156 50580 4165
rect 50712 4156 50764 4208
rect 55220 4156 55272 4208
rect 58808 4156 58860 4208
rect 51356 4088 51408 4140
rect 52276 4088 52328 4140
rect 56876 4088 56928 4140
rect 57336 4131 57388 4140
rect 57336 4097 57345 4131
rect 57345 4097 57379 4131
rect 57379 4097 57388 4131
rect 57336 4088 57388 4097
rect 58072 4131 58124 4140
rect 58072 4097 58081 4131
rect 58081 4097 58115 4131
rect 58115 4097 58124 4131
rect 58072 4088 58124 4097
rect 52920 4020 52972 4072
rect 53748 4020 53800 4072
rect 48320 3952 48372 4004
rect 46664 3884 46716 3936
rect 56324 4063 56376 4072
rect 56324 4029 56333 4063
rect 56333 4029 56367 4063
rect 56367 4029 56376 4063
rect 56324 4020 56376 4029
rect 49516 3884 49568 3936
rect 50528 3884 50580 3936
rect 50620 3927 50672 3936
rect 50620 3893 50629 3927
rect 50629 3893 50663 3927
rect 50663 3893 50672 3927
rect 50620 3884 50672 3893
rect 51448 3884 51500 3936
rect 54852 3884 54904 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 8484 3723 8536 3732
rect 8484 3689 8493 3723
rect 8493 3689 8527 3723
rect 8527 3689 8536 3723
rect 8484 3680 8536 3689
rect 9588 3680 9640 3732
rect 9772 3680 9824 3732
rect 9404 3612 9456 3664
rect 7656 3544 7708 3596
rect 13544 3680 13596 3732
rect 14464 3723 14516 3732
rect 14464 3689 14473 3723
rect 14473 3689 14507 3723
rect 14507 3689 14516 3723
rect 14464 3680 14516 3689
rect 15292 3723 15344 3732
rect 15292 3689 15301 3723
rect 15301 3689 15335 3723
rect 15335 3689 15344 3723
rect 15292 3680 15344 3689
rect 16028 3723 16080 3732
rect 16028 3689 16037 3723
rect 16037 3689 16071 3723
rect 16071 3689 16080 3723
rect 16028 3680 16080 3689
rect 16672 3680 16724 3732
rect 20444 3680 20496 3732
rect 20720 3680 20772 3732
rect 27620 3680 27672 3732
rect 27896 3680 27948 3732
rect 17132 3612 17184 3664
rect 17316 3612 17368 3664
rect 21180 3612 21232 3664
rect 22100 3612 22152 3664
rect 23020 3612 23072 3664
rect 9680 3544 9732 3596
rect 10048 3587 10100 3596
rect 10048 3553 10057 3587
rect 10057 3553 10091 3587
rect 10091 3553 10100 3587
rect 10048 3544 10100 3553
rect 12716 3544 12768 3596
rect 9772 3476 9824 3528
rect 7564 3408 7616 3460
rect 8208 3408 8260 3460
rect 8668 3408 8720 3460
rect 10048 3340 10100 3392
rect 10876 3340 10928 3392
rect 12072 3340 12124 3392
rect 12624 3340 12676 3392
rect 12808 3451 12860 3460
rect 12808 3417 12817 3451
rect 12817 3417 12851 3451
rect 12851 3417 12860 3451
rect 12808 3408 12860 3417
rect 13360 3408 13412 3460
rect 14188 3408 14240 3460
rect 15292 3408 15344 3460
rect 16120 3408 16172 3460
rect 16672 3476 16724 3528
rect 17960 3476 18012 3528
rect 18512 3476 18564 3528
rect 16764 3408 16816 3460
rect 16948 3408 17000 3460
rect 17592 3408 17644 3460
rect 18696 3451 18748 3460
rect 18696 3417 18705 3451
rect 18705 3417 18739 3451
rect 18739 3417 18748 3451
rect 18696 3408 18748 3417
rect 20536 3476 20588 3528
rect 21916 3519 21968 3528
rect 21916 3485 21925 3519
rect 21925 3485 21959 3519
rect 21959 3485 21968 3519
rect 21916 3476 21968 3485
rect 20168 3408 20220 3460
rect 20352 3451 20404 3460
rect 20352 3417 20361 3451
rect 20361 3417 20395 3451
rect 20395 3417 20404 3451
rect 20352 3408 20404 3417
rect 23480 3544 23532 3596
rect 23848 3612 23900 3664
rect 25320 3612 25372 3664
rect 29368 3612 29420 3664
rect 31576 3680 31628 3732
rect 32220 3680 32272 3732
rect 35808 3680 35860 3732
rect 22560 3476 22612 3528
rect 22744 3408 22796 3460
rect 23020 3451 23072 3460
rect 23020 3417 23029 3451
rect 23029 3417 23063 3451
rect 23063 3417 23072 3451
rect 23020 3408 23072 3417
rect 23112 3451 23164 3460
rect 23112 3417 23131 3451
rect 23131 3417 23164 3451
rect 24952 3519 25004 3528
rect 24952 3485 24961 3519
rect 24961 3485 24995 3519
rect 24995 3485 25004 3519
rect 24952 3476 25004 3485
rect 25872 3587 25924 3596
rect 25872 3553 25881 3587
rect 25881 3553 25915 3587
rect 25915 3553 25924 3587
rect 25872 3544 25924 3553
rect 26976 3544 27028 3596
rect 30380 3544 30432 3596
rect 30472 3587 30524 3596
rect 30472 3553 30481 3587
rect 30481 3553 30515 3587
rect 30515 3553 30524 3587
rect 30472 3544 30524 3553
rect 25964 3476 26016 3528
rect 27160 3476 27212 3528
rect 28908 3476 28960 3528
rect 30288 3519 30340 3528
rect 30288 3485 30297 3519
rect 30297 3485 30331 3519
rect 30331 3485 30340 3519
rect 30288 3476 30340 3485
rect 31024 3519 31076 3528
rect 31024 3485 31033 3519
rect 31033 3485 31067 3519
rect 31067 3485 31076 3519
rect 31024 3476 31076 3485
rect 32128 3612 32180 3664
rect 31300 3519 31352 3528
rect 31300 3485 31309 3519
rect 31309 3485 31343 3519
rect 31343 3485 31352 3519
rect 31300 3476 31352 3485
rect 31484 3544 31536 3596
rect 32404 3544 32456 3596
rect 34060 3544 34112 3596
rect 23112 3408 23164 3417
rect 12992 3340 13044 3392
rect 16580 3340 16632 3392
rect 19432 3340 19484 3392
rect 20444 3340 20496 3392
rect 23296 3340 23348 3392
rect 23940 3383 23992 3392
rect 23940 3349 23949 3383
rect 23949 3349 23983 3383
rect 23983 3349 23992 3383
rect 23940 3340 23992 3349
rect 25780 3408 25832 3460
rect 26240 3408 26292 3460
rect 27160 3340 27212 3392
rect 28816 3340 28868 3392
rect 29736 3340 29788 3392
rect 30012 3340 30064 3392
rect 30288 3340 30340 3392
rect 32036 3476 32088 3528
rect 32128 3340 32180 3392
rect 32956 3519 33008 3528
rect 32956 3485 32965 3519
rect 32965 3485 32999 3519
rect 32999 3485 33008 3519
rect 32956 3476 33008 3485
rect 33968 3476 34020 3528
rect 36544 3680 36596 3732
rect 37464 3680 37516 3732
rect 37924 3680 37976 3732
rect 38936 3680 38988 3732
rect 38200 3612 38252 3664
rect 42708 3680 42760 3732
rect 42984 3680 43036 3732
rect 44088 3680 44140 3732
rect 44180 3723 44232 3732
rect 44180 3689 44189 3723
rect 44189 3689 44223 3723
rect 44223 3689 44232 3723
rect 44180 3680 44232 3689
rect 36176 3544 36228 3596
rect 37372 3544 37424 3596
rect 41788 3612 41840 3664
rect 36360 3476 36412 3528
rect 32864 3408 32916 3460
rect 33232 3408 33284 3460
rect 39212 3476 39264 3528
rect 38476 3408 38528 3460
rect 39120 3408 39172 3460
rect 39396 3519 39448 3528
rect 39396 3485 39405 3519
rect 39405 3485 39439 3519
rect 39439 3485 39448 3519
rect 43444 3544 43496 3596
rect 39396 3476 39448 3485
rect 40040 3408 40092 3460
rect 41052 3408 41104 3460
rect 35992 3340 36044 3392
rect 40960 3383 41012 3392
rect 40960 3349 40969 3383
rect 40969 3349 41003 3383
rect 41003 3349 41012 3383
rect 40960 3340 41012 3349
rect 42800 3476 42852 3528
rect 42892 3519 42944 3528
rect 42892 3485 42901 3519
rect 42901 3485 42935 3519
rect 42935 3485 42944 3519
rect 42892 3476 42944 3485
rect 42984 3519 43036 3528
rect 42984 3485 42993 3519
rect 42993 3485 43027 3519
rect 43027 3485 43036 3519
rect 42984 3476 43036 3485
rect 43076 3476 43128 3528
rect 43720 3519 43772 3528
rect 43720 3485 43727 3519
rect 43727 3485 43772 3519
rect 43720 3476 43772 3485
rect 43904 3519 43956 3528
rect 43904 3485 43913 3519
rect 43913 3485 43947 3519
rect 43947 3485 43956 3519
rect 43904 3476 43956 3485
rect 44180 3476 44232 3528
rect 47308 3612 47360 3664
rect 47584 3723 47636 3732
rect 47584 3689 47593 3723
rect 47593 3689 47627 3723
rect 47627 3689 47636 3723
rect 47584 3680 47636 3689
rect 49976 3680 50028 3732
rect 53472 3723 53524 3732
rect 53472 3689 53481 3723
rect 53481 3689 53515 3723
rect 53515 3689 53524 3723
rect 53472 3680 53524 3689
rect 54208 3723 54260 3732
rect 54208 3689 54217 3723
rect 54217 3689 54251 3723
rect 54251 3689 54260 3723
rect 54208 3680 54260 3689
rect 50620 3612 50672 3664
rect 52184 3612 52236 3664
rect 53656 3612 53708 3664
rect 41880 3451 41932 3460
rect 41880 3417 41889 3451
rect 41889 3417 41923 3451
rect 41923 3417 41932 3451
rect 41880 3408 41932 3417
rect 44456 3408 44508 3460
rect 45468 3408 45520 3460
rect 57336 3544 57388 3596
rect 47400 3519 47452 3528
rect 47400 3485 47414 3519
rect 47414 3485 47448 3519
rect 47448 3485 47452 3519
rect 47400 3476 47452 3485
rect 47952 3476 48004 3528
rect 48596 3519 48648 3528
rect 48596 3485 48605 3519
rect 48605 3485 48639 3519
rect 48639 3485 48648 3519
rect 48596 3476 48648 3485
rect 48780 3519 48832 3528
rect 48780 3485 48789 3519
rect 48789 3485 48823 3519
rect 48823 3485 48832 3519
rect 48780 3476 48832 3485
rect 47216 3451 47268 3460
rect 47216 3417 47225 3451
rect 47225 3417 47259 3451
rect 47259 3417 47268 3451
rect 47216 3408 47268 3417
rect 47308 3451 47360 3460
rect 47308 3417 47317 3451
rect 47317 3417 47351 3451
rect 47351 3417 47360 3451
rect 47308 3408 47360 3417
rect 49240 3519 49292 3528
rect 49240 3485 49249 3519
rect 49249 3485 49283 3519
rect 49283 3485 49292 3519
rect 49240 3476 49292 3485
rect 49976 3476 50028 3528
rect 50436 3476 50488 3528
rect 51448 3476 51500 3528
rect 53104 3476 53156 3528
rect 54760 3519 54812 3528
rect 54760 3485 54769 3519
rect 54769 3485 54803 3519
rect 54803 3485 54812 3519
rect 54760 3476 54812 3485
rect 55496 3476 55548 3528
rect 56416 3476 56468 3528
rect 42984 3340 43036 3392
rect 43628 3340 43680 3392
rect 44088 3340 44140 3392
rect 49792 3408 49844 3460
rect 50068 3340 50120 3392
rect 52000 3408 52052 3460
rect 56876 3408 56928 3460
rect 56784 3340 56836 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 50294 3238 50346 3290
rect 50358 3238 50410 3290
rect 50422 3238 50474 3290
rect 50486 3238 50538 3290
rect 50550 3238 50602 3290
rect 7656 3179 7708 3188
rect 7656 3145 7665 3179
rect 7665 3145 7699 3179
rect 7699 3145 7708 3179
rect 7656 3136 7708 3145
rect 12072 3136 12124 3188
rect 9588 3068 9640 3120
rect 10048 3068 10100 3120
rect 5908 3000 5960 3052
rect 6828 3043 6880 3052
rect 6828 3009 6837 3043
rect 6837 3009 6871 3043
rect 6871 3009 6880 3043
rect 6828 3000 6880 3009
rect 7932 3000 7984 3052
rect 9036 3043 9088 3052
rect 9036 3009 9045 3043
rect 9045 3009 9079 3043
rect 9079 3009 9088 3043
rect 9036 3000 9088 3009
rect 9128 3000 9180 3052
rect 11980 3068 12032 3120
rect 13820 3179 13872 3188
rect 13820 3145 13829 3179
rect 13829 3145 13863 3179
rect 13863 3145 13872 3179
rect 13820 3136 13872 3145
rect 18604 3136 18656 3188
rect 17960 3068 18012 3120
rect 21916 3136 21968 3188
rect 10968 3043 11020 3052
rect 10968 3009 10977 3043
rect 10977 3009 11011 3043
rect 11011 3009 11020 3043
rect 10968 3000 11020 3009
rect 10232 2932 10284 2984
rect 10876 2932 10928 2984
rect 13636 3000 13688 3052
rect 13728 3043 13780 3052
rect 13728 3009 13737 3043
rect 13737 3009 13771 3043
rect 13771 3009 13780 3043
rect 13728 3000 13780 3009
rect 15016 3000 15068 3052
rect 15752 3000 15804 3052
rect 15844 3043 15896 3052
rect 15844 3009 15853 3043
rect 15853 3009 15887 3043
rect 15887 3009 15896 3043
rect 15844 3000 15896 3009
rect 18236 3000 18288 3052
rect 22100 3068 22152 3120
rect 13084 2932 13136 2984
rect 13912 2932 13964 2984
rect 8300 2864 8352 2916
rect 11888 2864 11940 2916
rect 16488 2932 16540 2984
rect 17868 2932 17920 2984
rect 21180 3000 21232 3052
rect 21456 3000 21508 3052
rect 19432 2932 19484 2984
rect 20352 2932 20404 2984
rect 23756 3136 23808 3188
rect 25688 3136 25740 3188
rect 25964 3136 26016 3188
rect 27160 3136 27212 3188
rect 33600 3136 33652 3188
rect 38476 3136 38528 3188
rect 41328 3136 41380 3188
rect 41696 3136 41748 3188
rect 43904 3179 43956 3188
rect 43904 3145 43913 3179
rect 43913 3145 43947 3179
rect 43947 3145 43956 3179
rect 43904 3136 43956 3145
rect 44640 3179 44692 3188
rect 44640 3145 44649 3179
rect 44649 3145 44683 3179
rect 44683 3145 44692 3179
rect 44640 3136 44692 3145
rect 22376 3068 22428 3120
rect 23940 3068 23992 3120
rect 25228 3068 25280 3120
rect 25320 3068 25372 3120
rect 27896 3068 27948 3120
rect 29828 3068 29880 3120
rect 23388 3000 23440 3052
rect 17316 2864 17368 2916
rect 18144 2864 18196 2916
rect 20996 2864 21048 2916
rect 15660 2796 15712 2848
rect 17040 2839 17092 2848
rect 17040 2805 17049 2839
rect 17049 2805 17083 2839
rect 17083 2805 17092 2839
rect 17040 2796 17092 2805
rect 20812 2796 20864 2848
rect 21548 2864 21600 2916
rect 22836 2975 22888 2984
rect 22836 2941 22845 2975
rect 22845 2941 22879 2975
rect 22879 2941 22888 2975
rect 22836 2932 22888 2941
rect 24492 3000 24544 3052
rect 26240 3043 26292 3052
rect 23756 2975 23808 2984
rect 23756 2941 23765 2975
rect 23765 2941 23799 2975
rect 23799 2941 23808 2975
rect 23756 2932 23808 2941
rect 24216 2864 24268 2916
rect 22652 2796 22704 2848
rect 22744 2796 22796 2848
rect 26240 3009 26249 3043
rect 26249 3009 26283 3043
rect 26283 3009 26292 3043
rect 26240 3000 26292 3009
rect 26516 2932 26568 2984
rect 29368 3000 29420 3052
rect 29736 3000 29788 3052
rect 32680 3068 32732 3120
rect 39120 3068 39172 3120
rect 31852 3000 31904 3052
rect 33048 3000 33100 3052
rect 34152 3043 34204 3052
rect 34152 3009 34161 3043
rect 34161 3009 34195 3043
rect 34195 3009 34204 3043
rect 34152 3000 34204 3009
rect 34244 3000 34296 3052
rect 35992 3043 36044 3052
rect 35992 3009 36001 3043
rect 36001 3009 36035 3043
rect 36035 3009 36044 3043
rect 35992 3000 36044 3009
rect 38292 3000 38344 3052
rect 38384 3043 38436 3052
rect 38384 3009 38393 3043
rect 38393 3009 38427 3043
rect 38427 3009 38436 3043
rect 38384 3000 38436 3009
rect 38660 3043 38712 3052
rect 38660 3009 38669 3043
rect 38669 3009 38703 3043
rect 38703 3009 38712 3043
rect 38660 3000 38712 3009
rect 39396 3000 39448 3052
rect 42800 3111 42852 3120
rect 42800 3077 42809 3111
rect 42809 3077 42843 3111
rect 42843 3077 42852 3111
rect 42800 3068 42852 3077
rect 46112 3136 46164 3188
rect 46296 3136 46348 3188
rect 44916 3068 44968 3120
rect 46388 3068 46440 3120
rect 40868 3000 40920 3052
rect 41512 3000 41564 3052
rect 42708 3000 42760 3052
rect 29092 2932 29144 2984
rect 29644 2932 29696 2984
rect 30196 2975 30248 2984
rect 30196 2941 30205 2975
rect 30205 2941 30239 2975
rect 30239 2941 30248 2975
rect 30196 2932 30248 2941
rect 30748 2932 30800 2984
rect 31576 2932 31628 2984
rect 31484 2864 31536 2916
rect 32128 2864 32180 2916
rect 33508 2864 33560 2916
rect 36176 2975 36228 2984
rect 36176 2941 36185 2975
rect 36185 2941 36219 2975
rect 36219 2941 36228 2975
rect 36176 2932 36228 2941
rect 37280 2932 37332 2984
rect 39672 2975 39724 2984
rect 39672 2941 39681 2975
rect 39681 2941 39715 2975
rect 39715 2941 39724 2975
rect 39672 2932 39724 2941
rect 43260 3000 43312 3052
rect 44088 3000 44140 3052
rect 45284 3043 45336 3052
rect 45284 3009 45293 3043
rect 45293 3009 45327 3043
rect 45327 3009 45336 3043
rect 45284 3000 45336 3009
rect 45376 3000 45428 3052
rect 46296 3000 46348 3052
rect 44180 2932 44232 2984
rect 48412 3136 48464 3188
rect 48504 3179 48556 3188
rect 48504 3145 48513 3179
rect 48513 3145 48547 3179
rect 48547 3145 48556 3179
rect 48504 3136 48556 3145
rect 48596 3136 48648 3188
rect 47308 3068 47360 3120
rect 52828 3136 52880 3188
rect 54576 3179 54628 3188
rect 54576 3145 54585 3179
rect 54585 3145 54619 3179
rect 54619 3145 54628 3179
rect 54576 3136 54628 3145
rect 55312 3179 55364 3188
rect 55312 3145 55321 3179
rect 55321 3145 55355 3179
rect 55355 3145 55364 3179
rect 55312 3136 55364 3145
rect 56968 3179 57020 3188
rect 56968 3145 56977 3179
rect 56977 3145 57011 3179
rect 57011 3145 57020 3179
rect 56968 3136 57020 3145
rect 58348 3068 58400 3120
rect 47860 3043 47912 3052
rect 47860 3009 47869 3043
rect 47869 3009 47903 3043
rect 47903 3009 47912 3043
rect 47860 3000 47912 3009
rect 48044 3043 48096 3052
rect 48044 3009 48051 3043
rect 48051 3009 48096 3043
rect 48044 3000 48096 3009
rect 47216 2932 47268 2984
rect 47768 2932 47820 2984
rect 48228 3043 48280 3052
rect 48228 3009 48237 3043
rect 48237 3009 48271 3043
rect 48271 3009 48280 3043
rect 48228 3000 48280 3009
rect 48412 3000 48464 3052
rect 48504 3000 48556 3052
rect 49424 3000 49476 3052
rect 50804 3043 50856 3052
rect 50804 3009 50813 3043
rect 50813 3009 50847 3043
rect 50847 3009 50856 3043
rect 50804 3000 50856 3009
rect 51540 3043 51592 3052
rect 51540 3009 51549 3043
rect 51549 3009 51583 3043
rect 51583 3009 51592 3043
rect 51540 3000 51592 3009
rect 52644 3000 52696 3052
rect 53012 3000 53064 3052
rect 54392 3043 54444 3052
rect 54392 3009 54401 3043
rect 54401 3009 54435 3043
rect 54435 3009 54444 3043
rect 54392 3000 54444 3009
rect 55220 3043 55272 3052
rect 55220 3009 55229 3043
rect 55229 3009 55263 3043
rect 55263 3009 55272 3043
rect 55220 3000 55272 3009
rect 55956 3043 56008 3052
rect 55956 3009 55965 3043
rect 55965 3009 55999 3043
rect 55999 3009 56008 3043
rect 55956 3000 56008 3009
rect 56140 3000 56192 3052
rect 56784 3043 56836 3052
rect 56784 3009 56793 3043
rect 56793 3009 56827 3043
rect 56827 3009 56836 3043
rect 56784 3000 56836 3009
rect 56968 3000 57020 3052
rect 48780 2932 48832 2984
rect 49056 2932 49108 2984
rect 38844 2864 38896 2916
rect 40592 2864 40644 2916
rect 43720 2864 43772 2916
rect 25964 2796 26016 2848
rect 28724 2796 28776 2848
rect 42892 2796 42944 2848
rect 45284 2796 45336 2848
rect 49240 2839 49292 2848
rect 49240 2805 49249 2839
rect 49249 2805 49283 2839
rect 49283 2805 49292 2839
rect 49240 2796 49292 2805
rect 49884 2796 49936 2848
rect 52460 2796 52512 2848
rect 56048 2839 56100 2848
rect 56048 2805 56057 2839
rect 56057 2805 56091 2839
rect 56091 2805 56100 2839
rect 56048 2796 56100 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 8392 2592 8444 2644
rect 8300 2524 8352 2576
rect 8760 2524 8812 2576
rect 10600 2524 10652 2576
rect 13176 2592 13228 2644
rect 13268 2592 13320 2644
rect 12532 2524 12584 2576
rect 13452 2524 13504 2576
rect 17776 2524 17828 2576
rect 5816 2363 5868 2372
rect 5816 2329 5825 2363
rect 5825 2329 5859 2363
rect 5859 2329 5868 2363
rect 5816 2320 5868 2329
rect 8024 2320 8076 2372
rect 8392 2363 8444 2372
rect 8392 2329 8401 2363
rect 8401 2329 8435 2363
rect 8435 2329 8444 2363
rect 8392 2320 8444 2329
rect 10048 2320 10100 2372
rect 10232 2363 10284 2372
rect 10232 2329 10241 2363
rect 10241 2329 10275 2363
rect 10275 2329 10284 2363
rect 10232 2320 10284 2329
rect 12532 2388 12584 2440
rect 11704 2320 11756 2372
rect 12072 2363 12124 2372
rect 12072 2329 12081 2363
rect 12081 2329 12115 2363
rect 12115 2329 12124 2363
rect 12072 2320 12124 2329
rect 13268 2320 13320 2372
rect 13544 2363 13596 2372
rect 13544 2329 13553 2363
rect 13553 2329 13587 2363
rect 13587 2329 13596 2363
rect 13544 2320 13596 2329
rect 16396 2456 16448 2508
rect 19432 2592 19484 2644
rect 27528 2592 27580 2644
rect 39764 2592 39816 2644
rect 41420 2635 41472 2644
rect 41420 2601 41429 2635
rect 41429 2601 41463 2635
rect 41463 2601 41472 2635
rect 41420 2592 41472 2601
rect 43812 2592 43864 2644
rect 44456 2635 44508 2644
rect 44456 2601 44465 2635
rect 44465 2601 44499 2635
rect 44499 2601 44508 2635
rect 44456 2592 44508 2601
rect 14924 2431 14976 2440
rect 14924 2397 14933 2431
rect 14933 2397 14967 2431
rect 14967 2397 14976 2431
rect 14924 2388 14976 2397
rect 15844 2431 15896 2440
rect 15844 2397 15853 2431
rect 15853 2397 15887 2431
rect 15887 2397 15896 2431
rect 15844 2388 15896 2397
rect 17408 2388 17460 2440
rect 20812 2456 20864 2508
rect 18236 2388 18288 2440
rect 18420 2431 18472 2440
rect 18420 2397 18429 2431
rect 18429 2397 18463 2431
rect 18463 2397 18472 2431
rect 18420 2388 18472 2397
rect 19340 2388 19392 2440
rect 20076 2431 20128 2440
rect 20076 2397 20085 2431
rect 20085 2397 20119 2431
rect 20119 2397 20128 2431
rect 20076 2388 20128 2397
rect 39212 2524 39264 2576
rect 46112 2635 46164 2644
rect 46112 2601 46121 2635
rect 46121 2601 46155 2635
rect 46155 2601 46164 2635
rect 46112 2592 46164 2601
rect 47124 2592 47176 2644
rect 49148 2592 49200 2644
rect 49332 2635 49384 2644
rect 49332 2601 49341 2635
rect 49341 2601 49375 2635
rect 49375 2601 49384 2635
rect 49332 2592 49384 2601
rect 49700 2592 49752 2644
rect 51632 2635 51684 2644
rect 51632 2601 51641 2635
rect 51641 2601 51675 2635
rect 51675 2601 51684 2635
rect 51632 2592 51684 2601
rect 52736 2592 52788 2644
rect 24124 2456 24176 2508
rect 21824 2388 21876 2440
rect 22652 2431 22704 2440
rect 22652 2397 22661 2431
rect 22661 2397 22695 2431
rect 22695 2397 22704 2431
rect 22652 2388 22704 2397
rect 15936 2252 15988 2304
rect 18604 2320 18656 2372
rect 19432 2252 19484 2304
rect 23296 2388 23348 2440
rect 23572 2431 23624 2440
rect 23572 2397 23581 2431
rect 23581 2397 23615 2431
rect 23615 2397 23624 2431
rect 23572 2388 23624 2397
rect 25228 2431 25280 2440
rect 25228 2397 25237 2431
rect 25237 2397 25271 2431
rect 25271 2397 25280 2431
rect 25228 2388 25280 2397
rect 44824 2456 44876 2508
rect 47032 2524 47084 2576
rect 48044 2524 48096 2576
rect 56876 2524 56928 2576
rect 48872 2456 48924 2508
rect 54300 2499 54352 2508
rect 54300 2465 54309 2499
rect 54309 2465 54343 2499
rect 54343 2465 54352 2499
rect 54300 2456 54352 2465
rect 26976 2388 27028 2440
rect 28724 2431 28776 2440
rect 28724 2397 28733 2431
rect 28733 2397 28767 2431
rect 28767 2397 28776 2431
rect 28724 2388 28776 2397
rect 30288 2388 30340 2440
rect 30840 2388 30892 2440
rect 31944 2388 31996 2440
rect 22468 2252 22520 2304
rect 24768 2320 24820 2372
rect 26056 2320 26108 2372
rect 26608 2320 26660 2372
rect 26884 2320 26936 2372
rect 29920 2320 29972 2372
rect 30472 2363 30524 2372
rect 30472 2329 30481 2363
rect 30481 2329 30515 2363
rect 30515 2329 30524 2363
rect 30472 2320 30524 2329
rect 31024 2320 31076 2372
rect 31760 2320 31812 2372
rect 33692 2388 33744 2440
rect 36728 2388 36780 2440
rect 32588 2363 32640 2372
rect 32588 2329 32597 2363
rect 32597 2329 32631 2363
rect 32631 2329 32640 2363
rect 32588 2320 32640 2329
rect 33140 2320 33192 2372
rect 34520 2320 34572 2372
rect 36084 2363 36136 2372
rect 36084 2329 36093 2363
rect 36093 2329 36127 2363
rect 36127 2329 36136 2363
rect 36084 2320 36136 2329
rect 24952 2252 25004 2304
rect 28908 2252 28960 2304
rect 37556 2388 37608 2440
rect 37740 2363 37792 2372
rect 37740 2329 37749 2363
rect 37749 2329 37783 2363
rect 37783 2329 37792 2363
rect 37740 2320 37792 2329
rect 37832 2320 37884 2372
rect 38660 2363 38712 2372
rect 38660 2329 38669 2363
rect 38669 2329 38703 2363
rect 38703 2329 38712 2363
rect 38660 2320 38712 2329
rect 39304 2388 39356 2440
rect 40316 2363 40368 2372
rect 40316 2329 40325 2363
rect 40325 2329 40359 2363
rect 40359 2329 40368 2363
rect 40316 2320 40368 2329
rect 40960 2320 41012 2372
rect 40868 2252 40920 2304
rect 41420 2388 41472 2440
rect 47952 2431 48004 2440
rect 47952 2397 47961 2431
rect 47961 2397 47995 2431
rect 47995 2397 48004 2431
rect 47952 2388 48004 2397
rect 48136 2431 48188 2440
rect 48136 2397 48143 2431
rect 48143 2397 48188 2431
rect 48136 2388 48188 2397
rect 48320 2431 48372 2440
rect 48320 2397 48329 2431
rect 48329 2397 48363 2431
rect 48363 2397 48372 2431
rect 48320 2388 48372 2397
rect 48596 2388 48648 2440
rect 51080 2388 51132 2440
rect 53932 2388 53984 2440
rect 58256 2524 58308 2576
rect 58348 2567 58400 2576
rect 58348 2533 58357 2567
rect 58357 2533 58391 2567
rect 58391 2533 58400 2567
rect 58348 2524 58400 2533
rect 58900 2456 58952 2508
rect 41788 2320 41840 2372
rect 43812 2320 43864 2372
rect 44456 2320 44508 2372
rect 46020 2363 46072 2372
rect 46020 2329 46029 2363
rect 46029 2329 46063 2363
rect 46063 2329 46072 2363
rect 46020 2320 46072 2329
rect 46112 2320 46164 2372
rect 47768 2320 47820 2372
rect 48504 2320 48556 2372
rect 49884 2320 49936 2372
rect 51264 2320 51316 2372
rect 55588 2363 55640 2372
rect 55588 2329 55597 2363
rect 55597 2329 55631 2363
rect 55631 2329 55640 2363
rect 55588 2320 55640 2329
rect 58992 2388 59044 2440
rect 57336 2320 57388 2372
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 50294 2150 50346 2202
rect 50358 2150 50410 2202
rect 50422 2150 50474 2202
rect 50486 2150 50538 2202
rect 50550 2150 50602 2202
rect 18604 2048 18656 2100
rect 22376 2048 22428 2100
rect 48136 2048 48188 2100
rect 56048 2048 56100 2100
rect 18236 1980 18288 2032
rect 20628 1980 20680 2032
rect 23572 1980 23624 2032
rect 44640 1980 44692 2032
rect 15844 1912 15896 1964
rect 30564 1912 30616 1964
rect 22652 1776 22704 1828
rect 39488 1776 39540 1828
rect 22836 1504 22888 1556
rect 24400 1504 24452 1556
rect 36268 1232 36320 1284
rect 39672 1232 39724 1284
rect 50344 1232 50396 1284
rect 54392 1232 54444 1284
rect 34336 1164 34388 1216
rect 36176 1164 36228 1216
rect 36820 1164 36872 1216
rect 38752 1164 38804 1216
rect 39028 1164 39080 1216
rect 43352 1164 43404 1216
rect 47032 1164 47084 1216
rect 51540 1164 51592 1216
rect 53656 1164 53708 1216
rect 56968 1164 57020 1216
rect 7932 1096 7984 1148
rect 9220 1096 9272 1148
rect 35716 1096 35768 1148
rect 38660 1096 38712 1148
rect 39856 1096 39908 1148
rect 44088 1096 44140 1148
rect 47584 1096 47636 1148
rect 49976 1096 50028 1148
rect 52552 1096 52604 1148
rect 55956 1096 56008 1148
rect 8392 1028 8444 1080
rect 10876 1028 10928 1080
rect 13268 1028 13320 1080
rect 13912 1028 13964 1080
rect 17868 1028 17920 1080
rect 19984 1028 20036 1080
rect 20536 1028 20588 1080
rect 22192 1028 22244 1080
rect 34888 1028 34940 1080
rect 37740 1028 37792 1080
rect 39304 1028 39356 1080
rect 43260 1028 43312 1080
rect 43720 1028 43772 1080
rect 46296 1028 46348 1080
rect 47308 1028 47360 1080
rect 51264 1028 51316 1080
rect 51724 1028 51776 1080
rect 55220 1028 55272 1080
rect 6828 960 6880 1012
rect 7840 960 7892 1012
rect 9036 960 9088 1012
rect 10600 960 10652 1012
rect 10968 960 11020 1012
rect 12256 960 12308 1012
rect 13544 960 13596 1012
rect 14740 960 14792 1012
rect 17408 960 17460 1012
rect 18880 960 18932 1012
rect 20444 960 20496 1012
rect 20812 960 20864 1012
rect 21180 960 21232 1012
rect 22744 960 22796 1012
rect 23756 960 23808 1012
rect 25228 960 25280 1012
rect 31852 960 31904 1012
rect 33140 960 33192 1012
rect 33784 960 33836 1012
rect 36084 960 36136 1012
rect 36544 960 36596 1012
rect 40316 960 40368 1012
rect 42340 960 42392 1012
rect 46020 960 46072 1012
rect 48964 960 49016 1012
rect 52644 960 52696 1012
rect 52828 960 52880 1012
rect 57336 960 57388 1012
rect 5816 892 5868 944
rect 7288 892 7340 944
rect 8024 892 8076 944
rect 9496 892 9548 944
rect 10232 892 10284 944
rect 11980 892 12032 944
rect 12072 892 12124 944
rect 13084 892 13136 944
rect 13728 892 13780 944
rect 14464 892 14516 944
rect 17040 892 17092 944
rect 18604 892 18656 944
rect 18696 892 18748 944
rect 20536 892 20588 944
rect 20628 892 20680 944
rect 21640 892 21692 944
rect 24768 892 24820 944
rect 25504 892 25556 944
rect 27528 892 27580 944
rect 27988 892 28040 944
rect 31300 892 31352 944
rect 32588 892 32640 944
rect 32956 892 33008 944
rect 34520 892 34572 944
rect 35440 892 35492 944
rect 37280 892 37332 944
rect 37648 892 37700 944
rect 23204 824 23256 876
rect 23756 824 23808 876
rect 38752 892 38804 944
rect 40684 892 40736 944
rect 44456 892 44508 944
rect 44824 892 44876 944
rect 46112 892 46164 944
rect 47860 892 47912 944
rect 48504 892 48556 944
rect 49240 892 49292 944
rect 49884 892 49936 944
rect 50896 892 50948 944
rect 53012 892 53064 944
rect 53380 892 53432 944
rect 55588 892 55640 944
rect 43812 824 43864 876
rect 48780 824 48832 876
rect 51080 824 51132 876
rect 41420 756 41472 808
rect 46664 756 46716 808
rect 50804 756 50856 808
rect 44088 76 44140 128
rect 49424 76 49476 128
<< metal2 >>
rect 2226 59200 2282 60000
rect 3514 59200 3570 60000
rect 4802 59200 4858 60000
rect 6090 59200 6146 60000
rect 7378 59200 7434 60000
rect 8666 59200 8722 60000
rect 9954 59200 10010 60000
rect 11242 59200 11298 60000
rect 12530 59200 12586 60000
rect 13818 59200 13874 60000
rect 15106 59200 15162 60000
rect 16394 59200 16450 60000
rect 17682 59200 17738 60000
rect 18970 59200 19026 60000
rect 20258 59200 20314 60000
rect 21546 59200 21602 60000
rect 22834 59200 22890 60000
rect 24122 59200 24178 60000
rect 25410 59200 25466 60000
rect 26698 59200 26754 60000
rect 27986 59200 28042 60000
rect 29274 59200 29330 60000
rect 30562 59200 30618 60000
rect 31850 59200 31906 60000
rect 33138 59200 33194 60000
rect 34426 59200 34482 60000
rect 35714 59200 35770 60000
rect 37002 59200 37058 60000
rect 38290 59200 38346 60000
rect 39578 59200 39634 60000
rect 40866 59200 40922 60000
rect 42154 59200 42210 60000
rect 43442 59200 43498 60000
rect 44730 59200 44786 60000
rect 46018 59200 46074 60000
rect 47306 59200 47362 60000
rect 48594 59200 48650 60000
rect 49882 59200 49938 60000
rect 51170 59200 51226 60000
rect 52458 59200 52514 60000
rect 53746 59200 53802 60000
rect 55034 59200 55090 60000
rect 56322 59200 56378 60000
rect 57610 59200 57666 60000
rect 2240 57526 2268 59200
rect 3528 57526 3556 59200
rect 4816 57526 4844 59200
rect 2228 57520 2280 57526
rect 2228 57462 2280 57468
rect 3516 57520 3568 57526
rect 3516 57462 3568 57468
rect 4804 57520 4856 57526
rect 4804 57462 4856 57468
rect 6104 57458 6132 59200
rect 7392 57526 7420 59200
rect 8680 57526 8708 59200
rect 9968 57526 9996 59200
rect 7380 57520 7432 57526
rect 7380 57462 7432 57468
rect 8668 57520 8720 57526
rect 8668 57462 8720 57468
rect 9956 57520 10008 57526
rect 9956 57462 10008 57468
rect 11256 57458 11284 59200
rect 12544 57526 12572 59200
rect 12532 57520 12584 57526
rect 12532 57462 12584 57468
rect 13832 57458 13860 59200
rect 15120 59140 15148 59200
rect 16408 59158 16436 59200
rect 16396 59152 16448 59158
rect 15120 59112 15240 59140
rect 15212 57458 15240 59112
rect 16396 59094 16448 59100
rect 16948 59152 17000 59158
rect 16948 59094 17000 59100
rect 16960 57526 16988 59094
rect 17696 57526 17724 59200
rect 18984 59158 19012 59200
rect 18972 59152 19024 59158
rect 18972 59094 19024 59100
rect 19432 59152 19484 59158
rect 19432 59094 19484 59100
rect 16948 57520 17000 57526
rect 16948 57462 17000 57468
rect 17684 57520 17736 57526
rect 17684 57462 17736 57468
rect 19444 57458 19472 59094
rect 19574 57692 19882 57701
rect 19574 57690 19580 57692
rect 19636 57690 19660 57692
rect 19716 57690 19740 57692
rect 19796 57690 19820 57692
rect 19876 57690 19882 57692
rect 19636 57638 19638 57690
rect 19818 57638 19820 57690
rect 19574 57636 19580 57638
rect 19636 57636 19660 57638
rect 19716 57636 19740 57638
rect 19796 57636 19820 57638
rect 19876 57636 19882 57638
rect 19574 57627 19882 57636
rect 20272 57526 20300 59200
rect 21560 59158 21588 59200
rect 21548 59152 21600 59158
rect 21548 59094 21600 59100
rect 22100 59152 22152 59158
rect 22100 59094 22152 59100
rect 22112 57526 22140 59094
rect 22848 57526 22876 59200
rect 20260 57520 20312 57526
rect 20260 57462 20312 57468
rect 22100 57520 22152 57526
rect 22100 57462 22152 57468
rect 22836 57520 22888 57526
rect 22836 57462 22888 57468
rect 24136 57458 24164 59200
rect 25424 57526 25452 59200
rect 26712 57526 26740 59200
rect 28000 57526 28028 59200
rect 29288 57526 29316 59200
rect 30576 57526 30604 59200
rect 31864 57526 31892 59200
rect 33152 57526 33180 59200
rect 34440 59106 34468 59200
rect 35728 59106 35756 59200
rect 37016 59158 37044 59200
rect 37004 59152 37056 59158
rect 34440 59078 34560 59106
rect 35728 59078 35940 59106
rect 37004 59094 37056 59100
rect 37556 59152 37608 59158
rect 37556 59094 37608 59100
rect 34532 57526 34560 59078
rect 35912 57526 35940 59078
rect 37568 57526 37596 59094
rect 38304 57526 38332 59200
rect 39592 59158 39620 59200
rect 39580 59152 39632 59158
rect 39580 59094 39632 59100
rect 40040 59152 40092 59158
rect 40040 59094 40092 59100
rect 25412 57520 25464 57526
rect 25412 57462 25464 57468
rect 26700 57520 26752 57526
rect 26700 57462 26752 57468
rect 27988 57520 28040 57526
rect 27988 57462 28040 57468
rect 29276 57520 29328 57526
rect 29276 57462 29328 57468
rect 30564 57520 30616 57526
rect 30564 57462 30616 57468
rect 31852 57520 31904 57526
rect 31852 57462 31904 57468
rect 33140 57520 33192 57526
rect 33140 57462 33192 57468
rect 34520 57520 34572 57526
rect 34520 57462 34572 57468
rect 35900 57520 35952 57526
rect 35900 57462 35952 57468
rect 37556 57520 37608 57526
rect 37556 57462 37608 57468
rect 38292 57520 38344 57526
rect 38292 57462 38344 57468
rect 40052 57458 40080 59094
rect 40880 57526 40908 59200
rect 42168 57526 42196 59200
rect 43456 57526 43484 59200
rect 44744 57526 44772 59200
rect 40868 57520 40920 57526
rect 40868 57462 40920 57468
rect 42156 57520 42208 57526
rect 42156 57462 42208 57468
rect 43444 57520 43496 57526
rect 43444 57462 43496 57468
rect 44732 57520 44784 57526
rect 44732 57462 44784 57468
rect 46032 57458 46060 59200
rect 47320 57526 47348 59200
rect 47308 57520 47360 57526
rect 47308 57462 47360 57468
rect 48608 57458 48636 59200
rect 49896 57526 49924 59200
rect 50294 57692 50602 57701
rect 50294 57690 50300 57692
rect 50356 57690 50380 57692
rect 50436 57690 50460 57692
rect 50516 57690 50540 57692
rect 50596 57690 50602 57692
rect 50356 57638 50358 57690
rect 50538 57638 50540 57690
rect 50294 57636 50300 57638
rect 50356 57636 50380 57638
rect 50436 57636 50460 57638
rect 50516 57636 50540 57638
rect 50596 57636 50602 57638
rect 50294 57627 50602 57636
rect 49884 57520 49936 57526
rect 49884 57462 49936 57468
rect 51184 57458 51212 59200
rect 52472 57458 52500 59200
rect 53760 59140 53788 59200
rect 55048 59158 55076 59200
rect 55036 59152 55088 59158
rect 53760 59112 53880 59140
rect 53852 57526 53880 59112
rect 55036 59094 55088 59100
rect 55588 59152 55640 59158
rect 55588 59094 55640 59100
rect 55600 57526 55628 59094
rect 56336 57526 56364 59200
rect 56784 57996 56836 58002
rect 56784 57938 56836 57944
rect 53840 57520 53892 57526
rect 53840 57462 53892 57468
rect 55588 57520 55640 57526
rect 55588 57462 55640 57468
rect 56324 57520 56376 57526
rect 56324 57462 56376 57468
rect 6092 57452 6144 57458
rect 6092 57394 6144 57400
rect 11244 57452 11296 57458
rect 11244 57394 11296 57400
rect 13820 57452 13872 57458
rect 13820 57394 13872 57400
rect 15200 57452 15252 57458
rect 15200 57394 15252 57400
rect 19432 57452 19484 57458
rect 19432 57394 19484 57400
rect 24124 57452 24176 57458
rect 24124 57394 24176 57400
rect 40040 57452 40092 57458
rect 40040 57394 40092 57400
rect 46020 57452 46072 57458
rect 46020 57394 46072 57400
rect 48596 57452 48648 57458
rect 48596 57394 48648 57400
rect 51172 57452 51224 57458
rect 51172 57394 51224 57400
rect 52460 57452 52512 57458
rect 52460 57394 52512 57400
rect 26884 57384 26936 57390
rect 26884 57326 26936 57332
rect 3424 57316 3476 57322
rect 3424 57258 3476 57264
rect 17132 57316 17184 57322
rect 17132 57258 17184 57264
rect 940 56364 992 56370
rect 940 56306 992 56312
rect 952 55865 980 56306
rect 938 55856 994 55865
rect 938 55791 994 55800
rect 940 55752 992 55758
rect 940 55694 992 55700
rect 952 55321 980 55694
rect 938 55312 994 55321
rect 938 55247 994 55256
rect 1032 55276 1084 55282
rect 1032 55218 1084 55224
rect 1044 54777 1072 55218
rect 1952 55072 2004 55078
rect 1952 55014 2004 55020
rect 1030 54768 1086 54777
rect 1030 54703 1086 54712
rect 940 54596 992 54602
rect 940 54538 992 54544
rect 952 54233 980 54538
rect 938 54224 994 54233
rect 938 54159 994 54168
rect 1032 54188 1084 54194
rect 1032 54130 1084 54136
rect 1044 53689 1072 54130
rect 1030 53680 1086 53689
rect 1030 53615 1086 53624
rect 940 53508 992 53514
rect 940 53450 992 53456
rect 952 53145 980 53450
rect 1964 53242 1992 55014
rect 2688 54596 2740 54602
rect 2688 54538 2740 54544
rect 2596 53984 2648 53990
rect 2596 53926 2648 53932
rect 1952 53236 2004 53242
rect 1952 53178 2004 53184
rect 938 53136 994 53145
rect 938 53071 994 53080
rect 1032 53100 1084 53106
rect 1032 53042 1084 53048
rect 1044 52601 1072 53042
rect 1030 52592 1086 52601
rect 1030 52527 1086 52536
rect 940 52420 992 52426
rect 940 52362 992 52368
rect 2044 52420 2096 52426
rect 2044 52362 2096 52368
rect 952 52057 980 52362
rect 938 52048 994 52057
rect 938 51983 994 51992
rect 1032 52012 1084 52018
rect 1032 51954 1084 51960
rect 1044 51513 1072 51954
rect 2056 51950 2084 52362
rect 2044 51944 2096 51950
rect 2044 51886 2096 51892
rect 1030 51504 1086 51513
rect 1030 51439 1086 51448
rect 940 51332 992 51338
rect 940 51274 992 51280
rect 2044 51332 2096 51338
rect 2044 51274 2096 51280
rect 952 50969 980 51274
rect 938 50960 994 50969
rect 938 50895 994 50904
rect 1032 50924 1084 50930
rect 1032 50866 1084 50872
rect 1044 50425 1072 50866
rect 2056 50862 2084 51274
rect 2044 50856 2096 50862
rect 2044 50798 2096 50804
rect 2608 50726 2636 53926
rect 2700 51610 2728 54538
rect 2688 51604 2740 51610
rect 2688 51546 2740 51552
rect 2412 50720 2464 50726
rect 2412 50662 2464 50668
rect 2596 50720 2648 50726
rect 2596 50662 2648 50668
rect 1030 50416 1086 50425
rect 1030 50351 1086 50360
rect 940 50244 992 50250
rect 940 50186 992 50192
rect 952 49881 980 50186
rect 938 49872 994 49881
rect 938 49807 994 49816
rect 1032 49836 1084 49842
rect 1032 49778 1084 49784
rect 1044 49337 1072 49778
rect 1860 49768 1912 49774
rect 1860 49710 1912 49716
rect 1030 49328 1086 49337
rect 1030 49263 1086 49272
rect 940 49156 992 49162
rect 940 49098 992 49104
rect 952 48793 980 49098
rect 938 48784 994 48793
rect 938 48719 994 48728
rect 1032 48748 1084 48754
rect 1032 48690 1084 48696
rect 1044 48249 1072 48690
rect 1030 48240 1086 48249
rect 1030 48175 1086 48184
rect 940 48068 992 48074
rect 940 48010 992 48016
rect 952 47705 980 48010
rect 938 47696 994 47705
rect 938 47631 994 47640
rect 1032 47660 1084 47666
rect 1032 47602 1084 47608
rect 1044 47161 1072 47602
rect 1030 47152 1086 47161
rect 1030 47087 1086 47096
rect 940 46980 992 46986
rect 940 46922 992 46928
rect 952 46617 980 46922
rect 938 46608 994 46617
rect 938 46543 994 46552
rect 1032 46572 1084 46578
rect 1032 46514 1084 46520
rect 1044 46073 1072 46514
rect 1030 46064 1086 46073
rect 1030 45999 1086 46008
rect 940 45960 992 45966
rect 940 45902 992 45908
rect 952 45529 980 45902
rect 1768 45824 1820 45830
rect 1768 45766 1820 45772
rect 938 45520 994 45529
rect 938 45455 994 45464
rect 1032 45484 1084 45490
rect 1032 45426 1084 45432
rect 1044 44985 1072 45426
rect 1780 45422 1808 45766
rect 1768 45416 1820 45422
rect 1768 45358 1820 45364
rect 1030 44976 1086 44985
rect 1030 44911 1086 44920
rect 940 44804 992 44810
rect 940 44746 992 44752
rect 952 44441 980 44746
rect 938 44432 994 44441
rect 938 44367 994 44376
rect 1032 44396 1084 44402
rect 1032 44338 1084 44344
rect 1044 43897 1072 44338
rect 1030 43888 1086 43897
rect 1030 43823 1086 43832
rect 940 43716 992 43722
rect 940 43658 992 43664
rect 952 43353 980 43658
rect 938 43344 994 43353
rect 938 43279 994 43288
rect 1032 43308 1084 43314
rect 1032 43250 1084 43256
rect 1044 42809 1072 43250
rect 1030 42800 1086 42809
rect 1030 42735 1086 42744
rect 940 42628 992 42634
rect 940 42570 992 42576
rect 952 42265 980 42570
rect 938 42256 994 42265
rect 938 42191 994 42200
rect 1032 42220 1084 42226
rect 1032 42162 1084 42168
rect 1044 41721 1072 42162
rect 1030 41712 1086 41721
rect 1030 41647 1086 41656
rect 940 41608 992 41614
rect 940 41550 992 41556
rect 952 41177 980 41550
rect 938 41168 994 41177
rect 938 41103 994 41112
rect 1032 41132 1084 41138
rect 1032 41074 1084 41080
rect 1044 40633 1072 41074
rect 1030 40624 1086 40633
rect 1030 40559 1086 40568
rect 940 40452 992 40458
rect 940 40394 992 40400
rect 952 40089 980 40394
rect 1032 40112 1084 40118
rect 938 40080 994 40089
rect 1032 40054 1084 40060
rect 938 40015 994 40024
rect 1044 39545 1072 40054
rect 1030 39536 1086 39545
rect 1030 39471 1086 39480
rect 940 39364 992 39370
rect 940 39306 992 39312
rect 952 39001 980 39306
rect 938 38992 994 39001
rect 938 38927 994 38936
rect 1032 38956 1084 38962
rect 1032 38898 1084 38904
rect 1044 38457 1072 38898
rect 1030 38448 1086 38457
rect 1030 38383 1086 38392
rect 940 38276 992 38282
rect 940 38218 992 38224
rect 952 37913 980 38218
rect 938 37904 994 37913
rect 938 37839 994 37848
rect 1032 37868 1084 37874
rect 1032 37810 1084 37816
rect 1044 37369 1072 37810
rect 1030 37360 1086 37369
rect 1030 37295 1086 37304
rect 940 37188 992 37194
rect 940 37130 992 37136
rect 952 36825 980 37130
rect 938 36816 994 36825
rect 938 36751 994 36760
rect 1032 36780 1084 36786
rect 1032 36722 1084 36728
rect 1044 36281 1072 36722
rect 1030 36272 1086 36281
rect 1030 36207 1086 36216
rect 940 36168 992 36174
rect 940 36110 992 36116
rect 952 35737 980 36110
rect 938 35728 994 35737
rect 938 35663 994 35672
rect 1032 35692 1084 35698
rect 1032 35634 1084 35640
rect 1044 35193 1072 35634
rect 1768 35284 1820 35290
rect 1768 35226 1820 35232
rect 1030 35184 1086 35193
rect 1030 35119 1086 35128
rect 940 35012 992 35018
rect 940 34954 992 34960
rect 952 34649 980 34954
rect 1780 34746 1808 35226
rect 1768 34740 1820 34746
rect 1768 34682 1820 34688
rect 938 34640 994 34649
rect 938 34575 994 34584
rect 1032 34604 1084 34610
rect 1032 34546 1084 34552
rect 1044 34105 1072 34546
rect 1030 34096 1086 34105
rect 1030 34031 1086 34040
rect 940 33924 992 33930
rect 940 33866 992 33872
rect 952 33561 980 33866
rect 938 33552 994 33561
rect 938 33487 994 33496
rect 1032 33516 1084 33522
rect 1032 33458 1084 33464
rect 1044 33017 1072 33458
rect 1030 33008 1086 33017
rect 1030 32943 1086 32952
rect 940 32836 992 32842
rect 940 32778 992 32784
rect 952 32473 980 32778
rect 938 32464 994 32473
rect 938 32399 994 32408
rect 938 31920 994 31929
rect 938 31855 994 31864
rect 1032 31884 1084 31890
rect 952 31822 980 31855
rect 1032 31826 1084 31832
rect 940 31816 992 31822
rect 940 31758 992 31764
rect 1044 31385 1072 31826
rect 1030 31376 1086 31385
rect 1030 31311 1086 31320
rect 938 30832 994 30841
rect 938 30767 994 30776
rect 952 30734 980 30767
rect 940 30728 992 30734
rect 940 30670 992 30676
rect 1768 30592 1820 30598
rect 1768 30534 1820 30540
rect 1780 30394 1808 30534
rect 1768 30388 1820 30394
rect 1768 30330 1820 30336
rect 940 30320 992 30326
rect 938 30288 940 30297
rect 992 30288 994 30297
rect 938 30223 994 30232
rect 938 29744 994 29753
rect 938 29679 994 29688
rect 952 29646 980 29679
rect 940 29640 992 29646
rect 940 29582 992 29588
rect 1032 29572 1084 29578
rect 1032 29514 1084 29520
rect 1044 29209 1072 29514
rect 1030 29200 1086 29209
rect 1030 29135 1086 29144
rect 938 28656 994 28665
rect 938 28591 994 28600
rect 952 28558 980 28591
rect 940 28552 992 28558
rect 940 28494 992 28500
rect 940 28144 992 28150
rect 938 28112 940 28121
rect 992 28112 994 28121
rect 938 28047 994 28056
rect 938 27568 994 27577
rect 938 27503 994 27512
rect 952 27470 980 27503
rect 940 27464 992 27470
rect 940 27406 992 27412
rect 1872 27062 1900 49710
rect 1952 49088 2004 49094
rect 1952 49030 2004 49036
rect 1964 35630 1992 49030
rect 2228 48680 2280 48686
rect 2228 48622 2280 48628
rect 2136 44804 2188 44810
rect 2136 44746 2188 44752
rect 2044 36644 2096 36650
rect 2044 36586 2096 36592
rect 1952 35624 2004 35630
rect 1952 35566 2004 35572
rect 1952 33108 2004 33114
rect 1952 33050 2004 33056
rect 940 27056 992 27062
rect 938 27024 940 27033
rect 1860 27056 1912 27062
rect 992 27024 994 27033
rect 1860 26998 1912 27004
rect 938 26959 994 26968
rect 1032 26988 1084 26994
rect 1032 26930 1084 26936
rect 1044 26489 1072 26930
rect 1030 26480 1086 26489
rect 1030 26415 1086 26424
rect 1964 26314 1992 33050
rect 2056 31346 2084 36586
rect 2148 32434 2176 44746
rect 2240 32978 2268 48622
rect 2320 43716 2372 43722
rect 2320 43658 2372 43664
rect 2228 32972 2280 32978
rect 2228 32914 2280 32920
rect 2332 32858 2360 43658
rect 2424 33114 2452 50662
rect 3436 36922 3464 57258
rect 3976 57248 4028 57254
rect 3976 57190 4028 57196
rect 4712 57248 4764 57254
rect 4712 57190 4764 57196
rect 6736 57248 6788 57254
rect 6736 57190 6788 57196
rect 7380 57248 7432 57254
rect 7380 57190 7432 57196
rect 9128 57248 9180 57254
rect 9128 57190 9180 57196
rect 9956 57248 10008 57254
rect 9956 57190 10008 57196
rect 11888 57248 11940 57254
rect 11888 57190 11940 57196
rect 12808 57248 12860 57254
rect 12808 57190 12860 57196
rect 15384 57248 15436 57254
rect 15384 57190 15436 57196
rect 3608 38276 3660 38282
rect 3608 38218 3660 38224
rect 3424 36916 3476 36922
rect 3424 36858 3476 36864
rect 3620 36786 3648 38218
rect 3700 37732 3752 37738
rect 3700 37674 3752 37680
rect 3712 36786 3740 37674
rect 3148 36780 3200 36786
rect 3148 36722 3200 36728
rect 3608 36780 3660 36786
rect 3608 36722 3660 36728
rect 3700 36780 3752 36786
rect 3700 36722 3752 36728
rect 3884 36780 3936 36786
rect 3884 36722 3936 36728
rect 2872 35692 2924 35698
rect 2872 35634 2924 35640
rect 2964 35692 3016 35698
rect 2964 35634 3016 35640
rect 2412 33108 2464 33114
rect 2412 33050 2464 33056
rect 2412 32972 2464 32978
rect 2412 32914 2464 32920
rect 2240 32830 2360 32858
rect 2136 32428 2188 32434
rect 2136 32370 2188 32376
rect 2044 31340 2096 31346
rect 2044 31282 2096 31288
rect 2240 29186 2268 32830
rect 2320 32768 2372 32774
rect 2320 32710 2372 32716
rect 2332 32502 2360 32710
rect 2424 32570 2452 32914
rect 2884 32570 2912 35634
rect 2976 33590 3004 35634
rect 2964 33584 3016 33590
rect 2964 33526 3016 33532
rect 2412 32564 2464 32570
rect 2412 32506 2464 32512
rect 2872 32564 2924 32570
rect 2872 32506 2924 32512
rect 2320 32496 2372 32502
rect 2320 32438 2372 32444
rect 2320 31340 2372 31346
rect 2320 31282 2372 31288
rect 2332 29782 2360 31282
rect 2320 29776 2372 29782
rect 2320 29718 2372 29724
rect 2320 29504 2372 29510
rect 2320 29446 2372 29452
rect 2332 29238 2360 29446
rect 2424 29306 2452 32506
rect 2504 32428 2556 32434
rect 2504 32370 2556 32376
rect 2412 29300 2464 29306
rect 2412 29242 2464 29248
rect 2148 29170 2268 29186
rect 2320 29232 2372 29238
rect 2320 29174 2372 29180
rect 2136 29164 2268 29170
rect 2188 29158 2268 29164
rect 2136 29106 2188 29112
rect 2136 29028 2188 29034
rect 2136 28970 2188 28976
rect 940 26308 992 26314
rect 940 26250 992 26256
rect 1952 26308 2004 26314
rect 1952 26250 2004 26256
rect 952 25945 980 26250
rect 938 25936 994 25945
rect 938 25871 994 25880
rect 1584 25900 1636 25906
rect 1584 25842 1636 25848
rect 940 25832 992 25838
rect 940 25774 992 25780
rect 952 25401 980 25774
rect 1596 25498 1624 25842
rect 1584 25492 1636 25498
rect 1584 25434 1636 25440
rect 938 25392 994 25401
rect 938 25327 994 25336
rect 940 25220 992 25226
rect 940 25162 992 25168
rect 952 24857 980 25162
rect 938 24848 994 24857
rect 938 24783 994 24792
rect 1584 24812 1636 24818
rect 1584 24754 1636 24760
rect 940 24744 992 24750
rect 940 24686 992 24692
rect 952 24313 980 24686
rect 1596 24410 1624 24754
rect 2148 24750 2176 28970
rect 2424 26234 2452 29242
rect 2516 29050 2544 32370
rect 2596 32224 2648 32230
rect 2596 32166 2648 32172
rect 2608 30258 2636 32166
rect 2688 31340 2740 31346
rect 2688 31282 2740 31288
rect 2700 30258 2728 31282
rect 2596 30252 2648 30258
rect 2596 30194 2648 30200
rect 2688 30252 2740 30258
rect 2688 30194 2740 30200
rect 2700 29170 2728 30194
rect 2688 29164 2740 29170
rect 2688 29106 2740 29112
rect 2516 29022 2728 29050
rect 2424 26206 2636 26234
rect 2504 25288 2556 25294
rect 2504 25230 2556 25236
rect 2516 24970 2544 25230
rect 2424 24954 2544 24970
rect 2424 24948 2556 24954
rect 2424 24942 2504 24948
rect 2424 24818 2452 24942
rect 2504 24890 2556 24896
rect 2412 24812 2464 24818
rect 2412 24754 2464 24760
rect 2136 24744 2188 24750
rect 2136 24686 2188 24692
rect 1584 24404 1636 24410
rect 1584 24346 1636 24352
rect 938 24304 994 24313
rect 938 24239 994 24248
rect 2424 24206 2452 24754
rect 2412 24200 2464 24206
rect 2412 24142 2464 24148
rect 940 24132 992 24138
rect 940 24074 992 24080
rect 952 23769 980 24074
rect 938 23760 994 23769
rect 938 23695 994 23704
rect 940 23656 992 23662
rect 940 23598 992 23604
rect 952 23225 980 23598
rect 938 23216 994 23225
rect 2424 23186 2452 24142
rect 938 23151 994 23160
rect 2412 23180 2464 23186
rect 2412 23122 2464 23128
rect 940 23044 992 23050
rect 940 22986 992 22992
rect 952 22681 980 22986
rect 2424 22778 2452 23122
rect 2412 22772 2464 22778
rect 2412 22714 2464 22720
rect 938 22672 994 22681
rect 2424 22658 2452 22714
rect 2424 22630 2544 22658
rect 938 22607 994 22616
rect 938 22128 994 22137
rect 938 22063 940 22072
rect 992 22063 994 22072
rect 940 22034 992 22040
rect 2516 22030 2544 22630
rect 2608 22030 2636 26206
rect 2700 24206 2728 29022
rect 3160 25294 3188 36722
rect 3424 36032 3476 36038
rect 3424 35974 3476 35980
rect 3436 35894 3464 35974
rect 3436 35866 3556 35894
rect 3424 32768 3476 32774
rect 3424 32710 3476 32716
rect 3240 32564 3292 32570
rect 3240 32506 3292 32512
rect 3252 29102 3280 32506
rect 3436 32434 3464 32710
rect 3332 32428 3384 32434
rect 3332 32370 3384 32376
rect 3424 32428 3476 32434
rect 3424 32370 3476 32376
rect 3344 31482 3372 32370
rect 3332 31476 3384 31482
rect 3332 31418 3384 31424
rect 3240 29096 3292 29102
rect 3240 29038 3292 29044
rect 3252 26234 3280 29038
rect 3252 26206 3464 26234
rect 3148 25288 3200 25294
rect 3148 25230 3200 25236
rect 2964 24676 3016 24682
rect 2964 24618 3016 24624
rect 2688 24200 2740 24206
rect 2688 24142 2740 24148
rect 2872 23724 2924 23730
rect 2872 23666 2924 23672
rect 2884 23254 2912 23666
rect 2872 23248 2924 23254
rect 2872 23190 2924 23196
rect 2780 23044 2832 23050
rect 2780 22986 2832 22992
rect 2792 22234 2820 22986
rect 2780 22228 2832 22234
rect 2780 22170 2832 22176
rect 2504 22024 2556 22030
rect 2504 21966 2556 21972
rect 2596 22024 2648 22030
rect 2596 21966 2648 21972
rect 938 21584 994 21593
rect 938 21519 994 21528
rect 952 21486 980 21519
rect 940 21480 992 21486
rect 940 21422 992 21428
rect 938 21040 994 21049
rect 938 20975 940 20984
rect 992 20975 994 20984
rect 940 20946 992 20952
rect 938 20496 994 20505
rect 2976 20466 3004 24618
rect 3436 23118 3464 26206
rect 3424 23112 3476 23118
rect 3424 23054 3476 23060
rect 938 20431 994 20440
rect 2964 20460 3016 20466
rect 952 20398 980 20431
rect 2964 20402 3016 20408
rect 940 20392 992 20398
rect 940 20334 992 20340
rect 938 19952 994 19961
rect 938 19887 940 19896
rect 992 19887 994 19896
rect 940 19858 992 19864
rect 940 19712 992 19718
rect 940 19654 992 19660
rect 952 19417 980 19654
rect 1032 19440 1084 19446
rect 938 19408 994 19417
rect 1032 19382 1084 19388
rect 938 19343 994 19352
rect 1044 18873 1072 19382
rect 1030 18864 1086 18873
rect 1030 18799 1086 18808
rect 940 18692 992 18698
rect 940 18634 992 18640
rect 952 18329 980 18634
rect 938 18320 994 18329
rect 938 18255 994 18264
rect 940 18216 992 18222
rect 940 18158 992 18164
rect 952 17785 980 18158
rect 938 17776 994 17785
rect 938 17711 994 17720
rect 940 17604 992 17610
rect 940 17546 992 17552
rect 952 17241 980 17546
rect 3528 17270 3556 35866
rect 3896 35834 3924 36722
rect 3884 35828 3936 35834
rect 3884 35770 3936 35776
rect 3988 33998 4016 57190
rect 4214 57148 4522 57157
rect 4214 57146 4220 57148
rect 4276 57146 4300 57148
rect 4356 57146 4380 57148
rect 4436 57146 4460 57148
rect 4516 57146 4522 57148
rect 4276 57094 4278 57146
rect 4458 57094 4460 57146
rect 4214 57092 4220 57094
rect 4276 57092 4300 57094
rect 4356 57092 4380 57094
rect 4436 57092 4460 57094
rect 4516 57092 4522 57094
rect 4214 57083 4522 57092
rect 4214 56060 4522 56069
rect 4214 56058 4220 56060
rect 4276 56058 4300 56060
rect 4356 56058 4380 56060
rect 4436 56058 4460 56060
rect 4516 56058 4522 56060
rect 4276 56006 4278 56058
rect 4458 56006 4460 56058
rect 4214 56004 4220 56006
rect 4276 56004 4300 56006
rect 4356 56004 4380 56006
rect 4436 56004 4460 56006
rect 4516 56004 4522 56006
rect 4214 55995 4522 56004
rect 4214 54972 4522 54981
rect 4214 54970 4220 54972
rect 4276 54970 4300 54972
rect 4356 54970 4380 54972
rect 4436 54970 4460 54972
rect 4516 54970 4522 54972
rect 4276 54918 4278 54970
rect 4458 54918 4460 54970
rect 4214 54916 4220 54918
rect 4276 54916 4300 54918
rect 4356 54916 4380 54918
rect 4436 54916 4460 54918
rect 4516 54916 4522 54918
rect 4214 54907 4522 54916
rect 4214 53884 4522 53893
rect 4214 53882 4220 53884
rect 4276 53882 4300 53884
rect 4356 53882 4380 53884
rect 4436 53882 4460 53884
rect 4516 53882 4522 53884
rect 4276 53830 4278 53882
rect 4458 53830 4460 53882
rect 4214 53828 4220 53830
rect 4276 53828 4300 53830
rect 4356 53828 4380 53830
rect 4436 53828 4460 53830
rect 4516 53828 4522 53830
rect 4214 53819 4522 53828
rect 4214 52796 4522 52805
rect 4214 52794 4220 52796
rect 4276 52794 4300 52796
rect 4356 52794 4380 52796
rect 4436 52794 4460 52796
rect 4516 52794 4522 52796
rect 4276 52742 4278 52794
rect 4458 52742 4460 52794
rect 4214 52740 4220 52742
rect 4276 52740 4300 52742
rect 4356 52740 4380 52742
rect 4436 52740 4460 52742
rect 4516 52740 4522 52742
rect 4214 52731 4522 52740
rect 4214 51708 4522 51717
rect 4214 51706 4220 51708
rect 4276 51706 4300 51708
rect 4356 51706 4380 51708
rect 4436 51706 4460 51708
rect 4516 51706 4522 51708
rect 4276 51654 4278 51706
rect 4458 51654 4460 51706
rect 4214 51652 4220 51654
rect 4276 51652 4300 51654
rect 4356 51652 4380 51654
rect 4436 51652 4460 51654
rect 4516 51652 4522 51654
rect 4214 51643 4522 51652
rect 4214 50620 4522 50629
rect 4214 50618 4220 50620
rect 4276 50618 4300 50620
rect 4356 50618 4380 50620
rect 4436 50618 4460 50620
rect 4516 50618 4522 50620
rect 4276 50566 4278 50618
rect 4458 50566 4460 50618
rect 4214 50564 4220 50566
rect 4276 50564 4300 50566
rect 4356 50564 4380 50566
rect 4436 50564 4460 50566
rect 4516 50564 4522 50566
rect 4214 50555 4522 50564
rect 4214 49532 4522 49541
rect 4214 49530 4220 49532
rect 4276 49530 4300 49532
rect 4356 49530 4380 49532
rect 4436 49530 4460 49532
rect 4516 49530 4522 49532
rect 4276 49478 4278 49530
rect 4458 49478 4460 49530
rect 4214 49476 4220 49478
rect 4276 49476 4300 49478
rect 4356 49476 4380 49478
rect 4436 49476 4460 49478
rect 4516 49476 4522 49478
rect 4214 49467 4522 49476
rect 4214 48444 4522 48453
rect 4214 48442 4220 48444
rect 4276 48442 4300 48444
rect 4356 48442 4380 48444
rect 4436 48442 4460 48444
rect 4516 48442 4522 48444
rect 4276 48390 4278 48442
rect 4458 48390 4460 48442
rect 4214 48388 4220 48390
rect 4276 48388 4300 48390
rect 4356 48388 4380 48390
rect 4436 48388 4460 48390
rect 4516 48388 4522 48390
rect 4214 48379 4522 48388
rect 4214 47356 4522 47365
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47291 4522 47300
rect 4214 46268 4522 46277
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46203 4522 46212
rect 4214 45180 4522 45189
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45115 4522 45124
rect 4214 44092 4522 44101
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44027 4522 44036
rect 4214 43004 4522 43013
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42939 4522 42948
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 4724 38350 4752 57190
rect 6748 45082 6776 57190
rect 7196 45280 7248 45286
rect 7196 45222 7248 45228
rect 6736 45076 6788 45082
rect 6736 45018 6788 45024
rect 4896 39364 4948 39370
rect 4896 39306 4948 39312
rect 4908 38350 4936 39306
rect 4988 38820 5040 38826
rect 4988 38762 5040 38768
rect 5000 38350 5028 38762
rect 5264 38480 5316 38486
rect 5264 38422 5316 38428
rect 4712 38344 4764 38350
rect 4712 38286 4764 38292
rect 4896 38344 4948 38350
rect 4896 38286 4948 38292
rect 4988 38344 5040 38350
rect 4988 38286 5040 38292
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 4908 36718 4936 38286
rect 4620 36712 4672 36718
rect 4620 36654 4672 36660
rect 4896 36712 4948 36718
rect 4896 36654 4948 36660
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4068 35692 4120 35698
rect 4068 35634 4120 35640
rect 4080 34134 4108 35634
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4068 34128 4120 34134
rect 4068 34070 4120 34076
rect 3976 33992 4028 33998
rect 3976 33934 4028 33940
rect 4080 32434 4108 34070
rect 4632 33930 4660 36654
rect 5276 34678 5304 38422
rect 7208 37942 7236 45222
rect 7392 39438 7420 57190
rect 9140 40526 9168 57190
rect 9968 48754 9996 57190
rect 11704 52896 11756 52902
rect 11704 52838 11756 52844
rect 9956 48748 10008 48754
rect 9956 48690 10008 48696
rect 10140 48748 10192 48754
rect 10140 48690 10192 48696
rect 9220 40928 9272 40934
rect 9220 40870 9272 40876
rect 9128 40520 9180 40526
rect 9128 40462 9180 40468
rect 7656 39840 7708 39846
rect 7656 39782 7708 39788
rect 7668 39438 7696 39782
rect 7932 39568 7984 39574
rect 7932 39510 7984 39516
rect 7380 39432 7432 39438
rect 7380 39374 7432 39380
rect 7656 39432 7708 39438
rect 7656 39374 7708 39380
rect 7840 39432 7892 39438
rect 7840 39374 7892 39380
rect 7852 38554 7880 39374
rect 7840 38548 7892 38554
rect 7840 38490 7892 38496
rect 7852 38350 7880 38490
rect 7840 38344 7892 38350
rect 7840 38286 7892 38292
rect 7196 37936 7248 37942
rect 7196 37878 7248 37884
rect 5264 34672 5316 34678
rect 5264 34614 5316 34620
rect 4620 33924 4672 33930
rect 4620 33866 4672 33872
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 3700 32428 3752 32434
rect 3700 32370 3752 32376
rect 4068 32428 4120 32434
rect 4068 32370 4120 32376
rect 3712 31958 3740 32370
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 3700 31952 3752 31958
rect 3700 31894 3752 31900
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 7944 29782 7972 39510
rect 9232 39438 9260 40870
rect 9588 40520 9640 40526
rect 9588 40462 9640 40468
rect 9312 40452 9364 40458
rect 9312 40394 9364 40400
rect 9220 39432 9272 39438
rect 9220 39374 9272 39380
rect 9324 39370 9352 40394
rect 9312 39364 9364 39370
rect 9312 39306 9364 39312
rect 9600 38554 9628 40462
rect 10152 40458 10180 48690
rect 10508 48544 10560 48550
rect 10508 48486 10560 48492
rect 10520 48210 10548 48486
rect 10508 48204 10560 48210
rect 10508 48146 10560 48152
rect 11716 43450 11744 52838
rect 11900 52494 11928 57190
rect 11888 52488 11940 52494
rect 11888 52430 11940 52436
rect 11704 43444 11756 43450
rect 11704 43386 11756 43392
rect 11704 43104 11756 43110
rect 11704 43046 11756 43052
rect 10140 40452 10192 40458
rect 10140 40394 10192 40400
rect 9588 38548 9640 38554
rect 9588 38490 9640 38496
rect 10152 34746 10180 40394
rect 11716 39370 11744 43046
rect 11704 39364 11756 39370
rect 11704 39306 11756 39312
rect 11428 38548 11480 38554
rect 11428 38490 11480 38496
rect 11440 36718 11468 38490
rect 11428 36712 11480 36718
rect 11428 36654 11480 36660
rect 10140 34740 10192 34746
rect 10140 34682 10192 34688
rect 7932 29776 7984 29782
rect 7932 29718 7984 29724
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 10508 22636 10560 22642
rect 10508 22578 10560 22584
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 10520 22030 10548 22578
rect 10140 22024 10192 22030
rect 10140 21966 10192 21972
rect 10508 22024 10560 22030
rect 10508 21966 10560 21972
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 3516 17264 3568 17270
rect 938 17232 994 17241
rect 3516 17206 3568 17212
rect 938 17167 994 17176
rect 940 17128 992 17134
rect 940 17070 992 17076
rect 952 16697 980 17070
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 938 16688 994 16697
rect 938 16623 994 16632
rect 1584 16584 1636 16590
rect 1584 16526 1636 16532
rect 940 16516 992 16522
rect 940 16458 992 16464
rect 952 16153 980 16458
rect 938 16144 994 16153
rect 938 16079 994 16088
rect 940 16040 992 16046
rect 940 15982 992 15988
rect 952 15609 980 15982
rect 938 15600 994 15609
rect 938 15535 994 15544
rect 940 15428 992 15434
rect 940 15370 992 15376
rect 952 15065 980 15370
rect 938 15056 994 15065
rect 938 14991 994 15000
rect 940 14952 992 14958
rect 940 14894 992 14900
rect 952 14521 980 14894
rect 938 14512 994 14521
rect 938 14447 994 14456
rect 940 14340 992 14346
rect 940 14282 992 14288
rect 952 13977 980 14282
rect 938 13968 994 13977
rect 938 13903 994 13912
rect 940 13864 992 13870
rect 940 13806 992 13812
rect 952 13433 980 13806
rect 938 13424 994 13433
rect 938 13359 994 13368
rect 940 13252 992 13258
rect 940 13194 992 13200
rect 952 12889 980 13194
rect 938 12880 994 12889
rect 938 12815 994 12824
rect 940 12776 992 12782
rect 940 12718 992 12724
rect 952 12345 980 12718
rect 938 12336 994 12345
rect 938 12271 994 12280
rect 940 12164 992 12170
rect 940 12106 992 12112
rect 952 11801 980 12106
rect 1596 11898 1624 16526
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 2688 15496 2740 15502
rect 2688 15438 2740 15444
rect 1584 11892 1636 11898
rect 1584 11834 1636 11840
rect 938 11792 994 11801
rect 938 11727 994 11736
rect 940 11688 992 11694
rect 940 11630 992 11636
rect 952 11257 980 11630
rect 938 11248 994 11257
rect 938 11183 994 11192
rect 940 11076 992 11082
rect 940 11018 992 11024
rect 952 10713 980 11018
rect 2700 10742 2728 15438
rect 5448 15088 5500 15094
rect 5448 15030 5500 15036
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 5460 14414 5488 15030
rect 5448 14408 5500 14414
rect 5448 14350 5500 14356
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4252 13320 4304 13326
rect 4252 13262 4304 13268
rect 8484 13320 8536 13326
rect 8484 13262 8536 13268
rect 4264 12918 4292 13262
rect 4252 12912 4304 12918
rect 4252 12854 4304 12860
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 2688 10736 2740 10742
rect 938 10704 994 10713
rect 2688 10678 2740 10684
rect 938 10639 994 10648
rect 940 10600 992 10606
rect 940 10542 992 10548
rect 952 10169 980 10542
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 938 10160 994 10169
rect 938 10095 994 10104
rect 940 9988 992 9994
rect 940 9930 992 9936
rect 952 9625 980 9930
rect 938 9616 994 9625
rect 938 9551 994 9560
rect 940 9512 992 9518
rect 940 9454 992 9460
rect 952 9081 980 9454
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 938 9072 994 9081
rect 938 9007 994 9016
rect 940 8900 992 8906
rect 940 8842 992 8848
rect 952 8537 980 8842
rect 938 8528 994 8537
rect 938 8463 994 8472
rect 940 8424 992 8430
rect 940 8366 992 8372
rect 952 7993 980 8366
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 938 7984 994 7993
rect 938 7919 994 7928
rect 940 7812 992 7818
rect 940 7754 992 7760
rect 952 7449 980 7754
rect 938 7440 994 7449
rect 938 7375 994 7384
rect 940 7336 992 7342
rect 940 7278 992 7284
rect 952 6905 980 7278
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 938 6896 994 6905
rect 938 6831 994 6840
rect 940 6724 992 6730
rect 940 6666 992 6672
rect 952 6361 980 6666
rect 938 6352 994 6361
rect 938 6287 994 6296
rect 940 6248 992 6254
rect 940 6190 992 6196
rect 952 5817 980 6190
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 8392 5840 8444 5846
rect 938 5808 994 5817
rect 8392 5782 8444 5788
rect 938 5743 994 5752
rect 4620 5704 4672 5710
rect 4620 5646 4672 5652
rect 940 5636 992 5642
rect 940 5578 992 5584
rect 952 5273 980 5578
rect 938 5264 994 5273
rect 938 5199 994 5208
rect 940 5160 992 5166
rect 940 5102 992 5108
rect 952 4729 980 5102
rect 1584 5092 1636 5098
rect 1584 5034 1636 5040
rect 938 4720 994 4729
rect 938 4655 994 4664
rect 1596 4622 1624 5034
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 1584 4616 1636 4622
rect 1584 4558 1636 4564
rect 940 4548 992 4554
rect 940 4490 992 4496
rect 952 4185 980 4490
rect 938 4176 994 4185
rect 938 4111 994 4120
rect 4632 4010 4660 5646
rect 8116 4140 8168 4146
rect 8116 4082 8168 4088
rect 4620 4004 4672 4010
rect 4620 3946 4672 3952
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 7656 3596 7708 3602
rect 7656 3538 7708 3544
rect 7564 3460 7616 3466
rect 7564 3402 7616 3408
rect 5908 3052 5960 3058
rect 5908 2994 5960 3000
rect 6828 3052 6880 3058
rect 6828 2994 6880 3000
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 5816 2372 5868 2378
rect 5816 2314 5868 2320
rect 5828 950 5856 2314
rect 5816 944 5868 950
rect 5816 886 5868 892
rect 5920 800 5948 2994
rect 6840 1018 6868 2994
rect 6828 1012 6880 1018
rect 6828 954 6880 960
rect 7288 944 7340 950
rect 7288 886 7340 892
rect 7300 800 7328 886
rect 7576 800 7604 3402
rect 7668 3194 7696 3538
rect 7656 3188 7708 3194
rect 7656 3130 7708 3136
rect 7932 3052 7984 3058
rect 7932 2994 7984 3000
rect 7944 1154 7972 2994
rect 8024 2372 8076 2378
rect 8024 2314 8076 2320
rect 7932 1148 7984 1154
rect 7932 1090 7984 1096
rect 7840 1012 7892 1018
rect 7840 954 7892 960
rect 7852 800 7880 954
rect 8036 950 8064 2314
rect 8024 944 8076 950
rect 8024 886 8076 892
rect 8128 800 8156 4082
rect 8208 3460 8260 3466
rect 8208 3402 8260 3408
rect 8220 898 8248 3402
rect 8300 2916 8352 2922
rect 8300 2858 8352 2864
rect 8312 2582 8340 2858
rect 8404 2650 8432 5782
rect 8496 3738 8524 13262
rect 8760 8016 8812 8022
rect 8760 7958 8812 7964
rect 8484 3732 8536 3738
rect 8484 3674 8536 3680
rect 8668 3460 8720 3466
rect 8668 3402 8720 3408
rect 8392 2644 8444 2650
rect 8392 2586 8444 2592
rect 8300 2576 8352 2582
rect 8300 2518 8352 2524
rect 8392 2372 8444 2378
rect 8392 2314 8444 2320
rect 8404 1086 8432 2314
rect 8392 1080 8444 1086
rect 8392 1022 8444 1028
rect 8220 870 8432 898
rect 8404 800 8432 870
rect 8680 800 8708 3402
rect 8772 2582 8800 7958
rect 9128 7268 9180 7274
rect 9128 7210 9180 7216
rect 8944 4208 8996 4214
rect 8944 4150 8996 4156
rect 8760 2576 8812 2582
rect 8760 2518 8812 2524
rect 8956 800 8984 4150
rect 9140 3058 9168 7210
rect 9494 5808 9550 5817
rect 10152 5778 10180 21966
rect 11336 16176 11388 16182
rect 11336 16118 11388 16124
rect 11348 15502 11376 16118
rect 11440 15570 11468 36654
rect 11796 32428 11848 32434
rect 11796 32370 11848 32376
rect 11808 29578 11836 32370
rect 11796 29572 11848 29578
rect 11796 29514 11848 29520
rect 11704 21548 11756 21554
rect 11704 21490 11756 21496
rect 11716 19310 11744 21490
rect 11704 19304 11756 19310
rect 11704 19246 11756 19252
rect 11704 17264 11756 17270
rect 11704 17206 11756 17212
rect 11428 15564 11480 15570
rect 11428 15506 11480 15512
rect 11716 15502 11744 17206
rect 11808 15570 11836 29514
rect 12820 24342 12848 57190
rect 14464 47456 14516 47462
rect 14464 47398 14516 47404
rect 14476 42090 14504 47398
rect 14464 42084 14516 42090
rect 14464 42026 14516 42032
rect 13820 30252 13872 30258
rect 13820 30194 13872 30200
rect 13832 28422 13860 30194
rect 13912 29504 13964 29510
rect 13912 29446 13964 29452
rect 15016 29504 15068 29510
rect 15016 29446 15068 29452
rect 13924 29102 13952 29446
rect 13912 29096 13964 29102
rect 13912 29038 13964 29044
rect 13820 28416 13872 28422
rect 13820 28358 13872 28364
rect 12808 24336 12860 24342
rect 12808 24278 12860 24284
rect 12256 18760 12308 18766
rect 12256 18702 12308 18708
rect 11796 15564 11848 15570
rect 11796 15506 11848 15512
rect 11336 15496 11388 15502
rect 11336 15438 11388 15444
rect 11704 15496 11756 15502
rect 11704 15438 11756 15444
rect 10508 15428 10560 15434
rect 10508 15370 10560 15376
rect 10416 6792 10468 6798
rect 10416 6734 10468 6740
rect 10428 6458 10456 6734
rect 10416 6452 10468 6458
rect 10416 6394 10468 6400
rect 10520 6254 10548 15370
rect 11348 8634 11376 15438
rect 12268 15366 12296 18702
rect 12348 17196 12400 17202
rect 12348 17138 12400 17144
rect 12256 15360 12308 15366
rect 12256 15302 12308 15308
rect 12360 15162 12388 17138
rect 14924 16992 14976 16998
rect 14924 16934 14976 16940
rect 14556 16108 14608 16114
rect 14556 16050 14608 16056
rect 14568 15706 14596 16050
rect 14556 15700 14608 15706
rect 14556 15642 14608 15648
rect 12348 15156 12400 15162
rect 12348 15098 12400 15104
rect 12440 15020 12492 15026
rect 12440 14962 12492 14968
rect 12452 13297 12480 14962
rect 13360 14544 13412 14550
rect 13360 14486 13412 14492
rect 12532 14340 12584 14346
rect 12532 14282 12584 14288
rect 12438 13288 12494 13297
rect 12438 13223 12494 13232
rect 12348 12844 12400 12850
rect 12348 12786 12400 12792
rect 12360 12442 12388 12786
rect 12348 12436 12400 12442
rect 12348 12378 12400 12384
rect 11704 11892 11756 11898
rect 11704 11834 11756 11840
rect 11152 8628 11204 8634
rect 11152 8570 11204 8576
rect 11336 8628 11388 8634
rect 11336 8570 11388 8576
rect 10968 8424 11020 8430
rect 10968 8366 11020 8372
rect 11060 8424 11112 8430
rect 11060 8366 11112 8372
rect 10876 8356 10928 8362
rect 10876 8298 10928 8304
rect 10600 8016 10652 8022
rect 10600 7958 10652 7964
rect 10508 6248 10560 6254
rect 10508 6190 10560 6196
rect 9494 5743 9550 5752
rect 10140 5772 10192 5778
rect 9508 5710 9536 5743
rect 10140 5714 10192 5720
rect 9404 5704 9456 5710
rect 9404 5646 9456 5652
rect 9496 5704 9548 5710
rect 9496 5646 9548 5652
rect 9416 3670 9444 5646
rect 10140 5636 10192 5642
rect 10140 5578 10192 5584
rect 9588 5228 9640 5234
rect 9588 5170 9640 5176
rect 9600 3738 9628 5170
rect 10152 4146 10180 5578
rect 10324 4548 10376 4554
rect 10324 4490 10376 4496
rect 10140 4140 10192 4146
rect 10140 4082 10192 4088
rect 9680 4072 9732 4078
rect 10048 4072 10100 4078
rect 9680 4014 9732 4020
rect 10046 4040 10048 4049
rect 10100 4040 10102 4049
rect 9588 3732 9640 3738
rect 9588 3674 9640 3680
rect 9404 3664 9456 3670
rect 9404 3606 9456 3612
rect 9692 3602 9720 4014
rect 10046 3975 10102 3984
rect 10152 3890 10180 4082
rect 10232 4072 10284 4078
rect 10232 4014 10284 4020
rect 10060 3862 10180 3890
rect 9772 3732 9824 3738
rect 9772 3674 9824 3680
rect 9680 3596 9732 3602
rect 9680 3538 9732 3544
rect 9784 3534 9812 3674
rect 10060 3602 10088 3862
rect 10048 3596 10100 3602
rect 10048 3538 10100 3544
rect 9772 3528 9824 3534
rect 9772 3470 9824 3476
rect 10060 3398 10088 3538
rect 10048 3392 10100 3398
rect 10048 3334 10100 3340
rect 10060 3126 10088 3334
rect 9588 3120 9640 3126
rect 9588 3062 9640 3068
rect 10048 3120 10100 3126
rect 10048 3062 10100 3068
rect 9036 3052 9088 3058
rect 9036 2994 9088 3000
rect 9128 3052 9180 3058
rect 9128 2994 9180 3000
rect 9048 1018 9076 2994
rect 9220 1148 9272 1154
rect 9220 1090 9272 1096
rect 9036 1012 9088 1018
rect 9036 954 9088 960
rect 9232 800 9260 1090
rect 9496 944 9548 950
rect 9496 886 9548 892
rect 9600 898 9628 3062
rect 10244 2990 10272 4014
rect 10232 2984 10284 2990
rect 10232 2926 10284 2932
rect 10048 2372 10100 2378
rect 10048 2314 10100 2320
rect 10232 2372 10284 2378
rect 10232 2314 10284 2320
rect 9508 800 9536 886
rect 9600 870 9812 898
rect 9784 800 9812 870
rect 10060 800 10088 2314
rect 10244 950 10272 2314
rect 10232 944 10284 950
rect 10232 886 10284 892
rect 10336 800 10364 4490
rect 10612 2582 10640 7958
rect 10888 6914 10916 8298
rect 10980 7818 11008 8366
rect 11072 8090 11100 8366
rect 11060 8084 11112 8090
rect 11060 8026 11112 8032
rect 11164 7954 11192 8570
rect 11152 7948 11204 7954
rect 11152 7890 11204 7896
rect 11244 7948 11296 7954
rect 11244 7890 11296 7896
rect 10968 7812 11020 7818
rect 10968 7754 11020 7760
rect 10980 7478 11008 7754
rect 11256 7750 11284 7890
rect 11428 7880 11480 7886
rect 11428 7822 11480 7828
rect 11520 7880 11572 7886
rect 11520 7822 11572 7828
rect 11244 7744 11296 7750
rect 11244 7686 11296 7692
rect 11440 7546 11468 7822
rect 11428 7540 11480 7546
rect 11428 7482 11480 7488
rect 10968 7472 11020 7478
rect 10968 7414 11020 7420
rect 10796 6886 10916 6914
rect 10692 6384 10744 6390
rect 10692 6326 10744 6332
rect 10704 6254 10732 6326
rect 10796 6254 10824 6886
rect 10692 6248 10744 6254
rect 10692 6190 10744 6196
rect 10784 6248 10836 6254
rect 10784 6190 10836 6196
rect 11060 6248 11112 6254
rect 11060 6190 11112 6196
rect 10796 5778 10824 6190
rect 11072 5914 11100 6190
rect 11060 5908 11112 5914
rect 11060 5850 11112 5856
rect 10784 5772 10836 5778
rect 10784 5714 10836 5720
rect 11428 4548 11480 4554
rect 11428 4490 11480 4496
rect 11060 4208 11112 4214
rect 11060 4150 11112 4156
rect 10876 3392 10928 3398
rect 10876 3334 10928 3340
rect 10888 2990 10916 3334
rect 10968 3052 11020 3058
rect 10968 2994 11020 3000
rect 10876 2984 10928 2990
rect 10876 2926 10928 2932
rect 10600 2576 10652 2582
rect 10600 2518 10652 2524
rect 10876 1080 10928 1086
rect 10876 1022 10928 1028
rect 10600 1012 10652 1018
rect 10600 954 10652 960
rect 10612 800 10640 954
rect 10888 800 10916 1022
rect 10980 1018 11008 2994
rect 11072 2122 11100 4150
rect 11072 2094 11192 2122
rect 10968 1012 11020 1018
rect 10968 954 11020 960
rect 11164 800 11192 2094
rect 11440 800 11468 4490
rect 11532 4146 11560 7822
rect 11716 7449 11744 11834
rect 12440 11076 12492 11082
rect 12440 11018 12492 11024
rect 12452 10674 12480 11018
rect 12348 10668 12400 10674
rect 12348 10610 12400 10616
rect 12440 10668 12492 10674
rect 12440 10610 12492 10616
rect 12360 10266 12388 10610
rect 12348 10260 12400 10266
rect 12348 10202 12400 10208
rect 12452 10062 12480 10610
rect 12544 10130 12572 14282
rect 13372 12434 13400 14486
rect 14464 14272 14516 14278
rect 14464 14214 14516 14220
rect 13280 12406 13400 12434
rect 13084 12232 13136 12238
rect 13084 12174 13136 12180
rect 13096 11898 13124 12174
rect 13176 12164 13228 12170
rect 13176 12106 13228 12112
rect 13084 11892 13136 11898
rect 13084 11834 13136 11840
rect 13188 11694 13216 12106
rect 13176 11688 13228 11694
rect 13176 11630 13228 11636
rect 13176 11280 13228 11286
rect 13176 11222 13228 11228
rect 13084 10532 13136 10538
rect 13084 10474 13136 10480
rect 12622 10160 12678 10169
rect 12532 10124 12584 10130
rect 12622 10095 12624 10104
rect 12532 10066 12584 10072
rect 12676 10095 12678 10104
rect 12624 10066 12676 10072
rect 12348 10056 12400 10062
rect 12348 9998 12400 10004
rect 12440 10056 12492 10062
rect 12440 9998 12492 10004
rect 12256 9580 12308 9586
rect 12256 9522 12308 9528
rect 12268 9178 12296 9522
rect 12360 9518 12388 9998
rect 12544 9586 12572 10066
rect 12532 9580 12584 9586
rect 12532 9522 12584 9528
rect 12348 9512 12400 9518
rect 12348 9454 12400 9460
rect 12808 9512 12860 9518
rect 12808 9454 12860 9460
rect 12624 9444 12676 9450
rect 12624 9386 12676 9392
rect 12256 9172 12308 9178
rect 12256 9114 12308 9120
rect 12636 8974 12664 9386
rect 12164 8968 12216 8974
rect 12624 8968 12676 8974
rect 12164 8910 12216 8916
rect 12544 8928 12624 8956
rect 12176 8634 12204 8910
rect 12348 8900 12400 8906
rect 12348 8842 12400 8848
rect 12164 8628 12216 8634
rect 12164 8570 12216 8576
rect 12360 8498 12388 8842
rect 12440 8832 12492 8838
rect 12440 8774 12492 8780
rect 12452 8498 12480 8774
rect 12544 8566 12572 8928
rect 12624 8910 12676 8916
rect 12716 8968 12768 8974
rect 12716 8910 12768 8916
rect 12532 8560 12584 8566
rect 12532 8502 12584 8508
rect 12348 8492 12400 8498
rect 12348 8434 12400 8440
rect 12440 8492 12492 8498
rect 12440 8434 12492 8440
rect 12544 8430 12572 8502
rect 12532 8424 12584 8430
rect 12452 8372 12532 8378
rect 12452 8366 12584 8372
rect 12624 8424 12676 8430
rect 12624 8366 12676 8372
rect 12452 8350 12572 8366
rect 12452 7954 12480 8350
rect 12636 8090 12664 8366
rect 12624 8084 12676 8090
rect 12624 8026 12676 8032
rect 12440 7948 12492 7954
rect 12440 7890 12492 7896
rect 12728 7546 12756 8910
rect 12820 8022 12848 9454
rect 12900 9376 12952 9382
rect 12900 9318 12952 9324
rect 12808 8016 12860 8022
rect 12808 7958 12860 7964
rect 12716 7540 12768 7546
rect 12716 7482 12768 7488
rect 11702 7440 11758 7449
rect 11702 7375 11758 7384
rect 12348 7404 12400 7410
rect 12348 7346 12400 7352
rect 12072 7268 12124 7274
rect 12072 7210 12124 7216
rect 12084 4758 12112 7210
rect 12360 5914 12388 7346
rect 12912 6338 12940 9318
rect 12544 6310 12940 6338
rect 12348 5908 12400 5914
rect 12348 5850 12400 5856
rect 12072 4752 12124 4758
rect 12072 4694 12124 4700
rect 11520 4140 11572 4146
rect 11520 4082 11572 4088
rect 11980 4004 12032 4010
rect 11980 3946 12032 3952
rect 11888 3936 11940 3942
rect 11888 3878 11940 3884
rect 11900 2922 11928 3878
rect 11992 3126 12020 3946
rect 12072 3392 12124 3398
rect 12072 3334 12124 3340
rect 12084 3194 12112 3334
rect 12072 3188 12124 3194
rect 12072 3130 12124 3136
rect 11980 3120 12032 3126
rect 11980 3062 12032 3068
rect 11888 2916 11940 2922
rect 11888 2858 11940 2864
rect 12544 2582 12572 6310
rect 12716 4072 12768 4078
rect 12636 4020 12716 4026
rect 12636 4014 12768 4020
rect 12636 3998 12756 4014
rect 12636 3398 12664 3998
rect 12716 3936 12768 3942
rect 12716 3878 12768 3884
rect 12992 3936 13044 3942
rect 12992 3878 13044 3884
rect 12728 3602 12756 3878
rect 12716 3596 12768 3602
rect 12716 3538 12768 3544
rect 12808 3460 12860 3466
rect 12808 3402 12860 3408
rect 12624 3392 12676 3398
rect 12624 3334 12676 3340
rect 12532 2576 12584 2582
rect 12532 2518 12584 2524
rect 12532 2440 12584 2446
rect 12532 2382 12584 2388
rect 11704 2372 11756 2378
rect 11704 2314 11756 2320
rect 12072 2372 12124 2378
rect 12072 2314 12124 2320
rect 11716 800 11744 2314
rect 12084 950 12112 2314
rect 12256 1012 12308 1018
rect 12256 954 12308 960
rect 11980 944 12032 950
rect 11980 886 12032 892
rect 12072 944 12124 950
rect 12072 886 12124 892
rect 11992 800 12020 886
rect 12268 800 12296 954
rect 12544 800 12572 2382
rect 12820 800 12848 3402
rect 13004 3398 13032 3878
rect 12992 3392 13044 3398
rect 12992 3334 13044 3340
rect 13096 2990 13124 10474
rect 13084 2984 13136 2990
rect 13084 2926 13136 2932
rect 13188 2650 13216 11222
rect 13280 2650 13308 12406
rect 13544 12300 13596 12306
rect 13544 12242 13596 12248
rect 13452 12232 13504 12238
rect 13452 12174 13504 12180
rect 13464 11898 13492 12174
rect 13452 11892 13504 11898
rect 13452 11834 13504 11840
rect 13556 11778 13584 12242
rect 13636 12232 13688 12238
rect 13636 12174 13688 12180
rect 13464 11750 13584 11778
rect 13464 11694 13492 11750
rect 13452 11688 13504 11694
rect 13452 11630 13504 11636
rect 13544 11688 13596 11694
rect 13544 11630 13596 11636
rect 13464 11150 13492 11630
rect 13452 11144 13504 11150
rect 13452 11086 13504 11092
rect 13464 10674 13492 11086
rect 13556 10810 13584 11630
rect 13648 11354 13676 12174
rect 13636 11348 13688 11354
rect 13636 11290 13688 11296
rect 14476 11218 14504 14214
rect 14554 11248 14610 11257
rect 14464 11212 14516 11218
rect 14554 11183 14556 11192
rect 14464 11154 14516 11160
rect 14608 11183 14610 11192
rect 14556 11154 14608 11160
rect 14740 11144 14792 11150
rect 14740 11086 14792 11092
rect 14752 10810 14780 11086
rect 13544 10804 13596 10810
rect 13544 10746 13596 10752
rect 14740 10804 14792 10810
rect 14740 10746 14792 10752
rect 13452 10668 13504 10674
rect 13452 10610 13504 10616
rect 13544 10464 13596 10470
rect 13544 10406 13596 10412
rect 13360 9988 13412 9994
rect 13360 9930 13412 9936
rect 13372 7954 13400 9930
rect 13360 7948 13412 7954
rect 13360 7890 13412 7896
rect 13372 3942 13400 7890
rect 13452 7268 13504 7274
rect 13452 7210 13504 7216
rect 13360 3936 13412 3942
rect 13360 3878 13412 3884
rect 13360 3460 13412 3466
rect 13360 3402 13412 3408
rect 13176 2644 13228 2650
rect 13176 2586 13228 2592
rect 13268 2644 13320 2650
rect 13268 2586 13320 2592
rect 13268 2372 13320 2378
rect 13268 2314 13320 2320
rect 13280 1086 13308 2314
rect 13268 1080 13320 1086
rect 13268 1022 13320 1028
rect 13084 944 13136 950
rect 13084 886 13136 892
rect 13096 800 13124 886
rect 13372 800 13400 3402
rect 13464 2582 13492 7210
rect 13556 3738 13584 10406
rect 13820 10056 13872 10062
rect 13820 9998 13872 10004
rect 13832 9518 13860 9998
rect 13820 9512 13872 9518
rect 13820 9454 13872 9460
rect 14464 6860 14516 6866
rect 14464 6802 14516 6808
rect 13912 6792 13964 6798
rect 13912 6734 13964 6740
rect 13820 5840 13872 5846
rect 13820 5782 13872 5788
rect 13544 3732 13596 3738
rect 13544 3674 13596 3680
rect 13832 3194 13860 5782
rect 13820 3188 13872 3194
rect 13820 3130 13872 3136
rect 13636 3052 13688 3058
rect 13636 2994 13688 3000
rect 13728 3052 13780 3058
rect 13728 2994 13780 3000
rect 13452 2576 13504 2582
rect 13452 2518 13504 2524
rect 13544 2372 13596 2378
rect 13544 2314 13596 2320
rect 13556 1018 13584 2314
rect 13544 1012 13596 1018
rect 13544 954 13596 960
rect 13648 800 13676 2994
rect 13740 950 13768 2994
rect 13924 2990 13952 6734
rect 14476 3738 14504 6802
rect 14464 3732 14516 3738
rect 14464 3674 14516 3680
rect 14188 3460 14240 3466
rect 14188 3402 14240 3408
rect 13912 2984 13964 2990
rect 13912 2926 13964 2932
rect 13912 1080 13964 1086
rect 13912 1022 13964 1028
rect 13728 944 13780 950
rect 13728 886 13780 892
rect 13924 800 13952 1022
rect 14200 800 14228 3402
rect 14936 2446 14964 16934
rect 15028 14414 15056 29446
rect 15396 28150 15424 57190
rect 17144 30326 17172 57258
rect 17960 57248 18012 57254
rect 17960 57190 18012 57196
rect 19984 57248 20036 57254
rect 19984 57190 20036 57196
rect 20168 57248 20220 57254
rect 20168 57190 20220 57196
rect 22192 57248 22244 57254
rect 22192 57190 22244 57196
rect 22652 57248 22704 57254
rect 22652 57190 22704 57196
rect 24768 57248 24820 57254
rect 24768 57190 24820 57196
rect 25688 57248 25740 57254
rect 25688 57190 25740 57196
rect 26700 57248 26752 57254
rect 26700 57190 26752 57196
rect 17972 56914 18000 57190
rect 17960 56908 18012 56914
rect 17960 56850 18012 56856
rect 19574 56604 19882 56613
rect 19574 56602 19580 56604
rect 19636 56602 19660 56604
rect 19716 56602 19740 56604
rect 19796 56602 19820 56604
rect 19876 56602 19882 56604
rect 19636 56550 19638 56602
rect 19818 56550 19820 56602
rect 19574 56548 19580 56550
rect 19636 56548 19660 56550
rect 19716 56548 19740 56550
rect 19796 56548 19820 56550
rect 19876 56548 19882 56550
rect 19574 56539 19882 56548
rect 18604 56296 18656 56302
rect 18604 56238 18656 56244
rect 17132 30320 17184 30326
rect 17132 30262 17184 30268
rect 17224 30252 17276 30258
rect 17224 30194 17276 30200
rect 15384 28144 15436 28150
rect 15384 28086 15436 28092
rect 15752 24812 15804 24818
rect 15752 24754 15804 24760
rect 15764 23730 15792 24754
rect 17236 24342 17264 30194
rect 17224 24336 17276 24342
rect 17224 24278 17276 24284
rect 17776 24336 17828 24342
rect 17776 24278 17828 24284
rect 16120 24268 16172 24274
rect 16120 24210 16172 24216
rect 16132 23866 16160 24210
rect 16120 23860 16172 23866
rect 16120 23802 16172 23808
rect 17788 23730 17816 24278
rect 15752 23724 15804 23730
rect 15752 23666 15804 23672
rect 17776 23724 17828 23730
rect 17776 23666 17828 23672
rect 18512 22772 18564 22778
rect 18512 22714 18564 22720
rect 17408 20256 17460 20262
rect 17408 20198 17460 20204
rect 17224 19780 17276 19786
rect 17224 19722 17276 19728
rect 17236 16658 17264 19722
rect 17420 16998 17448 20198
rect 17960 17672 18012 17678
rect 17960 17614 18012 17620
rect 18420 17672 18472 17678
rect 18420 17614 18472 17620
rect 17592 17196 17644 17202
rect 17592 17138 17644 17144
rect 17408 16992 17460 16998
rect 17408 16934 17460 16940
rect 17500 16992 17552 16998
rect 17500 16934 17552 16940
rect 17224 16652 17276 16658
rect 17224 16594 17276 16600
rect 16212 16584 16264 16590
rect 16212 16526 16264 16532
rect 16224 16250 16252 16526
rect 16212 16244 16264 16250
rect 16212 16186 16264 16192
rect 17236 16046 17264 16594
rect 17512 16590 17540 16934
rect 17604 16794 17632 17138
rect 17868 16992 17920 16998
rect 17868 16934 17920 16940
rect 17592 16788 17644 16794
rect 17592 16730 17644 16736
rect 17500 16584 17552 16590
rect 17500 16526 17552 16532
rect 17776 16108 17828 16114
rect 17776 16050 17828 16056
rect 17224 16040 17276 16046
rect 17224 15982 17276 15988
rect 17684 16040 17736 16046
rect 17684 15982 17736 15988
rect 15476 15632 15528 15638
rect 15476 15574 15528 15580
rect 15842 15600 15898 15609
rect 15488 14958 15516 15574
rect 15842 15535 15844 15544
rect 15896 15535 15898 15544
rect 15844 15506 15896 15512
rect 15660 15496 15712 15502
rect 15660 15438 15712 15444
rect 15752 15496 15804 15502
rect 15752 15438 15804 15444
rect 16212 15496 16264 15502
rect 16212 15438 16264 15444
rect 15476 14952 15528 14958
rect 15476 14894 15528 14900
rect 15568 14952 15620 14958
rect 15568 14894 15620 14900
rect 15108 14476 15160 14482
rect 15108 14418 15160 14424
rect 15016 14408 15068 14414
rect 15016 14350 15068 14356
rect 15120 14278 15148 14418
rect 15108 14272 15160 14278
rect 15108 14214 15160 14220
rect 15488 14006 15516 14894
rect 15580 14074 15608 14894
rect 15672 14618 15700 15438
rect 15764 15162 15792 15438
rect 15752 15156 15804 15162
rect 15752 15098 15804 15104
rect 15764 15026 15792 15098
rect 15752 15020 15804 15026
rect 15752 14962 15804 14968
rect 15660 14612 15712 14618
rect 15660 14554 15712 14560
rect 15844 14340 15896 14346
rect 15844 14282 15896 14288
rect 15568 14068 15620 14074
rect 15568 14010 15620 14016
rect 15476 14000 15528 14006
rect 15476 13942 15528 13948
rect 15292 13796 15344 13802
rect 15292 13738 15344 13744
rect 15108 11008 15160 11014
rect 15108 10950 15160 10956
rect 15120 4146 15148 10950
rect 15108 4140 15160 4146
rect 15108 4082 15160 4088
rect 15304 3738 15332 13738
rect 15488 13394 15516 13942
rect 15476 13388 15528 13394
rect 15476 13330 15528 13336
rect 15488 12306 15516 13330
rect 15476 12300 15528 12306
rect 15476 12242 15528 12248
rect 15488 11354 15516 12242
rect 15476 11348 15528 11354
rect 15476 11290 15528 11296
rect 15856 11150 15884 14282
rect 16224 13530 16252 15438
rect 17408 15156 17460 15162
rect 17408 15098 17460 15104
rect 17420 14482 17448 15098
rect 17500 14816 17552 14822
rect 17500 14758 17552 14764
rect 17316 14476 17368 14482
rect 17316 14418 17368 14424
rect 17408 14476 17460 14482
rect 17408 14418 17460 14424
rect 17328 14006 17356 14418
rect 17512 14414 17540 14758
rect 17696 14550 17724 15982
rect 17788 15638 17816 16050
rect 17776 15632 17828 15638
rect 17776 15574 17828 15580
rect 17880 15570 17908 16934
rect 17868 15564 17920 15570
rect 17868 15506 17920 15512
rect 17880 15094 17908 15506
rect 17972 15434 18000 17614
rect 18328 17536 18380 17542
rect 18328 17478 18380 17484
rect 18340 17202 18368 17478
rect 18328 17196 18380 17202
rect 18328 17138 18380 17144
rect 18432 16046 18460 17614
rect 18420 16040 18472 16046
rect 18420 15982 18472 15988
rect 18236 15904 18288 15910
rect 18236 15846 18288 15852
rect 17960 15428 18012 15434
rect 17960 15370 18012 15376
rect 17868 15088 17920 15094
rect 17868 15030 17920 15036
rect 17684 14544 17736 14550
rect 17684 14486 17736 14492
rect 17500 14408 17552 14414
rect 17500 14350 17552 14356
rect 17316 14000 17368 14006
rect 17316 13942 17368 13948
rect 16212 13524 16264 13530
rect 16212 13466 16264 13472
rect 16028 13456 16080 13462
rect 16028 13398 16080 13404
rect 15936 11280 15988 11286
rect 15936 11222 15988 11228
rect 15844 11144 15896 11150
rect 15844 11086 15896 11092
rect 15844 4820 15896 4826
rect 15844 4762 15896 4768
rect 15568 4208 15620 4214
rect 15568 4150 15620 4156
rect 15292 3732 15344 3738
rect 15292 3674 15344 3680
rect 15292 3460 15344 3466
rect 15292 3402 15344 3408
rect 15016 3052 15068 3058
rect 15016 2994 15068 3000
rect 14924 2440 14976 2446
rect 14924 2382 14976 2388
rect 14740 1012 14792 1018
rect 14740 954 14792 960
rect 14464 944 14516 950
rect 14464 886 14516 892
rect 14476 800 14504 886
rect 14752 800 14780 954
rect 15028 800 15056 2994
rect 15304 800 15332 3402
rect 15580 800 15608 4150
rect 15660 4140 15712 4146
rect 15660 4082 15712 4088
rect 15672 2854 15700 4082
rect 15856 3058 15884 4762
rect 15752 3052 15804 3058
rect 15752 2994 15804 3000
rect 15844 3052 15896 3058
rect 15844 2994 15896 3000
rect 15660 2848 15712 2854
rect 15660 2790 15712 2796
rect 15764 1578 15792 2994
rect 15844 2440 15896 2446
rect 15844 2382 15896 2388
rect 15856 1970 15884 2382
rect 15948 2310 15976 11222
rect 16040 3738 16068 13398
rect 18052 11688 18104 11694
rect 18052 11630 18104 11636
rect 18144 11688 18196 11694
rect 18144 11630 18196 11636
rect 16120 11212 16172 11218
rect 16120 11154 16172 11160
rect 16132 4078 16160 11154
rect 18064 11082 18092 11630
rect 18156 11354 18184 11630
rect 18144 11348 18196 11354
rect 18144 11290 18196 11296
rect 18052 11076 18104 11082
rect 18052 11018 18104 11024
rect 17040 10464 17092 10470
rect 17040 10406 17092 10412
rect 16580 6180 16632 6186
rect 16580 6122 16632 6128
rect 16120 4072 16172 4078
rect 16120 4014 16172 4020
rect 16028 3732 16080 3738
rect 16028 3674 16080 3680
rect 16120 3460 16172 3466
rect 16120 3402 16172 3408
rect 15936 2304 15988 2310
rect 15936 2246 15988 2252
rect 15844 1964 15896 1970
rect 15844 1906 15896 1912
rect 15764 1550 15884 1578
rect 15856 800 15884 1550
rect 16132 800 16160 3402
rect 16592 3398 16620 6122
rect 17052 4146 17080 10406
rect 17960 9716 18012 9722
rect 17960 9658 18012 9664
rect 17316 9580 17368 9586
rect 17316 9522 17368 9528
rect 17328 8906 17356 9522
rect 17316 8900 17368 8906
rect 17316 8842 17368 8848
rect 17316 8288 17368 8294
rect 17316 8230 17368 8236
rect 17132 4480 17184 4486
rect 17132 4422 17184 4428
rect 17040 4140 17092 4146
rect 17040 4082 17092 4088
rect 16672 3732 16724 3738
rect 16672 3674 16724 3680
rect 16684 3534 16712 3674
rect 17144 3670 17172 4422
rect 17328 4146 17356 8230
rect 17316 4140 17368 4146
rect 17316 4082 17368 4088
rect 17224 4072 17276 4078
rect 17224 4014 17276 4020
rect 17132 3664 17184 3670
rect 17132 3606 17184 3612
rect 16672 3528 16724 3534
rect 16672 3470 16724 3476
rect 16762 3496 16818 3505
rect 16762 3431 16764 3440
rect 16816 3431 16818 3440
rect 16948 3460 17000 3466
rect 16764 3402 16816 3408
rect 16948 3402 17000 3408
rect 16580 3392 16632 3398
rect 16580 3334 16632 3340
rect 16488 2984 16540 2990
rect 16488 2926 16540 2932
rect 16396 2508 16448 2514
rect 16396 2450 16448 2456
rect 16408 800 16436 2450
rect 16500 898 16528 2926
rect 16500 870 16712 898
rect 16684 800 16712 870
rect 16960 800 16988 3402
rect 17040 2848 17092 2854
rect 17040 2790 17092 2796
rect 17052 950 17080 2790
rect 17040 944 17092 950
rect 17040 886 17092 892
rect 17236 800 17264 4014
rect 17316 3664 17368 3670
rect 17316 3606 17368 3612
rect 17328 2922 17356 3606
rect 17972 3534 18000 9658
rect 18248 8294 18276 15846
rect 18432 15434 18460 15982
rect 18420 15428 18472 15434
rect 18420 15370 18472 15376
rect 18420 8968 18472 8974
rect 18420 8910 18472 8916
rect 18236 8288 18288 8294
rect 18236 8230 18288 8236
rect 18328 6452 18380 6458
rect 18328 6394 18380 6400
rect 18144 5704 18196 5710
rect 18144 5646 18196 5652
rect 18236 5704 18288 5710
rect 18236 5646 18288 5652
rect 18156 4690 18184 5646
rect 18248 4826 18276 5646
rect 18236 4820 18288 4826
rect 18236 4762 18288 4768
rect 18340 4706 18368 6394
rect 18144 4684 18196 4690
rect 18144 4626 18196 4632
rect 18248 4678 18368 4706
rect 18052 4616 18104 4622
rect 18052 4558 18104 4564
rect 17960 3528 18012 3534
rect 17960 3470 18012 3476
rect 17592 3460 17644 3466
rect 17592 3402 17644 3408
rect 17316 2916 17368 2922
rect 17316 2858 17368 2864
rect 17408 2440 17460 2446
rect 17408 2382 17460 2388
rect 17420 1018 17448 2382
rect 17604 1714 17632 3402
rect 17960 3120 18012 3126
rect 17958 3088 17960 3097
rect 18012 3088 18014 3097
rect 17958 3023 18014 3032
rect 17868 2984 17920 2990
rect 17868 2926 17920 2932
rect 17776 2576 17828 2582
rect 17776 2518 17828 2524
rect 17512 1686 17632 1714
rect 17408 1012 17460 1018
rect 17408 954 17460 960
rect 17512 800 17540 1686
rect 17788 800 17816 2518
rect 17880 1086 17908 2926
rect 17868 1080 17920 1086
rect 17868 1022 17920 1028
rect 18064 800 18092 4558
rect 18144 3936 18196 3942
rect 18144 3878 18196 3884
rect 18156 2922 18184 3878
rect 18248 3058 18276 4678
rect 18328 3936 18380 3942
rect 18328 3878 18380 3884
rect 18236 3052 18288 3058
rect 18236 2994 18288 3000
rect 18144 2916 18196 2922
rect 18144 2858 18196 2864
rect 18236 2440 18288 2446
rect 18236 2382 18288 2388
rect 18248 2038 18276 2382
rect 18236 2032 18288 2038
rect 18236 1974 18288 1980
rect 18340 800 18368 3878
rect 18432 2446 18460 8910
rect 18524 3534 18552 22714
rect 18616 18086 18644 56238
rect 19574 55516 19882 55525
rect 19574 55514 19580 55516
rect 19636 55514 19660 55516
rect 19716 55514 19740 55516
rect 19796 55514 19820 55516
rect 19876 55514 19882 55516
rect 19636 55462 19638 55514
rect 19818 55462 19820 55514
rect 19574 55460 19580 55462
rect 19636 55460 19660 55462
rect 19716 55460 19740 55462
rect 19796 55460 19820 55462
rect 19876 55460 19882 55462
rect 19574 55451 19882 55460
rect 19574 54428 19882 54437
rect 19574 54426 19580 54428
rect 19636 54426 19660 54428
rect 19716 54426 19740 54428
rect 19796 54426 19820 54428
rect 19876 54426 19882 54428
rect 19636 54374 19638 54426
rect 19818 54374 19820 54426
rect 19574 54372 19580 54374
rect 19636 54372 19660 54374
rect 19716 54372 19740 54374
rect 19796 54372 19820 54374
rect 19876 54372 19882 54374
rect 19574 54363 19882 54372
rect 19574 53340 19882 53349
rect 19574 53338 19580 53340
rect 19636 53338 19660 53340
rect 19716 53338 19740 53340
rect 19796 53338 19820 53340
rect 19876 53338 19882 53340
rect 19636 53286 19638 53338
rect 19818 53286 19820 53338
rect 19574 53284 19580 53286
rect 19636 53284 19660 53286
rect 19716 53284 19740 53286
rect 19796 53284 19820 53286
rect 19876 53284 19882 53286
rect 19574 53275 19882 53284
rect 19574 52252 19882 52261
rect 19574 52250 19580 52252
rect 19636 52250 19660 52252
rect 19716 52250 19740 52252
rect 19796 52250 19820 52252
rect 19876 52250 19882 52252
rect 19636 52198 19638 52250
rect 19818 52198 19820 52250
rect 19574 52196 19580 52198
rect 19636 52196 19660 52198
rect 19716 52196 19740 52198
rect 19796 52196 19820 52198
rect 19876 52196 19882 52198
rect 19574 52187 19882 52196
rect 19574 51164 19882 51173
rect 19574 51162 19580 51164
rect 19636 51162 19660 51164
rect 19716 51162 19740 51164
rect 19796 51162 19820 51164
rect 19876 51162 19882 51164
rect 19636 51110 19638 51162
rect 19818 51110 19820 51162
rect 19574 51108 19580 51110
rect 19636 51108 19660 51110
rect 19716 51108 19740 51110
rect 19796 51108 19820 51110
rect 19876 51108 19882 51110
rect 19574 51099 19882 51108
rect 19574 50076 19882 50085
rect 19574 50074 19580 50076
rect 19636 50074 19660 50076
rect 19716 50074 19740 50076
rect 19796 50074 19820 50076
rect 19876 50074 19882 50076
rect 19636 50022 19638 50074
rect 19818 50022 19820 50074
rect 19574 50020 19580 50022
rect 19636 50020 19660 50022
rect 19716 50020 19740 50022
rect 19796 50020 19820 50022
rect 19876 50020 19882 50022
rect 19574 50011 19882 50020
rect 19574 48988 19882 48997
rect 19574 48986 19580 48988
rect 19636 48986 19660 48988
rect 19716 48986 19740 48988
rect 19796 48986 19820 48988
rect 19876 48986 19882 48988
rect 19636 48934 19638 48986
rect 19818 48934 19820 48986
rect 19574 48932 19580 48934
rect 19636 48932 19660 48934
rect 19716 48932 19740 48934
rect 19796 48932 19820 48934
rect 19876 48932 19882 48934
rect 19574 48923 19882 48932
rect 19574 47900 19882 47909
rect 19574 47898 19580 47900
rect 19636 47898 19660 47900
rect 19716 47898 19740 47900
rect 19796 47898 19820 47900
rect 19876 47898 19882 47900
rect 19636 47846 19638 47898
rect 19818 47846 19820 47898
rect 19574 47844 19580 47846
rect 19636 47844 19660 47846
rect 19716 47844 19740 47846
rect 19796 47844 19820 47846
rect 19876 47844 19882 47846
rect 19574 47835 19882 47844
rect 19574 46812 19882 46821
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46747 19882 46756
rect 19574 45724 19882 45733
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45659 19882 45668
rect 19574 44636 19882 44645
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44571 19882 44580
rect 19574 43548 19882 43557
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43483 19882 43492
rect 19574 42460 19882 42469
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42395 19882 42404
rect 19574 41372 19882 41381
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41307 19882 41316
rect 19574 40284 19882 40293
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40219 19882 40228
rect 19574 39196 19882 39205
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39131 19882 39140
rect 19574 38108 19882 38117
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38043 19882 38052
rect 19432 37324 19484 37330
rect 19432 37266 19484 37272
rect 19340 36780 19392 36786
rect 19340 36722 19392 36728
rect 19352 35894 19380 36722
rect 19444 36174 19472 37266
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 19432 36168 19484 36174
rect 19432 36110 19484 36116
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19352 35866 19472 35894
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19444 31278 19472 35866
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19996 32502 20024 57190
rect 20180 36174 20208 57190
rect 22204 57050 22232 57190
rect 22192 57044 22244 57050
rect 22192 56986 22244 56992
rect 21364 55684 21416 55690
rect 21364 55626 21416 55632
rect 21272 41472 21324 41478
rect 21272 41414 21324 41420
rect 21284 38350 21312 41414
rect 21272 38344 21324 38350
rect 21272 38286 21324 38292
rect 20168 36168 20220 36174
rect 20168 36110 20220 36116
rect 19984 32496 20036 32502
rect 19984 32438 20036 32444
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19432 31272 19484 31278
rect 19432 31214 19484 31220
rect 19444 28626 19472 31214
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19432 28620 19484 28626
rect 19432 28562 19484 28568
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 18972 28212 19024 28218
rect 18972 28154 19024 28160
rect 18984 27334 19012 28154
rect 18972 27328 19024 27334
rect 18972 27270 19024 27276
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 20168 26376 20220 26382
rect 20168 26318 20220 26324
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 20180 25974 20208 26318
rect 20168 25968 20220 25974
rect 20168 25910 20220 25916
rect 20996 25900 21048 25906
rect 20996 25842 21048 25848
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 21008 24818 21036 25842
rect 20996 24812 21048 24818
rect 20996 24754 21048 24760
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 21008 23798 21036 24754
rect 20996 23792 21048 23798
rect 20996 23734 21048 23740
rect 21376 23322 21404 55626
rect 21456 36712 21508 36718
rect 21456 36654 21508 36660
rect 21468 36106 21496 36654
rect 21456 36100 21508 36106
rect 21456 36042 21508 36048
rect 22468 30252 22520 30258
rect 22468 30194 22520 30200
rect 22376 30184 22428 30190
rect 22376 30126 22428 30132
rect 22284 30048 22336 30054
rect 22282 30016 22284 30025
rect 22336 30016 22338 30025
rect 22282 29951 22338 29960
rect 22282 29336 22338 29345
rect 22282 29271 22284 29280
rect 22336 29271 22338 29280
rect 22284 29242 22336 29248
rect 22284 28212 22336 28218
rect 22284 28154 22336 28160
rect 22296 28014 22324 28154
rect 22284 28008 22336 28014
rect 22284 27950 22336 27956
rect 22388 27674 22416 30126
rect 22480 29306 22508 30194
rect 22468 29300 22520 29306
rect 22468 29242 22520 29248
rect 22468 28212 22520 28218
rect 22468 28154 22520 28160
rect 22376 27668 22428 27674
rect 22376 27610 22428 27616
rect 22100 27464 22152 27470
rect 22100 27406 22152 27412
rect 21364 23316 21416 23322
rect 21364 23258 21416 23264
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 22008 22024 22060 22030
rect 22008 21966 22060 21972
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 22020 20942 22048 21966
rect 22112 21554 22140 27406
rect 22388 25906 22416 27610
rect 22376 25900 22428 25906
rect 22376 25842 22428 25848
rect 22284 25152 22336 25158
rect 22284 25094 22336 25100
rect 22296 24886 22324 25094
rect 22284 24880 22336 24886
rect 22284 24822 22336 24828
rect 22192 24812 22244 24818
rect 22192 24754 22244 24760
rect 22100 21548 22152 21554
rect 22100 21490 22152 21496
rect 22008 20936 22060 20942
rect 22008 20878 22060 20884
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 22204 19922 22232 24754
rect 22480 22710 22508 28154
rect 22468 22704 22520 22710
rect 22468 22646 22520 22652
rect 22664 22094 22692 57190
rect 22744 42084 22796 42090
rect 22744 42026 22796 42032
rect 22756 29306 22784 42026
rect 23204 35488 23256 35494
rect 23204 35430 23256 35436
rect 23020 32972 23072 32978
rect 23020 32914 23072 32920
rect 22836 30320 22888 30326
rect 22836 30262 22888 30268
rect 22848 30054 22876 30262
rect 22928 30252 22980 30258
rect 22928 30194 22980 30200
rect 22836 30048 22888 30054
rect 22836 29990 22888 29996
rect 22940 29306 22968 30194
rect 22744 29300 22796 29306
rect 22744 29242 22796 29248
rect 22928 29300 22980 29306
rect 22928 29242 22980 29248
rect 22756 29170 22784 29242
rect 22744 29164 22796 29170
rect 22744 29106 22796 29112
rect 23032 27538 23060 32914
rect 23216 30258 23244 35430
rect 24400 34740 24452 34746
rect 24400 34682 24452 34688
rect 24412 34626 24440 34682
rect 24412 34610 24624 34626
rect 24308 34604 24360 34610
rect 24412 34604 24636 34610
rect 24412 34598 24584 34604
rect 24308 34546 24360 34552
rect 24584 34546 24636 34552
rect 24320 31754 24348 34546
rect 24780 31754 24808 57190
rect 24320 31726 24440 31754
rect 23112 30252 23164 30258
rect 23112 30194 23164 30200
rect 23204 30252 23256 30258
rect 23204 30194 23256 30200
rect 23296 30252 23348 30258
rect 23296 30194 23348 30200
rect 24216 30252 24268 30258
rect 24216 30194 24268 30200
rect 23124 29714 23152 30194
rect 23112 29708 23164 29714
rect 23112 29650 23164 29656
rect 23308 29646 23336 30194
rect 23756 30048 23808 30054
rect 23756 29990 23808 29996
rect 23296 29640 23348 29646
rect 23296 29582 23348 29588
rect 23570 29336 23626 29345
rect 23388 29300 23440 29306
rect 23570 29271 23626 29280
rect 23388 29242 23440 29248
rect 23204 29164 23256 29170
rect 23204 29106 23256 29112
rect 23216 29073 23244 29106
rect 23202 29064 23258 29073
rect 23202 28999 23258 29008
rect 23296 28552 23348 28558
rect 23296 28494 23348 28500
rect 23308 28082 23336 28494
rect 23400 28490 23428 29242
rect 23584 29238 23612 29271
rect 23572 29232 23624 29238
rect 23572 29174 23624 29180
rect 23768 29170 23796 29990
rect 23756 29164 23808 29170
rect 23756 29106 23808 29112
rect 23662 29064 23718 29073
rect 23662 28999 23718 29008
rect 23676 28626 23704 28999
rect 23664 28620 23716 28626
rect 23664 28562 23716 28568
rect 23388 28484 23440 28490
rect 23388 28426 23440 28432
rect 23400 28082 23428 28426
rect 23296 28076 23348 28082
rect 23296 28018 23348 28024
rect 23388 28076 23440 28082
rect 23440 28036 23612 28064
rect 23388 28018 23440 28024
rect 23308 27826 23336 28018
rect 23308 27798 23428 27826
rect 23020 27532 23072 27538
rect 23020 27474 23072 27480
rect 23296 27464 23348 27470
rect 23296 27406 23348 27412
rect 23018 27024 23074 27033
rect 23018 26959 23020 26968
rect 23072 26959 23074 26968
rect 23020 26930 23072 26936
rect 22928 26920 22980 26926
rect 22928 26862 22980 26868
rect 22940 26586 22968 26862
rect 22928 26580 22980 26586
rect 22928 26522 22980 26528
rect 22940 25974 22968 26522
rect 23032 26042 23060 26930
rect 23204 26308 23256 26314
rect 23204 26250 23256 26256
rect 23020 26036 23072 26042
rect 23020 25978 23072 25984
rect 22928 25968 22980 25974
rect 22928 25910 22980 25916
rect 22940 25362 22968 25910
rect 23112 25764 23164 25770
rect 23112 25706 23164 25712
rect 22928 25356 22980 25362
rect 22928 25298 22980 25304
rect 23124 24206 23152 25706
rect 23216 24614 23244 26250
rect 23308 25906 23336 27406
rect 23400 26994 23428 27798
rect 23584 27470 23612 28036
rect 23676 27606 23704 28562
rect 23768 28558 23796 29106
rect 23756 28552 23808 28558
rect 23756 28494 23808 28500
rect 23768 28082 23796 28494
rect 23756 28076 23808 28082
rect 23756 28018 23808 28024
rect 23664 27600 23716 27606
rect 23664 27542 23716 27548
rect 23572 27464 23624 27470
rect 23572 27406 23624 27412
rect 23664 27464 23716 27470
rect 23664 27406 23716 27412
rect 23584 27130 23612 27406
rect 23572 27124 23624 27130
rect 23572 27066 23624 27072
rect 23388 26988 23440 26994
rect 23388 26930 23440 26936
rect 23400 26602 23428 26930
rect 23400 26574 23520 26602
rect 23296 25900 23348 25906
rect 23296 25842 23348 25848
rect 23308 25226 23336 25842
rect 23492 25362 23520 26574
rect 23676 25974 23704 27406
rect 23768 27334 23796 28018
rect 23756 27328 23808 27334
rect 23756 27270 23808 27276
rect 23664 25968 23716 25974
rect 23664 25910 23716 25916
rect 23940 25968 23992 25974
rect 23940 25910 23992 25916
rect 23572 25832 23624 25838
rect 23572 25774 23624 25780
rect 23480 25356 23532 25362
rect 23480 25298 23532 25304
rect 23584 25294 23612 25774
rect 23676 25430 23704 25910
rect 23664 25424 23716 25430
rect 23664 25366 23716 25372
rect 23572 25288 23624 25294
rect 23572 25230 23624 25236
rect 23296 25220 23348 25226
rect 23296 25162 23348 25168
rect 23308 24954 23336 25162
rect 23296 24948 23348 24954
rect 23296 24890 23348 24896
rect 23204 24608 23256 24614
rect 23204 24550 23256 24556
rect 23112 24200 23164 24206
rect 23112 24142 23164 24148
rect 23216 24138 23244 24550
rect 23308 24206 23336 24890
rect 23676 24886 23704 25366
rect 23664 24880 23716 24886
rect 23664 24822 23716 24828
rect 23480 24676 23532 24682
rect 23480 24618 23532 24624
rect 23296 24200 23348 24206
rect 23296 24142 23348 24148
rect 23204 24132 23256 24138
rect 23204 24074 23256 24080
rect 23216 23866 23244 24074
rect 23204 23860 23256 23866
rect 23204 23802 23256 23808
rect 22664 22066 22784 22094
rect 22284 21548 22336 21554
rect 22284 21490 22336 21496
rect 22192 19916 22244 19922
rect 22192 19858 22244 19864
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 18788 19372 18840 19378
rect 18788 19314 18840 19320
rect 20536 19372 20588 19378
rect 20536 19314 20588 19320
rect 18604 18080 18656 18086
rect 18604 18022 18656 18028
rect 18696 16448 18748 16454
rect 18696 16390 18748 16396
rect 18604 15360 18656 15366
rect 18604 15302 18656 15308
rect 18616 15026 18644 15302
rect 18604 15020 18656 15026
rect 18604 14962 18656 14968
rect 18708 10674 18736 16390
rect 18800 14550 18828 19314
rect 20548 19258 20576 19314
rect 20548 19230 20760 19258
rect 20732 18970 20760 19230
rect 22100 19168 22152 19174
rect 22100 19110 22152 19116
rect 20720 18964 20772 18970
rect 20720 18906 20772 18912
rect 22112 18834 22140 19110
rect 22100 18828 22152 18834
rect 22100 18770 22152 18776
rect 20812 18760 20864 18766
rect 20812 18702 20864 18708
rect 21548 18760 21600 18766
rect 21548 18702 21600 18708
rect 21732 18760 21784 18766
rect 21732 18702 21784 18708
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 20536 18352 20588 18358
rect 20536 18294 20588 18300
rect 20352 17536 20404 17542
rect 20352 17478 20404 17484
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19432 16652 19484 16658
rect 19432 16594 19484 16600
rect 19444 16114 19472 16594
rect 20364 16590 20392 17478
rect 20352 16584 20404 16590
rect 20548 16574 20576 18294
rect 20352 16526 20404 16532
rect 20456 16546 20576 16574
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 20456 16130 20484 16546
rect 19432 16108 19484 16114
rect 19432 16050 19484 16056
rect 20088 16102 20484 16130
rect 20720 16108 20772 16114
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 18788 14544 18840 14550
rect 18788 14486 18840 14492
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 18696 10668 18748 10674
rect 18696 10610 18748 10616
rect 18708 9722 18736 10610
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 18696 9716 18748 9722
rect 18696 9658 18748 9664
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19156 7948 19208 7954
rect 19156 7890 19208 7896
rect 19168 4146 19196 7890
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19798 5264 19854 5273
rect 19798 5199 19800 5208
rect 19852 5199 19854 5208
rect 19800 5170 19852 5176
rect 19984 5160 20036 5166
rect 19984 5102 20036 5108
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19890 4176 19946 4185
rect 19156 4140 19208 4146
rect 19156 4082 19208 4088
rect 19432 4140 19484 4146
rect 19890 4111 19946 4120
rect 19432 4082 19484 4088
rect 18696 3936 18748 3942
rect 18696 3878 18748 3884
rect 18708 3754 18736 3878
rect 18616 3726 18736 3754
rect 18512 3528 18564 3534
rect 18512 3470 18564 3476
rect 18616 3194 18644 3726
rect 18696 3460 18748 3466
rect 18696 3402 18748 3408
rect 18604 3188 18656 3194
rect 18604 3130 18656 3136
rect 18420 2440 18472 2446
rect 18420 2382 18472 2388
rect 18604 2372 18656 2378
rect 18604 2314 18656 2320
rect 18616 2106 18644 2314
rect 18604 2100 18656 2106
rect 18604 2042 18656 2048
rect 18708 950 18736 3402
rect 19444 3398 19472 4082
rect 19904 4010 19932 4111
rect 19892 4004 19944 4010
rect 19892 3946 19944 3952
rect 19432 3392 19484 3398
rect 19432 3334 19484 3340
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 19432 2984 19484 2990
rect 19432 2926 19484 2932
rect 19444 2650 19472 2926
rect 19432 2644 19484 2650
rect 19432 2586 19484 2592
rect 19340 2440 19392 2446
rect 19340 2382 19392 2388
rect 18880 1012 18932 1018
rect 18880 954 18932 960
rect 18604 944 18656 950
rect 18604 886 18656 892
rect 18696 944 18748 950
rect 18696 886 18748 892
rect 18616 800 18644 886
rect 18892 800 18920 954
rect 19352 898 19380 2382
rect 19432 2304 19484 2310
rect 19432 2246 19484 2252
rect 19168 870 19380 898
rect 19168 800 19196 870
rect 19444 800 19472 2246
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 19996 1986 20024 5102
rect 20088 2446 20116 16102
rect 20720 16050 20772 16056
rect 20352 16040 20404 16046
rect 20352 15982 20404 15988
rect 20628 16040 20680 16046
rect 20628 15982 20680 15988
rect 20166 15872 20222 15881
rect 20166 15807 20222 15816
rect 20180 3466 20208 15807
rect 20260 15360 20312 15366
rect 20260 15302 20312 15308
rect 20272 15026 20300 15302
rect 20364 15162 20392 15982
rect 20640 15434 20668 15982
rect 20732 15502 20760 16050
rect 20720 15496 20772 15502
rect 20720 15438 20772 15444
rect 20628 15428 20680 15434
rect 20628 15370 20680 15376
rect 20352 15156 20404 15162
rect 20352 15098 20404 15104
rect 20260 15020 20312 15026
rect 20260 14962 20312 14968
rect 20444 14340 20496 14346
rect 20444 14282 20496 14288
rect 20628 14340 20680 14346
rect 20628 14282 20680 14288
rect 20456 11082 20484 14282
rect 20536 13252 20588 13258
rect 20536 13194 20588 13200
rect 20444 11076 20496 11082
rect 20444 11018 20496 11024
rect 20548 8838 20576 13194
rect 20640 11354 20668 14282
rect 20732 14074 20760 15438
rect 20824 15162 20852 18702
rect 20904 18420 20956 18426
rect 20904 18362 20956 18368
rect 20812 15156 20864 15162
rect 20812 15098 20864 15104
rect 20720 14068 20772 14074
rect 20720 14010 20772 14016
rect 20812 12640 20864 12646
rect 20812 12582 20864 12588
rect 20718 12200 20774 12209
rect 20718 12135 20774 12144
rect 20732 11626 20760 12135
rect 20720 11620 20772 11626
rect 20720 11562 20772 11568
rect 20628 11348 20680 11354
rect 20628 11290 20680 11296
rect 20536 8832 20588 8838
rect 20536 8774 20588 8780
rect 20444 7336 20496 7342
rect 20444 7278 20496 7284
rect 20456 6730 20484 7278
rect 20444 6724 20496 6730
rect 20444 6666 20496 6672
rect 20456 6254 20484 6666
rect 20444 6248 20496 6254
rect 20444 6190 20496 6196
rect 20456 5710 20484 6190
rect 20444 5704 20496 5710
rect 20444 5646 20496 5652
rect 20352 5092 20404 5098
rect 20352 5034 20404 5040
rect 20364 4622 20392 5034
rect 20352 4616 20404 4622
rect 20352 4558 20404 4564
rect 20260 4548 20312 4554
rect 20260 4490 20312 4496
rect 20168 3460 20220 3466
rect 20168 3402 20220 3408
rect 20076 2440 20128 2446
rect 20076 2382 20128 2388
rect 19720 1958 20024 1986
rect 19720 800 19748 1958
rect 19984 1080 20036 1086
rect 19984 1022 20036 1028
rect 19996 800 20024 1022
rect 20272 800 20300 4490
rect 20456 4146 20484 5646
rect 20824 5234 20852 12582
rect 20812 5228 20864 5234
rect 20812 5170 20864 5176
rect 20916 4622 20944 18362
rect 21180 17672 21232 17678
rect 21180 17614 21232 17620
rect 21192 17338 21220 17614
rect 21364 17536 21416 17542
rect 21364 17478 21416 17484
rect 21180 17332 21232 17338
rect 21180 17274 21232 17280
rect 21376 17134 21404 17478
rect 21364 17128 21416 17134
rect 21364 17070 21416 17076
rect 21560 16658 21588 18702
rect 21640 17604 21692 17610
rect 21640 17546 21692 17552
rect 21548 16652 21600 16658
rect 21548 16594 21600 16600
rect 21364 15972 21416 15978
rect 21364 15914 21416 15920
rect 21180 15904 21232 15910
rect 21180 15846 21232 15852
rect 20996 15360 21048 15366
rect 20996 15302 21048 15308
rect 21008 15026 21036 15302
rect 20996 15020 21048 15026
rect 20996 14962 21048 14968
rect 21088 14816 21140 14822
rect 21088 14758 21140 14764
rect 21100 14414 21128 14758
rect 21088 14408 21140 14414
rect 21088 14350 21140 14356
rect 21192 8430 21220 15846
rect 21272 15564 21324 15570
rect 21272 15506 21324 15512
rect 21284 14550 21312 15506
rect 21272 14544 21324 14550
rect 21272 14486 21324 14492
rect 21376 13530 21404 15914
rect 21456 15496 21508 15502
rect 21456 15438 21508 15444
rect 21468 15162 21496 15438
rect 21652 15434 21680 17546
rect 21640 15428 21692 15434
rect 21640 15370 21692 15376
rect 21456 15156 21508 15162
rect 21456 15098 21508 15104
rect 21652 14550 21680 15370
rect 21744 14958 21772 18702
rect 22296 18290 22324 21490
rect 22468 21412 22520 21418
rect 22468 21354 22520 21360
rect 22480 20942 22508 21354
rect 22468 20936 22520 20942
rect 22468 20878 22520 20884
rect 22376 19848 22428 19854
rect 22376 19790 22428 19796
rect 22388 19514 22416 19790
rect 22376 19508 22428 19514
rect 22376 19450 22428 19456
rect 22284 18284 22336 18290
rect 22284 18226 22336 18232
rect 22756 17746 22784 22066
rect 23216 21622 23244 23802
rect 23308 23662 23336 24142
rect 23296 23656 23348 23662
rect 23296 23598 23348 23604
rect 23492 22098 23520 24618
rect 23676 24206 23704 24822
rect 23664 24200 23716 24206
rect 23664 24142 23716 24148
rect 23676 23730 23704 24142
rect 23664 23724 23716 23730
rect 23664 23666 23716 23672
rect 23848 23248 23900 23254
rect 23848 23190 23900 23196
rect 23480 22092 23532 22098
rect 23480 22034 23532 22040
rect 23294 21992 23350 22001
rect 23294 21927 23350 21936
rect 23204 21616 23256 21622
rect 23204 21558 23256 21564
rect 23216 21146 23244 21558
rect 23204 21140 23256 21146
rect 23204 21082 23256 21088
rect 23112 19916 23164 19922
rect 23112 19858 23164 19864
rect 23124 19378 23152 19858
rect 23112 19372 23164 19378
rect 23112 19314 23164 19320
rect 22928 19236 22980 19242
rect 22928 19178 22980 19184
rect 22744 17740 22796 17746
rect 22744 17682 22796 17688
rect 22652 17672 22704 17678
rect 22652 17614 22704 17620
rect 21914 17368 21970 17377
rect 21914 17303 21970 17312
rect 21732 14952 21784 14958
rect 21732 14894 21784 14900
rect 21640 14544 21692 14550
rect 21640 14486 21692 14492
rect 21364 13524 21416 13530
rect 21364 13466 21416 13472
rect 21456 13524 21508 13530
rect 21456 13466 21508 13472
rect 21180 8424 21232 8430
rect 21180 8366 21232 8372
rect 20996 8288 21048 8294
rect 20996 8230 21048 8236
rect 21008 7002 21036 8230
rect 20996 6996 21048 7002
rect 20996 6938 21048 6944
rect 21180 6928 21232 6934
rect 21180 6870 21232 6876
rect 20994 6488 21050 6497
rect 20994 6423 21050 6432
rect 20904 4616 20956 4622
rect 20904 4558 20956 4564
rect 20812 4548 20864 4554
rect 20812 4490 20864 4496
rect 20444 4140 20496 4146
rect 20444 4082 20496 4088
rect 20718 4040 20774 4049
rect 20444 4004 20496 4010
rect 20718 3975 20774 3984
rect 20444 3946 20496 3952
rect 20456 3738 20484 3946
rect 20732 3738 20760 3975
rect 20444 3732 20496 3738
rect 20444 3674 20496 3680
rect 20720 3732 20772 3738
rect 20720 3674 20772 3680
rect 20536 3528 20588 3534
rect 20536 3470 20588 3476
rect 20352 3460 20404 3466
rect 20352 3402 20404 3408
rect 20364 2990 20392 3402
rect 20444 3392 20496 3398
rect 20444 3334 20496 3340
rect 20352 2984 20404 2990
rect 20352 2926 20404 2932
rect 20456 1018 20484 3334
rect 20548 1086 20576 3470
rect 20824 2938 20852 4490
rect 20904 4480 20956 4486
rect 20902 4448 20904 4457
rect 20956 4448 20958 4457
rect 20902 4383 20958 4392
rect 20824 2910 20944 2938
rect 21008 2922 21036 6423
rect 21192 3670 21220 6870
rect 21272 5160 21324 5166
rect 21272 5102 21324 5108
rect 21180 3664 21232 3670
rect 21180 3606 21232 3612
rect 21180 3052 21232 3058
rect 21180 2994 21232 3000
rect 20812 2848 20864 2854
rect 20812 2790 20864 2796
rect 20824 2514 20852 2790
rect 20916 2774 20944 2910
rect 20996 2916 21048 2922
rect 20996 2858 21048 2864
rect 20916 2746 21128 2774
rect 20812 2508 20864 2514
rect 20812 2450 20864 2456
rect 20628 2032 20680 2038
rect 20628 1974 20680 1980
rect 20536 1080 20588 1086
rect 20536 1022 20588 1028
rect 20444 1012 20496 1018
rect 20444 954 20496 960
rect 20640 950 20668 1974
rect 20812 1012 20864 1018
rect 20812 954 20864 960
rect 20536 944 20588 950
rect 20536 886 20588 892
rect 20628 944 20680 950
rect 20628 886 20680 892
rect 20548 800 20576 886
rect 20824 800 20852 954
rect 21100 800 21128 2746
rect 21192 1018 21220 2994
rect 21284 2774 21312 5102
rect 21364 4548 21416 4554
rect 21364 4490 21416 4496
rect 21376 4214 21404 4490
rect 21364 4208 21416 4214
rect 21364 4150 21416 4156
rect 21468 3058 21496 13466
rect 21822 13152 21878 13161
rect 21822 13087 21878 13096
rect 21548 8424 21600 8430
rect 21548 8366 21600 8372
rect 21560 4010 21588 8366
rect 21732 5160 21784 5166
rect 21732 5102 21784 5108
rect 21744 4826 21772 5102
rect 21732 4820 21784 4826
rect 21732 4762 21784 4768
rect 21548 4004 21600 4010
rect 21548 3946 21600 3952
rect 21456 3052 21508 3058
rect 21456 2994 21508 3000
rect 21560 2922 21588 3946
rect 21548 2916 21600 2922
rect 21548 2858 21600 2864
rect 21284 2746 21404 2774
rect 21180 1012 21232 1018
rect 21180 954 21232 960
rect 21376 800 21404 2746
rect 21836 2446 21864 13087
rect 21928 3534 21956 17303
rect 22468 16992 22520 16998
rect 22468 16934 22520 16940
rect 22480 16590 22508 16934
rect 22468 16584 22520 16590
rect 22468 16526 22520 16532
rect 22284 16040 22336 16046
rect 22284 15982 22336 15988
rect 22192 15428 22244 15434
rect 22296 15416 22324 15982
rect 22376 15428 22428 15434
rect 22296 15388 22376 15416
rect 22192 15370 22244 15376
rect 22376 15370 22428 15376
rect 22008 14952 22060 14958
rect 22204 14940 22232 15370
rect 22468 15360 22520 15366
rect 22468 15302 22520 15308
rect 22560 15360 22612 15366
rect 22560 15302 22612 15308
rect 22376 14952 22428 14958
rect 22204 14912 22376 14940
rect 22008 14894 22060 14900
rect 22376 14894 22428 14900
rect 22020 10577 22048 14894
rect 22388 14482 22416 14894
rect 22284 14476 22336 14482
rect 22284 14418 22336 14424
rect 22376 14476 22428 14482
rect 22376 14418 22428 14424
rect 22296 14074 22324 14418
rect 22284 14068 22336 14074
rect 22284 14010 22336 14016
rect 22480 13938 22508 15302
rect 22192 13932 22244 13938
rect 22192 13874 22244 13880
rect 22468 13932 22520 13938
rect 22468 13874 22520 13880
rect 22100 13864 22152 13870
rect 22100 13806 22152 13812
rect 22112 10713 22140 13806
rect 22204 11286 22232 13874
rect 22572 13326 22600 15302
rect 22664 15094 22692 17614
rect 22940 17082 22968 19178
rect 23020 17128 23072 17134
rect 22940 17076 23020 17082
rect 22940 17070 23072 17076
rect 22940 17054 23060 17070
rect 22836 16584 22888 16590
rect 22836 16526 22888 16532
rect 22744 15428 22796 15434
rect 22744 15370 22796 15376
rect 22756 15094 22784 15370
rect 22652 15088 22704 15094
rect 22652 15030 22704 15036
rect 22744 15088 22796 15094
rect 22744 15030 22796 15036
rect 22664 14822 22692 15030
rect 22652 14816 22704 14822
rect 22652 14758 22704 14764
rect 22744 13796 22796 13802
rect 22744 13738 22796 13744
rect 22560 13320 22612 13326
rect 22560 13262 22612 13268
rect 22572 12442 22600 13262
rect 22756 12646 22784 13738
rect 22744 12640 22796 12646
rect 22744 12582 22796 12588
rect 22560 12436 22612 12442
rect 22560 12378 22612 12384
rect 22744 11824 22796 11830
rect 22744 11766 22796 11772
rect 22756 11665 22784 11766
rect 22742 11656 22798 11665
rect 22742 11591 22798 11600
rect 22192 11280 22244 11286
rect 22192 11222 22244 11228
rect 22098 10704 22154 10713
rect 22098 10639 22154 10648
rect 22006 10568 22062 10577
rect 22006 10503 22062 10512
rect 22744 9580 22796 9586
rect 22744 9522 22796 9528
rect 22098 9480 22154 9489
rect 22098 9415 22154 9424
rect 22112 8362 22140 9415
rect 22756 8786 22784 9522
rect 22848 8974 22876 16526
rect 22940 9058 22968 17054
rect 23112 16040 23164 16046
rect 23112 15982 23164 15988
rect 23124 15434 23152 15982
rect 23202 15736 23258 15745
rect 23202 15671 23204 15680
rect 23256 15671 23258 15680
rect 23204 15642 23256 15648
rect 23112 15428 23164 15434
rect 23112 15370 23164 15376
rect 23204 15020 23256 15026
rect 23204 14962 23256 14968
rect 23216 14822 23244 14962
rect 23204 14816 23256 14822
rect 23204 14758 23256 14764
rect 23216 14521 23244 14758
rect 23202 14512 23258 14521
rect 23202 14447 23258 14456
rect 23112 13456 23164 13462
rect 23112 13398 23164 13404
rect 23020 12912 23072 12918
rect 23020 12854 23072 12860
rect 23032 12374 23060 12854
rect 23020 12368 23072 12374
rect 23020 12310 23072 12316
rect 23032 11558 23060 12310
rect 23020 11552 23072 11558
rect 23020 11494 23072 11500
rect 23032 9586 23060 11494
rect 23020 9580 23072 9586
rect 23020 9522 23072 9528
rect 23018 9072 23074 9081
rect 22940 9030 23018 9058
rect 23018 9007 23074 9016
rect 23032 8974 23060 9007
rect 23124 8974 23152 13398
rect 23308 13274 23336 21927
rect 23492 21622 23520 22034
rect 23480 21616 23532 21622
rect 23480 21558 23532 21564
rect 23662 21040 23718 21049
rect 23662 20975 23718 20984
rect 23676 20534 23704 20975
rect 23756 20936 23808 20942
rect 23756 20878 23808 20884
rect 23664 20528 23716 20534
rect 23664 20470 23716 20476
rect 23676 20262 23704 20470
rect 23664 20256 23716 20262
rect 23664 20198 23716 20204
rect 23768 17610 23796 20878
rect 23756 17604 23808 17610
rect 23756 17546 23808 17552
rect 23860 17218 23888 23190
rect 23952 21894 23980 25910
rect 24032 25900 24084 25906
rect 24032 25842 24084 25848
rect 24044 24818 24072 25842
rect 24228 24954 24256 30194
rect 24308 28688 24360 28694
rect 24308 28630 24360 28636
rect 24320 28218 24348 28630
rect 24308 28212 24360 28218
rect 24308 28154 24360 28160
rect 24216 24948 24268 24954
rect 24216 24890 24268 24896
rect 24032 24812 24084 24818
rect 24032 24754 24084 24760
rect 24044 24070 24072 24754
rect 24308 24676 24360 24682
rect 24308 24618 24360 24624
rect 24032 24064 24084 24070
rect 24032 24006 24084 24012
rect 24044 23730 24072 24006
rect 24032 23724 24084 23730
rect 24032 23666 24084 23672
rect 23940 21888 23992 21894
rect 23940 21830 23992 21836
rect 23952 20534 23980 21830
rect 24044 21690 24072 23666
rect 24124 22704 24176 22710
rect 24124 22646 24176 22652
rect 24136 22030 24164 22646
rect 24320 22094 24348 24618
rect 24412 23866 24440 31726
rect 24688 31726 24808 31754
rect 24492 28960 24544 28966
rect 24492 28902 24544 28908
rect 24504 28082 24532 28902
rect 24584 28552 24636 28558
rect 24584 28494 24636 28500
rect 24492 28076 24544 28082
rect 24492 28018 24544 28024
rect 24504 26926 24532 28018
rect 24596 26994 24624 28494
rect 24584 26988 24636 26994
rect 24584 26930 24636 26936
rect 24492 26920 24544 26926
rect 24492 26862 24544 26868
rect 24596 26042 24624 26930
rect 24584 26036 24636 26042
rect 24584 25978 24636 25984
rect 24596 25838 24624 25978
rect 24584 25832 24636 25838
rect 24584 25774 24636 25780
rect 24688 25650 24716 31726
rect 24952 29096 25004 29102
rect 24952 29038 25004 29044
rect 24964 28082 24992 29038
rect 25504 28620 25556 28626
rect 25504 28562 25556 28568
rect 25412 28416 25464 28422
rect 25412 28358 25464 28364
rect 24952 28076 25004 28082
rect 24952 28018 25004 28024
rect 24964 27470 24992 28018
rect 25044 27940 25096 27946
rect 25044 27882 25096 27888
rect 24952 27464 25004 27470
rect 24952 27406 25004 27412
rect 24860 27328 24912 27334
rect 24860 27270 24912 27276
rect 24872 26994 24900 27270
rect 25056 27130 25084 27882
rect 25424 27470 25452 28358
rect 25516 28082 25544 28562
rect 25504 28076 25556 28082
rect 25504 28018 25556 28024
rect 25596 28076 25648 28082
rect 25596 28018 25648 28024
rect 25228 27464 25280 27470
rect 25228 27406 25280 27412
rect 25412 27464 25464 27470
rect 25412 27406 25464 27412
rect 25504 27464 25556 27470
rect 25504 27406 25556 27412
rect 25044 27124 25096 27130
rect 25044 27066 25096 27072
rect 25056 26994 25084 27066
rect 25240 26994 25268 27406
rect 25320 27124 25372 27130
rect 25320 27066 25372 27072
rect 24860 26988 24912 26994
rect 24860 26930 24912 26936
rect 25044 26988 25096 26994
rect 25044 26930 25096 26936
rect 25136 26988 25188 26994
rect 25136 26930 25188 26936
rect 25228 26988 25280 26994
rect 25228 26930 25280 26936
rect 24872 26314 24900 26930
rect 24952 26920 25004 26926
rect 25148 26874 25176 26930
rect 25004 26868 25176 26874
rect 24952 26862 25176 26868
rect 24964 26846 25176 26862
rect 24860 26308 24912 26314
rect 24860 26250 24912 26256
rect 24768 26240 24820 26246
rect 24768 26182 24820 26188
rect 24596 25622 24716 25650
rect 24596 25362 24624 25622
rect 24584 25356 24636 25362
rect 24584 25298 24636 25304
rect 24492 25288 24544 25294
rect 24492 25230 24544 25236
rect 24400 23860 24452 23866
rect 24400 23802 24452 23808
rect 24412 22642 24440 23802
rect 24400 22636 24452 22642
rect 24400 22578 24452 22584
rect 24320 22066 24440 22094
rect 24124 22024 24176 22030
rect 24124 21966 24176 21972
rect 24032 21684 24084 21690
rect 24032 21626 24084 21632
rect 24136 21026 24164 21966
rect 24044 20998 24164 21026
rect 23940 20528 23992 20534
rect 23940 20470 23992 20476
rect 24044 17542 24072 20998
rect 24124 20868 24176 20874
rect 24124 20810 24176 20816
rect 24136 19786 24164 20810
rect 24308 20596 24360 20602
rect 24308 20538 24360 20544
rect 24124 19780 24176 19786
rect 24124 19722 24176 19728
rect 24136 19378 24164 19722
rect 24124 19372 24176 19378
rect 24124 19314 24176 19320
rect 24320 18290 24348 20538
rect 24412 20466 24440 22066
rect 24504 21486 24532 25230
rect 24676 23316 24728 23322
rect 24676 23258 24728 23264
rect 24584 21548 24636 21554
rect 24584 21490 24636 21496
rect 24492 21480 24544 21486
rect 24492 21422 24544 21428
rect 24400 20460 24452 20466
rect 24400 20402 24452 20408
rect 24504 19854 24532 21422
rect 24492 19848 24544 19854
rect 24492 19790 24544 19796
rect 24400 19440 24452 19446
rect 24400 19382 24452 19388
rect 24412 18834 24440 19382
rect 24596 19378 24624 21490
rect 24688 20466 24716 23258
rect 24780 22710 24808 26182
rect 25148 24818 25176 26846
rect 25332 26364 25360 27066
rect 25424 26586 25452 27406
rect 25516 27062 25544 27406
rect 25608 27402 25636 28018
rect 25596 27396 25648 27402
rect 25596 27338 25648 27344
rect 25504 27056 25556 27062
rect 25504 26998 25556 27004
rect 25596 26852 25648 26858
rect 25596 26794 25648 26800
rect 25412 26580 25464 26586
rect 25412 26522 25464 26528
rect 25608 26382 25636 26794
rect 25412 26376 25464 26382
rect 25332 26336 25412 26364
rect 25412 26318 25464 26324
rect 25596 26376 25648 26382
rect 25596 26318 25648 26324
rect 25700 24818 25728 57190
rect 26148 43444 26200 43450
rect 26148 43386 26200 43392
rect 25872 28552 25924 28558
rect 25872 28494 25924 28500
rect 25884 28082 25912 28494
rect 25872 28076 25924 28082
rect 25872 28018 25924 28024
rect 26056 27940 26108 27946
rect 26056 27882 26108 27888
rect 26068 27334 26096 27882
rect 26056 27328 26108 27334
rect 26056 27270 26108 27276
rect 26054 27160 26110 27169
rect 26054 27095 26056 27104
rect 26108 27095 26110 27104
rect 26056 27066 26108 27072
rect 26160 27062 26188 43386
rect 26424 42016 26476 42022
rect 26424 41958 26476 41964
rect 26436 41614 26464 41958
rect 26712 41614 26740 57190
rect 26792 55888 26844 55894
rect 26792 55830 26844 55836
rect 26424 41608 26476 41614
rect 26424 41550 26476 41556
rect 26700 41608 26752 41614
rect 26700 41550 26752 41556
rect 26700 35284 26752 35290
rect 26700 35226 26752 35232
rect 26712 34542 26740 35226
rect 26700 34536 26752 34542
rect 26700 34478 26752 34484
rect 26240 30728 26292 30734
rect 26240 30670 26292 30676
rect 26252 30190 26280 30670
rect 26240 30184 26292 30190
rect 26240 30126 26292 30132
rect 26332 27600 26384 27606
rect 26332 27542 26384 27548
rect 26240 27396 26292 27402
rect 26240 27338 26292 27344
rect 26252 27130 26280 27338
rect 26344 27334 26372 27542
rect 26332 27328 26384 27334
rect 26332 27270 26384 27276
rect 26516 27328 26568 27334
rect 26516 27270 26568 27276
rect 26608 27328 26660 27334
rect 26608 27270 26660 27276
rect 26344 27130 26372 27270
rect 26240 27124 26292 27130
rect 26240 27066 26292 27072
rect 26332 27124 26384 27130
rect 26332 27066 26384 27072
rect 26424 27124 26476 27130
rect 26424 27066 26476 27072
rect 26148 27056 26200 27062
rect 26436 27033 26464 27066
rect 26148 26998 26200 27004
rect 26422 27024 26478 27033
rect 26422 26959 26478 26968
rect 26528 26382 26556 27270
rect 26620 26926 26648 27270
rect 26608 26920 26660 26926
rect 26608 26862 26660 26868
rect 26516 26376 26568 26382
rect 26516 26318 26568 26324
rect 26332 26308 26384 26314
rect 26332 26250 26384 26256
rect 26700 26308 26752 26314
rect 26700 26250 26752 26256
rect 26344 25702 26372 26250
rect 26332 25696 26384 25702
rect 26332 25638 26384 25644
rect 24860 24812 24912 24818
rect 24860 24754 24912 24760
rect 25136 24812 25188 24818
rect 25136 24754 25188 24760
rect 25688 24812 25740 24818
rect 25688 24754 25740 24760
rect 24768 22704 24820 22710
rect 24768 22646 24820 22652
rect 24872 21622 24900 24754
rect 26712 23254 26740 26250
rect 26700 23248 26752 23254
rect 26700 23190 26752 23196
rect 26608 22024 26660 22030
rect 26608 21966 26660 21972
rect 25228 21888 25280 21894
rect 25228 21830 25280 21836
rect 24860 21616 24912 21622
rect 24860 21558 24912 21564
rect 24872 21146 24900 21558
rect 24860 21140 24912 21146
rect 24860 21082 24912 21088
rect 25240 20942 25268 21830
rect 25412 21548 25464 21554
rect 25412 21490 25464 21496
rect 25424 21146 25452 21490
rect 26240 21344 26292 21350
rect 26240 21286 26292 21292
rect 25412 21140 25464 21146
rect 25412 21082 25464 21088
rect 25228 20936 25280 20942
rect 25228 20878 25280 20884
rect 26252 20874 26280 21286
rect 26240 20868 26292 20874
rect 26240 20810 26292 20816
rect 26332 20868 26384 20874
rect 26332 20810 26384 20816
rect 24676 20460 24728 20466
rect 24676 20402 24728 20408
rect 24676 20324 24728 20330
rect 24676 20266 24728 20272
rect 24688 19718 24716 20266
rect 26344 19854 26372 20810
rect 26620 20602 26648 21966
rect 26608 20596 26660 20602
rect 26608 20538 26660 20544
rect 24768 19848 24820 19854
rect 24768 19790 24820 19796
rect 25320 19848 25372 19854
rect 25320 19790 25372 19796
rect 26332 19848 26384 19854
rect 26332 19790 26384 19796
rect 24676 19712 24728 19718
rect 24676 19654 24728 19660
rect 24584 19372 24636 19378
rect 24584 19314 24636 19320
rect 24400 18828 24452 18834
rect 24400 18770 24452 18776
rect 24584 18760 24636 18766
rect 24584 18702 24636 18708
rect 24308 18284 24360 18290
rect 24308 18226 24360 18232
rect 24124 18080 24176 18086
rect 24124 18022 24176 18028
rect 24032 17536 24084 17542
rect 24032 17478 24084 17484
rect 24136 17338 24164 18022
rect 24216 17604 24268 17610
rect 24216 17546 24268 17552
rect 24124 17332 24176 17338
rect 24124 17274 24176 17280
rect 23572 17196 23624 17202
rect 23860 17190 24072 17218
rect 23572 17138 23624 17144
rect 23480 16992 23532 16998
rect 23480 16934 23532 16940
rect 23492 16130 23520 16934
rect 23584 16250 23612 17138
rect 23940 17128 23992 17134
rect 23940 17070 23992 17076
rect 23664 17060 23716 17066
rect 23664 17002 23716 17008
rect 23572 16244 23624 16250
rect 23572 16186 23624 16192
rect 23492 16102 23612 16130
rect 23388 15972 23440 15978
rect 23388 15914 23440 15920
rect 23400 15706 23428 15914
rect 23480 15904 23532 15910
rect 23480 15846 23532 15852
rect 23388 15700 23440 15706
rect 23388 15642 23440 15648
rect 23492 15502 23520 15846
rect 23480 15496 23532 15502
rect 23480 15438 23532 15444
rect 23584 15348 23612 16102
rect 23492 15320 23612 15348
rect 23386 14920 23442 14929
rect 23386 14855 23442 14864
rect 23400 14278 23428 14855
rect 23388 14272 23440 14278
rect 23388 14214 23440 14220
rect 23216 13246 23336 13274
rect 23216 10010 23244 13246
rect 23296 13184 23348 13190
rect 23296 13126 23348 13132
rect 23308 12986 23336 13126
rect 23296 12980 23348 12986
rect 23296 12922 23348 12928
rect 23388 12776 23440 12782
rect 23388 12718 23440 12724
rect 23294 12336 23350 12345
rect 23294 12271 23350 12280
rect 23308 11898 23336 12271
rect 23296 11892 23348 11898
rect 23296 11834 23348 11840
rect 23400 11354 23428 12718
rect 23492 12238 23520 15320
rect 23676 14278 23704 17002
rect 23848 16040 23900 16046
rect 23848 15982 23900 15988
rect 23756 15428 23808 15434
rect 23756 15370 23808 15376
rect 23664 14272 23716 14278
rect 23664 14214 23716 14220
rect 23572 13728 23624 13734
rect 23572 13670 23624 13676
rect 23480 12232 23532 12238
rect 23480 12174 23532 12180
rect 23478 12064 23534 12073
rect 23478 11999 23534 12008
rect 23388 11348 23440 11354
rect 23388 11290 23440 11296
rect 23388 10804 23440 10810
rect 23388 10746 23440 10752
rect 23400 10470 23428 10746
rect 23388 10464 23440 10470
rect 23388 10406 23440 10412
rect 23216 9982 23428 10010
rect 23296 9920 23348 9926
rect 23296 9862 23348 9868
rect 23204 9512 23256 9518
rect 23204 9454 23256 9460
rect 22836 8968 22888 8974
rect 22836 8910 22888 8916
rect 23020 8968 23072 8974
rect 23020 8910 23072 8916
rect 23112 8968 23164 8974
rect 23112 8910 23164 8916
rect 22756 8758 22876 8786
rect 22100 8356 22152 8362
rect 22100 8298 22152 8304
rect 22468 7744 22520 7750
rect 22468 7686 22520 7692
rect 22100 5024 22152 5030
rect 22100 4966 22152 4972
rect 22008 4752 22060 4758
rect 22006 4720 22008 4729
rect 22060 4720 22062 4729
rect 22006 4655 22062 4664
rect 22112 3670 22140 4966
rect 22284 4684 22336 4690
rect 22284 4626 22336 4632
rect 22296 4146 22324 4626
rect 22284 4140 22336 4146
rect 22284 4082 22336 4088
rect 22100 3664 22152 3670
rect 22100 3606 22152 3612
rect 21916 3528 21968 3534
rect 21916 3470 21968 3476
rect 21916 3188 21968 3194
rect 21916 3130 21968 3136
rect 21824 2440 21876 2446
rect 21824 2382 21876 2388
rect 21640 944 21692 950
rect 21640 886 21692 892
rect 21652 800 21680 886
rect 21928 800 21956 3130
rect 22100 3120 22152 3126
rect 22376 3120 22428 3126
rect 22152 3068 22376 3074
rect 22100 3062 22428 3068
rect 22112 3046 22416 3062
rect 22480 2394 22508 7686
rect 22848 5166 22876 8758
rect 23124 5914 23152 8910
rect 23216 8090 23244 9454
rect 23308 8634 23336 9862
rect 23296 8628 23348 8634
rect 23296 8570 23348 8576
rect 23204 8084 23256 8090
rect 23204 8026 23256 8032
rect 23112 5908 23164 5914
rect 23112 5850 23164 5856
rect 23124 5370 23152 5850
rect 23112 5364 23164 5370
rect 23112 5306 23164 5312
rect 22836 5160 22888 5166
rect 22836 5102 22888 5108
rect 23296 4684 23348 4690
rect 23296 4626 23348 4632
rect 23308 4486 23336 4626
rect 22560 4480 22612 4486
rect 22558 4448 22560 4457
rect 23296 4480 23348 4486
rect 22612 4448 22614 4457
rect 23296 4422 23348 4428
rect 22558 4383 22614 4392
rect 22928 4208 22980 4214
rect 22558 4176 22614 4185
rect 22928 4150 22980 4156
rect 22558 4111 22560 4120
rect 22612 4111 22614 4120
rect 22560 4082 22612 4088
rect 22836 3936 22888 3942
rect 22836 3878 22888 3884
rect 22560 3528 22612 3534
rect 22560 3470 22612 3476
rect 22572 3097 22600 3470
rect 22744 3460 22796 3466
rect 22744 3402 22796 3408
rect 22558 3088 22614 3097
rect 22558 3023 22614 3032
rect 22650 2952 22706 2961
rect 22650 2887 22706 2896
rect 22664 2854 22692 2887
rect 22756 2854 22784 3402
rect 22848 3233 22876 3878
rect 22834 3224 22890 3233
rect 22834 3159 22890 3168
rect 22836 2984 22888 2990
rect 22836 2926 22888 2932
rect 22652 2848 22704 2854
rect 22652 2790 22704 2796
rect 22744 2848 22796 2854
rect 22744 2790 22796 2796
rect 22388 2366 22508 2394
rect 22652 2440 22704 2446
rect 22652 2382 22704 2388
rect 22388 2106 22416 2366
rect 22468 2304 22520 2310
rect 22468 2246 22520 2252
rect 22376 2100 22428 2106
rect 22376 2042 22428 2048
rect 22192 1080 22244 1086
rect 22192 1022 22244 1028
rect 22204 800 22232 1022
rect 22480 800 22508 2246
rect 22664 1834 22692 2382
rect 22652 1828 22704 1834
rect 22652 1770 22704 1776
rect 22848 1562 22876 2926
rect 22940 2258 22968 4150
rect 23204 4072 23256 4078
rect 23204 4014 23256 4020
rect 23020 3664 23072 3670
rect 23020 3606 23072 3612
rect 23032 3466 23060 3606
rect 23020 3460 23072 3466
rect 23020 3402 23072 3408
rect 23112 3460 23164 3466
rect 23112 3402 23164 3408
rect 23124 3369 23152 3402
rect 23110 3360 23166 3369
rect 23110 3295 23166 3304
rect 22940 2230 23060 2258
rect 22836 1556 22888 1562
rect 22836 1498 22888 1504
rect 22744 1012 22796 1018
rect 22744 954 22796 960
rect 22756 800 22784 954
rect 23032 800 23060 2230
rect 23216 882 23244 4014
rect 23308 3398 23336 4422
rect 23296 3392 23348 3398
rect 23296 3334 23348 3340
rect 23400 3058 23428 9982
rect 23492 5098 23520 11999
rect 23584 10198 23612 13670
rect 23768 13394 23796 15370
rect 23756 13388 23808 13394
rect 23756 13330 23808 13336
rect 23664 13320 23716 13326
rect 23664 13262 23716 13268
rect 23676 12986 23704 13262
rect 23664 12980 23716 12986
rect 23664 12922 23716 12928
rect 23664 12436 23716 12442
rect 23664 12378 23716 12384
rect 23676 12238 23704 12378
rect 23664 12232 23716 12238
rect 23664 12174 23716 12180
rect 23676 11898 23704 12174
rect 23756 12096 23808 12102
rect 23756 12038 23808 12044
rect 23664 11892 23716 11898
rect 23664 11834 23716 11840
rect 23664 11008 23716 11014
rect 23664 10950 23716 10956
rect 23676 10538 23704 10950
rect 23768 10810 23796 12038
rect 23860 11370 23888 15982
rect 23952 15162 23980 17070
rect 23940 15156 23992 15162
rect 23940 15098 23992 15104
rect 23940 15020 23992 15026
rect 23940 14962 23992 14968
rect 23952 13938 23980 14962
rect 23940 13932 23992 13938
rect 23940 13874 23992 13880
rect 23952 12442 23980 13874
rect 23940 12436 23992 12442
rect 23940 12378 23992 12384
rect 23940 12096 23992 12102
rect 23940 12038 23992 12044
rect 23952 11830 23980 12038
rect 23940 11824 23992 11830
rect 23940 11766 23992 11772
rect 23860 11342 23980 11370
rect 23848 11212 23900 11218
rect 23848 11154 23900 11160
rect 23860 11082 23888 11154
rect 23848 11076 23900 11082
rect 23848 11018 23900 11024
rect 23952 10962 23980 11342
rect 23860 10934 23980 10962
rect 23756 10804 23808 10810
rect 23756 10746 23808 10752
rect 23664 10532 23716 10538
rect 23664 10474 23716 10480
rect 23572 10192 23624 10198
rect 23572 10134 23624 10140
rect 23584 9654 23612 10134
rect 23572 9648 23624 9654
rect 23572 9590 23624 9596
rect 23584 9042 23612 9590
rect 23572 9036 23624 9042
rect 23572 8978 23624 8984
rect 23676 8922 23704 10474
rect 23584 8894 23704 8922
rect 23584 7954 23612 8894
rect 23572 7948 23624 7954
rect 23572 7890 23624 7896
rect 23480 5092 23532 5098
rect 23480 5034 23532 5040
rect 23584 4554 23612 7890
rect 23572 4548 23624 4554
rect 23572 4490 23624 4496
rect 23584 4078 23612 4490
rect 23572 4072 23624 4078
rect 23572 4014 23624 4020
rect 23480 3596 23532 3602
rect 23480 3538 23532 3544
rect 23388 3052 23440 3058
rect 23388 2994 23440 3000
rect 23296 2440 23348 2446
rect 23296 2382 23348 2388
rect 23204 876 23256 882
rect 23204 818 23256 824
rect 23308 800 23336 2382
rect 23492 1714 23520 3538
rect 23584 2961 23612 4014
rect 23756 3936 23808 3942
rect 23756 3878 23808 3884
rect 23768 3194 23796 3878
rect 23860 3670 23888 10934
rect 23940 10600 23992 10606
rect 23940 10542 23992 10548
rect 23952 10266 23980 10542
rect 23940 10260 23992 10266
rect 23940 10202 23992 10208
rect 24044 4010 24072 17190
rect 24124 17196 24176 17202
rect 24124 17138 24176 17144
rect 24136 16114 24164 17138
rect 24124 16108 24176 16114
rect 24124 16050 24176 16056
rect 24124 15156 24176 15162
rect 24124 15098 24176 15104
rect 24136 14822 24164 15098
rect 24124 14816 24176 14822
rect 24124 14758 24176 14764
rect 24124 14000 24176 14006
rect 24124 13942 24176 13948
rect 24136 13462 24164 13942
rect 24228 13734 24256 17546
rect 24320 17202 24348 18226
rect 24400 18216 24452 18222
rect 24400 18158 24452 18164
rect 24308 17196 24360 17202
rect 24308 17138 24360 17144
rect 24412 16114 24440 18158
rect 24596 17678 24624 18702
rect 24688 17814 24716 19654
rect 24780 18902 24808 19790
rect 25332 19378 25360 19790
rect 25504 19780 25556 19786
rect 25504 19722 25556 19728
rect 25320 19372 25372 19378
rect 25320 19314 25372 19320
rect 24768 18896 24820 18902
rect 24768 18838 24820 18844
rect 24860 18692 24912 18698
rect 24860 18634 24912 18640
rect 24768 18216 24820 18222
rect 24768 18158 24820 18164
rect 24780 18086 24808 18158
rect 24768 18080 24820 18086
rect 24768 18022 24820 18028
rect 24676 17808 24728 17814
rect 24676 17750 24728 17756
rect 24584 17672 24636 17678
rect 24584 17614 24636 17620
rect 24768 17672 24820 17678
rect 24768 17614 24820 17620
rect 24490 17232 24546 17241
rect 24596 17202 24624 17614
rect 24780 17542 24808 17614
rect 24768 17536 24820 17542
rect 24768 17478 24820 17484
rect 24780 17338 24808 17478
rect 24768 17332 24820 17338
rect 24768 17274 24820 17280
rect 24490 17167 24546 17176
rect 24584 17196 24636 17202
rect 24400 16108 24452 16114
rect 24400 16050 24452 16056
rect 24308 16040 24360 16046
rect 24308 15982 24360 15988
rect 24320 13870 24348 15982
rect 24504 15348 24532 17167
rect 24584 17138 24636 17144
rect 24872 16590 24900 18634
rect 25044 16788 25096 16794
rect 25044 16730 25096 16736
rect 24860 16584 24912 16590
rect 24860 16526 24912 16532
rect 24768 16448 24820 16454
rect 24768 16390 24820 16396
rect 24412 15320 24532 15348
rect 24308 13864 24360 13870
rect 24308 13806 24360 13812
rect 24412 13818 24440 15320
rect 24674 15192 24730 15201
rect 24674 15127 24730 15136
rect 24584 15088 24636 15094
rect 24584 15030 24636 15036
rect 24492 14816 24544 14822
rect 24492 14758 24544 14764
rect 24504 13938 24532 14758
rect 24596 14618 24624 15030
rect 24688 14890 24716 15127
rect 24676 14884 24728 14890
rect 24676 14826 24728 14832
rect 24584 14612 24636 14618
rect 24584 14554 24636 14560
rect 24492 13932 24544 13938
rect 24492 13874 24544 13880
rect 24412 13790 24716 13818
rect 24216 13728 24268 13734
rect 24216 13670 24268 13676
rect 24124 13456 24176 13462
rect 24124 13398 24176 13404
rect 24584 13388 24636 13394
rect 24584 13330 24636 13336
rect 24596 12918 24624 13330
rect 24584 12912 24636 12918
rect 24584 12854 24636 12860
rect 24596 12306 24624 12854
rect 24584 12300 24636 12306
rect 24584 12242 24636 12248
rect 24584 10056 24636 10062
rect 24584 9998 24636 10004
rect 24596 9654 24624 9998
rect 24584 9648 24636 9654
rect 24584 9590 24636 9596
rect 24308 9376 24360 9382
rect 24308 9318 24360 9324
rect 24320 9178 24348 9318
rect 24308 9172 24360 9178
rect 24308 9114 24360 9120
rect 24214 8936 24270 8945
rect 24214 8871 24270 8880
rect 24124 8492 24176 8498
rect 24124 8434 24176 8440
rect 24136 7410 24164 8434
rect 24124 7404 24176 7410
rect 24124 7346 24176 7352
rect 24124 5228 24176 5234
rect 24124 5170 24176 5176
rect 24136 4690 24164 5170
rect 24124 4684 24176 4690
rect 24124 4626 24176 4632
rect 24032 4004 24084 4010
rect 24032 3946 24084 3952
rect 23848 3664 23900 3670
rect 23848 3606 23900 3612
rect 23940 3392 23992 3398
rect 23940 3334 23992 3340
rect 23756 3188 23808 3194
rect 23756 3130 23808 3136
rect 23952 3126 23980 3334
rect 23940 3120 23992 3126
rect 23940 3062 23992 3068
rect 23756 2984 23808 2990
rect 23570 2952 23626 2961
rect 23756 2926 23808 2932
rect 23570 2887 23626 2896
rect 23572 2440 23624 2446
rect 23572 2382 23624 2388
rect 23584 2038 23612 2382
rect 23572 2032 23624 2038
rect 23572 1974 23624 1980
rect 23492 1686 23612 1714
rect 23584 800 23612 1686
rect 23768 1018 23796 2926
rect 24228 2922 24256 8871
rect 24596 8566 24624 9590
rect 24584 8560 24636 8566
rect 24584 8502 24636 8508
rect 24688 8276 24716 13790
rect 24780 12442 24808 16390
rect 24872 14006 24900 16526
rect 25056 15978 25084 16730
rect 25332 16590 25360 19314
rect 25516 16658 25544 19722
rect 26424 18964 26476 18970
rect 26424 18906 26476 18912
rect 26332 18624 26384 18630
rect 26332 18566 26384 18572
rect 26344 18290 26372 18566
rect 26332 18284 26384 18290
rect 26332 18226 26384 18232
rect 26148 17672 26200 17678
rect 26148 17614 26200 17620
rect 26240 17672 26292 17678
rect 26240 17614 26292 17620
rect 25872 17536 25924 17542
rect 25872 17478 25924 17484
rect 25688 17196 25740 17202
rect 25688 17138 25740 17144
rect 25504 16652 25556 16658
rect 25424 16612 25504 16640
rect 25320 16584 25372 16590
rect 25320 16526 25372 16532
rect 24952 15972 25004 15978
rect 24952 15914 25004 15920
rect 25044 15972 25096 15978
rect 25044 15914 25096 15920
rect 24964 14618 24992 15914
rect 25056 15706 25084 15914
rect 25044 15700 25096 15706
rect 25044 15642 25096 15648
rect 25044 15564 25096 15570
rect 25044 15506 25096 15512
rect 25056 15042 25084 15506
rect 25056 15014 25268 15042
rect 24952 14612 25004 14618
rect 24952 14554 25004 14560
rect 24950 14512 25006 14521
rect 24950 14447 25006 14456
rect 24860 14000 24912 14006
rect 24860 13942 24912 13948
rect 24768 12436 24820 12442
rect 24768 12378 24820 12384
rect 24964 11898 24992 14447
rect 25056 14414 25084 15014
rect 25136 14952 25188 14958
rect 25136 14894 25188 14900
rect 25044 14408 25096 14414
rect 25044 14350 25096 14356
rect 25148 12850 25176 14894
rect 25240 14346 25268 15014
rect 25332 14958 25360 16526
rect 25424 15026 25452 16612
rect 25504 16594 25556 16600
rect 25700 16590 25728 17138
rect 25780 17128 25832 17134
rect 25780 17070 25832 17076
rect 25688 16584 25740 16590
rect 25688 16526 25740 16532
rect 25596 16516 25648 16522
rect 25596 16458 25648 16464
rect 25504 16040 25556 16046
rect 25504 15982 25556 15988
rect 25516 15434 25544 15982
rect 25608 15706 25636 16458
rect 25596 15700 25648 15706
rect 25596 15642 25648 15648
rect 25504 15428 25556 15434
rect 25504 15370 25556 15376
rect 25412 15020 25464 15026
rect 25412 14962 25464 14968
rect 25700 14958 25728 16526
rect 25792 15008 25820 17070
rect 25884 16538 25912 17478
rect 26160 17134 26188 17614
rect 26252 17542 26280 17614
rect 26240 17536 26292 17542
rect 26240 17478 26292 17484
rect 26148 17128 26200 17134
rect 26148 17070 26200 17076
rect 26332 16992 26384 16998
rect 26332 16934 26384 16940
rect 26344 16590 26372 16934
rect 26332 16584 26384 16590
rect 25884 16510 26096 16538
rect 26332 16526 26384 16532
rect 25872 16448 25924 16454
rect 25872 16390 25924 16396
rect 25884 16182 25912 16390
rect 25872 16176 25924 16182
rect 25872 16118 25924 16124
rect 25964 16040 26016 16046
rect 25964 15982 26016 15988
rect 25872 15020 25924 15026
rect 25792 14980 25872 15008
rect 25872 14962 25924 14968
rect 25320 14952 25372 14958
rect 25320 14894 25372 14900
rect 25688 14952 25740 14958
rect 25688 14894 25740 14900
rect 25228 14340 25280 14346
rect 25228 14282 25280 14288
rect 25228 13932 25280 13938
rect 25228 13874 25280 13880
rect 25240 13394 25268 13874
rect 25228 13388 25280 13394
rect 25228 13330 25280 13336
rect 25332 13190 25360 14894
rect 25884 14890 25912 14962
rect 25872 14884 25924 14890
rect 25872 14826 25924 14832
rect 25412 14476 25464 14482
rect 25412 14418 25464 14424
rect 25320 13184 25372 13190
rect 25320 13126 25372 13132
rect 25136 12844 25188 12850
rect 25136 12786 25188 12792
rect 25424 11898 25452 14418
rect 25884 12782 25912 14826
rect 25976 14006 26004 15982
rect 25964 14000 26016 14006
rect 25964 13942 26016 13948
rect 25964 12844 26016 12850
rect 25964 12786 26016 12792
rect 25872 12776 25924 12782
rect 25872 12718 25924 12724
rect 25872 12640 25924 12646
rect 25872 12582 25924 12588
rect 24952 11892 25004 11898
rect 24952 11834 25004 11840
rect 25412 11892 25464 11898
rect 25412 11834 25464 11840
rect 25136 11756 25188 11762
rect 25136 11698 25188 11704
rect 25148 9178 25176 11698
rect 25412 10668 25464 10674
rect 25412 10610 25464 10616
rect 25320 10464 25372 10470
rect 25320 10406 25372 10412
rect 25332 10062 25360 10406
rect 25320 10056 25372 10062
rect 25320 9998 25372 10004
rect 25228 9988 25280 9994
rect 25228 9930 25280 9936
rect 25240 9722 25268 9930
rect 25228 9716 25280 9722
rect 25228 9658 25280 9664
rect 25136 9172 25188 9178
rect 25136 9114 25188 9120
rect 25424 8974 25452 10610
rect 25780 10600 25832 10606
rect 25780 10542 25832 10548
rect 25792 9926 25820 10542
rect 25780 9920 25832 9926
rect 25780 9862 25832 9868
rect 25884 9110 25912 12582
rect 25976 12434 26004 12786
rect 26068 12646 26096 16510
rect 26148 15360 26200 15366
rect 26148 15302 26200 15308
rect 26160 12986 26188 15302
rect 26240 14272 26292 14278
rect 26240 14214 26292 14220
rect 26252 13938 26280 14214
rect 26332 14068 26384 14074
rect 26332 14010 26384 14016
rect 26240 13932 26292 13938
rect 26240 13874 26292 13880
rect 26344 13870 26372 14010
rect 26332 13864 26384 13870
rect 26332 13806 26384 13812
rect 26148 12980 26200 12986
rect 26148 12922 26200 12928
rect 26056 12640 26108 12646
rect 26056 12582 26108 12588
rect 25976 12406 26096 12434
rect 25964 10600 26016 10606
rect 25964 10542 26016 10548
rect 25976 10130 26004 10542
rect 26068 10198 26096 12406
rect 26148 12232 26200 12238
rect 26148 12174 26200 12180
rect 26056 10192 26108 10198
rect 26056 10134 26108 10140
rect 25964 10124 26016 10130
rect 25964 10066 26016 10072
rect 26160 9450 26188 12174
rect 26332 9580 26384 9586
rect 26332 9522 26384 9528
rect 26344 9489 26372 9522
rect 26330 9480 26386 9489
rect 26148 9444 26200 9450
rect 26330 9415 26386 9424
rect 26148 9386 26200 9392
rect 25872 9104 25924 9110
rect 25872 9046 25924 9052
rect 25688 9036 25740 9042
rect 25688 8978 25740 8984
rect 25412 8968 25464 8974
rect 25412 8910 25464 8916
rect 25044 8832 25096 8838
rect 25044 8774 25096 8780
rect 25596 8832 25648 8838
rect 25596 8774 25648 8780
rect 24768 8560 24820 8566
rect 24768 8502 24820 8508
rect 24504 8248 24716 8276
rect 24308 5364 24360 5370
rect 24308 5306 24360 5312
rect 24320 4758 24348 5306
rect 24308 4752 24360 4758
rect 24308 4694 24360 4700
rect 24504 4146 24532 8248
rect 24584 6112 24636 6118
rect 24584 6054 24636 6060
rect 24676 6112 24728 6118
rect 24676 6054 24728 6060
rect 24596 5914 24624 6054
rect 24584 5908 24636 5914
rect 24584 5850 24636 5856
rect 24688 5302 24716 6054
rect 24780 5846 24808 8502
rect 25056 8498 25084 8774
rect 25044 8492 25096 8498
rect 25044 8434 25096 8440
rect 25608 8362 25636 8774
rect 25596 8356 25648 8362
rect 25596 8298 25648 8304
rect 25608 7818 25636 8298
rect 25596 7812 25648 7818
rect 25596 7754 25648 7760
rect 24952 7404 25004 7410
rect 24952 7346 25004 7352
rect 24964 7002 24992 7346
rect 25044 7200 25096 7206
rect 25044 7142 25096 7148
rect 25136 7200 25188 7206
rect 25136 7142 25188 7148
rect 24952 6996 25004 7002
rect 24952 6938 25004 6944
rect 24768 5840 24820 5846
rect 24768 5782 24820 5788
rect 24768 5636 24820 5642
rect 24768 5578 24820 5584
rect 24676 5296 24728 5302
rect 24676 5238 24728 5244
rect 24584 4616 24636 4622
rect 24584 4558 24636 4564
rect 24492 4140 24544 4146
rect 24492 4082 24544 4088
rect 24596 4010 24624 4558
rect 24780 4486 24808 5578
rect 25056 5370 25084 7142
rect 25148 6730 25176 7142
rect 25700 6866 25728 8978
rect 26436 8974 26464 18906
rect 26700 18216 26752 18222
rect 26700 18158 26752 18164
rect 26608 17604 26660 17610
rect 26608 17546 26660 17552
rect 26516 17536 26568 17542
rect 26516 17478 26568 17484
rect 26528 16658 26556 17478
rect 26620 17202 26648 17546
rect 26608 17196 26660 17202
rect 26608 17138 26660 17144
rect 26712 16658 26740 18158
rect 26804 17134 26832 55830
rect 26896 18193 26924 57326
rect 52644 57316 52696 57322
rect 52644 57258 52696 57264
rect 56692 57316 56744 57322
rect 56692 57258 56744 57264
rect 27988 57248 28040 57254
rect 27988 57190 28040 57196
rect 29920 57248 29972 57254
rect 29920 57190 29972 57196
rect 30840 57248 30892 57254
rect 30840 57190 30892 57196
rect 31208 57248 31260 57254
rect 31208 57190 31260 57196
rect 33416 57248 33468 57254
rect 33416 57190 33468 57196
rect 34796 57248 34848 57254
rect 34796 57190 34848 57196
rect 35624 57248 35676 57254
rect 35624 57190 35676 57196
rect 37096 57248 37148 57254
rect 37096 57190 37148 57196
rect 37924 57248 37976 57254
rect 37924 57190 37976 57196
rect 39304 57248 39356 57254
rect 39304 57190 39356 57196
rect 40316 57248 40368 57254
rect 40316 57190 40368 57196
rect 41696 57248 41748 57254
rect 41696 57190 41748 57196
rect 43628 57248 43680 57254
rect 43628 57190 43680 57196
rect 45376 57248 45428 57254
rect 45376 57190 45428 57196
rect 46296 57248 46348 57254
rect 46296 57190 46348 57196
rect 46388 57248 46440 57254
rect 46388 57190 46440 57196
rect 48872 57248 48924 57254
rect 48872 57190 48924 57196
rect 49056 57248 49108 57254
rect 49056 57190 49108 57196
rect 51448 57248 51500 57254
rect 51448 57190 51500 57196
rect 51724 57248 51776 57254
rect 51724 57190 51776 57196
rect 28000 55214 28028 57190
rect 28000 55186 28212 55214
rect 26976 46368 27028 46374
rect 26976 46310 27028 46316
rect 26988 45966 27016 46310
rect 26976 45960 27028 45966
rect 26976 45902 27028 45908
rect 26976 44192 27028 44198
rect 26976 44134 27028 44140
rect 26988 31890 27016 44134
rect 27896 42560 27948 42566
rect 27896 42502 27948 42508
rect 27908 42226 27936 42502
rect 28184 42294 28212 55186
rect 29932 51074 29960 57190
rect 30472 56908 30524 56914
rect 30472 56850 30524 56856
rect 29932 51046 30052 51074
rect 28356 49088 28408 49094
rect 28356 49030 28408 49036
rect 28080 42288 28132 42294
rect 28080 42230 28132 42236
rect 28172 42288 28224 42294
rect 28172 42230 28224 42236
rect 27896 42220 27948 42226
rect 27896 42162 27948 42168
rect 28092 41546 28120 42230
rect 28264 42220 28316 42226
rect 28264 42162 28316 42168
rect 28276 41614 28304 42162
rect 28264 41608 28316 41614
rect 28264 41550 28316 41556
rect 28080 41540 28132 41546
rect 28080 41482 28132 41488
rect 27160 38344 27212 38350
rect 27160 38286 27212 38292
rect 26976 31884 27028 31890
rect 26976 31826 27028 31832
rect 26976 27464 27028 27470
rect 26974 27432 26976 27441
rect 27068 27464 27120 27470
rect 27028 27432 27030 27441
rect 27068 27406 27120 27412
rect 26974 27367 27030 27376
rect 26988 27062 27016 27367
rect 26976 27056 27028 27062
rect 26976 26998 27028 27004
rect 27080 26858 27108 27406
rect 27068 26852 27120 26858
rect 27068 26794 27120 26800
rect 27172 25294 27200 38286
rect 27804 36168 27856 36174
rect 27804 36110 27856 36116
rect 27712 32836 27764 32842
rect 27712 32778 27764 32784
rect 27618 32464 27674 32473
rect 27618 32399 27674 32408
rect 27632 32366 27660 32399
rect 27620 32360 27672 32366
rect 27620 32302 27672 32308
rect 27620 32020 27672 32026
rect 27620 31962 27672 31968
rect 27632 30938 27660 31962
rect 27724 31822 27752 32778
rect 27816 32337 27844 36110
rect 27988 35488 28040 35494
rect 27988 35430 28040 35436
rect 27896 32428 27948 32434
rect 27896 32370 27948 32376
rect 27802 32328 27858 32337
rect 27802 32263 27858 32272
rect 27712 31816 27764 31822
rect 27712 31758 27764 31764
rect 27620 30932 27672 30938
rect 27620 30874 27672 30880
rect 27724 30598 27752 31758
rect 27712 30592 27764 30598
rect 27712 30534 27764 30540
rect 27344 28008 27396 28014
rect 27344 27950 27396 27956
rect 27528 28008 27580 28014
rect 27528 27950 27580 27956
rect 27356 27606 27384 27950
rect 27344 27600 27396 27606
rect 27344 27542 27396 27548
rect 27540 25294 27568 27950
rect 27712 27464 27764 27470
rect 27712 27406 27764 27412
rect 27724 27062 27752 27406
rect 27712 27056 27764 27062
rect 27712 26998 27764 27004
rect 27712 25832 27764 25838
rect 27712 25774 27764 25780
rect 27724 25362 27752 25774
rect 27712 25356 27764 25362
rect 27712 25298 27764 25304
rect 27160 25288 27212 25294
rect 27160 25230 27212 25236
rect 27528 25288 27580 25294
rect 27528 25230 27580 25236
rect 27620 25288 27672 25294
rect 27620 25230 27672 25236
rect 27436 25220 27488 25226
rect 27436 25162 27488 25168
rect 27344 21344 27396 21350
rect 27344 21286 27396 21292
rect 27356 21146 27384 21286
rect 27344 21140 27396 21146
rect 27344 21082 27396 21088
rect 27068 19780 27120 19786
rect 27068 19722 27120 19728
rect 27080 18970 27108 19722
rect 27068 18964 27120 18970
rect 27068 18906 27120 18912
rect 26882 18184 26938 18193
rect 26882 18119 26938 18128
rect 26884 18080 26936 18086
rect 26884 18022 26936 18028
rect 26792 17128 26844 17134
rect 26792 17070 26844 17076
rect 26896 16946 26924 18022
rect 26804 16918 26924 16946
rect 27160 16992 27212 16998
rect 27160 16934 27212 16940
rect 27252 16992 27304 16998
rect 27252 16934 27304 16940
rect 26516 16652 26568 16658
rect 26516 16594 26568 16600
rect 26700 16652 26752 16658
rect 26700 16594 26752 16600
rect 26700 15428 26752 15434
rect 26700 15370 26752 15376
rect 26516 14952 26568 14958
rect 26516 14894 26568 14900
rect 26528 14414 26556 14894
rect 26516 14408 26568 14414
rect 26516 14350 26568 14356
rect 26608 14408 26660 14414
rect 26608 14350 26660 14356
rect 26528 12986 26556 14350
rect 26620 14074 26648 14350
rect 26608 14068 26660 14074
rect 26608 14010 26660 14016
rect 26516 12980 26568 12986
rect 26516 12922 26568 12928
rect 26620 9382 26648 14010
rect 26608 9376 26660 9382
rect 26608 9318 26660 9324
rect 26424 8968 26476 8974
rect 26424 8910 26476 8916
rect 25688 6860 25740 6866
rect 25688 6802 25740 6808
rect 25136 6724 25188 6730
rect 25136 6666 25188 6672
rect 25148 6390 25176 6666
rect 25136 6384 25188 6390
rect 25228 6384 25280 6390
rect 25136 6326 25188 6332
rect 25226 6352 25228 6361
rect 25280 6352 25282 6361
rect 25226 6287 25282 6296
rect 25700 6254 25728 6802
rect 26056 6316 26108 6322
rect 26056 6258 26108 6264
rect 25320 6248 25372 6254
rect 25688 6248 25740 6254
rect 25320 6190 25372 6196
rect 25686 6216 25688 6225
rect 25740 6216 25742 6225
rect 25332 5778 25360 6190
rect 25742 6174 25820 6202
rect 25686 6151 25742 6160
rect 25688 6112 25740 6118
rect 25688 6054 25740 6060
rect 25320 5772 25372 5778
rect 25320 5714 25372 5720
rect 25332 5370 25360 5714
rect 25700 5642 25728 6054
rect 25688 5636 25740 5642
rect 25688 5578 25740 5584
rect 25044 5364 25096 5370
rect 25044 5306 25096 5312
rect 25320 5364 25372 5370
rect 25320 5306 25372 5312
rect 24860 5024 24912 5030
rect 24860 4966 24912 4972
rect 25044 5024 25096 5030
rect 25044 4966 25096 4972
rect 24872 4622 24900 4966
rect 24860 4616 24912 4622
rect 24860 4558 24912 4564
rect 24768 4480 24820 4486
rect 24768 4422 24820 4428
rect 25056 4282 25084 4966
rect 25596 4752 25648 4758
rect 25594 4720 25596 4729
rect 25648 4720 25650 4729
rect 25594 4655 25650 4664
rect 25044 4276 25096 4282
rect 25044 4218 25096 4224
rect 25228 4276 25280 4282
rect 25228 4218 25280 4224
rect 24676 4140 24728 4146
rect 24676 4082 24728 4088
rect 24584 4004 24636 4010
rect 24584 3946 24636 3952
rect 24492 3052 24544 3058
rect 24596 3040 24624 3946
rect 24544 3012 24624 3040
rect 24492 2994 24544 3000
rect 24216 2916 24268 2922
rect 24216 2858 24268 2864
rect 24124 2508 24176 2514
rect 24124 2450 24176 2456
rect 23756 1012 23808 1018
rect 23756 954 23808 960
rect 23768 882 23888 898
rect 23756 876 23888 882
rect 23808 870 23888 876
rect 23756 818 23808 824
rect 23860 800 23888 870
rect 24136 800 24164 2450
rect 24400 1556 24452 1562
rect 24400 1498 24452 1504
rect 24412 800 24440 1498
rect 24688 800 24716 4082
rect 24950 3632 25006 3641
rect 24950 3567 25006 3576
rect 24964 3534 24992 3567
rect 24952 3528 25004 3534
rect 24952 3470 25004 3476
rect 25240 3126 25268 4218
rect 25792 4214 25820 6174
rect 25872 5636 25924 5642
rect 25872 5578 25924 5584
rect 25780 4208 25832 4214
rect 25780 4150 25832 4156
rect 25792 4078 25820 4150
rect 25688 4072 25740 4078
rect 25688 4014 25740 4020
rect 25780 4072 25832 4078
rect 25780 4014 25832 4020
rect 25320 3664 25372 3670
rect 25320 3606 25372 3612
rect 25332 3126 25360 3606
rect 25700 3369 25728 4014
rect 25884 4010 25912 5578
rect 26068 5302 26096 6258
rect 26332 6248 26384 6254
rect 26332 6190 26384 6196
rect 26344 5370 26372 6190
rect 26436 5642 26464 8910
rect 26608 8288 26660 8294
rect 26608 8230 26660 8236
rect 26620 8022 26648 8230
rect 26608 8016 26660 8022
rect 26608 7958 26660 7964
rect 26424 5636 26476 5642
rect 26424 5578 26476 5584
rect 26712 5522 26740 15370
rect 26804 11665 26832 16918
rect 27172 16658 27200 16934
rect 27264 16794 27292 16934
rect 27252 16788 27304 16794
rect 27252 16730 27304 16736
rect 27160 16652 27212 16658
rect 27160 16594 27212 16600
rect 27252 16516 27304 16522
rect 27252 16458 27304 16464
rect 27068 14884 27120 14890
rect 27068 14826 27120 14832
rect 26884 14476 26936 14482
rect 26884 14418 26936 14424
rect 26896 13394 26924 14418
rect 26884 13388 26936 13394
rect 26884 13330 26936 13336
rect 26896 13274 26924 13330
rect 26896 13246 27016 13274
rect 26884 12980 26936 12986
rect 26884 12922 26936 12928
rect 26790 11656 26846 11665
rect 26790 11591 26846 11600
rect 26792 8288 26844 8294
rect 26792 8230 26844 8236
rect 26804 8090 26832 8230
rect 26792 8084 26844 8090
rect 26792 8026 26844 8032
rect 26792 6248 26844 6254
rect 26792 6190 26844 6196
rect 26804 5914 26832 6190
rect 26792 5908 26844 5914
rect 26792 5850 26844 5856
rect 26436 5494 26740 5522
rect 26436 5370 26464 5494
rect 26332 5364 26384 5370
rect 26332 5306 26384 5312
rect 26424 5364 26476 5370
rect 26424 5306 26476 5312
rect 26056 5296 26108 5302
rect 26056 5238 26108 5244
rect 26608 5228 26660 5234
rect 26608 5170 26660 5176
rect 26620 5030 26648 5170
rect 26712 5030 26740 5494
rect 26608 5024 26660 5030
rect 26608 4966 26660 4972
rect 26700 5024 26752 5030
rect 26700 4966 26752 4972
rect 25872 4004 25924 4010
rect 25872 3946 25924 3952
rect 25884 3602 25912 3946
rect 25872 3596 25924 3602
rect 25872 3538 25924 3544
rect 25964 3528 26016 3534
rect 25964 3470 26016 3476
rect 25780 3460 25832 3466
rect 25780 3402 25832 3408
rect 25686 3360 25742 3369
rect 25686 3295 25742 3304
rect 25700 3194 25728 3295
rect 25688 3188 25740 3194
rect 25688 3130 25740 3136
rect 25228 3120 25280 3126
rect 25228 3062 25280 3068
rect 25320 3120 25372 3126
rect 25320 3062 25372 3068
rect 25228 2440 25280 2446
rect 25226 2408 25228 2417
rect 25280 2408 25282 2417
rect 24768 2372 24820 2378
rect 25226 2343 25282 2352
rect 24768 2314 24820 2320
rect 24780 950 24808 2314
rect 24952 2304 25004 2310
rect 24952 2246 25004 2252
rect 24768 944 24820 950
rect 24768 886 24820 892
rect 24964 800 24992 2246
rect 25228 1012 25280 1018
rect 25228 954 25280 960
rect 25240 800 25268 954
rect 25504 944 25556 950
rect 25504 886 25556 892
rect 25516 800 25544 886
rect 25792 800 25820 3402
rect 25976 3194 26004 3470
rect 26240 3460 26292 3466
rect 26240 3402 26292 3408
rect 25964 3188 26016 3194
rect 25964 3130 26016 3136
rect 25976 2854 26004 3130
rect 26252 3058 26280 3402
rect 26240 3052 26292 3058
rect 26240 2994 26292 3000
rect 26516 2984 26568 2990
rect 26516 2926 26568 2932
rect 25964 2848 26016 2854
rect 25964 2790 26016 2796
rect 26528 2774 26556 2926
rect 26344 2746 26556 2774
rect 26896 2774 26924 12922
rect 26988 9217 27016 13246
rect 26974 9208 27030 9217
rect 26974 9143 27030 9152
rect 26988 9042 27016 9143
rect 26976 9036 27028 9042
rect 26976 8978 27028 8984
rect 27080 8498 27108 14826
rect 27160 13456 27212 13462
rect 27160 13398 27212 13404
rect 27172 12345 27200 13398
rect 27158 12336 27214 12345
rect 27158 12271 27214 12280
rect 27264 9674 27292 16458
rect 27264 9646 27384 9674
rect 27160 9580 27212 9586
rect 27160 9522 27212 9528
rect 27172 9042 27200 9522
rect 27250 9480 27306 9489
rect 27250 9415 27306 9424
rect 27160 9036 27212 9042
rect 27160 8978 27212 8984
rect 27068 8492 27120 8498
rect 27068 8434 27120 8440
rect 27172 6866 27200 8978
rect 27264 7818 27292 9415
rect 27356 9178 27384 9646
rect 27344 9172 27396 9178
rect 27344 9114 27396 9120
rect 27252 7812 27304 7818
rect 27252 7754 27304 7760
rect 27264 7206 27292 7754
rect 27252 7200 27304 7206
rect 27252 7142 27304 7148
rect 27160 6860 27212 6866
rect 27160 6802 27212 6808
rect 27448 5148 27476 25162
rect 27632 24818 27660 25230
rect 27620 24812 27672 24818
rect 27620 24754 27672 24760
rect 27724 24070 27752 25298
rect 27816 24410 27844 32263
rect 27908 32026 27936 32370
rect 27896 32020 27948 32026
rect 27896 31962 27948 31968
rect 28000 29782 28028 35430
rect 28092 35018 28120 41482
rect 28368 36174 28396 49030
rect 29736 45552 29788 45558
rect 29736 45494 29788 45500
rect 28540 42016 28592 42022
rect 28540 41958 28592 41964
rect 28356 36168 28408 36174
rect 28356 36110 28408 36116
rect 28264 35828 28316 35834
rect 28264 35770 28316 35776
rect 28276 35698 28304 35770
rect 28264 35692 28316 35698
rect 28264 35634 28316 35640
rect 28448 35692 28500 35698
rect 28448 35634 28500 35640
rect 28460 35494 28488 35634
rect 28448 35488 28500 35494
rect 28448 35430 28500 35436
rect 28080 35012 28132 35018
rect 28080 34954 28132 34960
rect 28092 32842 28120 34954
rect 28264 32904 28316 32910
rect 28264 32846 28316 32852
rect 28080 32836 28132 32842
rect 28080 32778 28132 32784
rect 28172 32564 28224 32570
rect 28172 32506 28224 32512
rect 28080 32292 28132 32298
rect 28080 32234 28132 32240
rect 28092 32201 28120 32234
rect 28078 32192 28134 32201
rect 28078 32127 28134 32136
rect 28184 31890 28212 32506
rect 28172 31884 28224 31890
rect 28172 31826 28224 31832
rect 28080 31816 28132 31822
rect 28080 31758 28132 31764
rect 27988 29776 28040 29782
rect 27988 29718 28040 29724
rect 27988 28416 28040 28422
rect 27988 28358 28040 28364
rect 27896 27396 27948 27402
rect 27896 27338 27948 27344
rect 27908 26586 27936 27338
rect 28000 26994 28028 28358
rect 27988 26988 28040 26994
rect 27988 26930 28040 26936
rect 27896 26580 27948 26586
rect 27896 26522 27948 26528
rect 27908 25770 27936 26522
rect 27896 25764 27948 25770
rect 27896 25706 27948 25712
rect 27896 25356 27948 25362
rect 27896 25298 27948 25304
rect 27804 24404 27856 24410
rect 27804 24346 27856 24352
rect 27712 24064 27764 24070
rect 27712 24006 27764 24012
rect 27816 23798 27844 24346
rect 27804 23792 27856 23798
rect 27804 23734 27856 23740
rect 27712 21616 27764 21622
rect 27712 21558 27764 21564
rect 27620 20800 27672 20806
rect 27620 20742 27672 20748
rect 27632 20398 27660 20742
rect 27620 20392 27672 20398
rect 27620 20334 27672 20340
rect 27620 19508 27672 19514
rect 27620 19450 27672 19456
rect 27632 18766 27660 19450
rect 27620 18760 27672 18766
rect 27620 18702 27672 18708
rect 27724 18578 27752 21558
rect 27908 20482 27936 25298
rect 28092 25242 28120 31758
rect 28172 30660 28224 30666
rect 28172 30602 28224 30608
rect 28184 30054 28212 30602
rect 28172 30048 28224 30054
rect 28172 29990 28224 29996
rect 28172 27328 28224 27334
rect 28172 27270 28224 27276
rect 28184 26450 28212 27270
rect 28172 26444 28224 26450
rect 28172 26386 28224 26392
rect 28172 25900 28224 25906
rect 28172 25842 28224 25848
rect 28184 25498 28212 25842
rect 28276 25838 28304 32846
rect 28448 32428 28500 32434
rect 28448 32370 28500 32376
rect 28460 32337 28488 32370
rect 28446 32328 28502 32337
rect 28446 32263 28502 32272
rect 28356 30048 28408 30054
rect 28356 29990 28408 29996
rect 28446 30016 28502 30025
rect 28368 26450 28396 29990
rect 28446 29951 28502 29960
rect 28460 29646 28488 29951
rect 28448 29640 28500 29646
rect 28448 29582 28500 29588
rect 28448 28756 28500 28762
rect 28448 28698 28500 28704
rect 28460 27674 28488 28698
rect 28552 28558 28580 41958
rect 28724 41608 28776 41614
rect 28724 41550 28776 41556
rect 28632 36032 28684 36038
rect 28632 35974 28684 35980
rect 28644 35698 28672 35974
rect 28632 35692 28684 35698
rect 28632 35634 28684 35640
rect 28736 35630 28764 41550
rect 29552 39432 29604 39438
rect 29552 39374 29604 39380
rect 29368 39364 29420 39370
rect 29368 39306 29420 39312
rect 29092 35692 29144 35698
rect 29092 35634 29144 35640
rect 28724 35624 28776 35630
rect 28724 35566 28776 35572
rect 29104 35222 29132 35634
rect 29092 35216 29144 35222
rect 29092 35158 29144 35164
rect 28632 32224 28684 32230
rect 28630 32192 28632 32201
rect 28684 32192 28686 32201
rect 28630 32127 28686 32136
rect 28724 30728 28776 30734
rect 28724 30670 28776 30676
rect 28632 30660 28684 30666
rect 28632 30602 28684 30608
rect 28644 30394 28672 30602
rect 28632 30388 28684 30394
rect 28632 30330 28684 30336
rect 28736 30258 28764 30670
rect 28724 30252 28776 30258
rect 28724 30194 28776 30200
rect 28722 29744 28778 29753
rect 28722 29679 28778 29688
rect 28736 29646 28764 29679
rect 28724 29640 28776 29646
rect 28724 29582 28776 29588
rect 28632 29504 28684 29510
rect 28632 29446 28684 29452
rect 28644 29170 28672 29446
rect 28908 29300 28960 29306
rect 28908 29242 28960 29248
rect 28632 29164 28684 29170
rect 28632 29106 28684 29112
rect 28724 29164 28776 29170
rect 28724 29106 28776 29112
rect 28816 29164 28868 29170
rect 28816 29106 28868 29112
rect 28736 28642 28764 29106
rect 28828 28762 28856 29106
rect 28816 28756 28868 28762
rect 28816 28698 28868 28704
rect 28644 28614 28764 28642
rect 28540 28552 28592 28558
rect 28540 28494 28592 28500
rect 28540 28076 28592 28082
rect 28540 28018 28592 28024
rect 28448 27668 28500 27674
rect 28448 27610 28500 27616
rect 28448 27464 28500 27470
rect 28446 27432 28448 27441
rect 28500 27432 28502 27441
rect 28446 27367 28502 27376
rect 28448 27328 28500 27334
rect 28448 27270 28500 27276
rect 28356 26444 28408 26450
rect 28356 26386 28408 26392
rect 28264 25832 28316 25838
rect 28264 25774 28316 25780
rect 28172 25492 28224 25498
rect 28172 25434 28224 25440
rect 28264 25288 28316 25294
rect 28092 25214 28212 25242
rect 28264 25230 28316 25236
rect 28080 25152 28132 25158
rect 28080 25094 28132 25100
rect 28092 24818 28120 25094
rect 28080 24812 28132 24818
rect 28080 24754 28132 24760
rect 28080 24676 28132 24682
rect 28080 24618 28132 24624
rect 27988 24132 28040 24138
rect 27988 24074 28040 24080
rect 28000 20618 28028 24074
rect 28092 22098 28120 24618
rect 28184 24342 28212 25214
rect 28276 24410 28304 25230
rect 28368 25226 28396 26386
rect 28460 25294 28488 27270
rect 28448 25288 28500 25294
rect 28448 25230 28500 25236
rect 28356 25220 28408 25226
rect 28356 25162 28408 25168
rect 28368 24886 28396 25162
rect 28356 24880 28408 24886
rect 28356 24822 28408 24828
rect 28264 24404 28316 24410
rect 28264 24346 28316 24352
rect 28172 24336 28224 24342
rect 28172 24278 28224 24284
rect 28172 24200 28224 24206
rect 28172 24142 28224 24148
rect 28184 23866 28212 24142
rect 28172 23860 28224 23866
rect 28172 23802 28224 23808
rect 28080 22092 28132 22098
rect 28080 22034 28132 22040
rect 28092 21622 28120 22034
rect 28264 22024 28316 22030
rect 28264 21966 28316 21972
rect 28172 21888 28224 21894
rect 28172 21830 28224 21836
rect 28080 21616 28132 21622
rect 28080 21558 28132 21564
rect 28000 20590 28120 20618
rect 27908 20454 28028 20482
rect 27896 20392 27948 20398
rect 27896 20334 27948 20340
rect 27908 19854 27936 20334
rect 27896 19848 27948 19854
rect 27802 19816 27858 19825
rect 27896 19790 27948 19796
rect 27802 19751 27858 19760
rect 27816 19718 27844 19751
rect 27804 19712 27856 19718
rect 27804 19654 27856 19660
rect 27632 18550 27752 18578
rect 27896 18624 27948 18630
rect 27896 18566 27948 18572
rect 27528 17808 27580 17814
rect 27528 17750 27580 17756
rect 27540 17202 27568 17750
rect 27632 17202 27660 18550
rect 27908 18290 27936 18566
rect 27896 18284 27948 18290
rect 27896 18226 27948 18232
rect 27528 17196 27580 17202
rect 27528 17138 27580 17144
rect 27620 17196 27672 17202
rect 27620 17138 27672 17144
rect 27528 11144 27580 11150
rect 27528 11086 27580 11092
rect 27540 10198 27568 11086
rect 27632 11014 27660 17138
rect 27804 16176 27856 16182
rect 27804 16118 27856 16124
rect 27712 14340 27764 14346
rect 27712 14282 27764 14288
rect 27724 14074 27752 14282
rect 27712 14068 27764 14074
rect 27712 14010 27764 14016
rect 27620 11008 27672 11014
rect 27620 10950 27672 10956
rect 27620 10532 27672 10538
rect 27620 10474 27672 10480
rect 27712 10532 27764 10538
rect 27712 10474 27764 10480
rect 27528 10192 27580 10198
rect 27528 10134 27580 10140
rect 27632 8401 27660 10474
rect 27724 10441 27752 10474
rect 27710 10432 27766 10441
rect 27710 10367 27766 10376
rect 27712 9580 27764 9586
rect 27712 9522 27764 9528
rect 27724 8634 27752 9522
rect 27816 9489 27844 16118
rect 27896 16040 27948 16046
rect 27896 15982 27948 15988
rect 27908 15366 27936 15982
rect 27896 15360 27948 15366
rect 27896 15302 27948 15308
rect 27896 15156 27948 15162
rect 27896 15098 27948 15104
rect 27908 13394 27936 15098
rect 27896 13388 27948 13394
rect 27896 13330 27948 13336
rect 28000 12434 28028 20454
rect 27908 12406 28028 12434
rect 28092 12434 28120 20590
rect 28184 20534 28212 21830
rect 28276 21690 28304 21966
rect 28264 21684 28316 21690
rect 28264 21626 28316 21632
rect 28368 21570 28396 24822
rect 28552 24342 28580 28018
rect 28644 27878 28672 28614
rect 28816 28552 28868 28558
rect 28816 28494 28868 28500
rect 28724 28484 28776 28490
rect 28724 28426 28776 28432
rect 28736 28218 28764 28426
rect 28828 28218 28856 28494
rect 28724 28212 28776 28218
rect 28724 28154 28776 28160
rect 28816 28212 28868 28218
rect 28816 28154 28868 28160
rect 28920 28082 28948 29242
rect 29000 28960 29052 28966
rect 29000 28902 29052 28908
rect 29012 28762 29040 28902
rect 29000 28756 29052 28762
rect 29000 28698 29052 28704
rect 28908 28076 28960 28082
rect 28908 28018 28960 28024
rect 28632 27872 28684 27878
rect 28632 27814 28684 27820
rect 28632 27532 28684 27538
rect 28632 27474 28684 27480
rect 28644 27169 28672 27474
rect 28630 27160 28686 27169
rect 28630 27095 28686 27104
rect 28920 24818 28948 28018
rect 29000 28008 29052 28014
rect 29000 27950 29052 27956
rect 29012 27878 29040 27950
rect 29000 27872 29052 27878
rect 29000 27814 29052 27820
rect 29104 26994 29132 35158
rect 29380 30802 29408 39306
rect 29460 38752 29512 38758
rect 29460 38694 29512 38700
rect 29368 30796 29420 30802
rect 29368 30738 29420 30744
rect 29184 29572 29236 29578
rect 29184 29514 29236 29520
rect 29092 26988 29144 26994
rect 29092 26930 29144 26936
rect 29104 26382 29132 26930
rect 29092 26376 29144 26382
rect 29092 26318 29144 26324
rect 29104 25974 29132 26318
rect 29092 25968 29144 25974
rect 29092 25910 29144 25916
rect 28908 24812 28960 24818
rect 28908 24754 28960 24760
rect 28632 24744 28684 24750
rect 28632 24686 28684 24692
rect 28448 24336 28500 24342
rect 28448 24278 28500 24284
rect 28540 24336 28592 24342
rect 28540 24278 28592 24284
rect 28460 24206 28488 24278
rect 28644 24206 28672 24686
rect 28448 24200 28500 24206
rect 28448 24142 28500 24148
rect 28632 24200 28684 24206
rect 28632 24142 28684 24148
rect 29090 24168 29146 24177
rect 28276 21542 28396 21570
rect 28172 20528 28224 20534
rect 28172 20470 28224 20476
rect 28276 20346 28304 21542
rect 28460 21486 28488 24142
rect 28644 23798 28672 24142
rect 29090 24103 29092 24112
rect 29144 24103 29146 24112
rect 29092 24074 29144 24080
rect 28632 23792 28684 23798
rect 28632 23734 28684 23740
rect 28448 21480 28500 21486
rect 28448 21422 28500 21428
rect 28356 21412 28408 21418
rect 28356 21354 28408 21360
rect 29092 21412 29144 21418
rect 29092 21354 29144 21360
rect 28184 20318 28304 20346
rect 28184 17762 28212 20318
rect 28264 20256 28316 20262
rect 28264 20198 28316 20204
rect 28276 19378 28304 20198
rect 28368 19514 28396 21354
rect 29104 21078 29132 21354
rect 29092 21072 29144 21078
rect 29092 21014 29144 21020
rect 28632 21004 28684 21010
rect 28632 20946 28684 20952
rect 28540 20936 28592 20942
rect 28540 20878 28592 20884
rect 28448 20460 28500 20466
rect 28448 20402 28500 20408
rect 28460 20058 28488 20402
rect 28448 20052 28500 20058
rect 28448 19994 28500 20000
rect 28552 19786 28580 20878
rect 28644 20058 28672 20946
rect 28816 20596 28868 20602
rect 28816 20538 28868 20544
rect 28724 20460 28776 20466
rect 28724 20402 28776 20408
rect 28632 20052 28684 20058
rect 28632 19994 28684 20000
rect 28540 19780 28592 19786
rect 28540 19722 28592 19728
rect 28552 19689 28580 19722
rect 28538 19680 28594 19689
rect 28538 19615 28594 19624
rect 28644 19514 28672 19994
rect 28736 19718 28764 20402
rect 28828 20058 28856 20538
rect 28908 20256 28960 20262
rect 28908 20198 28960 20204
rect 28816 20052 28868 20058
rect 28816 19994 28868 20000
rect 28828 19922 28856 19994
rect 28920 19922 28948 20198
rect 28816 19916 28868 19922
rect 28816 19858 28868 19864
rect 28908 19916 28960 19922
rect 28908 19858 28960 19864
rect 28814 19816 28870 19825
rect 28814 19751 28816 19760
rect 28868 19751 28870 19760
rect 28816 19722 28868 19728
rect 28724 19712 28776 19718
rect 29000 19712 29052 19718
rect 28724 19654 28776 19660
rect 28906 19680 28962 19689
rect 28356 19508 28408 19514
rect 28356 19450 28408 19456
rect 28632 19508 28684 19514
rect 28632 19450 28684 19456
rect 28264 19372 28316 19378
rect 28264 19314 28316 19320
rect 28644 19242 28672 19450
rect 28632 19236 28684 19242
rect 28632 19178 28684 19184
rect 28184 17746 28304 17762
rect 28184 17740 28316 17746
rect 28184 17734 28264 17740
rect 28264 17682 28316 17688
rect 28356 17740 28408 17746
rect 28356 17682 28408 17688
rect 28276 17134 28304 17682
rect 28264 17128 28316 17134
rect 28264 17070 28316 17076
rect 28368 16946 28396 17682
rect 28540 17672 28592 17678
rect 28540 17614 28592 17620
rect 28276 16918 28396 16946
rect 28172 16448 28224 16454
rect 28172 16390 28224 16396
rect 28184 16114 28212 16390
rect 28276 16114 28304 16918
rect 28356 16584 28408 16590
rect 28356 16526 28408 16532
rect 28368 16250 28396 16526
rect 28552 16454 28580 17614
rect 28632 17332 28684 17338
rect 28632 17274 28684 17280
rect 28540 16448 28592 16454
rect 28540 16390 28592 16396
rect 28356 16244 28408 16250
rect 28356 16186 28408 16192
rect 28172 16108 28224 16114
rect 28172 16050 28224 16056
rect 28264 16108 28316 16114
rect 28264 16050 28316 16056
rect 28276 15910 28304 16050
rect 28356 16040 28408 16046
rect 28356 15982 28408 15988
rect 28264 15904 28316 15910
rect 28264 15846 28316 15852
rect 28368 15366 28396 15982
rect 28264 15360 28316 15366
rect 28264 15302 28316 15308
rect 28356 15360 28408 15366
rect 28356 15302 28408 15308
rect 28172 13524 28224 13530
rect 28172 13466 28224 13472
rect 28184 13190 28212 13466
rect 28172 13184 28224 13190
rect 28172 13126 28224 13132
rect 28092 12406 28212 12434
rect 27802 9480 27858 9489
rect 27802 9415 27858 9424
rect 27804 8900 27856 8906
rect 27804 8842 27856 8848
rect 27712 8628 27764 8634
rect 27712 8570 27764 8576
rect 27618 8392 27674 8401
rect 27618 8327 27674 8336
rect 27816 8090 27844 8842
rect 27804 8084 27856 8090
rect 27804 8026 27856 8032
rect 27712 7948 27764 7954
rect 27712 7890 27764 7896
rect 27528 7744 27580 7750
rect 27528 7686 27580 7692
rect 27540 7342 27568 7686
rect 27528 7336 27580 7342
rect 27528 7278 27580 7284
rect 27528 6860 27580 6866
rect 27528 6802 27580 6808
rect 27540 5710 27568 6802
rect 27620 6792 27672 6798
rect 27620 6734 27672 6740
rect 27528 5704 27580 5710
rect 27632 5681 27660 6734
rect 27724 5846 27752 7890
rect 27908 6798 27936 12406
rect 27988 11008 28040 11014
rect 27988 10950 28040 10956
rect 28000 9586 28028 10950
rect 28080 10736 28132 10742
rect 28080 10678 28132 10684
rect 28092 10062 28120 10678
rect 28080 10056 28132 10062
rect 28080 9998 28132 10004
rect 28184 9874 28212 12406
rect 28092 9846 28212 9874
rect 27988 9580 28040 9586
rect 27988 9522 28040 9528
rect 27988 8900 28040 8906
rect 27988 8842 28040 8848
rect 28000 8566 28028 8842
rect 27988 8560 28040 8566
rect 27988 8502 28040 8508
rect 28092 7562 28120 9846
rect 28276 8838 28304 15302
rect 28552 15162 28580 16390
rect 28540 15156 28592 15162
rect 28540 15098 28592 15104
rect 28448 15020 28500 15026
rect 28448 14962 28500 14968
rect 28460 14618 28488 14962
rect 28448 14612 28500 14618
rect 28448 14554 28500 14560
rect 28540 11552 28592 11558
rect 28540 11494 28592 11500
rect 28552 11286 28580 11494
rect 28540 11280 28592 11286
rect 28540 11222 28592 11228
rect 28552 10674 28580 11222
rect 28644 11121 28672 17274
rect 28736 17134 28764 19654
rect 28962 19660 29000 19666
rect 28962 19654 29052 19660
rect 28962 19638 29040 19654
rect 28906 19615 28962 19624
rect 29000 18284 29052 18290
rect 29000 18226 29052 18232
rect 29092 18284 29144 18290
rect 29092 18226 29144 18232
rect 29012 17814 29040 18226
rect 29000 17808 29052 17814
rect 29000 17750 29052 17756
rect 28724 17128 28776 17134
rect 28724 17070 28776 17076
rect 28736 16658 28764 17070
rect 28724 16652 28776 16658
rect 28724 16594 28776 16600
rect 28736 16046 28764 16594
rect 29104 16454 29132 18226
rect 29092 16448 29144 16454
rect 29092 16390 29144 16396
rect 28724 16040 28776 16046
rect 28724 15982 28776 15988
rect 28722 15736 28778 15745
rect 29196 15706 29224 29514
rect 29368 28076 29420 28082
rect 29368 28018 29420 28024
rect 29276 22024 29328 22030
rect 29276 21966 29328 21972
rect 29288 21486 29316 21966
rect 29276 21480 29328 21486
rect 29276 21422 29328 21428
rect 29380 19446 29408 28018
rect 29472 22094 29500 38694
rect 29564 32994 29592 39374
rect 29748 33114 29776 45494
rect 29736 33108 29788 33114
rect 29736 33050 29788 33056
rect 29564 32966 29776 32994
rect 29552 32360 29604 32366
rect 29552 32302 29604 32308
rect 29564 32065 29592 32302
rect 29550 32056 29606 32065
rect 29550 31991 29606 32000
rect 29748 31754 29776 32966
rect 29828 32972 29880 32978
rect 29828 32914 29880 32920
rect 29840 32366 29868 32914
rect 29828 32360 29880 32366
rect 29828 32302 29880 32308
rect 30024 32042 30052 51046
rect 30484 49230 30512 56850
rect 30852 49298 30880 57190
rect 30840 49292 30892 49298
rect 30840 49234 30892 49240
rect 30472 49224 30524 49230
rect 30472 49166 30524 49172
rect 30380 49156 30432 49162
rect 30380 49098 30432 49104
rect 30392 48226 30420 49098
rect 30932 49088 30984 49094
rect 30932 49030 30984 49036
rect 30656 48544 30708 48550
rect 30656 48486 30708 48492
rect 30392 48198 30512 48226
rect 30380 48136 30432 48142
rect 30380 48078 30432 48084
rect 30392 47666 30420 48078
rect 30380 47660 30432 47666
rect 30380 47602 30432 47608
rect 30392 36174 30420 47602
rect 30484 47054 30512 48198
rect 30472 47048 30524 47054
rect 30472 46990 30524 46996
rect 30484 42226 30512 46990
rect 30472 42220 30524 42226
rect 30472 42162 30524 42168
rect 30564 37936 30616 37942
rect 30564 37878 30616 37884
rect 30380 36168 30432 36174
rect 30380 36110 30432 36116
rect 30104 35488 30156 35494
rect 30104 35430 30156 35436
rect 30116 33522 30144 35430
rect 30104 33516 30156 33522
rect 30104 33458 30156 33464
rect 29932 32014 30052 32042
rect 29748 31726 29868 31754
rect 29644 30728 29696 30734
rect 29644 30670 29696 30676
rect 29656 30394 29684 30670
rect 29736 30592 29788 30598
rect 29736 30534 29788 30540
rect 29644 30388 29696 30394
rect 29644 30330 29696 30336
rect 29748 30326 29776 30534
rect 29736 30320 29788 30326
rect 29736 30262 29788 30268
rect 29748 29646 29776 30262
rect 29736 29640 29788 29646
rect 29736 29582 29788 29588
rect 29644 29164 29696 29170
rect 29644 29106 29696 29112
rect 29656 28121 29684 29106
rect 29642 28112 29698 28121
rect 29642 28047 29698 28056
rect 29736 24744 29788 24750
rect 29736 24686 29788 24692
rect 29748 24614 29776 24686
rect 29736 24608 29788 24614
rect 29736 24550 29788 24556
rect 29748 24206 29776 24550
rect 29840 24206 29868 31726
rect 29932 30870 29960 32014
rect 29920 30864 29972 30870
rect 29920 30806 29972 30812
rect 30116 30394 30144 33458
rect 30196 33108 30248 33114
rect 30196 33050 30248 33056
rect 30208 32230 30236 33050
rect 30196 32224 30248 32230
rect 30196 32166 30248 32172
rect 30208 31754 30236 32166
rect 30392 31754 30420 36110
rect 30472 36032 30524 36038
rect 30470 36000 30472 36009
rect 30524 36000 30526 36009
rect 30470 35935 30526 35944
rect 30576 35086 30604 37878
rect 30668 36174 30696 48486
rect 30840 48000 30892 48006
rect 30840 47942 30892 47948
rect 30852 47666 30880 47942
rect 30840 47660 30892 47666
rect 30840 47602 30892 47608
rect 30656 36168 30708 36174
rect 30656 36110 30708 36116
rect 30840 35692 30892 35698
rect 30840 35634 30892 35640
rect 30852 35086 30880 35634
rect 30564 35080 30616 35086
rect 30564 35022 30616 35028
rect 30840 35080 30892 35086
rect 30840 35022 30892 35028
rect 30748 35012 30800 35018
rect 30748 34954 30800 34960
rect 30760 34649 30788 34954
rect 30746 34640 30802 34649
rect 30746 34575 30802 34584
rect 30852 31822 30880 35022
rect 30840 31816 30892 31822
rect 30840 31758 30892 31764
rect 30208 31726 30328 31754
rect 30392 31726 30512 31754
rect 30300 30734 30328 31726
rect 30288 30728 30340 30734
rect 30288 30670 30340 30676
rect 30104 30388 30156 30394
rect 30104 30330 30156 30336
rect 30012 30184 30064 30190
rect 30012 30126 30064 30132
rect 30024 29646 30052 30126
rect 30012 29640 30064 29646
rect 30012 29582 30064 29588
rect 30196 29504 30248 29510
rect 30196 29446 30248 29452
rect 30012 28484 30064 28490
rect 30012 28426 30064 28432
rect 29918 28112 29974 28121
rect 30024 28082 30052 28426
rect 30104 28212 30156 28218
rect 30104 28154 30156 28160
rect 29918 28047 29974 28056
rect 30012 28076 30064 28082
rect 29932 26586 29960 28047
rect 30012 28018 30064 28024
rect 30116 27606 30144 28154
rect 30104 27600 30156 27606
rect 30104 27542 30156 27548
rect 30012 26784 30064 26790
rect 30012 26726 30064 26732
rect 29920 26580 29972 26586
rect 29920 26522 29972 26528
rect 29932 26382 29960 26522
rect 30024 26382 30052 26726
rect 30116 26382 30144 27542
rect 29920 26376 29972 26382
rect 29920 26318 29972 26324
rect 30012 26376 30064 26382
rect 30012 26318 30064 26324
rect 30104 26376 30156 26382
rect 30104 26318 30156 26324
rect 30104 25900 30156 25906
rect 30104 25842 30156 25848
rect 30116 25498 30144 25842
rect 30104 25492 30156 25498
rect 30104 25434 30156 25440
rect 29736 24200 29788 24206
rect 29736 24142 29788 24148
rect 29828 24200 29880 24206
rect 29828 24142 29880 24148
rect 29736 23112 29788 23118
rect 29736 23054 29788 23060
rect 29552 22976 29604 22982
rect 29552 22918 29604 22924
rect 29564 22642 29592 22918
rect 29552 22636 29604 22642
rect 29552 22578 29604 22584
rect 29748 22234 29776 23054
rect 29828 23044 29880 23050
rect 29828 22986 29880 22992
rect 29736 22228 29788 22234
rect 29736 22170 29788 22176
rect 29472 22066 29592 22094
rect 29368 19440 29420 19446
rect 29368 19382 29420 19388
rect 28722 15671 28778 15680
rect 29000 15700 29052 15706
rect 28736 15638 28764 15671
rect 29000 15642 29052 15648
rect 29184 15700 29236 15706
rect 29184 15642 29236 15648
rect 28724 15632 28776 15638
rect 28724 15574 28776 15580
rect 28908 15496 28960 15502
rect 28908 15438 28960 15444
rect 28920 14958 28948 15438
rect 28908 14952 28960 14958
rect 28828 14912 28908 14940
rect 28828 14414 28856 14912
rect 28908 14894 28960 14900
rect 28816 14408 28868 14414
rect 28816 14350 28868 14356
rect 28814 13968 28870 13977
rect 28814 13903 28870 13912
rect 28908 13932 28960 13938
rect 28724 13864 28776 13870
rect 28724 13806 28776 13812
rect 28630 11112 28686 11121
rect 28630 11047 28686 11056
rect 28540 10668 28592 10674
rect 28540 10610 28592 10616
rect 28632 10668 28684 10674
rect 28632 10610 28684 10616
rect 28354 9888 28410 9897
rect 28354 9823 28410 9832
rect 28368 8974 28396 9823
rect 28552 9722 28580 10610
rect 28644 10441 28672 10610
rect 28630 10432 28686 10441
rect 28630 10367 28686 10376
rect 28540 9716 28592 9722
rect 28540 9658 28592 9664
rect 28538 9480 28594 9489
rect 28538 9415 28540 9424
rect 28592 9415 28594 9424
rect 28632 9444 28684 9450
rect 28540 9386 28592 9392
rect 28632 9386 28684 9392
rect 28356 8968 28408 8974
rect 28356 8910 28408 8916
rect 28264 8832 28316 8838
rect 28264 8774 28316 8780
rect 28276 7818 28304 8774
rect 28448 8628 28500 8634
rect 28552 8616 28580 9386
rect 28500 8588 28580 8616
rect 28448 8570 28500 8576
rect 28538 8528 28594 8537
rect 28538 8463 28594 8472
rect 28356 8424 28408 8430
rect 28356 8366 28408 8372
rect 28264 7812 28316 7818
rect 28264 7754 28316 7760
rect 28092 7534 28304 7562
rect 28172 6860 28224 6866
rect 28172 6802 28224 6808
rect 27896 6792 27948 6798
rect 27896 6734 27948 6740
rect 27804 6248 27856 6254
rect 27802 6216 27804 6225
rect 27856 6216 27858 6225
rect 27802 6151 27858 6160
rect 27712 5840 27764 5846
rect 27712 5782 27764 5788
rect 27724 5710 27752 5782
rect 27712 5704 27764 5710
rect 27528 5646 27580 5652
rect 27618 5672 27674 5681
rect 27540 5216 27568 5646
rect 27712 5646 27764 5652
rect 27618 5607 27674 5616
rect 27908 5273 27936 6734
rect 28184 6458 28212 6802
rect 28172 6452 28224 6458
rect 28172 6394 28224 6400
rect 28080 6248 28132 6254
rect 28080 6190 28132 6196
rect 27894 5264 27950 5273
rect 27620 5228 27672 5234
rect 27540 5188 27620 5216
rect 27894 5199 27950 5208
rect 27620 5170 27672 5176
rect 27712 5160 27764 5166
rect 27448 5120 27568 5148
rect 27068 4616 27120 4622
rect 27068 4558 27120 4564
rect 26976 3936 27028 3942
rect 26976 3878 27028 3884
rect 26988 3602 27016 3878
rect 26976 3596 27028 3602
rect 26976 3538 27028 3544
rect 26896 2746 27016 2774
rect 26056 2372 26108 2378
rect 26056 2314 26108 2320
rect 26068 800 26096 2314
rect 26344 800 26372 2746
rect 26988 2446 27016 2746
rect 26976 2440 27028 2446
rect 26976 2382 27028 2388
rect 26608 2372 26660 2378
rect 26608 2314 26660 2320
rect 26884 2372 26936 2378
rect 27080 2360 27108 4558
rect 27436 4004 27488 4010
rect 27436 3946 27488 3952
rect 27160 3936 27212 3942
rect 27160 3878 27212 3884
rect 27172 3534 27200 3878
rect 27160 3528 27212 3534
rect 27160 3470 27212 3476
rect 27160 3392 27212 3398
rect 27160 3334 27212 3340
rect 27172 3194 27200 3334
rect 27160 3188 27212 3194
rect 27160 3130 27212 3136
rect 27080 2332 27200 2360
rect 26884 2314 26936 2320
rect 26620 800 26648 2314
rect 26896 800 26924 2314
rect 27172 800 27200 2332
rect 27448 800 27476 3946
rect 27540 3913 27568 5120
rect 27712 5102 27764 5108
rect 27724 4826 27752 5102
rect 27712 4820 27764 4826
rect 27712 4762 27764 4768
rect 27804 4820 27856 4826
rect 27804 4762 27856 4768
rect 27712 4616 27764 4622
rect 27712 4558 27764 4564
rect 27620 4072 27672 4078
rect 27620 4014 27672 4020
rect 27526 3904 27582 3913
rect 27526 3839 27582 3848
rect 27632 3738 27660 4014
rect 27620 3732 27672 3738
rect 27620 3674 27672 3680
rect 27528 2644 27580 2650
rect 27528 2586 27580 2592
rect 27540 950 27568 2586
rect 27528 944 27580 950
rect 27528 886 27580 892
rect 27724 800 27752 4558
rect 27816 4554 27844 4762
rect 27896 4684 27948 4690
rect 27896 4626 27948 4632
rect 27804 4548 27856 4554
rect 27804 4490 27856 4496
rect 27908 4214 27936 4626
rect 28092 4622 28120 6190
rect 28172 5568 28224 5574
rect 28172 5510 28224 5516
rect 28184 4622 28212 5510
rect 27988 4616 28040 4622
rect 27988 4558 28040 4564
rect 28080 4616 28132 4622
rect 28080 4558 28132 4564
rect 28172 4616 28224 4622
rect 28276 4593 28304 7534
rect 28368 7313 28396 8366
rect 28448 8356 28500 8362
rect 28552 8344 28580 8463
rect 28644 8430 28672 9386
rect 28632 8424 28684 8430
rect 28632 8366 28684 8372
rect 28500 8316 28580 8344
rect 28448 8298 28500 8304
rect 28448 7744 28500 7750
rect 28448 7686 28500 7692
rect 28354 7304 28410 7313
rect 28354 7239 28410 7248
rect 28368 6322 28396 7239
rect 28356 6316 28408 6322
rect 28356 6258 28408 6264
rect 28460 4690 28488 7686
rect 28552 6254 28580 8316
rect 28644 7954 28672 8366
rect 28632 7948 28684 7954
rect 28632 7890 28684 7896
rect 28540 6248 28592 6254
rect 28540 6190 28592 6196
rect 28736 6118 28764 13806
rect 28828 13802 28856 13903
rect 28908 13874 28960 13880
rect 28816 13796 28868 13802
rect 28816 13738 28868 13744
rect 28828 13258 28856 13738
rect 28816 13252 28868 13258
rect 28816 13194 28868 13200
rect 28920 12442 28948 13874
rect 28908 12436 28960 12442
rect 28908 12378 28960 12384
rect 28816 11552 28868 11558
rect 28816 11494 28868 11500
rect 28828 11150 28856 11494
rect 29012 11393 29040 15642
rect 29276 15564 29328 15570
rect 29276 15506 29328 15512
rect 29092 14272 29144 14278
rect 29092 14214 29144 14220
rect 29184 14272 29236 14278
rect 29184 14214 29236 14220
rect 29104 13841 29132 14214
rect 29196 14074 29224 14214
rect 29184 14068 29236 14074
rect 29184 14010 29236 14016
rect 29090 13832 29146 13841
rect 29090 13767 29146 13776
rect 29288 13530 29316 15506
rect 29276 13524 29328 13530
rect 29276 13466 29328 13472
rect 29090 13016 29146 13025
rect 29090 12951 29146 12960
rect 29104 11626 29132 12951
rect 29276 12708 29328 12714
rect 29276 12650 29328 12656
rect 29184 12436 29236 12442
rect 29184 12378 29236 12384
rect 29092 11620 29144 11626
rect 29092 11562 29144 11568
rect 28998 11384 29054 11393
rect 28998 11319 29054 11328
rect 29196 11218 29224 12378
rect 29184 11212 29236 11218
rect 29184 11154 29236 11160
rect 28816 11144 28868 11150
rect 28816 11086 28868 11092
rect 28908 11144 28960 11150
rect 28908 11086 28960 11092
rect 28920 10996 28948 11086
rect 28828 10968 28948 10996
rect 29092 11008 29144 11014
rect 28828 10538 28856 10968
rect 29092 10950 29144 10956
rect 29104 10742 29132 10950
rect 29092 10736 29144 10742
rect 29092 10678 29144 10684
rect 29000 10600 29052 10606
rect 29000 10542 29052 10548
rect 28816 10532 28868 10538
rect 28816 10474 28868 10480
rect 28828 8537 28856 10474
rect 28908 9988 28960 9994
rect 28908 9930 28960 9936
rect 28920 8634 28948 9930
rect 29012 9654 29040 10542
rect 29288 9926 29316 12650
rect 29276 9920 29328 9926
rect 29276 9862 29328 9868
rect 29000 9648 29052 9654
rect 29000 9590 29052 9596
rect 28908 8628 28960 8634
rect 28908 8570 28960 8576
rect 28814 8528 28870 8537
rect 28814 8463 28870 8472
rect 29012 8430 29040 9590
rect 29184 9580 29236 9586
rect 29184 9522 29236 9528
rect 29092 8832 29144 8838
rect 29092 8774 29144 8780
rect 29000 8424 29052 8430
rect 29000 8366 29052 8372
rect 29104 7954 29132 8774
rect 29092 7948 29144 7954
rect 29092 7890 29144 7896
rect 28816 7880 28868 7886
rect 28816 7822 28868 7828
rect 28828 6322 28856 7822
rect 29196 7818 29224 9522
rect 29276 8492 29328 8498
rect 29276 8434 29328 8440
rect 29184 7812 29236 7818
rect 29184 7754 29236 7760
rect 29000 7744 29052 7750
rect 29000 7686 29052 7692
rect 29012 7206 29040 7686
rect 29000 7200 29052 7206
rect 29000 7142 29052 7148
rect 29012 6866 29040 7142
rect 29000 6860 29052 6866
rect 29000 6802 29052 6808
rect 29090 6760 29146 6769
rect 29090 6695 29146 6704
rect 28816 6316 28868 6322
rect 28816 6258 28868 6264
rect 28998 6216 29054 6225
rect 28998 6151 29000 6160
rect 29052 6151 29054 6160
rect 29000 6122 29052 6128
rect 28724 6112 28776 6118
rect 28724 6054 28776 6060
rect 28448 4684 28500 4690
rect 28448 4626 28500 4632
rect 28172 4558 28224 4564
rect 28262 4584 28318 4593
rect 28000 4486 28028 4558
rect 28262 4519 28318 4528
rect 27988 4480 28040 4486
rect 27988 4422 28040 4428
rect 28264 4480 28316 4486
rect 28264 4422 28316 4428
rect 28000 4282 28028 4422
rect 27988 4276 28040 4282
rect 27988 4218 28040 4224
rect 27896 4208 27948 4214
rect 27896 4150 27948 4156
rect 27896 3732 27948 3738
rect 27896 3674 27948 3680
rect 27908 3126 27936 3674
rect 27896 3120 27948 3126
rect 27896 3062 27948 3068
rect 27988 944 28040 950
rect 27988 886 28040 892
rect 28000 800 28028 886
rect 28276 800 28304 4422
rect 28540 4208 28592 4214
rect 28540 4150 28592 4156
rect 28552 800 28580 4150
rect 28908 3528 28960 3534
rect 28906 3496 28908 3505
rect 28960 3496 28962 3505
rect 28906 3431 28962 3440
rect 28816 3392 28868 3398
rect 28816 3334 28868 3340
rect 28724 2848 28776 2854
rect 28724 2790 28776 2796
rect 28736 2446 28764 2790
rect 28724 2440 28776 2446
rect 28724 2382 28776 2388
rect 28828 800 28856 3334
rect 29104 2990 29132 6695
rect 29196 6458 29224 7754
rect 29288 6866 29316 8434
rect 29276 6860 29328 6866
rect 29276 6802 29328 6808
rect 29184 6452 29236 6458
rect 29184 6394 29236 6400
rect 29184 5704 29236 5710
rect 29184 5646 29236 5652
rect 29196 5574 29224 5646
rect 29184 5568 29236 5574
rect 29184 5510 29236 5516
rect 29196 5370 29224 5510
rect 29184 5364 29236 5370
rect 29184 5306 29236 5312
rect 29184 5228 29236 5234
rect 29184 5170 29236 5176
rect 29196 4146 29224 5170
rect 29184 4140 29236 4146
rect 29184 4082 29236 4088
rect 29380 3670 29408 19382
rect 29564 18698 29592 22066
rect 29734 21584 29790 21593
rect 29734 21519 29736 21528
rect 29788 21519 29790 21528
rect 29736 21490 29788 21496
rect 29840 21486 29868 22986
rect 30208 22778 30236 29446
rect 30300 28490 30328 30670
rect 30380 30592 30432 30598
rect 30380 30534 30432 30540
rect 30392 30258 30420 30534
rect 30380 30252 30432 30258
rect 30380 30194 30432 30200
rect 30392 29782 30420 30194
rect 30380 29776 30432 29782
rect 30380 29718 30432 29724
rect 30380 28688 30432 28694
rect 30380 28630 30432 28636
rect 30288 28484 30340 28490
rect 30288 28426 30340 28432
rect 30300 28014 30328 28426
rect 30288 28008 30340 28014
rect 30288 27950 30340 27956
rect 30392 27606 30420 28630
rect 30484 28626 30512 31726
rect 30748 30932 30800 30938
rect 30748 30874 30800 30880
rect 30564 30048 30616 30054
rect 30564 29990 30616 29996
rect 30576 29578 30604 29990
rect 30564 29572 30616 29578
rect 30564 29514 30616 29520
rect 30472 28620 30524 28626
rect 30472 28562 30524 28568
rect 30484 28082 30512 28562
rect 30472 28076 30524 28082
rect 30472 28018 30524 28024
rect 30484 27674 30512 28018
rect 30472 27668 30524 27674
rect 30472 27610 30524 27616
rect 30380 27600 30432 27606
rect 30380 27542 30432 27548
rect 30656 27464 30708 27470
rect 30656 27406 30708 27412
rect 30668 27130 30696 27406
rect 30656 27124 30708 27130
rect 30656 27066 30708 27072
rect 30564 27056 30616 27062
rect 30562 27024 30564 27033
rect 30616 27024 30618 27033
rect 30668 26994 30696 27066
rect 30760 26994 30788 30874
rect 30840 30388 30892 30394
rect 30840 30330 30892 30336
rect 30562 26959 30618 26968
rect 30656 26988 30708 26994
rect 30656 26930 30708 26936
rect 30748 26988 30800 26994
rect 30748 26930 30800 26936
rect 30668 26382 30696 26930
rect 30852 26738 30880 30330
rect 30944 28966 30972 49030
rect 31220 48142 31248 57190
rect 31576 57044 31628 57050
rect 31576 56986 31628 56992
rect 31392 49156 31444 49162
rect 31392 49098 31444 49104
rect 31404 48754 31432 49098
rect 31588 48754 31616 56986
rect 31392 48748 31444 48754
rect 31392 48690 31444 48696
rect 31576 48748 31628 48754
rect 31576 48690 31628 48696
rect 33048 48680 33100 48686
rect 33048 48622 33100 48628
rect 31484 48612 31536 48618
rect 31484 48554 31536 48560
rect 31392 48272 31444 48278
rect 31392 48214 31444 48220
rect 31404 48142 31432 48214
rect 31496 48142 31524 48554
rect 31208 48136 31260 48142
rect 31208 48078 31260 48084
rect 31392 48136 31444 48142
rect 31392 48078 31444 48084
rect 31484 48136 31536 48142
rect 31484 48078 31536 48084
rect 31300 48068 31352 48074
rect 31300 48010 31352 48016
rect 31024 47660 31076 47666
rect 31024 47602 31076 47608
rect 31036 46510 31064 47602
rect 31312 47054 31340 48010
rect 31496 47666 31524 48078
rect 31668 48000 31720 48006
rect 31668 47942 31720 47948
rect 31484 47660 31536 47666
rect 31484 47602 31536 47608
rect 31392 47456 31444 47462
rect 31392 47398 31444 47404
rect 31300 47048 31352 47054
rect 31300 46990 31352 46996
rect 31024 46504 31076 46510
rect 31024 46446 31076 46452
rect 31036 42362 31064 46446
rect 31024 42356 31076 42362
rect 31024 42298 31076 42304
rect 31404 40526 31432 47398
rect 31392 40520 31444 40526
rect 31392 40462 31444 40468
rect 31484 40384 31536 40390
rect 31484 40326 31536 40332
rect 31496 38758 31524 40326
rect 31484 38752 31536 38758
rect 31484 38694 31536 38700
rect 31680 36938 31708 47942
rect 33060 47666 33088 48622
rect 32956 47660 33008 47666
rect 32956 47602 33008 47608
rect 33048 47660 33100 47666
rect 33048 47602 33100 47608
rect 32680 47048 32732 47054
rect 32680 46990 32732 46996
rect 32312 46980 32364 46986
rect 32312 46922 32364 46928
rect 32324 46578 32352 46922
rect 32692 46578 32720 46990
rect 32312 46572 32364 46578
rect 32312 46514 32364 46520
rect 32680 46572 32732 46578
rect 32680 46514 32732 46520
rect 32312 46368 32364 46374
rect 32312 46310 32364 46316
rect 32324 45490 32352 46310
rect 32968 45554 32996 47602
rect 32678 45520 32734 45529
rect 32968 45526 33088 45554
rect 32312 45484 32364 45490
rect 32312 45426 32364 45432
rect 32404 45484 32456 45490
rect 32404 45426 32456 45432
rect 32588 45484 32640 45490
rect 32678 45455 32680 45464
rect 32588 45426 32640 45432
rect 32732 45455 32734 45464
rect 32680 45426 32732 45432
rect 32416 45082 32444 45426
rect 32600 45354 32628 45426
rect 32588 45348 32640 45354
rect 32588 45290 32640 45296
rect 32404 45076 32456 45082
rect 32404 45018 32456 45024
rect 31852 41744 31904 41750
rect 31852 41686 31904 41692
rect 31496 36910 31708 36938
rect 31024 36644 31076 36650
rect 31024 36586 31076 36592
rect 31036 36174 31064 36586
rect 31024 36168 31076 36174
rect 31024 36110 31076 36116
rect 31392 36168 31444 36174
rect 31392 36110 31444 36116
rect 31300 36100 31352 36106
rect 31300 36042 31352 36048
rect 31208 30252 31260 30258
rect 31208 30194 31260 30200
rect 31024 29164 31076 29170
rect 31024 29106 31076 29112
rect 30932 28960 30984 28966
rect 30932 28902 30984 28908
rect 30932 27464 30984 27470
rect 30932 27406 30984 27412
rect 30944 26926 30972 27406
rect 31036 27130 31064 29106
rect 31114 28112 31170 28121
rect 31114 28047 31170 28056
rect 31128 28014 31156 28047
rect 31116 28008 31168 28014
rect 31116 27950 31168 27956
rect 31024 27124 31076 27130
rect 31024 27066 31076 27072
rect 30932 26920 30984 26926
rect 30932 26862 30984 26868
rect 30852 26710 31064 26738
rect 30656 26376 30708 26382
rect 30656 26318 30708 26324
rect 30748 26308 30800 26314
rect 30748 26250 30800 26256
rect 30288 26240 30340 26246
rect 30288 26182 30340 26188
rect 30300 25906 30328 26182
rect 30288 25900 30340 25906
rect 30288 25842 30340 25848
rect 30380 25900 30432 25906
rect 30380 25842 30432 25848
rect 30392 24410 30420 25842
rect 30564 25832 30616 25838
rect 30564 25774 30616 25780
rect 30380 24404 30432 24410
rect 30380 24346 30432 24352
rect 30288 24200 30340 24206
rect 30286 24168 30288 24177
rect 30340 24168 30342 24177
rect 30286 24103 30342 24112
rect 30196 22772 30248 22778
rect 30196 22714 30248 22720
rect 30288 22636 30340 22642
rect 30288 22578 30340 22584
rect 30012 22432 30064 22438
rect 30012 22374 30064 22380
rect 29828 21480 29880 21486
rect 29828 21422 29880 21428
rect 29736 20936 29788 20942
rect 29736 20878 29788 20884
rect 29748 20466 29776 20878
rect 30024 20874 30052 22374
rect 30300 21690 30328 22578
rect 30380 22432 30432 22438
rect 30380 22374 30432 22380
rect 30288 21684 30340 21690
rect 30288 21626 30340 21632
rect 30286 21448 30342 21457
rect 30286 21383 30342 21392
rect 30300 21350 30328 21383
rect 30288 21344 30340 21350
rect 30288 21286 30340 21292
rect 30012 20868 30064 20874
rect 30012 20810 30064 20816
rect 29736 20460 29788 20466
rect 29736 20402 29788 20408
rect 30392 19938 30420 22374
rect 30470 21856 30526 21865
rect 30470 21791 30526 21800
rect 30300 19910 30420 19938
rect 30300 19854 30328 19910
rect 30288 19848 30340 19854
rect 30288 19790 30340 19796
rect 30484 19786 30512 21791
rect 30472 19780 30524 19786
rect 30472 19722 30524 19728
rect 29552 18692 29604 18698
rect 29552 18634 29604 18640
rect 29564 18426 29592 18634
rect 29552 18420 29604 18426
rect 29552 18362 29604 18368
rect 29644 18420 29696 18426
rect 29644 18362 29696 18368
rect 29656 18290 29684 18362
rect 29644 18284 29696 18290
rect 29644 18226 29696 18232
rect 30380 18284 30432 18290
rect 30380 18226 30432 18232
rect 30104 18080 30156 18086
rect 30104 18022 30156 18028
rect 30116 17678 30144 18022
rect 30104 17672 30156 17678
rect 30104 17614 30156 17620
rect 30012 17536 30064 17542
rect 30012 17478 30064 17484
rect 30024 17270 30052 17478
rect 30012 17264 30064 17270
rect 30012 17206 30064 17212
rect 29736 16992 29788 16998
rect 29736 16934 29788 16940
rect 29552 14816 29604 14822
rect 29550 14784 29552 14793
rect 29644 14816 29696 14822
rect 29604 14784 29606 14793
rect 29644 14758 29696 14764
rect 29550 14719 29606 14728
rect 29656 14550 29684 14758
rect 29644 14544 29696 14550
rect 29644 14486 29696 14492
rect 29460 14408 29512 14414
rect 29460 14350 29512 14356
rect 29472 12986 29500 14350
rect 29552 14340 29604 14346
rect 29552 14282 29604 14288
rect 29564 13938 29592 14282
rect 29656 13938 29684 14486
rect 29552 13932 29604 13938
rect 29552 13874 29604 13880
rect 29644 13932 29696 13938
rect 29644 13874 29696 13880
rect 29460 12980 29512 12986
rect 29460 12922 29512 12928
rect 29748 12850 29776 16934
rect 30104 16516 30156 16522
rect 30104 16458 30156 16464
rect 30012 15700 30064 15706
rect 30012 15642 30064 15648
rect 29828 15360 29880 15366
rect 29828 15302 29880 15308
rect 29920 15360 29972 15366
rect 29920 15302 29972 15308
rect 29840 14498 29868 15302
rect 29932 15026 29960 15302
rect 29920 15020 29972 15026
rect 29920 14962 29972 14968
rect 29840 14470 29960 14498
rect 29828 14340 29880 14346
rect 29828 14282 29880 14288
rect 29840 14006 29868 14282
rect 29828 14000 29880 14006
rect 29828 13942 29880 13948
rect 29736 12844 29788 12850
rect 29736 12786 29788 12792
rect 29840 12434 29868 13942
rect 29932 13938 29960 14470
rect 29920 13932 29972 13938
rect 29920 13874 29972 13880
rect 30024 13734 30052 15642
rect 30116 15162 30144 16458
rect 30392 15910 30420 18226
rect 30288 15904 30340 15910
rect 30288 15846 30340 15852
rect 30380 15904 30432 15910
rect 30380 15846 30432 15852
rect 30196 15496 30248 15502
rect 30196 15438 30248 15444
rect 30104 15156 30156 15162
rect 30104 15098 30156 15104
rect 30208 14346 30236 15438
rect 30104 14340 30156 14346
rect 30104 14282 30156 14288
rect 30196 14340 30248 14346
rect 30196 14282 30248 14288
rect 30116 13870 30144 14282
rect 30208 14074 30236 14282
rect 30196 14068 30248 14074
rect 30196 14010 30248 14016
rect 30104 13864 30156 13870
rect 30104 13806 30156 13812
rect 30012 13728 30064 13734
rect 30012 13670 30064 13676
rect 30024 12986 30052 13670
rect 30116 13433 30144 13806
rect 30102 13424 30158 13433
rect 30102 13359 30158 13368
rect 30300 13326 30328 15846
rect 30378 15056 30434 15065
rect 30378 14991 30434 15000
rect 30392 13802 30420 14991
rect 30380 13796 30432 13802
rect 30380 13738 30432 13744
rect 30288 13320 30340 13326
rect 30288 13262 30340 13268
rect 30392 13190 30420 13738
rect 30380 13184 30432 13190
rect 30380 13126 30432 13132
rect 30012 12980 30064 12986
rect 30012 12922 30064 12928
rect 30288 12844 30340 12850
rect 30288 12786 30340 12792
rect 30380 12844 30432 12850
rect 30380 12786 30432 12792
rect 29564 12406 29868 12434
rect 29564 11694 29592 12406
rect 30300 12102 30328 12786
rect 30392 12238 30420 12786
rect 30380 12232 30432 12238
rect 30380 12174 30432 12180
rect 30288 12096 30340 12102
rect 30288 12038 30340 12044
rect 29644 11824 29696 11830
rect 29644 11766 29696 11772
rect 29552 11688 29604 11694
rect 29552 11630 29604 11636
rect 29564 10674 29592 11630
rect 29552 10668 29604 10674
rect 29552 10610 29604 10616
rect 29460 9648 29512 9654
rect 29460 9590 29512 9596
rect 29472 6322 29500 9590
rect 29656 9110 29684 11766
rect 29828 11756 29880 11762
rect 29828 11698 29880 11704
rect 29840 11354 29868 11698
rect 30300 11370 30328 12038
rect 29828 11348 29880 11354
rect 29828 11290 29880 11296
rect 29932 11342 30328 11370
rect 29828 11212 29880 11218
rect 29828 11154 29880 11160
rect 29840 10985 29868 11154
rect 29932 11082 29960 11342
rect 30104 11280 30156 11286
rect 30104 11222 30156 11228
rect 30012 11144 30064 11150
rect 30012 11086 30064 11092
rect 29920 11076 29972 11082
rect 29920 11018 29972 11024
rect 29826 10976 29882 10985
rect 29826 10911 29882 10920
rect 30024 10810 30052 11086
rect 30012 10804 30064 10810
rect 30012 10746 30064 10752
rect 30012 9512 30064 9518
rect 30012 9454 30064 9460
rect 29920 9444 29972 9450
rect 29920 9386 29972 9392
rect 29644 9104 29696 9110
rect 29644 9046 29696 9052
rect 29552 9036 29604 9042
rect 29552 8978 29604 8984
rect 29736 9036 29788 9042
rect 29736 8978 29788 8984
rect 29564 8242 29592 8978
rect 29644 8968 29696 8974
rect 29644 8910 29696 8916
rect 29656 8634 29684 8910
rect 29644 8628 29696 8634
rect 29644 8570 29696 8576
rect 29748 8362 29776 8978
rect 29828 8968 29880 8974
rect 29828 8910 29880 8916
rect 29840 8673 29868 8910
rect 29826 8664 29882 8673
rect 29826 8599 29882 8608
rect 29736 8356 29788 8362
rect 29736 8298 29788 8304
rect 29564 8214 29776 8242
rect 29644 6452 29696 6458
rect 29644 6394 29696 6400
rect 29656 6322 29684 6394
rect 29460 6316 29512 6322
rect 29460 6258 29512 6264
rect 29644 6316 29696 6322
rect 29748 6304 29776 8214
rect 29840 6730 29868 8599
rect 29932 8537 29960 9386
rect 29918 8528 29974 8537
rect 29918 8463 29974 8472
rect 29920 8424 29972 8430
rect 29920 8366 29972 8372
rect 29932 7546 29960 8366
rect 29920 7540 29972 7546
rect 29920 7482 29972 7488
rect 30024 7290 30052 9454
rect 30116 7886 30144 11222
rect 30300 10810 30328 11342
rect 30472 11348 30524 11354
rect 30472 11290 30524 11296
rect 30484 11150 30512 11290
rect 30472 11144 30524 11150
rect 30472 11086 30524 11092
rect 30288 10804 30340 10810
rect 30288 10746 30340 10752
rect 30472 10804 30524 10810
rect 30472 10746 30524 10752
rect 30484 10470 30512 10746
rect 30472 10464 30524 10470
rect 30472 10406 30524 10412
rect 30380 10056 30432 10062
rect 30380 9998 30432 10004
rect 30196 9648 30248 9654
rect 30196 9590 30248 9596
rect 30208 8974 30236 9590
rect 30288 9580 30340 9586
rect 30288 9522 30340 9528
rect 30300 9042 30328 9522
rect 30288 9036 30340 9042
rect 30288 8978 30340 8984
rect 30196 8968 30248 8974
rect 30196 8910 30248 8916
rect 30392 8838 30420 9998
rect 30470 9344 30526 9353
rect 30470 9279 30526 9288
rect 30484 8974 30512 9279
rect 30472 8968 30524 8974
rect 30472 8910 30524 8916
rect 30288 8832 30340 8838
rect 30288 8774 30340 8780
rect 30380 8832 30432 8838
rect 30380 8774 30432 8780
rect 30300 8498 30328 8774
rect 30288 8492 30340 8498
rect 30288 8434 30340 8440
rect 30380 8492 30432 8498
rect 30380 8434 30432 8440
rect 30104 7880 30156 7886
rect 30104 7822 30156 7828
rect 29932 7262 30052 7290
rect 29828 6724 29880 6730
rect 29828 6666 29880 6672
rect 29828 6316 29880 6322
rect 29748 6276 29828 6304
rect 29644 6258 29696 6264
rect 29828 6258 29880 6264
rect 29472 4622 29500 6258
rect 29840 5302 29868 6258
rect 29932 5914 29960 7262
rect 30012 7200 30064 7206
rect 30012 7142 30064 7148
rect 29920 5908 29972 5914
rect 29920 5850 29972 5856
rect 30024 5778 30052 7142
rect 30116 5778 30144 7822
rect 30392 7478 30420 8434
rect 30472 8084 30524 8090
rect 30472 8026 30524 8032
rect 30484 7818 30512 8026
rect 30472 7812 30524 7818
rect 30472 7754 30524 7760
rect 30380 7472 30432 7478
rect 30380 7414 30432 7420
rect 30484 7274 30512 7754
rect 30472 7268 30524 7274
rect 30472 7210 30524 7216
rect 30472 6860 30524 6866
rect 30472 6802 30524 6808
rect 30286 6624 30342 6633
rect 30286 6559 30342 6568
rect 30300 6186 30328 6559
rect 30484 6202 30512 6802
rect 30576 6254 30604 25774
rect 30760 25294 30788 26250
rect 30748 25288 30800 25294
rect 30748 25230 30800 25236
rect 31036 25158 31064 26710
rect 31024 25152 31076 25158
rect 31024 25094 31076 25100
rect 30748 24880 30800 24886
rect 30748 24822 30800 24828
rect 30656 23112 30708 23118
rect 30656 23054 30708 23060
rect 30668 21486 30696 23054
rect 30656 21480 30708 21486
rect 30656 21422 30708 21428
rect 30656 21140 30708 21146
rect 30656 21082 30708 21088
rect 30668 20466 30696 21082
rect 30656 20460 30708 20466
rect 30656 20402 30708 20408
rect 30656 19984 30708 19990
rect 30656 19926 30708 19932
rect 30668 19378 30696 19926
rect 30656 19372 30708 19378
rect 30656 19314 30708 19320
rect 30656 18080 30708 18086
rect 30656 18022 30708 18028
rect 30668 17202 30696 18022
rect 30656 17196 30708 17202
rect 30656 17138 30708 17144
rect 30656 15904 30708 15910
rect 30656 15846 30708 15852
rect 30668 15570 30696 15846
rect 30656 15564 30708 15570
rect 30656 15506 30708 15512
rect 30668 13870 30696 15506
rect 30656 13864 30708 13870
rect 30656 13806 30708 13812
rect 30656 13320 30708 13326
rect 30656 13262 30708 13268
rect 30668 12918 30696 13262
rect 30656 12912 30708 12918
rect 30656 12854 30708 12860
rect 30668 11898 30696 12854
rect 30656 11892 30708 11898
rect 30656 11834 30708 11840
rect 30760 11506 30788 24822
rect 31036 24750 31064 25094
rect 31024 24744 31076 24750
rect 31024 24686 31076 24692
rect 31036 24614 31064 24686
rect 31024 24608 31076 24614
rect 31024 24550 31076 24556
rect 30840 22228 30892 22234
rect 30840 22170 30892 22176
rect 30852 21622 30880 22170
rect 31116 22160 31168 22166
rect 31116 22102 31168 22108
rect 30932 22024 30984 22030
rect 30932 21966 30984 21972
rect 30944 21690 30972 21966
rect 31024 21956 31076 21962
rect 31024 21898 31076 21904
rect 31036 21690 31064 21898
rect 30932 21684 30984 21690
rect 30932 21626 30984 21632
rect 31024 21684 31076 21690
rect 31024 21626 31076 21632
rect 30840 21616 30892 21622
rect 30840 21558 30892 21564
rect 31128 21554 31156 22102
rect 31116 21548 31168 21554
rect 31116 21490 31168 21496
rect 30840 21344 30892 21350
rect 30840 21286 30892 21292
rect 30852 20058 30880 21286
rect 31220 21078 31248 30194
rect 31208 21072 31260 21078
rect 31208 21014 31260 21020
rect 31208 20392 31260 20398
rect 31208 20334 31260 20340
rect 31220 20058 31248 20334
rect 30840 20052 30892 20058
rect 30840 19994 30892 20000
rect 31208 20052 31260 20058
rect 31208 19994 31260 20000
rect 31312 19938 31340 36042
rect 31404 35290 31432 36110
rect 31392 35284 31444 35290
rect 31392 35226 31444 35232
rect 31496 32502 31524 36910
rect 31576 35012 31628 35018
rect 31576 34954 31628 34960
rect 31484 32496 31536 32502
rect 31484 32438 31536 32444
rect 31588 31754 31616 34954
rect 31404 31726 31616 31754
rect 31404 29714 31432 31726
rect 31392 29708 31444 29714
rect 31392 29650 31444 29656
rect 31404 26994 31432 29650
rect 31668 29096 31720 29102
rect 31668 29038 31720 29044
rect 31576 28416 31628 28422
rect 31576 28358 31628 28364
rect 31484 28212 31536 28218
rect 31484 28154 31536 28160
rect 31392 26988 31444 26994
rect 31392 26930 31444 26936
rect 31392 23180 31444 23186
rect 31392 23122 31444 23128
rect 31404 22166 31432 23122
rect 31392 22160 31444 22166
rect 31392 22102 31444 22108
rect 31404 22030 31432 22102
rect 31392 22024 31444 22030
rect 31392 21966 31444 21972
rect 31392 21888 31444 21894
rect 31392 21830 31444 21836
rect 31404 21593 31432 21830
rect 31390 21584 31446 21593
rect 31390 21519 31446 21528
rect 31392 21072 31444 21078
rect 31392 21014 31444 21020
rect 31220 19910 31340 19938
rect 30840 16992 30892 16998
rect 30840 16934 30892 16940
rect 30852 16182 30880 16934
rect 31116 16448 31168 16454
rect 31116 16390 31168 16396
rect 30840 16176 30892 16182
rect 30840 16118 30892 16124
rect 31024 16040 31076 16046
rect 31024 15982 31076 15988
rect 31036 15910 31064 15982
rect 31024 15904 31076 15910
rect 31024 15846 31076 15852
rect 31036 15706 31064 15846
rect 31024 15700 31076 15706
rect 31024 15642 31076 15648
rect 31036 15502 31064 15642
rect 30932 15496 30984 15502
rect 30932 15438 30984 15444
rect 31024 15496 31076 15502
rect 31024 15438 31076 15444
rect 30840 14816 30892 14822
rect 30840 14758 30892 14764
rect 30852 14550 30880 14758
rect 30944 14618 30972 15438
rect 31024 15360 31076 15366
rect 31024 15302 31076 15308
rect 30932 14612 30984 14618
rect 30932 14554 30984 14560
rect 30840 14544 30892 14550
rect 30840 14486 30892 14492
rect 31036 14074 31064 15302
rect 31128 14618 31156 16390
rect 31116 14612 31168 14618
rect 31116 14554 31168 14560
rect 31128 14414 31156 14554
rect 31116 14408 31168 14414
rect 31220 14396 31248 19910
rect 31404 19334 31432 21014
rect 31116 14350 31168 14356
rect 31198 14368 31248 14396
rect 31312 19306 31432 19334
rect 31198 14328 31226 14368
rect 31198 14300 31248 14328
rect 31116 14272 31168 14278
rect 31220 14260 31248 14300
rect 31312 14278 31340 19306
rect 31392 16176 31444 16182
rect 31392 16118 31444 16124
rect 31404 15366 31432 16118
rect 31392 15360 31444 15366
rect 31392 15302 31444 15308
rect 31392 14884 31444 14890
rect 31392 14826 31444 14832
rect 31116 14214 31168 14220
rect 31198 14232 31248 14260
rect 31300 14272 31352 14278
rect 31024 14068 31076 14074
rect 31024 14010 31076 14016
rect 31024 12912 31076 12918
rect 31024 12854 31076 12860
rect 31036 12306 31064 12854
rect 31024 12300 31076 12306
rect 31024 12242 31076 12248
rect 30932 12232 30984 12238
rect 30932 12174 30984 12180
rect 30944 12073 30972 12174
rect 31024 12164 31076 12170
rect 31024 12106 31076 12112
rect 30930 12064 30986 12073
rect 30930 11999 30986 12008
rect 31036 11898 31064 12106
rect 31024 11892 31076 11898
rect 31024 11834 31076 11840
rect 30932 11688 30984 11694
rect 30932 11630 30984 11636
rect 30668 11478 30788 11506
rect 30668 9568 30696 11478
rect 30746 11384 30802 11393
rect 30746 11319 30802 11328
rect 30760 9697 30788 11319
rect 30944 11218 30972 11630
rect 30932 11212 30984 11218
rect 30932 11154 30984 11160
rect 31024 9716 31076 9722
rect 30746 9688 30802 9697
rect 31024 9658 31076 9664
rect 30746 9623 30802 9632
rect 30932 9580 30984 9586
rect 30668 9540 30788 9568
rect 30760 9330 30788 9540
rect 30932 9522 30984 9528
rect 30840 9512 30892 9518
rect 30944 9489 30972 9522
rect 30840 9454 30892 9460
rect 30930 9480 30986 9489
rect 30852 9353 30880 9454
rect 30930 9415 30986 9424
rect 30673 9302 30788 9330
rect 30838 9344 30894 9353
rect 30673 9194 30701 9302
rect 30838 9279 30894 9288
rect 30668 9166 30701 9194
rect 30668 8786 30696 9166
rect 30668 8758 30788 8786
rect 30656 8628 30708 8634
rect 30656 8570 30708 8576
rect 30668 7886 30696 8570
rect 30656 7880 30708 7886
rect 30656 7822 30708 7828
rect 30760 7546 30788 8758
rect 30930 7576 30986 7585
rect 30748 7540 30800 7546
rect 30930 7511 30986 7520
rect 30748 7482 30800 7488
rect 30656 7472 30708 7478
rect 30656 7414 30708 7420
rect 30668 6866 30696 7414
rect 30944 7410 30972 7511
rect 30932 7404 30984 7410
rect 30932 7346 30984 7352
rect 30748 7336 30800 7342
rect 30748 7278 30800 7284
rect 30760 6882 30788 7278
rect 31036 7274 31064 9658
rect 31128 9450 31156 14214
rect 31198 14090 31226 14232
rect 31300 14214 31352 14220
rect 31198 14062 31340 14090
rect 31208 9988 31260 9994
rect 31208 9930 31260 9936
rect 31220 9568 31248 9930
rect 31312 9625 31340 14062
rect 31404 13938 31432 14826
rect 31392 13932 31444 13938
rect 31392 13874 31444 13880
rect 31496 11540 31524 28154
rect 31588 25242 31616 28358
rect 31680 27606 31708 29038
rect 31760 28960 31812 28966
rect 31760 28902 31812 28908
rect 31772 28694 31800 28902
rect 31760 28688 31812 28694
rect 31760 28630 31812 28636
rect 31668 27600 31720 27606
rect 31668 27542 31720 27548
rect 31668 26920 31720 26926
rect 31668 26862 31720 26868
rect 31680 26489 31708 26862
rect 31666 26480 31722 26489
rect 31666 26415 31668 26424
rect 31720 26415 31722 26424
rect 31668 26386 31720 26392
rect 31588 25214 31708 25242
rect 31576 22568 31628 22574
rect 31576 22510 31628 22516
rect 31588 22234 31616 22510
rect 31576 22228 31628 22234
rect 31576 22170 31628 22176
rect 31576 21616 31628 21622
rect 31576 21558 31628 21564
rect 31588 21418 31616 21558
rect 31576 21412 31628 21418
rect 31576 21354 31628 21360
rect 31576 17536 31628 17542
rect 31576 17478 31628 17484
rect 31588 17202 31616 17478
rect 31576 17196 31628 17202
rect 31576 17138 31628 17144
rect 31680 17082 31708 25214
rect 31760 17672 31812 17678
rect 31760 17614 31812 17620
rect 31772 17105 31800 17614
rect 31404 11512 31524 11540
rect 31588 17054 31708 17082
rect 31758 17096 31814 17105
rect 31404 9674 31432 11512
rect 31588 9692 31616 17054
rect 31758 17031 31814 17040
rect 31760 15020 31812 15026
rect 31760 14962 31812 14968
rect 31668 14816 31720 14822
rect 31668 14758 31720 14764
rect 31680 14074 31708 14758
rect 31772 14618 31800 14962
rect 31760 14612 31812 14618
rect 31760 14554 31812 14560
rect 31668 14068 31720 14074
rect 31668 14010 31720 14016
rect 31760 13728 31812 13734
rect 31864 13705 31892 41686
rect 32600 35894 32628 45290
rect 32772 45280 32824 45286
rect 32772 45222 32824 45228
rect 32680 39296 32732 39302
rect 32680 39238 32732 39244
rect 32692 38962 32720 39238
rect 32680 38956 32732 38962
rect 32680 38898 32732 38904
rect 32680 38208 32732 38214
rect 32680 38150 32732 38156
rect 32692 37874 32720 38150
rect 32680 37868 32732 37874
rect 32680 37810 32732 37816
rect 32416 35866 32628 35894
rect 32036 35012 32088 35018
rect 32036 34954 32088 34960
rect 32048 34898 32076 34954
rect 32220 34944 32272 34950
rect 32048 34892 32220 34898
rect 32048 34886 32272 34892
rect 32048 34870 32260 34886
rect 32048 29510 32076 34870
rect 32416 34610 32444 35866
rect 32784 35086 32812 45222
rect 33060 38962 33088 45526
rect 32864 38956 32916 38962
rect 32864 38898 32916 38904
rect 33048 38956 33100 38962
rect 33048 38898 33100 38904
rect 32876 37874 32904 38898
rect 33060 38418 33088 38898
rect 33048 38412 33100 38418
rect 33048 38354 33100 38360
rect 33060 37874 33088 38354
rect 33232 38344 33284 38350
rect 33232 38286 33284 38292
rect 32864 37868 32916 37874
rect 32864 37810 32916 37816
rect 33048 37868 33100 37874
rect 33048 37810 33100 37816
rect 32876 36106 32904 37810
rect 32864 36100 32916 36106
rect 32864 36042 32916 36048
rect 33244 35714 33272 38286
rect 33428 35834 33456 57190
rect 34808 48074 34836 57190
rect 34934 57148 35242 57157
rect 34934 57146 34940 57148
rect 34996 57146 35020 57148
rect 35076 57146 35100 57148
rect 35156 57146 35180 57148
rect 35236 57146 35242 57148
rect 34996 57094 34998 57146
rect 35178 57094 35180 57146
rect 34934 57092 34940 57094
rect 34996 57092 35020 57094
rect 35076 57092 35100 57094
rect 35156 57092 35180 57094
rect 35236 57092 35242 57094
rect 34934 57083 35242 57092
rect 34934 56060 35242 56069
rect 34934 56058 34940 56060
rect 34996 56058 35020 56060
rect 35076 56058 35100 56060
rect 35156 56058 35180 56060
rect 35236 56058 35242 56060
rect 34996 56006 34998 56058
rect 35178 56006 35180 56058
rect 34934 56004 34940 56006
rect 34996 56004 35020 56006
rect 35076 56004 35100 56006
rect 35156 56004 35180 56006
rect 35236 56004 35242 56006
rect 34934 55995 35242 56004
rect 34934 54972 35242 54981
rect 34934 54970 34940 54972
rect 34996 54970 35020 54972
rect 35076 54970 35100 54972
rect 35156 54970 35180 54972
rect 35236 54970 35242 54972
rect 34996 54918 34998 54970
rect 35178 54918 35180 54970
rect 34934 54916 34940 54918
rect 34996 54916 35020 54918
rect 35076 54916 35100 54918
rect 35156 54916 35180 54918
rect 35236 54916 35242 54918
rect 34934 54907 35242 54916
rect 34934 53884 35242 53893
rect 34934 53882 34940 53884
rect 34996 53882 35020 53884
rect 35076 53882 35100 53884
rect 35156 53882 35180 53884
rect 35236 53882 35242 53884
rect 34996 53830 34998 53882
rect 35178 53830 35180 53882
rect 34934 53828 34940 53830
rect 34996 53828 35020 53830
rect 35076 53828 35100 53830
rect 35156 53828 35180 53830
rect 35236 53828 35242 53830
rect 34934 53819 35242 53828
rect 34934 52796 35242 52805
rect 34934 52794 34940 52796
rect 34996 52794 35020 52796
rect 35076 52794 35100 52796
rect 35156 52794 35180 52796
rect 35236 52794 35242 52796
rect 34996 52742 34998 52794
rect 35178 52742 35180 52794
rect 34934 52740 34940 52742
rect 34996 52740 35020 52742
rect 35076 52740 35100 52742
rect 35156 52740 35180 52742
rect 35236 52740 35242 52742
rect 34934 52731 35242 52740
rect 34934 51708 35242 51717
rect 34934 51706 34940 51708
rect 34996 51706 35020 51708
rect 35076 51706 35100 51708
rect 35156 51706 35180 51708
rect 35236 51706 35242 51708
rect 34996 51654 34998 51706
rect 35178 51654 35180 51706
rect 34934 51652 34940 51654
rect 34996 51652 35020 51654
rect 35076 51652 35100 51654
rect 35156 51652 35180 51654
rect 35236 51652 35242 51654
rect 34934 51643 35242 51652
rect 34934 50620 35242 50629
rect 34934 50618 34940 50620
rect 34996 50618 35020 50620
rect 35076 50618 35100 50620
rect 35156 50618 35180 50620
rect 35236 50618 35242 50620
rect 34996 50566 34998 50618
rect 35178 50566 35180 50618
rect 34934 50564 34940 50566
rect 34996 50564 35020 50566
rect 35076 50564 35100 50566
rect 35156 50564 35180 50566
rect 35236 50564 35242 50566
rect 34934 50555 35242 50564
rect 34934 49532 35242 49541
rect 34934 49530 34940 49532
rect 34996 49530 35020 49532
rect 35076 49530 35100 49532
rect 35156 49530 35180 49532
rect 35236 49530 35242 49532
rect 34996 49478 34998 49530
rect 35178 49478 35180 49530
rect 34934 49476 34940 49478
rect 34996 49476 35020 49478
rect 35076 49476 35100 49478
rect 35156 49476 35180 49478
rect 35236 49476 35242 49478
rect 34934 49467 35242 49476
rect 34934 48444 35242 48453
rect 34934 48442 34940 48444
rect 34996 48442 35020 48444
rect 35076 48442 35100 48444
rect 35156 48442 35180 48444
rect 35236 48442 35242 48444
rect 34996 48390 34998 48442
rect 35178 48390 35180 48442
rect 34934 48388 34940 48390
rect 34996 48388 35020 48390
rect 35076 48388 35100 48390
rect 35156 48388 35180 48390
rect 35236 48388 35242 48390
rect 34934 48379 35242 48388
rect 34888 48136 34940 48142
rect 34888 48078 34940 48084
rect 34796 48068 34848 48074
rect 34796 48010 34848 48016
rect 34900 47802 34928 48078
rect 35440 48000 35492 48006
rect 35440 47942 35492 47948
rect 34888 47796 34940 47802
rect 34888 47738 34940 47744
rect 35348 47796 35400 47802
rect 35348 47738 35400 47744
rect 34934 47356 35242 47365
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47291 35242 47300
rect 34934 46268 35242 46277
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46203 35242 46212
rect 34934 45180 35242 45189
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45115 35242 45124
rect 34934 44092 35242 44101
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44027 35242 44036
rect 33784 43444 33836 43450
rect 33784 43386 33836 43392
rect 33508 42084 33560 42090
rect 33508 42026 33560 42032
rect 33416 35828 33468 35834
rect 33416 35770 33468 35776
rect 33060 35686 33272 35714
rect 33324 35692 33376 35698
rect 32772 35080 32824 35086
rect 32772 35022 32824 35028
rect 32956 35012 33008 35018
rect 32956 34954 33008 34960
rect 32772 34944 32824 34950
rect 32772 34886 32824 34892
rect 32784 34610 32812 34886
rect 32968 34610 32996 34954
rect 32404 34604 32456 34610
rect 32404 34546 32456 34552
rect 32496 34604 32548 34610
rect 32496 34546 32548 34552
rect 32772 34604 32824 34610
rect 32772 34546 32824 34552
rect 32956 34604 33008 34610
rect 32956 34546 33008 34552
rect 32128 30660 32180 30666
rect 32128 30602 32180 30608
rect 32140 30258 32168 30602
rect 32128 30252 32180 30258
rect 32128 30194 32180 30200
rect 32508 29594 32536 34546
rect 32784 33930 32812 34546
rect 32772 33924 32824 33930
rect 32772 33866 32824 33872
rect 33060 33402 33088 35686
rect 33324 35634 33376 35640
rect 33416 35692 33468 35698
rect 33416 35634 33468 35640
rect 33140 35488 33192 35494
rect 33140 35430 33192 35436
rect 33152 35086 33180 35430
rect 33232 35148 33284 35154
rect 33232 35090 33284 35096
rect 33140 35080 33192 35086
rect 33140 35022 33192 35028
rect 33244 34898 33272 35090
rect 33152 34870 33272 34898
rect 33152 33522 33180 34870
rect 33232 33652 33284 33658
rect 33232 33594 33284 33600
rect 33140 33516 33192 33522
rect 33140 33458 33192 33464
rect 33060 33374 33180 33402
rect 32588 30048 32640 30054
rect 32588 29990 32640 29996
rect 32600 29782 32628 29990
rect 32588 29776 32640 29782
rect 32588 29718 32640 29724
rect 32588 29640 32640 29646
rect 32508 29588 32588 29594
rect 32508 29582 32640 29588
rect 32508 29566 32628 29582
rect 32036 29504 32088 29510
rect 32036 29446 32088 29452
rect 31944 28416 31996 28422
rect 31944 28358 31996 28364
rect 31760 13670 31812 13676
rect 31850 13696 31906 13705
rect 31772 13002 31800 13670
rect 31850 13631 31906 13640
rect 31772 12974 31892 13002
rect 31668 12844 31720 12850
rect 31720 12804 31800 12832
rect 31668 12786 31720 12792
rect 31772 12238 31800 12804
rect 31760 12232 31812 12238
rect 31760 12174 31812 12180
rect 31864 11778 31892 12974
rect 31680 11750 31892 11778
rect 31576 9686 31628 9692
rect 31404 9646 31524 9674
rect 31198 9540 31248 9568
rect 31298 9616 31354 9625
rect 31496 9602 31524 9646
rect 31576 9628 31628 9634
rect 31680 9636 31708 11750
rect 31852 11688 31904 11694
rect 31852 11630 31904 11636
rect 31864 11558 31892 11630
rect 31852 11552 31904 11558
rect 31852 11494 31904 11500
rect 31956 11150 31984 28358
rect 32220 27464 32272 27470
rect 32220 27406 32272 27412
rect 32312 27464 32364 27470
rect 32312 27406 32364 27412
rect 32036 27056 32088 27062
rect 32034 27024 32036 27033
rect 32088 27024 32090 27033
rect 32034 26959 32090 26968
rect 32232 25770 32260 27406
rect 32220 25764 32272 25770
rect 32220 25706 32272 25712
rect 32324 24177 32352 27406
rect 32600 26858 32628 29566
rect 33152 27674 33180 33374
rect 33140 27668 33192 27674
rect 33140 27610 33192 27616
rect 32772 26988 32824 26994
rect 32772 26930 32824 26936
rect 32956 26988 33008 26994
rect 32956 26930 33008 26936
rect 33140 26988 33192 26994
rect 33140 26930 33192 26936
rect 32588 26852 32640 26858
rect 32588 26794 32640 26800
rect 32600 26042 32628 26794
rect 32588 26036 32640 26042
rect 32588 25978 32640 25984
rect 32784 24886 32812 26930
rect 32968 26450 32996 26930
rect 33152 26489 33180 26930
rect 33138 26480 33194 26489
rect 32956 26444 33008 26450
rect 33138 26415 33194 26424
rect 32956 26386 33008 26392
rect 32772 24880 32824 24886
rect 32772 24822 32824 24828
rect 33152 24342 33180 26415
rect 33140 24336 33192 24342
rect 33140 24278 33192 24284
rect 32310 24168 32366 24177
rect 32310 24103 32366 24112
rect 32036 24064 32088 24070
rect 32036 24006 32088 24012
rect 31944 11144 31996 11150
rect 31944 11086 31996 11092
rect 31680 9608 31892 9636
rect 31298 9551 31354 9560
rect 31404 9574 31524 9602
rect 31576 9580 31628 9586
rect 31116 9444 31168 9450
rect 31116 9386 31168 9392
rect 31198 9364 31226 9540
rect 31198 9336 31248 9364
rect 31116 8968 31168 8974
rect 31116 8910 31168 8916
rect 31128 8106 31156 8910
rect 31220 8498 31248 9336
rect 31298 8800 31354 8809
rect 31298 8735 31354 8744
rect 31208 8492 31260 8498
rect 31208 8434 31260 8440
rect 31128 8078 31248 8106
rect 31116 7336 31168 7342
rect 31116 7278 31168 7284
rect 30932 7268 30984 7274
rect 30932 7210 30984 7216
rect 31024 7268 31076 7274
rect 31024 7210 31076 7216
rect 30944 7177 30972 7210
rect 30930 7168 30986 7177
rect 30930 7103 30986 7112
rect 30656 6860 30708 6866
rect 30760 6854 30880 6882
rect 30656 6802 30708 6808
rect 30668 6322 30696 6802
rect 30748 6792 30800 6798
rect 30748 6734 30800 6740
rect 30760 6322 30788 6734
rect 30852 6458 30880 6854
rect 31036 6798 31064 7210
rect 31024 6792 31076 6798
rect 31024 6734 31076 6740
rect 31024 6656 31076 6662
rect 31024 6598 31076 6604
rect 30840 6452 30892 6458
rect 30840 6394 30892 6400
rect 30656 6316 30708 6322
rect 30656 6258 30708 6264
rect 30748 6316 30800 6322
rect 30748 6258 30800 6264
rect 30288 6180 30340 6186
rect 30288 6122 30340 6128
rect 30392 6174 30512 6202
rect 30564 6248 30616 6254
rect 30564 6190 30616 6196
rect 30012 5772 30064 5778
rect 30012 5714 30064 5720
rect 30104 5772 30156 5778
rect 30104 5714 30156 5720
rect 30104 5636 30156 5642
rect 30104 5578 30156 5584
rect 29828 5296 29880 5302
rect 29828 5238 29880 5244
rect 29460 4616 29512 4622
rect 29460 4558 29512 4564
rect 29552 4548 29604 4554
rect 29552 4490 29604 4496
rect 29564 4214 29592 4490
rect 29552 4208 29604 4214
rect 29552 4150 29604 4156
rect 29368 3664 29420 3670
rect 29368 3606 29420 3612
rect 29736 3392 29788 3398
rect 29736 3334 29788 3340
rect 29748 3058 29776 3334
rect 29840 3126 29868 5238
rect 30116 5166 30144 5578
rect 30392 5574 30420 6174
rect 30380 5568 30432 5574
rect 30380 5510 30432 5516
rect 30104 5160 30156 5166
rect 30104 5102 30156 5108
rect 30196 5024 30248 5030
rect 30196 4966 30248 4972
rect 30012 4140 30064 4146
rect 30012 4082 30064 4088
rect 30024 3398 30052 4082
rect 30012 3392 30064 3398
rect 30208 3380 30236 4966
rect 30392 4078 30420 5510
rect 30472 4276 30524 4282
rect 30472 4218 30524 4224
rect 30380 4072 30432 4078
rect 30380 4014 30432 4020
rect 30288 3936 30340 3942
rect 30288 3878 30340 3884
rect 30300 3534 30328 3878
rect 30392 3602 30420 4014
rect 30484 3602 30512 4218
rect 30380 3596 30432 3602
rect 30380 3538 30432 3544
rect 30472 3596 30524 3602
rect 30472 3538 30524 3544
rect 30288 3528 30340 3534
rect 30288 3470 30340 3476
rect 30288 3392 30340 3398
rect 30208 3352 30288 3380
rect 30012 3334 30064 3340
rect 30288 3334 30340 3340
rect 29828 3120 29880 3126
rect 29828 3062 29880 3068
rect 29368 3052 29420 3058
rect 29368 2994 29420 3000
rect 29736 3052 29788 3058
rect 29736 2994 29788 3000
rect 29092 2984 29144 2990
rect 29092 2926 29144 2932
rect 28908 2304 28960 2310
rect 28908 2246 28960 2252
rect 28920 864 28948 2246
rect 28920 836 29132 864
rect 29104 800 29132 836
rect 29380 800 29408 2994
rect 29644 2984 29696 2990
rect 29644 2926 29696 2932
rect 30196 2984 30248 2990
rect 30196 2926 30248 2932
rect 29656 800 29684 2926
rect 29920 2372 29972 2378
rect 29920 2314 29972 2320
rect 29932 800 29960 2314
rect 30208 800 30236 2926
rect 30300 2446 30328 3334
rect 30288 2440 30340 2446
rect 30288 2382 30340 2388
rect 30472 2372 30524 2378
rect 30472 2314 30524 2320
rect 30484 800 30512 2314
rect 30576 1970 30604 6190
rect 30668 5234 30696 6258
rect 30932 6248 30984 6254
rect 30932 6190 30984 6196
rect 30944 5914 30972 6190
rect 31036 5914 31064 6598
rect 31128 6390 31156 7278
rect 31116 6384 31168 6390
rect 31116 6326 31168 6332
rect 30840 5908 30892 5914
rect 30840 5850 30892 5856
rect 30932 5908 30984 5914
rect 30932 5850 30984 5856
rect 31024 5908 31076 5914
rect 31024 5850 31076 5856
rect 30656 5228 30708 5234
rect 30656 5170 30708 5176
rect 30748 2984 30800 2990
rect 30748 2926 30800 2932
rect 30564 1964 30616 1970
rect 30564 1906 30616 1912
rect 30760 800 30788 2926
rect 30852 2446 30880 5850
rect 31220 4758 31248 8078
rect 31312 5234 31340 8735
rect 31404 7002 31432 9574
rect 31576 9522 31628 9528
rect 31588 9353 31616 9522
rect 31864 9450 31892 9608
rect 31852 9444 31904 9450
rect 31852 9386 31904 9392
rect 31574 9344 31630 9353
rect 31574 9279 31630 9288
rect 31482 9208 31538 9217
rect 31482 9143 31484 9152
rect 31536 9143 31538 9152
rect 31484 9114 31536 9120
rect 31588 8956 31616 9279
rect 31668 8968 31720 8974
rect 31588 8928 31668 8956
rect 31668 8910 31720 8916
rect 31484 8900 31536 8906
rect 31484 8842 31536 8848
rect 31496 8809 31524 8842
rect 31576 8832 31628 8838
rect 31482 8800 31538 8809
rect 31576 8774 31628 8780
rect 31482 8735 31538 8744
rect 31588 8634 31616 8774
rect 31576 8628 31628 8634
rect 31576 8570 31628 8576
rect 31852 8560 31904 8566
rect 31852 8502 31904 8508
rect 31864 7954 31892 8502
rect 31956 8294 31984 11086
rect 31944 8288 31996 8294
rect 31944 8230 31996 8236
rect 31942 7984 31998 7993
rect 31852 7948 31904 7954
rect 31942 7919 31998 7928
rect 31852 7890 31904 7896
rect 31956 7886 31984 7919
rect 31576 7880 31628 7886
rect 31576 7822 31628 7828
rect 31760 7880 31812 7886
rect 31760 7822 31812 7828
rect 31944 7880 31996 7886
rect 31944 7822 31996 7828
rect 31484 7540 31536 7546
rect 31484 7482 31536 7488
rect 31392 6996 31444 7002
rect 31392 6938 31444 6944
rect 31392 5840 31444 5846
rect 31392 5782 31444 5788
rect 31300 5228 31352 5234
rect 31300 5170 31352 5176
rect 31208 4752 31260 4758
rect 31208 4694 31260 4700
rect 31404 4146 31432 5782
rect 31392 4140 31444 4146
rect 31392 4082 31444 4088
rect 31298 4040 31354 4049
rect 31298 3975 31354 3984
rect 31312 3534 31340 3975
rect 31496 3602 31524 7482
rect 31588 6934 31616 7822
rect 31772 7206 31800 7822
rect 31760 7200 31812 7206
rect 31760 7142 31812 7148
rect 31576 6928 31628 6934
rect 31576 6870 31628 6876
rect 31944 6928 31996 6934
rect 31944 6870 31996 6876
rect 31576 6792 31628 6798
rect 31576 6734 31628 6740
rect 31588 3738 31616 6734
rect 31760 6656 31812 6662
rect 31760 6598 31812 6604
rect 31772 6390 31800 6598
rect 31760 6384 31812 6390
rect 31760 6326 31812 6332
rect 31956 5710 31984 6870
rect 32048 6798 32076 24006
rect 32772 23044 32824 23050
rect 32772 22986 32824 22992
rect 32784 22642 32812 22986
rect 32772 22636 32824 22642
rect 32772 22578 32824 22584
rect 32220 22500 32272 22506
rect 32220 22442 32272 22448
rect 32232 22234 32260 22442
rect 32772 22432 32824 22438
rect 32772 22374 32824 22380
rect 32220 22228 32272 22234
rect 32220 22170 32272 22176
rect 32784 22030 32812 22374
rect 32956 22160 33008 22166
rect 32956 22102 33008 22108
rect 32772 22024 32824 22030
rect 32772 21966 32824 21972
rect 32864 21888 32916 21894
rect 32864 21830 32916 21836
rect 32312 21548 32364 21554
rect 32312 21490 32364 21496
rect 32324 20806 32352 21490
rect 32876 20874 32904 21830
rect 32968 21146 32996 22102
rect 33048 22024 33100 22030
rect 33048 21966 33100 21972
rect 33060 21622 33088 21966
rect 33048 21616 33100 21622
rect 33048 21558 33100 21564
rect 33048 21480 33100 21486
rect 33048 21422 33100 21428
rect 32956 21140 33008 21146
rect 32956 21082 33008 21088
rect 33060 21010 33088 21422
rect 33048 21004 33100 21010
rect 33048 20946 33100 20952
rect 32864 20868 32916 20874
rect 32864 20810 32916 20816
rect 32956 20868 33008 20874
rect 32956 20810 33008 20816
rect 32312 20800 32364 20806
rect 32312 20742 32364 20748
rect 32968 20398 32996 20810
rect 33060 20466 33088 20946
rect 33048 20460 33100 20466
rect 33048 20402 33100 20408
rect 32956 20392 33008 20398
rect 32956 20334 33008 20340
rect 33060 19854 33088 20402
rect 33048 19848 33100 19854
rect 33048 19790 33100 19796
rect 33060 19378 33088 19790
rect 33048 19372 33100 19378
rect 33048 19314 33100 19320
rect 32496 18760 32548 18766
rect 32496 18702 32548 18708
rect 32220 18624 32272 18630
rect 32220 18566 32272 18572
rect 32128 17672 32180 17678
rect 32128 17614 32180 17620
rect 32140 17338 32168 17614
rect 32128 17332 32180 17338
rect 32128 17274 32180 17280
rect 32232 17270 32260 18566
rect 32404 18284 32456 18290
rect 32404 18226 32456 18232
rect 32312 17536 32364 17542
rect 32312 17478 32364 17484
rect 32220 17264 32272 17270
rect 32220 17206 32272 17212
rect 32218 17096 32274 17105
rect 32218 17031 32274 17040
rect 32128 16176 32180 16182
rect 32128 16118 32180 16124
rect 32140 15366 32168 16118
rect 32232 15706 32260 17031
rect 32324 16522 32352 17478
rect 32416 17338 32444 18226
rect 32404 17332 32456 17338
rect 32404 17274 32456 17280
rect 32312 16516 32364 16522
rect 32312 16458 32364 16464
rect 32508 16250 32536 18702
rect 32588 18080 32640 18086
rect 32588 18022 32640 18028
rect 32680 18080 32732 18086
rect 32680 18022 32732 18028
rect 32496 16244 32548 16250
rect 32496 16186 32548 16192
rect 32600 16182 32628 18022
rect 32692 17746 32720 18022
rect 33060 17762 33088 19314
rect 32680 17740 32732 17746
rect 32680 17682 32732 17688
rect 32968 17734 33088 17762
rect 32968 17678 32996 17734
rect 32956 17672 33008 17678
rect 32956 17614 33008 17620
rect 32968 17202 32996 17614
rect 32956 17196 33008 17202
rect 32956 17138 33008 17144
rect 32968 16590 32996 17138
rect 32680 16584 32732 16590
rect 32680 16526 32732 16532
rect 32956 16584 33008 16590
rect 32956 16526 33008 16532
rect 32588 16176 32640 16182
rect 32588 16118 32640 16124
rect 32692 16114 32720 16526
rect 32772 16448 32824 16454
rect 32772 16390 32824 16396
rect 32680 16108 32732 16114
rect 32680 16050 32732 16056
rect 32220 15700 32272 15706
rect 32220 15642 32272 15648
rect 32128 15360 32180 15366
rect 32128 15302 32180 15308
rect 32140 14618 32168 15302
rect 32404 15156 32456 15162
rect 32404 15098 32456 15104
rect 32416 15026 32444 15098
rect 32404 15020 32456 15026
rect 32404 14962 32456 14968
rect 32128 14612 32180 14618
rect 32128 14554 32180 14560
rect 32680 14612 32732 14618
rect 32680 14554 32732 14560
rect 32588 14340 32640 14346
rect 32588 14282 32640 14288
rect 32600 13938 32628 14282
rect 32588 13932 32640 13938
rect 32588 13874 32640 13880
rect 32600 13530 32628 13874
rect 32692 13802 32720 14554
rect 32680 13796 32732 13802
rect 32680 13738 32732 13744
rect 32588 13524 32640 13530
rect 32588 13466 32640 13472
rect 32312 13252 32364 13258
rect 32312 13194 32364 13200
rect 32324 12646 32352 13194
rect 32312 12640 32364 12646
rect 32312 12582 32364 12588
rect 32128 11892 32180 11898
rect 32128 11834 32180 11840
rect 32140 11218 32168 11834
rect 32220 11688 32272 11694
rect 32220 11630 32272 11636
rect 32128 11212 32180 11218
rect 32128 11154 32180 11160
rect 32128 9648 32180 9654
rect 32128 9590 32180 9596
rect 32140 7886 32168 9590
rect 32128 7880 32180 7886
rect 32128 7822 32180 7828
rect 32036 6792 32088 6798
rect 32036 6734 32088 6740
rect 31944 5704 31996 5710
rect 31944 5646 31996 5652
rect 32036 5704 32088 5710
rect 32036 5646 32088 5652
rect 31760 5228 31812 5234
rect 31760 5170 31812 5176
rect 31772 4622 31800 5170
rect 31944 5160 31996 5166
rect 31944 5102 31996 5108
rect 31760 4616 31812 4622
rect 31760 4558 31812 4564
rect 31576 3732 31628 3738
rect 31576 3674 31628 3680
rect 31484 3596 31536 3602
rect 31484 3538 31536 3544
rect 31024 3528 31076 3534
rect 31024 3470 31076 3476
rect 31300 3528 31352 3534
rect 31300 3470 31352 3476
rect 31036 3097 31064 3470
rect 31022 3088 31078 3097
rect 31022 3023 31078 3032
rect 31496 2922 31524 3538
rect 31576 2984 31628 2990
rect 31576 2926 31628 2932
rect 31484 2916 31536 2922
rect 31484 2858 31536 2864
rect 30840 2440 30892 2446
rect 30840 2382 30892 2388
rect 31024 2372 31076 2378
rect 31024 2314 31076 2320
rect 31036 800 31064 2314
rect 31300 944 31352 950
rect 31300 886 31352 892
rect 31312 800 31340 886
rect 31588 800 31616 2926
rect 31772 2378 31800 4558
rect 31852 4548 31904 4554
rect 31852 4490 31904 4496
rect 31864 3058 31892 4490
rect 31852 3052 31904 3058
rect 31852 2994 31904 3000
rect 31956 2446 31984 5102
rect 32048 3534 32076 5646
rect 32128 5636 32180 5642
rect 32128 5578 32180 5584
rect 32140 4706 32168 5578
rect 32232 5234 32260 11630
rect 32324 5284 32352 12582
rect 32404 12368 32456 12374
rect 32404 12310 32456 12316
rect 32416 11150 32444 12310
rect 32680 12232 32732 12238
rect 32680 12174 32732 12180
rect 32496 12096 32548 12102
rect 32496 12038 32548 12044
rect 32508 11762 32536 12038
rect 32692 11762 32720 12174
rect 32784 11762 32812 16390
rect 32956 15496 33008 15502
rect 32956 15438 33008 15444
rect 32862 14784 32918 14793
rect 32862 14719 32918 14728
rect 32876 13938 32904 14719
rect 32864 13932 32916 13938
rect 32864 13874 32916 13880
rect 32968 12238 32996 15438
rect 33244 14414 33272 33594
rect 33336 29782 33364 35634
rect 33428 35154 33456 35634
rect 33416 35148 33468 35154
rect 33416 35090 33468 35096
rect 33416 34944 33468 34950
rect 33416 34886 33468 34892
rect 33324 29776 33376 29782
rect 33324 29718 33376 29724
rect 33428 22094 33456 34886
rect 33520 27470 33548 42026
rect 33692 38752 33744 38758
rect 33692 38694 33744 38700
rect 33600 37664 33652 37670
rect 33600 37606 33652 37612
rect 33612 33522 33640 37606
rect 33704 35698 33732 38694
rect 33692 35692 33744 35698
rect 33692 35634 33744 35640
rect 33692 35148 33744 35154
rect 33692 35090 33744 35096
rect 33704 34678 33732 35090
rect 33692 34672 33744 34678
rect 33692 34614 33744 34620
rect 33796 33930 33824 43386
rect 34934 43004 35242 43013
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42939 35242 42948
rect 34934 41916 35242 41925
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41851 35242 41860
rect 34934 40828 35242 40837
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40763 35242 40772
rect 34934 39740 35242 39749
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39675 35242 39684
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 35360 36553 35388 47738
rect 35452 47666 35480 47942
rect 35440 47660 35492 47666
rect 35440 47602 35492 47608
rect 35532 46436 35584 46442
rect 35532 46378 35584 46384
rect 35544 45898 35572 46378
rect 35532 45892 35584 45898
rect 35532 45834 35584 45840
rect 35544 45626 35572 45834
rect 35532 45620 35584 45626
rect 35532 45562 35584 45568
rect 35636 45558 35664 57190
rect 37108 51406 37136 57190
rect 37280 51876 37332 51882
rect 37280 51818 37332 51824
rect 37292 51406 37320 51818
rect 36912 51400 36964 51406
rect 36912 51342 36964 51348
rect 37096 51400 37148 51406
rect 37096 51342 37148 51348
rect 37280 51400 37332 51406
rect 37280 51342 37332 51348
rect 35716 48340 35768 48346
rect 35716 48282 35768 48288
rect 35900 48340 35952 48346
rect 35900 48282 35952 48288
rect 35728 47054 35756 48282
rect 35912 48142 35940 48282
rect 35900 48136 35952 48142
rect 35900 48078 35952 48084
rect 35900 48000 35952 48006
rect 35900 47942 35952 47948
rect 35716 47048 35768 47054
rect 35716 46990 35768 46996
rect 35624 45552 35676 45558
rect 35624 45494 35676 45500
rect 35728 45490 35756 46990
rect 35912 45558 35940 47942
rect 36924 46170 36952 51342
rect 37188 51332 37240 51338
rect 37188 51274 37240 51280
rect 37200 48142 37228 51274
rect 37556 51264 37608 51270
rect 37556 51206 37608 51212
rect 37188 48136 37240 48142
rect 37188 48078 37240 48084
rect 36912 46164 36964 46170
rect 36912 46106 36964 46112
rect 36820 45960 36872 45966
rect 36820 45902 36872 45908
rect 36832 45558 36860 45902
rect 35900 45552 35952 45558
rect 35900 45494 35952 45500
rect 36820 45552 36872 45558
rect 36820 45494 36872 45500
rect 35716 45484 35768 45490
rect 35716 45426 35768 45432
rect 36452 45280 36504 45286
rect 36452 45222 36504 45228
rect 35346 36544 35402 36553
rect 34934 36476 35242 36485
rect 35346 36479 35402 36488
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 34796 35692 34848 35698
rect 34796 35634 34848 35640
rect 33876 35624 33928 35630
rect 33876 35566 33928 35572
rect 33888 35290 33916 35566
rect 33876 35284 33928 35290
rect 33876 35226 33928 35232
rect 34060 34740 34112 34746
rect 34060 34682 34112 34688
rect 34072 34474 34100 34682
rect 34704 34604 34756 34610
rect 34704 34546 34756 34552
rect 34336 34536 34388 34542
rect 34336 34478 34388 34484
rect 34060 34468 34112 34474
rect 34060 34410 34112 34416
rect 33784 33924 33836 33930
rect 33784 33866 33836 33872
rect 33968 33856 34020 33862
rect 33968 33798 34020 33804
rect 33980 33590 34008 33798
rect 33968 33584 34020 33590
rect 33968 33526 34020 33532
rect 33600 33516 33652 33522
rect 33600 33458 33652 33464
rect 33968 29708 34020 29714
rect 33968 29650 34020 29656
rect 33784 27532 33836 27538
rect 33784 27474 33836 27480
rect 33508 27464 33560 27470
rect 33508 27406 33560 27412
rect 33600 27328 33652 27334
rect 33600 27270 33652 27276
rect 33508 22976 33560 22982
rect 33508 22918 33560 22924
rect 33336 22066 33456 22094
rect 33336 16998 33364 22066
rect 33520 20942 33548 22918
rect 33508 20936 33560 20942
rect 33508 20878 33560 20884
rect 33416 18896 33468 18902
rect 33416 18838 33468 18844
rect 33324 16992 33376 16998
rect 33324 16934 33376 16940
rect 33428 16658 33456 18838
rect 33416 16652 33468 16658
rect 33416 16594 33468 16600
rect 33232 14408 33284 14414
rect 33232 14350 33284 14356
rect 33244 13161 33272 14350
rect 33324 13932 33376 13938
rect 33324 13874 33376 13880
rect 33336 13433 33364 13874
rect 33322 13424 33378 13433
rect 33322 13359 33378 13368
rect 33428 13326 33456 16594
rect 33508 16108 33560 16114
rect 33508 16050 33560 16056
rect 33520 15434 33548 16050
rect 33508 15428 33560 15434
rect 33508 15370 33560 15376
rect 33416 13320 33468 13326
rect 33416 13262 33468 13268
rect 33230 13152 33286 13161
rect 33230 13087 33286 13096
rect 32956 12232 33008 12238
rect 32956 12174 33008 12180
rect 32496 11756 32548 11762
rect 32496 11698 32548 11704
rect 32680 11756 32732 11762
rect 32680 11698 32732 11704
rect 32772 11756 32824 11762
rect 32772 11698 32824 11704
rect 32404 11144 32456 11150
rect 32404 11086 32456 11092
rect 32416 10470 32444 11086
rect 32404 10464 32456 10470
rect 32404 10406 32456 10412
rect 32416 9722 32444 10406
rect 32404 9716 32456 9722
rect 32404 9658 32456 9664
rect 32508 9586 32536 11698
rect 32692 11642 32720 11698
rect 32692 11614 32812 11642
rect 32784 11150 32812 11614
rect 33232 11212 33284 11218
rect 33232 11154 33284 11160
rect 32772 11144 32824 11150
rect 32772 11086 32824 11092
rect 32680 10600 32732 10606
rect 32680 10542 32732 10548
rect 32692 10266 32720 10542
rect 32680 10260 32732 10266
rect 32680 10202 32732 10208
rect 32496 9580 32548 9586
rect 32548 9540 32628 9568
rect 32496 9522 32548 9528
rect 32404 9444 32456 9450
rect 32404 9386 32456 9392
rect 32416 8537 32444 9386
rect 32402 8528 32458 8537
rect 32402 8463 32458 8472
rect 32404 8084 32456 8090
rect 32404 8026 32456 8032
rect 32416 7410 32444 8026
rect 32404 7404 32456 7410
rect 32404 7346 32456 7352
rect 32496 6792 32548 6798
rect 32496 6734 32548 6740
rect 32508 5778 32536 6734
rect 32600 6322 32628 9540
rect 32784 7410 32812 11086
rect 32956 11076 33008 11082
rect 32956 11018 33008 11024
rect 32968 10985 32996 11018
rect 32954 10976 33010 10985
rect 32954 10911 33010 10920
rect 33138 10976 33194 10985
rect 33138 10911 33194 10920
rect 32864 9988 32916 9994
rect 32864 9930 32916 9936
rect 32876 9654 32904 9930
rect 32864 9648 32916 9654
rect 32864 9590 32916 9596
rect 32772 7404 32824 7410
rect 32772 7346 32824 7352
rect 32784 6934 32812 7346
rect 32772 6928 32824 6934
rect 32772 6870 32824 6876
rect 32784 6798 32812 6870
rect 32772 6792 32824 6798
rect 32772 6734 32824 6740
rect 32772 6656 32824 6662
rect 32772 6598 32824 6604
rect 32784 6322 32812 6598
rect 32588 6316 32640 6322
rect 32588 6258 32640 6264
rect 32772 6316 32824 6322
rect 32772 6258 32824 6264
rect 32600 5846 32628 6258
rect 32588 5840 32640 5846
rect 32588 5782 32640 5788
rect 32496 5772 32548 5778
rect 32496 5714 32548 5720
rect 32680 5704 32732 5710
rect 32680 5646 32732 5652
rect 32588 5568 32640 5574
rect 32588 5510 32640 5516
rect 32324 5256 32444 5284
rect 32220 5228 32272 5234
rect 32220 5170 32272 5176
rect 32312 5160 32364 5166
rect 32312 5102 32364 5108
rect 32140 4678 32260 4706
rect 32128 4616 32180 4622
rect 32128 4558 32180 4564
rect 32140 4282 32168 4558
rect 32232 4554 32260 4678
rect 32220 4548 32272 4554
rect 32220 4490 32272 4496
rect 32128 4276 32180 4282
rect 32128 4218 32180 4224
rect 32324 4146 32352 5102
rect 32416 4622 32444 5256
rect 32600 5234 32628 5510
rect 32692 5234 32720 5646
rect 32588 5228 32640 5234
rect 32588 5170 32640 5176
rect 32680 5228 32732 5234
rect 32680 5170 32732 5176
rect 32784 4758 32812 6258
rect 32968 6202 32996 10911
rect 33152 9466 33180 10911
rect 33244 10130 33272 11154
rect 33416 11008 33468 11014
rect 33416 10950 33468 10956
rect 33428 10742 33456 10950
rect 33416 10736 33468 10742
rect 33416 10678 33468 10684
rect 33232 10124 33284 10130
rect 33232 10066 33284 10072
rect 33244 9586 33272 10066
rect 33322 9616 33378 9625
rect 33232 9580 33284 9586
rect 33322 9551 33378 9560
rect 33232 9522 33284 9528
rect 33152 9438 33272 9466
rect 33046 9072 33102 9081
rect 33046 9007 33102 9016
rect 33060 8634 33088 9007
rect 33140 8832 33192 8838
rect 33140 8774 33192 8780
rect 33048 8628 33100 8634
rect 33048 8570 33100 8576
rect 33152 8498 33180 8774
rect 33140 8492 33192 8498
rect 33140 8434 33192 8440
rect 33140 8356 33192 8362
rect 33140 8298 33192 8304
rect 33152 6730 33180 8298
rect 33140 6724 33192 6730
rect 33140 6666 33192 6672
rect 33244 6361 33272 9438
rect 33336 8498 33364 9551
rect 33324 8492 33376 8498
rect 33324 8434 33376 8440
rect 33416 8492 33468 8498
rect 33416 8434 33468 8440
rect 33230 6352 33286 6361
rect 33230 6287 33286 6296
rect 33140 6248 33192 6254
rect 32968 6174 33088 6202
rect 33140 6190 33192 6196
rect 32956 6112 33008 6118
rect 32956 6054 33008 6060
rect 32968 5710 32996 6054
rect 33060 5778 33088 6174
rect 33048 5772 33100 5778
rect 33048 5714 33100 5720
rect 33152 5710 33180 6190
rect 32956 5704 33008 5710
rect 32956 5646 33008 5652
rect 33140 5704 33192 5710
rect 33140 5646 33192 5652
rect 32772 4752 32824 4758
rect 32772 4694 32824 4700
rect 32404 4616 32456 4622
rect 32404 4558 32456 4564
rect 32956 4616 33008 4622
rect 32956 4558 33008 4564
rect 32588 4480 32640 4486
rect 32588 4422 32640 4428
rect 32312 4140 32364 4146
rect 32312 4082 32364 4088
rect 32600 4078 32628 4422
rect 32588 4072 32640 4078
rect 32588 4014 32640 4020
rect 32220 4004 32272 4010
rect 32220 3946 32272 3952
rect 32232 3738 32260 3946
rect 32220 3732 32272 3738
rect 32220 3674 32272 3680
rect 32128 3664 32180 3670
rect 32128 3606 32180 3612
rect 32036 3528 32088 3534
rect 32036 3470 32088 3476
rect 32140 3398 32168 3606
rect 32404 3596 32456 3602
rect 32404 3538 32456 3544
rect 32128 3392 32180 3398
rect 32128 3334 32180 3340
rect 32128 2916 32180 2922
rect 32128 2858 32180 2864
rect 31944 2440 31996 2446
rect 31944 2382 31996 2388
rect 31760 2372 31812 2378
rect 31760 2314 31812 2320
rect 31852 1012 31904 1018
rect 31852 954 31904 960
rect 31864 800 31892 954
rect 32140 800 32168 2858
rect 32416 800 32444 3538
rect 32968 3534 32996 4558
rect 33048 4548 33100 4554
rect 33048 4490 33100 4496
rect 32956 3528 33008 3534
rect 32862 3496 32918 3505
rect 32956 3470 33008 3476
rect 32862 3431 32864 3440
rect 32916 3431 32918 3440
rect 32864 3402 32916 3408
rect 32680 3120 32732 3126
rect 32680 3062 32732 3068
rect 32588 2372 32640 2378
rect 32588 2314 32640 2320
rect 32600 950 32628 2314
rect 32588 944 32640 950
rect 32588 886 32640 892
rect 32692 800 32720 3062
rect 33060 3058 33088 4490
rect 33152 4486 33180 5646
rect 33428 5574 33456 8434
rect 33416 5568 33468 5574
rect 33416 5510 33468 5516
rect 33520 4622 33548 15370
rect 33612 15026 33640 27270
rect 33796 26353 33824 27474
rect 33980 27470 34008 29650
rect 34152 27668 34204 27674
rect 34152 27610 34204 27616
rect 33968 27464 34020 27470
rect 33968 27406 34020 27412
rect 34164 26926 34192 27610
rect 34152 26920 34204 26926
rect 34152 26862 34204 26868
rect 33782 26344 33838 26353
rect 33782 26279 33838 26288
rect 34152 23520 34204 23526
rect 34152 23462 34204 23468
rect 33784 23112 33836 23118
rect 33784 23054 33836 23060
rect 33692 22976 33744 22982
rect 33692 22918 33744 22924
rect 33704 22098 33732 22918
rect 33796 22778 33824 23054
rect 33784 22772 33836 22778
rect 33784 22714 33836 22720
rect 33692 22092 33744 22098
rect 33692 22034 33744 22040
rect 33692 21548 33744 21554
rect 33692 21490 33744 21496
rect 33704 21146 33732 21490
rect 34164 21486 34192 23462
rect 34348 22094 34376 34478
rect 34716 34202 34744 34546
rect 34704 34196 34756 34202
rect 34704 34138 34756 34144
rect 34808 33998 34836 35634
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34796 33992 34848 33998
rect 34796 33934 34848 33940
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 36464 31822 36492 45222
rect 37004 43716 37056 43722
rect 37004 43658 37056 43664
rect 37016 31822 37044 43658
rect 37568 34678 37596 51206
rect 37936 46510 37964 57190
rect 37924 46504 37976 46510
rect 37924 46446 37976 46452
rect 38292 45892 38344 45898
rect 38292 45834 38344 45840
rect 37924 43648 37976 43654
rect 37924 43590 37976 43596
rect 37740 42152 37792 42158
rect 37740 42094 37792 42100
rect 37556 34672 37608 34678
rect 37556 34614 37608 34620
rect 37096 33448 37148 33454
rect 37096 33390 37148 33396
rect 37108 32026 37136 33390
rect 37096 32020 37148 32026
rect 37096 31962 37148 31968
rect 36452 31816 36504 31822
rect 36452 31758 36504 31764
rect 36636 31816 36688 31822
rect 36820 31816 36872 31822
rect 36636 31758 36688 31764
rect 36818 31784 36820 31793
rect 37004 31816 37056 31822
rect 36872 31784 36874 31793
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 36544 30592 36596 30598
rect 36544 30534 36596 30540
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 36556 29073 36584 30534
rect 36648 29782 36676 31758
rect 37004 31758 37056 31764
rect 36818 31719 36874 31728
rect 36820 30252 36872 30258
rect 36820 30194 36872 30200
rect 36636 29776 36688 29782
rect 36636 29718 36688 29724
rect 36542 29064 36598 29073
rect 36542 28999 36598 29008
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 35348 27396 35400 27402
rect 35348 27338 35400 27344
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 35360 26450 35388 27338
rect 35348 26444 35400 26450
rect 35348 26386 35400 26392
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 36544 24608 36596 24614
rect 36544 24550 36596 24556
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 36556 24410 36584 24550
rect 36544 24404 36596 24410
rect 36544 24346 36596 24352
rect 36636 24132 36688 24138
rect 36636 24074 36688 24080
rect 36648 23866 36676 24074
rect 36636 23860 36688 23866
rect 36636 23802 36688 23808
rect 34428 23724 34480 23730
rect 34428 23666 34480 23672
rect 34256 22066 34376 22094
rect 34152 21480 34204 21486
rect 34152 21422 34204 21428
rect 33692 21140 33744 21146
rect 33692 21082 33744 21088
rect 34060 20256 34112 20262
rect 34060 20198 34112 20204
rect 33876 18828 33928 18834
rect 33876 18770 33928 18776
rect 33692 16584 33744 16590
rect 33692 16526 33744 16532
rect 33704 15706 33732 16526
rect 33888 16454 33916 18770
rect 33876 16448 33928 16454
rect 33876 16390 33928 16396
rect 33692 15700 33744 15706
rect 33692 15642 33744 15648
rect 33600 15020 33652 15026
rect 33600 14962 33652 14968
rect 33692 15020 33744 15026
rect 33692 14962 33744 14968
rect 33508 4616 33560 4622
rect 33508 4558 33560 4564
rect 33140 4480 33192 4486
rect 33140 4422 33192 4428
rect 33232 3460 33284 3466
rect 33232 3402 33284 3408
rect 33048 3052 33100 3058
rect 33048 2994 33100 3000
rect 33140 2372 33192 2378
rect 33140 2314 33192 2320
rect 33152 1018 33180 2314
rect 33140 1012 33192 1018
rect 33140 954 33192 960
rect 32956 944 33008 950
rect 32956 886 33008 892
rect 32968 800 32996 886
rect 33244 800 33272 3402
rect 33612 3194 33640 14962
rect 33704 14618 33732 14962
rect 33968 14884 34020 14890
rect 33968 14826 34020 14832
rect 33692 14612 33744 14618
rect 33692 14554 33744 14560
rect 33784 14612 33836 14618
rect 33784 14554 33836 14560
rect 33796 14414 33824 14554
rect 33784 14408 33836 14414
rect 33784 14350 33836 14356
rect 33796 13938 33824 14350
rect 33784 13932 33836 13938
rect 33784 13874 33836 13880
rect 33784 12912 33836 12918
rect 33784 12854 33836 12860
rect 33692 11144 33744 11150
rect 33692 11086 33744 11092
rect 33704 10985 33732 11086
rect 33690 10976 33746 10985
rect 33690 10911 33746 10920
rect 33692 10600 33744 10606
rect 33692 10542 33744 10548
rect 33704 9586 33732 10542
rect 33692 9580 33744 9586
rect 33692 9522 33744 9528
rect 33796 8838 33824 12854
rect 33874 11112 33930 11121
rect 33874 11047 33930 11056
rect 33784 8832 33836 8838
rect 33784 8774 33836 8780
rect 33692 8560 33744 8566
rect 33690 8528 33692 8537
rect 33744 8528 33746 8537
rect 33690 8463 33746 8472
rect 33796 7478 33824 8774
rect 33888 8498 33916 11047
rect 33876 8492 33928 8498
rect 33876 8434 33928 8440
rect 33784 7472 33836 7478
rect 33784 7414 33836 7420
rect 33692 5092 33744 5098
rect 33692 5034 33744 5040
rect 33704 4758 33732 5034
rect 33692 4752 33744 4758
rect 33692 4694 33744 4700
rect 33692 4616 33744 4622
rect 33692 4558 33744 4564
rect 33600 3188 33652 3194
rect 33600 3130 33652 3136
rect 33508 2916 33560 2922
rect 33508 2858 33560 2864
rect 33520 800 33548 2858
rect 33704 2446 33732 4558
rect 33980 3534 34008 14826
rect 34072 14278 34100 20198
rect 34256 16454 34284 22066
rect 34440 20754 34468 23666
rect 35900 23656 35952 23662
rect 35900 23598 35952 23604
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 35912 23118 35940 23598
rect 36728 23588 36780 23594
rect 36728 23530 36780 23536
rect 36360 23520 36412 23526
rect 36360 23462 36412 23468
rect 34888 23112 34940 23118
rect 34888 23054 34940 23060
rect 35900 23112 35952 23118
rect 35900 23054 35952 23060
rect 34900 22778 34928 23054
rect 35256 23044 35308 23050
rect 35256 22986 35308 22992
rect 36176 23044 36228 23050
rect 36176 22986 36228 22992
rect 35164 22976 35216 22982
rect 35164 22918 35216 22924
rect 34888 22772 34940 22778
rect 34888 22714 34940 22720
rect 35176 22420 35204 22918
rect 35268 22642 35296 22986
rect 35440 22704 35492 22710
rect 35492 22652 36124 22658
rect 35440 22646 36124 22652
rect 35452 22642 36124 22646
rect 35256 22636 35308 22642
rect 35452 22636 36136 22642
rect 35452 22630 36084 22636
rect 35256 22578 35308 22584
rect 36084 22578 36136 22584
rect 35348 22568 35400 22574
rect 35348 22510 35400 22516
rect 35440 22568 35492 22574
rect 35440 22510 35492 22516
rect 34808 22392 35204 22420
rect 34808 22030 34836 22392
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34796 22024 34848 22030
rect 34796 21966 34848 21972
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34348 20726 34468 20754
rect 34348 19786 34376 20726
rect 34426 20632 34482 20641
rect 34426 20567 34428 20576
rect 34480 20567 34482 20576
rect 34428 20538 34480 20544
rect 35254 20496 35310 20505
rect 34796 20460 34848 20466
rect 35254 20431 35256 20440
rect 34796 20402 34848 20408
rect 35308 20431 35310 20440
rect 35256 20402 35308 20408
rect 34704 20256 34756 20262
rect 34704 20198 34756 20204
rect 34716 19961 34744 20198
rect 34702 19952 34758 19961
rect 34702 19887 34758 19896
rect 34336 19780 34388 19786
rect 34336 19722 34388 19728
rect 34348 19514 34376 19722
rect 34426 19680 34482 19689
rect 34426 19615 34482 19624
rect 34336 19508 34388 19514
rect 34336 19450 34388 19456
rect 34440 18970 34468 19615
rect 34808 19514 34836 20402
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 35360 19530 35388 22510
rect 35452 22234 35480 22510
rect 35900 22432 35952 22438
rect 35900 22374 35952 22380
rect 35440 22228 35492 22234
rect 35440 22170 35492 22176
rect 35808 22160 35860 22166
rect 35808 22102 35860 22108
rect 35532 20460 35584 20466
rect 35532 20402 35584 20408
rect 35440 20256 35492 20262
rect 35440 20198 35492 20204
rect 35452 20058 35480 20198
rect 35440 20052 35492 20058
rect 35440 19994 35492 20000
rect 35544 19836 35572 20402
rect 35452 19808 35572 19836
rect 35452 19718 35480 19808
rect 35440 19712 35492 19718
rect 35440 19654 35492 19660
rect 35532 19712 35584 19718
rect 35532 19654 35584 19660
rect 34796 19508 34848 19514
rect 35360 19502 35480 19530
rect 34796 19450 34848 19456
rect 34612 19372 34664 19378
rect 34612 19314 34664 19320
rect 35348 19372 35400 19378
rect 35348 19314 35400 19320
rect 34428 18964 34480 18970
rect 34428 18906 34480 18912
rect 34624 18426 34652 19314
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 35360 18970 35388 19314
rect 35348 18964 35400 18970
rect 35348 18906 35400 18912
rect 34796 18896 34848 18902
rect 34796 18838 34848 18844
rect 34704 18624 34756 18630
rect 34704 18566 34756 18572
rect 34612 18420 34664 18426
rect 34612 18362 34664 18368
rect 34716 18290 34744 18566
rect 34612 18284 34664 18290
rect 34612 18226 34664 18232
rect 34704 18284 34756 18290
rect 34704 18226 34756 18232
rect 34520 16516 34572 16522
rect 34520 16458 34572 16464
rect 34244 16448 34296 16454
rect 34244 16390 34296 16396
rect 34256 15881 34284 16390
rect 34242 15872 34298 15881
rect 34242 15807 34298 15816
rect 34428 15020 34480 15026
rect 34428 14962 34480 14968
rect 34440 14550 34468 14962
rect 34428 14544 34480 14550
rect 34428 14486 34480 14492
rect 34532 14414 34560 16458
rect 34624 16250 34652 18226
rect 34808 17678 34836 18838
rect 34888 18760 34940 18766
rect 34888 18702 34940 18708
rect 34900 18408 34928 18702
rect 34980 18420 35032 18426
rect 34900 18380 34980 18408
rect 34980 18362 35032 18368
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34796 17672 34848 17678
rect 34796 17614 34848 17620
rect 34796 17196 34848 17202
rect 34796 17138 34848 17144
rect 34808 16590 34836 17138
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 34796 16584 34848 16590
rect 34796 16526 34848 16532
rect 34612 16244 34664 16250
rect 34612 16186 34664 16192
rect 34704 16108 34756 16114
rect 34704 16050 34756 16056
rect 34716 15910 34744 16050
rect 34704 15904 34756 15910
rect 34704 15846 34756 15852
rect 34716 15570 34744 15846
rect 34704 15564 34756 15570
rect 34704 15506 34756 15512
rect 34808 15502 34836 16526
rect 35164 16516 35216 16522
rect 35164 16458 35216 16464
rect 35176 15978 35204 16458
rect 35164 15972 35216 15978
rect 35164 15914 35216 15920
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34796 15496 34848 15502
rect 34796 15438 34848 15444
rect 34704 14816 34756 14822
rect 34704 14758 34756 14764
rect 34520 14408 34572 14414
rect 34520 14350 34572 14356
rect 34060 14272 34112 14278
rect 34060 14214 34112 14220
rect 34072 14056 34100 14214
rect 34072 14028 34284 14056
rect 34060 13932 34112 13938
rect 34060 13874 34112 13880
rect 34072 13530 34100 13874
rect 34152 13728 34204 13734
rect 34152 13670 34204 13676
rect 34060 13524 34112 13530
rect 34060 13466 34112 13472
rect 34058 13424 34114 13433
rect 34058 13359 34114 13368
rect 34072 13326 34100 13359
rect 34164 13326 34192 13670
rect 34256 13326 34284 14028
rect 34428 14000 34480 14006
rect 34428 13942 34480 13948
rect 34440 13841 34468 13942
rect 34426 13832 34482 13841
rect 34426 13767 34482 13776
rect 34440 13394 34468 13767
rect 34428 13388 34480 13394
rect 34428 13330 34480 13336
rect 34060 13320 34112 13326
rect 34060 13262 34112 13268
rect 34152 13320 34204 13326
rect 34152 13262 34204 13268
rect 34244 13320 34296 13326
rect 34244 13262 34296 13268
rect 34256 12434 34284 13262
rect 34612 12776 34664 12782
rect 34612 12718 34664 12724
rect 34256 12406 34376 12434
rect 34242 11656 34298 11665
rect 34242 11591 34298 11600
rect 34152 11076 34204 11082
rect 34152 11018 34204 11024
rect 34164 9994 34192 11018
rect 34152 9988 34204 9994
rect 34152 9930 34204 9936
rect 34152 7812 34204 7818
rect 34152 7754 34204 7760
rect 34164 6730 34192 7754
rect 34152 6724 34204 6730
rect 34152 6666 34204 6672
rect 34060 6656 34112 6662
rect 34060 6598 34112 6604
rect 34072 6186 34100 6598
rect 34060 6180 34112 6186
rect 34060 6122 34112 6128
rect 34072 4622 34100 6122
rect 34164 5710 34192 6666
rect 34152 5704 34204 5710
rect 34152 5646 34204 5652
rect 34060 4616 34112 4622
rect 34060 4558 34112 4564
rect 34152 4548 34204 4554
rect 34152 4490 34204 4496
rect 34060 3596 34112 3602
rect 34060 3538 34112 3544
rect 33968 3528 34020 3534
rect 33968 3470 34020 3476
rect 33692 2440 33744 2446
rect 33692 2382 33744 2388
rect 33784 1012 33836 1018
rect 33784 954 33836 960
rect 33796 800 33824 954
rect 34072 800 34100 3538
rect 34164 3058 34192 4490
rect 34256 3058 34284 11591
rect 34348 9994 34376 12406
rect 34520 11688 34572 11694
rect 34520 11630 34572 11636
rect 34336 9988 34388 9994
rect 34336 9930 34388 9936
rect 34532 9674 34560 11630
rect 34440 9646 34560 9674
rect 34440 9042 34468 9646
rect 34428 9036 34480 9042
rect 34428 8978 34480 8984
rect 34440 6186 34468 8978
rect 34624 8498 34652 12718
rect 34716 9897 34744 14758
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 35348 14408 35400 14414
rect 35348 14350 35400 14356
rect 35360 14074 35388 14350
rect 35348 14068 35400 14074
rect 35348 14010 35400 14016
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 34796 11756 34848 11762
rect 34796 11698 34848 11704
rect 35348 11756 35400 11762
rect 35348 11698 35400 11704
rect 34808 10810 34836 11698
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 35360 11234 35388 11698
rect 35452 11642 35480 19502
rect 35544 18290 35572 19654
rect 35716 18760 35768 18766
rect 35716 18702 35768 18708
rect 35532 18284 35584 18290
rect 35532 18226 35584 18232
rect 35544 17105 35572 18226
rect 35624 17876 35676 17882
rect 35624 17818 35676 17824
rect 35530 17096 35586 17105
rect 35530 17031 35586 17040
rect 35544 16114 35572 17031
rect 35532 16108 35584 16114
rect 35532 16050 35584 16056
rect 35636 13818 35664 17818
rect 35728 16794 35756 18702
rect 35820 17649 35848 22102
rect 35912 22030 35940 22374
rect 36188 22094 36216 22986
rect 36096 22066 36216 22094
rect 35900 22024 35952 22030
rect 35900 21966 35952 21972
rect 36096 21146 36124 22066
rect 36268 22024 36320 22030
rect 36268 21966 36320 21972
rect 36084 21140 36136 21146
rect 36084 21082 36136 21088
rect 35992 20392 36044 20398
rect 35992 20334 36044 20340
rect 35900 19712 35952 19718
rect 35900 19654 35952 19660
rect 35912 19446 35940 19654
rect 35900 19440 35952 19446
rect 35900 19382 35952 19388
rect 36004 19378 36032 20334
rect 36280 20330 36308 21966
rect 36372 21622 36400 23462
rect 36452 23316 36504 23322
rect 36452 23258 36504 23264
rect 36464 23186 36492 23258
rect 36452 23180 36504 23186
rect 36452 23122 36504 23128
rect 36636 21888 36688 21894
rect 36636 21830 36688 21836
rect 36360 21616 36412 21622
rect 36360 21558 36412 21564
rect 36648 20942 36676 21830
rect 36740 21690 36768 23530
rect 36832 23118 36860 30194
rect 37016 28762 37044 31758
rect 37004 28756 37056 28762
rect 37004 28698 37056 28704
rect 37016 25906 37044 28698
rect 37004 25900 37056 25906
rect 37004 25842 37056 25848
rect 37556 25832 37608 25838
rect 37556 25774 37608 25780
rect 37280 25288 37332 25294
rect 37280 25230 37332 25236
rect 37292 24954 37320 25230
rect 37568 25226 37596 25774
rect 37648 25424 37700 25430
rect 37648 25366 37700 25372
rect 37660 25294 37688 25366
rect 37648 25288 37700 25294
rect 37648 25230 37700 25236
rect 37556 25220 37608 25226
rect 37556 25162 37608 25168
rect 37280 24948 37332 24954
rect 37280 24890 37332 24896
rect 37372 24744 37424 24750
rect 37372 24686 37424 24692
rect 37096 24404 37148 24410
rect 37096 24346 37148 24352
rect 36912 23724 36964 23730
rect 36912 23666 36964 23672
rect 36820 23112 36872 23118
rect 36820 23054 36872 23060
rect 36728 21684 36780 21690
rect 36728 21626 36780 21632
rect 36728 21344 36780 21350
rect 36728 21286 36780 21292
rect 36740 20942 36768 21286
rect 36636 20936 36688 20942
rect 36636 20878 36688 20884
rect 36728 20936 36780 20942
rect 36728 20878 36780 20884
rect 36728 20460 36780 20466
rect 36728 20402 36780 20408
rect 36268 20324 36320 20330
rect 36268 20266 36320 20272
rect 36636 20324 36688 20330
rect 36636 20266 36688 20272
rect 36648 19854 36676 20266
rect 36176 19848 36228 19854
rect 36082 19816 36138 19825
rect 36176 19790 36228 19796
rect 36636 19848 36688 19854
rect 36636 19790 36688 19796
rect 36082 19751 36138 19760
rect 36096 19514 36124 19751
rect 36084 19508 36136 19514
rect 36084 19450 36136 19456
rect 35992 19372 36044 19378
rect 35992 19314 36044 19320
rect 36004 18902 36032 19314
rect 35992 18896 36044 18902
rect 35992 18838 36044 18844
rect 36188 18766 36216 19790
rect 36452 19712 36504 19718
rect 36452 19654 36504 19660
rect 36544 19712 36596 19718
rect 36544 19654 36596 19660
rect 36360 19236 36412 19242
rect 36360 19178 36412 19184
rect 36176 18760 36228 18766
rect 36176 18702 36228 18708
rect 36188 18358 36216 18702
rect 36176 18352 36228 18358
rect 36176 18294 36228 18300
rect 36188 17898 36216 18294
rect 36096 17870 36216 17898
rect 36096 17746 36124 17870
rect 36176 17808 36228 17814
rect 36176 17750 36228 17756
rect 36084 17740 36136 17746
rect 36084 17682 36136 17688
rect 35806 17640 35862 17649
rect 35806 17575 35862 17584
rect 35716 16788 35768 16794
rect 35716 16730 35768 16736
rect 35820 14634 35848 17575
rect 36082 17504 36138 17513
rect 36082 17439 36138 17448
rect 36096 17338 36124 17439
rect 36084 17332 36136 17338
rect 36084 17274 36136 17280
rect 36188 17202 36216 17750
rect 36268 17740 36320 17746
rect 36268 17682 36320 17688
rect 36176 17196 36228 17202
rect 36176 17138 36228 17144
rect 35900 17128 35952 17134
rect 35898 17096 35900 17105
rect 35952 17096 35954 17105
rect 35898 17031 35954 17040
rect 35900 16992 35952 16998
rect 35900 16934 35952 16940
rect 35912 16590 35940 16934
rect 36084 16720 36136 16726
rect 36084 16662 36136 16668
rect 35900 16584 35952 16590
rect 35900 16526 35952 16532
rect 36096 15910 36124 16662
rect 36280 16590 36308 17682
rect 36268 16584 36320 16590
rect 36268 16526 36320 16532
rect 36084 15904 36136 15910
rect 36084 15846 36136 15852
rect 36372 15094 36400 19178
rect 36464 18766 36492 19654
rect 36556 19446 36584 19654
rect 36544 19440 36596 19446
rect 36544 19382 36596 19388
rect 36544 18964 36596 18970
rect 36544 18906 36596 18912
rect 36452 18760 36504 18766
rect 36452 18702 36504 18708
rect 36556 17678 36584 18906
rect 36740 18630 36768 20402
rect 36832 20074 36860 23054
rect 36924 23050 36952 23666
rect 36912 23044 36964 23050
rect 36912 22986 36964 22992
rect 36924 22506 36952 22986
rect 36912 22500 36964 22506
rect 36912 22442 36964 22448
rect 36912 22024 36964 22030
rect 36912 21966 36964 21972
rect 36924 21146 36952 21966
rect 37108 21962 37136 24346
rect 37384 24206 37412 24686
rect 37280 24200 37332 24206
rect 37280 24142 37332 24148
rect 37372 24200 37424 24206
rect 37372 24142 37424 24148
rect 37096 21956 37148 21962
rect 37096 21898 37148 21904
rect 37004 21684 37056 21690
rect 37004 21626 37056 21632
rect 37016 21457 37044 21626
rect 37002 21448 37058 21457
rect 37002 21383 37058 21392
rect 36912 21140 36964 21146
rect 36912 21082 36964 21088
rect 37004 20256 37056 20262
rect 37004 20198 37056 20204
rect 36832 20046 36952 20074
rect 36820 19984 36872 19990
rect 36820 19926 36872 19932
rect 36832 19553 36860 19926
rect 36818 19544 36874 19553
rect 36818 19479 36874 19488
rect 36924 19242 36952 20046
rect 37016 19854 37044 20198
rect 37004 19848 37056 19854
rect 37004 19790 37056 19796
rect 36912 19236 36964 19242
rect 36912 19178 36964 19184
rect 36728 18624 36780 18630
rect 36728 18566 36780 18572
rect 36636 18080 36688 18086
rect 36636 18022 36688 18028
rect 36544 17672 36596 17678
rect 36544 17614 36596 17620
rect 36450 17504 36506 17513
rect 36450 17439 36506 17448
rect 36360 15088 36412 15094
rect 36360 15030 36412 15036
rect 35820 14606 35940 14634
rect 35808 14544 35860 14550
rect 35808 14486 35860 14492
rect 35820 13938 35848 14486
rect 35808 13932 35860 13938
rect 35808 13874 35860 13880
rect 35636 13790 35848 13818
rect 35624 12980 35676 12986
rect 35624 12922 35676 12928
rect 35452 11614 35572 11642
rect 35440 11552 35492 11558
rect 35440 11494 35492 11500
rect 35268 11206 35388 11234
rect 35268 11150 35296 11206
rect 35452 11150 35480 11494
rect 35256 11144 35308 11150
rect 35256 11086 35308 11092
rect 35440 11144 35492 11150
rect 35440 11086 35492 11092
rect 34796 10804 34848 10810
rect 34796 10746 34848 10752
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34702 9888 34758 9897
rect 34702 9823 34758 9832
rect 35440 9376 35492 9382
rect 35440 9318 35492 9324
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 35348 8968 35400 8974
rect 35348 8910 35400 8916
rect 34612 8492 34664 8498
rect 34612 8434 34664 8440
rect 35360 8430 35388 8910
rect 35348 8424 35400 8430
rect 35348 8366 35400 8372
rect 35452 8378 35480 9318
rect 35544 8566 35572 11614
rect 35636 10674 35664 12922
rect 35716 12436 35768 12442
rect 35716 12378 35768 12384
rect 35728 11150 35756 12378
rect 35716 11144 35768 11150
rect 35716 11086 35768 11092
rect 35728 10810 35756 11086
rect 35716 10804 35768 10810
rect 35716 10746 35768 10752
rect 35624 10668 35676 10674
rect 35624 10610 35676 10616
rect 35820 9674 35848 13790
rect 35912 13433 35940 14606
rect 35898 13424 35954 13433
rect 35898 13359 35954 13368
rect 36268 13320 36320 13326
rect 36082 13288 36138 13297
rect 36268 13262 36320 13268
rect 36082 13223 36138 13232
rect 35624 9648 35676 9654
rect 35624 9590 35676 9596
rect 35716 9648 35768 9654
rect 35820 9646 35940 9674
rect 35716 9590 35768 9596
rect 35532 8560 35584 8566
rect 35532 8502 35584 8508
rect 34520 8356 34572 8362
rect 34520 8298 34572 8304
rect 34532 7886 34560 8298
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 34520 7880 34572 7886
rect 35360 7868 35388 8366
rect 35452 8350 35572 8378
rect 35440 8288 35492 8294
rect 35440 8230 35492 8236
rect 35452 8090 35480 8230
rect 35440 8084 35492 8090
rect 35440 8026 35492 8032
rect 35440 7880 35492 7886
rect 35360 7840 35440 7868
rect 34520 7822 34572 7828
rect 35440 7822 35492 7828
rect 35348 7540 35400 7546
rect 35348 7482 35400 7488
rect 34796 7268 34848 7274
rect 34796 7210 34848 7216
rect 34808 7177 34836 7210
rect 34794 7168 34850 7177
rect 34794 7103 34850 7112
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34704 6724 34756 6730
rect 34704 6666 34756 6672
rect 34612 6656 34664 6662
rect 34612 6598 34664 6604
rect 34624 6458 34652 6598
rect 34716 6458 34744 6666
rect 34612 6452 34664 6458
rect 34612 6394 34664 6400
rect 34704 6452 34756 6458
rect 34704 6394 34756 6400
rect 35360 6322 35388 7482
rect 35348 6316 35400 6322
rect 35348 6258 35400 6264
rect 34612 6248 34664 6254
rect 34612 6190 34664 6196
rect 34428 6180 34480 6186
rect 34428 6122 34480 6128
rect 34624 5710 34652 6190
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34612 5704 34664 5710
rect 34612 5646 34664 5652
rect 34624 5302 34652 5646
rect 34612 5296 34664 5302
rect 34612 5238 34664 5244
rect 35360 5098 35388 6258
rect 35452 6202 35480 7822
rect 35544 6322 35572 8350
rect 35636 7342 35664 9590
rect 35728 9382 35756 9590
rect 35716 9376 35768 9382
rect 35716 9318 35768 9324
rect 35912 9058 35940 9646
rect 35912 9042 36032 9058
rect 35912 9036 36044 9042
rect 35912 9030 35992 9036
rect 35992 8978 36044 8984
rect 35808 8968 35860 8974
rect 35808 8910 35860 8916
rect 35820 8498 35848 8910
rect 35808 8492 35860 8498
rect 35808 8434 35860 8440
rect 35820 7886 35848 8434
rect 35900 8084 35952 8090
rect 35900 8026 35952 8032
rect 35808 7880 35860 7886
rect 35808 7822 35860 7828
rect 35820 7546 35848 7822
rect 35912 7818 35940 8026
rect 35990 7984 36046 7993
rect 35990 7919 35992 7928
rect 36044 7919 36046 7928
rect 35992 7890 36044 7896
rect 35900 7812 35952 7818
rect 35900 7754 35952 7760
rect 35808 7540 35860 7546
rect 35808 7482 35860 7488
rect 35624 7336 35676 7342
rect 35624 7278 35676 7284
rect 35636 6798 35664 7278
rect 35624 6792 35676 6798
rect 35624 6734 35676 6740
rect 35716 6792 35768 6798
rect 35716 6734 35768 6740
rect 35532 6316 35584 6322
rect 35532 6258 35584 6264
rect 35452 6174 35572 6202
rect 35544 5710 35572 6174
rect 35532 5704 35584 5710
rect 35532 5646 35584 5652
rect 35440 5636 35492 5642
rect 35440 5578 35492 5584
rect 35348 5092 35400 5098
rect 35348 5034 35400 5040
rect 34704 5024 34756 5030
rect 34704 4966 34756 4972
rect 34716 4146 34744 4966
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 35360 4758 35388 5034
rect 35348 4752 35400 4758
rect 35162 4720 35218 4729
rect 35348 4694 35400 4700
rect 35162 4655 35218 4664
rect 35176 4622 35204 4655
rect 35164 4616 35216 4622
rect 35164 4558 35216 4564
rect 35452 4146 35480 5578
rect 35544 5234 35572 5646
rect 35636 5302 35664 6734
rect 35728 6633 35756 6734
rect 35714 6624 35770 6633
rect 35714 6559 35770 6568
rect 35900 6316 35952 6322
rect 35900 6258 35952 6264
rect 35912 6225 35940 6258
rect 35898 6216 35954 6225
rect 35716 6180 35768 6186
rect 35898 6151 35954 6160
rect 35716 6122 35768 6128
rect 35624 5296 35676 5302
rect 35624 5238 35676 5244
rect 35532 5228 35584 5234
rect 35532 5170 35584 5176
rect 35728 4622 35756 6122
rect 35808 6112 35860 6118
rect 35808 6054 35860 6060
rect 35820 5710 35848 6054
rect 36096 5778 36124 13223
rect 36280 12782 36308 13262
rect 36268 12776 36320 12782
rect 36268 12718 36320 12724
rect 36280 12238 36308 12718
rect 36464 12434 36492 17439
rect 36556 17338 36584 17614
rect 36544 17332 36596 17338
rect 36544 17274 36596 17280
rect 36544 17060 36596 17066
rect 36544 17002 36596 17008
rect 36556 16017 36584 17002
rect 36648 16538 36676 18022
rect 36740 16726 36768 18566
rect 36820 18216 36872 18222
rect 36820 18158 36872 18164
rect 36832 17882 36860 18158
rect 36820 17876 36872 17882
rect 36820 17818 36872 17824
rect 36728 16720 36780 16726
rect 36728 16662 36780 16668
rect 36648 16510 36768 16538
rect 36542 16008 36598 16017
rect 36542 15943 36598 15952
rect 36636 12640 36688 12646
rect 36636 12582 36688 12588
rect 36464 12406 36584 12434
rect 36268 12232 36320 12238
rect 36268 12174 36320 12180
rect 36280 11830 36308 12174
rect 36268 11824 36320 11830
rect 36268 11766 36320 11772
rect 36452 9988 36504 9994
rect 36452 9930 36504 9936
rect 36268 9920 36320 9926
rect 36268 9862 36320 9868
rect 36280 9058 36308 9862
rect 36464 9518 36492 9930
rect 36452 9512 36504 9518
rect 36452 9454 36504 9460
rect 36464 9178 36492 9454
rect 36452 9172 36504 9178
rect 36452 9114 36504 9120
rect 36280 9030 36400 9058
rect 36268 8900 36320 8906
rect 36268 8842 36320 8848
rect 36174 8800 36230 8809
rect 36174 8735 36230 8744
rect 36188 8566 36216 8735
rect 36176 8560 36228 8566
rect 36176 8502 36228 8508
rect 36280 7936 36308 8842
rect 36188 7908 36308 7936
rect 36188 6497 36216 7908
rect 36268 7812 36320 7818
rect 36268 7754 36320 7760
rect 36280 7585 36308 7754
rect 36266 7576 36322 7585
rect 36266 7511 36322 7520
rect 36372 7290 36400 9030
rect 36450 8392 36506 8401
rect 36450 8327 36452 8336
rect 36504 8327 36506 8336
rect 36452 8298 36504 8304
rect 36280 7262 36400 7290
rect 36174 6488 36230 6497
rect 36174 6423 36230 6432
rect 36280 6186 36308 7262
rect 36360 6316 36412 6322
rect 36360 6258 36412 6264
rect 36268 6180 36320 6186
rect 36268 6122 36320 6128
rect 36084 5772 36136 5778
rect 36084 5714 36136 5720
rect 35808 5704 35860 5710
rect 35808 5646 35860 5652
rect 36266 5672 36322 5681
rect 35820 5234 35848 5646
rect 36266 5607 36268 5616
rect 36320 5607 36322 5616
rect 36268 5578 36320 5584
rect 36176 5296 36228 5302
rect 36176 5238 36228 5244
rect 35808 5228 35860 5234
rect 35808 5170 35860 5176
rect 35716 4616 35768 4622
rect 35716 4558 35768 4564
rect 34704 4140 34756 4146
rect 34704 4082 34756 4088
rect 35440 4140 35492 4146
rect 35440 4082 35492 4088
rect 34612 4072 34664 4078
rect 34612 4014 34664 4020
rect 35348 4072 35400 4078
rect 35348 4014 35400 4020
rect 34152 3052 34204 3058
rect 34152 2994 34204 3000
rect 34244 3052 34296 3058
rect 34244 2994 34296 3000
rect 34520 2372 34572 2378
rect 34520 2314 34572 2320
rect 34336 1216 34388 1222
rect 34336 1158 34388 1164
rect 34348 800 34376 1158
rect 34532 950 34560 2314
rect 34520 944 34572 950
rect 34520 886 34572 892
rect 34624 800 34652 4014
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 34888 1080 34940 1086
rect 34888 1022 34940 1028
rect 34900 800 34928 1022
rect 35360 898 35388 4014
rect 35820 3738 35848 5170
rect 35900 4616 35952 4622
rect 35900 4558 35952 4564
rect 35992 4616 36044 4622
rect 35992 4558 36044 4564
rect 35912 4321 35940 4558
rect 36004 4457 36032 4558
rect 35990 4448 36046 4457
rect 35990 4383 36046 4392
rect 35898 4312 35954 4321
rect 35898 4247 35954 4256
rect 36188 4214 36216 5238
rect 36268 5228 36320 5234
rect 36268 5170 36320 5176
rect 36176 4208 36228 4214
rect 36176 4150 36228 4156
rect 36084 4072 36136 4078
rect 36084 4014 36136 4020
rect 35808 3732 35860 3738
rect 35808 3674 35860 3680
rect 35992 3392 36044 3398
rect 35992 3334 36044 3340
rect 36004 3058 36032 3334
rect 35992 3052 36044 3058
rect 35992 2994 36044 3000
rect 36096 2774 36124 4014
rect 36188 3602 36216 4150
rect 36176 3596 36228 3602
rect 36176 3538 36228 3544
rect 36280 3233 36308 5170
rect 36372 4690 36400 6258
rect 36360 4684 36412 4690
rect 36360 4626 36412 4632
rect 36360 4480 36412 4486
rect 36360 4422 36412 4428
rect 36372 3534 36400 4422
rect 36556 4214 36584 12406
rect 36648 11762 36676 12582
rect 36636 11756 36688 11762
rect 36636 11698 36688 11704
rect 36634 9480 36690 9489
rect 36634 9415 36690 9424
rect 36648 9178 36676 9415
rect 36636 9172 36688 9178
rect 36636 9114 36688 9120
rect 36636 8016 36688 8022
rect 36636 7958 36688 7964
rect 36648 7818 36676 7958
rect 36636 7812 36688 7818
rect 36636 7754 36688 7760
rect 36740 5234 36768 16510
rect 36832 16114 36860 17818
rect 36912 17808 36964 17814
rect 36912 17750 36964 17756
rect 36924 17270 36952 17750
rect 36912 17264 36964 17270
rect 36912 17206 36964 17212
rect 36912 16584 36964 16590
rect 36912 16526 36964 16532
rect 36924 16250 36952 16526
rect 36912 16244 36964 16250
rect 36912 16186 36964 16192
rect 36820 16108 36872 16114
rect 36820 16050 36872 16056
rect 36912 13184 36964 13190
rect 36912 13126 36964 13132
rect 36924 8022 36952 13126
rect 37108 9654 37136 21898
rect 37188 21548 37240 21554
rect 37188 21490 37240 21496
rect 37200 21146 37228 21490
rect 37188 21140 37240 21146
rect 37188 21082 37240 21088
rect 37188 20460 37240 20466
rect 37188 20402 37240 20408
rect 37200 19854 37228 20402
rect 37188 19848 37240 19854
rect 37188 19790 37240 19796
rect 37188 19508 37240 19514
rect 37188 19450 37240 19456
rect 37200 17746 37228 19450
rect 37188 17740 37240 17746
rect 37188 17682 37240 17688
rect 37188 13388 37240 13394
rect 37188 13330 37240 13336
rect 37200 12850 37228 13330
rect 37188 12844 37240 12850
rect 37188 12786 37240 12792
rect 37096 9648 37148 9654
rect 37096 9590 37148 9596
rect 36912 8016 36964 8022
rect 36912 7958 36964 7964
rect 37292 7290 37320 24142
rect 37372 23792 37424 23798
rect 37372 23734 37424 23740
rect 37384 21554 37412 23734
rect 37464 23520 37516 23526
rect 37464 23462 37516 23468
rect 37476 22642 37504 23462
rect 37464 22636 37516 22642
rect 37464 22578 37516 22584
rect 37568 22094 37596 25162
rect 37752 24818 37780 42094
rect 37832 32224 37884 32230
rect 37832 32166 37884 32172
rect 37844 32026 37872 32166
rect 37832 32020 37884 32026
rect 37832 31962 37884 31968
rect 37936 28558 37964 43590
rect 38304 35894 38332 45834
rect 38304 35866 38424 35894
rect 37924 28552 37976 28558
rect 37924 28494 37976 28500
rect 37832 26444 37884 26450
rect 37832 26386 37884 26392
rect 37844 24818 37872 26386
rect 37740 24812 37792 24818
rect 37740 24754 37792 24760
rect 37832 24812 37884 24818
rect 37832 24754 37884 24760
rect 37648 24200 37700 24206
rect 37844 24188 37872 24754
rect 37700 24160 37872 24188
rect 37922 24168 37978 24177
rect 37648 24142 37700 24148
rect 37922 24103 37978 24112
rect 37936 24070 37964 24103
rect 37924 24064 37976 24070
rect 37924 24006 37976 24012
rect 37740 22772 37792 22778
rect 37740 22714 37792 22720
rect 37752 22234 37780 22714
rect 38200 22704 38252 22710
rect 38200 22646 38252 22652
rect 37740 22228 37792 22234
rect 37740 22170 37792 22176
rect 38108 22228 38160 22234
rect 38108 22170 38160 22176
rect 37568 22066 38056 22094
rect 37648 21888 37700 21894
rect 37648 21830 37700 21836
rect 37372 21548 37424 21554
rect 37372 21490 37424 21496
rect 37556 21344 37608 21350
rect 37556 21286 37608 21292
rect 37464 20936 37516 20942
rect 37464 20878 37516 20884
rect 37476 20602 37504 20878
rect 37464 20596 37516 20602
rect 37464 20538 37516 20544
rect 37464 20460 37516 20466
rect 37464 20402 37516 20408
rect 37372 20052 37424 20058
rect 37372 19994 37424 20000
rect 37384 19922 37412 19994
rect 37372 19916 37424 19922
rect 37372 19858 37424 19864
rect 37372 19712 37424 19718
rect 37372 19654 37424 19660
rect 37384 18290 37412 19654
rect 37476 19514 37504 20402
rect 37568 20058 37596 21286
rect 37556 20052 37608 20058
rect 37556 19994 37608 20000
rect 37464 19508 37516 19514
rect 37464 19450 37516 19456
rect 37568 19378 37596 19994
rect 37556 19372 37608 19378
rect 37556 19314 37608 19320
rect 37660 18358 37688 21830
rect 37740 21412 37792 21418
rect 37740 21354 37792 21360
rect 37752 21078 37780 21354
rect 37740 21072 37792 21078
rect 37740 21014 37792 21020
rect 37832 20868 37884 20874
rect 37832 20810 37884 20816
rect 37844 20330 37872 20810
rect 37832 20324 37884 20330
rect 37832 20266 37884 20272
rect 37740 20052 37792 20058
rect 37740 19994 37792 20000
rect 37648 18352 37700 18358
rect 37648 18294 37700 18300
rect 37372 18284 37424 18290
rect 37372 18226 37424 18232
rect 37464 18148 37516 18154
rect 37464 18090 37516 18096
rect 37372 17672 37424 17678
rect 37372 17614 37424 17620
rect 37384 16522 37412 17614
rect 37372 16516 37424 16522
rect 37372 16458 37424 16464
rect 37476 16250 37504 18090
rect 37556 18080 37608 18086
rect 37556 18022 37608 18028
rect 37568 16658 37596 18022
rect 37648 16992 37700 16998
rect 37648 16934 37700 16940
rect 37556 16652 37608 16658
rect 37556 16594 37608 16600
rect 37464 16244 37516 16250
rect 37464 16186 37516 16192
rect 37660 16182 37688 16934
rect 37752 16794 37780 19994
rect 37844 19514 37872 20266
rect 37832 19508 37884 19514
rect 37832 19450 37884 19456
rect 37924 18284 37976 18290
rect 37924 18226 37976 18232
rect 37832 18080 37884 18086
rect 37832 18022 37884 18028
rect 37844 17134 37872 18022
rect 37832 17128 37884 17134
rect 37832 17070 37884 17076
rect 37740 16788 37792 16794
rect 37740 16730 37792 16736
rect 37740 16516 37792 16522
rect 37740 16458 37792 16464
rect 37752 16250 37780 16458
rect 37740 16244 37792 16250
rect 37740 16186 37792 16192
rect 37648 16176 37700 16182
rect 37648 16118 37700 16124
rect 37832 16108 37884 16114
rect 37832 16050 37884 16056
rect 37740 15904 37792 15910
rect 37740 15846 37792 15852
rect 37648 15020 37700 15026
rect 37648 14962 37700 14968
rect 37464 13728 37516 13734
rect 37464 13670 37516 13676
rect 37476 13326 37504 13670
rect 37464 13320 37516 13326
rect 37464 13262 37516 13268
rect 37556 12776 37608 12782
rect 37556 12718 37608 12724
rect 37372 12368 37424 12374
rect 37372 12310 37424 12316
rect 37384 11014 37412 12310
rect 37464 12164 37516 12170
rect 37464 12106 37516 12112
rect 37476 11898 37504 12106
rect 37464 11892 37516 11898
rect 37464 11834 37516 11840
rect 37568 11558 37596 12718
rect 37660 12238 37688 14962
rect 37752 12434 37780 15846
rect 37844 15434 37872 16050
rect 37936 15978 37964 18226
rect 37924 15972 37976 15978
rect 37924 15914 37976 15920
rect 37832 15428 37884 15434
rect 37832 15370 37884 15376
rect 38028 14906 38056 22066
rect 38120 21962 38148 22170
rect 38108 21956 38160 21962
rect 38108 21898 38160 21904
rect 38120 21865 38148 21898
rect 38106 21856 38162 21865
rect 38106 21791 38162 21800
rect 38212 19378 38240 22646
rect 38396 22094 38424 35866
rect 39316 29510 39344 57190
rect 39396 45008 39448 45014
rect 39396 44950 39448 44956
rect 39304 29504 39356 29510
rect 39304 29446 39356 29452
rect 38476 25832 38528 25838
rect 38476 25774 38528 25780
rect 38844 25832 38896 25838
rect 38844 25774 38896 25780
rect 38488 25226 38516 25774
rect 38856 25294 38884 25774
rect 38844 25288 38896 25294
rect 38844 25230 38896 25236
rect 38476 25220 38528 25226
rect 38476 25162 38528 25168
rect 39304 24744 39356 24750
rect 39304 24686 39356 24692
rect 39120 23316 39172 23322
rect 39120 23258 39172 23264
rect 39132 23225 39160 23258
rect 39118 23216 39174 23225
rect 39118 23151 39174 23160
rect 39212 23112 39264 23118
rect 38948 23080 39212 23100
rect 39264 23080 39266 23089
rect 38948 23072 39210 23080
rect 38844 22976 38896 22982
rect 38844 22918 38896 22924
rect 38856 22710 38884 22918
rect 38844 22704 38896 22710
rect 38844 22646 38896 22652
rect 38844 22432 38896 22438
rect 38844 22374 38896 22380
rect 38750 22264 38806 22273
rect 38750 22199 38806 22208
rect 38764 22166 38792 22199
rect 38752 22160 38804 22166
rect 38752 22102 38804 22108
rect 38304 22066 38424 22094
rect 38304 19394 38332 22066
rect 38752 22024 38804 22030
rect 38672 21972 38752 21978
rect 38672 21966 38804 21972
rect 38672 21950 38792 21966
rect 38568 21888 38620 21894
rect 38672 21865 38700 21950
rect 38568 21830 38620 21836
rect 38658 21856 38714 21865
rect 38384 21140 38436 21146
rect 38384 21082 38436 21088
rect 38396 20942 38424 21082
rect 38580 20942 38608 21830
rect 38658 21791 38714 21800
rect 38856 21622 38884 22374
rect 38948 22166 38976 23072
rect 39210 23015 39266 23024
rect 39316 22250 39344 24686
rect 39408 24138 39436 44950
rect 40328 40526 40356 57190
rect 40960 48204 41012 48210
rect 40960 48146 41012 48152
rect 40972 47734 41000 48146
rect 41604 48068 41656 48074
rect 41604 48010 41656 48016
rect 41616 47734 41644 48010
rect 41708 47734 41736 57190
rect 42340 52488 42392 52494
rect 42340 52430 42392 52436
rect 42524 52488 42576 52494
rect 42524 52430 42576 52436
rect 41788 48136 41840 48142
rect 41788 48078 41840 48084
rect 40960 47728 41012 47734
rect 40960 47670 41012 47676
rect 41604 47728 41656 47734
rect 41604 47670 41656 47676
rect 41696 47728 41748 47734
rect 41696 47670 41748 47676
rect 41800 47666 41828 48078
rect 41788 47660 41840 47666
rect 41788 47602 41840 47608
rect 42156 47456 42208 47462
rect 42156 47398 42208 47404
rect 41696 44464 41748 44470
rect 41696 44406 41748 44412
rect 41420 44396 41472 44402
rect 41420 44338 41472 44344
rect 41328 43784 41380 43790
rect 41328 43726 41380 43732
rect 41340 42945 41368 43726
rect 41326 42936 41382 42945
rect 41326 42871 41382 42880
rect 40316 40520 40368 40526
rect 40316 40462 40368 40468
rect 40592 40520 40644 40526
rect 40592 40462 40644 40468
rect 39948 34060 40000 34066
rect 39948 34002 40000 34008
rect 39960 32434 39988 34002
rect 39948 32428 40000 32434
rect 39948 32370 40000 32376
rect 39488 25356 39540 25362
rect 39488 25298 39540 25304
rect 39396 24132 39448 24138
rect 39396 24074 39448 24080
rect 39040 22222 39344 22250
rect 38936 22160 38988 22166
rect 38936 22102 38988 22108
rect 38844 21616 38896 21622
rect 38844 21558 38896 21564
rect 38948 21434 38976 22102
rect 39040 22030 39068 22222
rect 39120 22160 39172 22166
rect 39120 22102 39172 22108
rect 39028 22024 39080 22030
rect 39028 21966 39080 21972
rect 39132 21894 39160 22102
rect 39120 21888 39172 21894
rect 39120 21830 39172 21836
rect 38764 21406 38976 21434
rect 38384 20936 38436 20942
rect 38384 20878 38436 20884
rect 38568 20936 38620 20942
rect 38568 20878 38620 20884
rect 38660 20868 38712 20874
rect 38660 20810 38712 20816
rect 38568 20392 38620 20398
rect 38568 20334 38620 20340
rect 38476 20052 38528 20058
rect 38476 19994 38528 20000
rect 38488 19854 38516 19994
rect 38476 19848 38528 19854
rect 38476 19790 38528 19796
rect 38476 19440 38528 19446
rect 38200 19372 38252 19378
rect 38304 19366 38424 19394
rect 38476 19382 38528 19388
rect 38200 19314 38252 19320
rect 38106 17640 38162 17649
rect 38106 17575 38162 17584
rect 38120 17542 38148 17575
rect 38108 17536 38160 17542
rect 38108 17478 38160 17484
rect 38212 17082 38240 19314
rect 38120 17054 38240 17082
rect 38120 16658 38148 17054
rect 38108 16652 38160 16658
rect 38108 16594 38160 16600
rect 38120 15094 38148 16594
rect 38198 16008 38254 16017
rect 38198 15943 38254 15952
rect 38212 15910 38240 15943
rect 38200 15904 38252 15910
rect 38200 15846 38252 15852
rect 38396 15858 38424 19366
rect 38488 18970 38516 19382
rect 38476 18964 38528 18970
rect 38476 18906 38528 18912
rect 38580 18136 38608 20334
rect 38672 19854 38700 20810
rect 38764 20398 38792 21406
rect 38844 20936 38896 20942
rect 38844 20878 38896 20884
rect 38856 20602 38884 20878
rect 39028 20868 39080 20874
rect 39028 20810 39080 20816
rect 38934 20768 38990 20777
rect 38934 20703 38990 20712
rect 38844 20596 38896 20602
rect 38844 20538 38896 20544
rect 38948 20466 38976 20703
rect 38844 20460 38896 20466
rect 38844 20402 38896 20408
rect 38936 20460 38988 20466
rect 38936 20402 38988 20408
rect 38752 20392 38804 20398
rect 38752 20334 38804 20340
rect 38660 19848 38712 19854
rect 38660 19790 38712 19796
rect 38672 18630 38700 19790
rect 38764 18766 38792 20334
rect 38856 19718 38884 20402
rect 38844 19712 38896 19718
rect 38844 19654 38896 19660
rect 38752 18760 38804 18766
rect 38752 18702 38804 18708
rect 38660 18624 38712 18630
rect 38660 18566 38712 18572
rect 38844 18624 38896 18630
rect 38844 18566 38896 18572
rect 38488 18108 38608 18136
rect 38488 17678 38516 18108
rect 38568 17808 38620 17814
rect 38568 17750 38620 17756
rect 38476 17672 38528 17678
rect 38476 17614 38528 17620
rect 38488 17066 38516 17614
rect 38580 17202 38608 17750
rect 38568 17196 38620 17202
rect 38568 17138 38620 17144
rect 38752 17196 38804 17202
rect 38752 17138 38804 17144
rect 38476 17060 38528 17066
rect 38476 17002 38528 17008
rect 38660 16992 38712 16998
rect 38660 16934 38712 16940
rect 38568 16516 38620 16522
rect 38568 16458 38620 16464
rect 38580 16046 38608 16458
rect 38672 16182 38700 16934
rect 38764 16794 38792 17138
rect 38752 16788 38804 16794
rect 38752 16730 38804 16736
rect 38764 16522 38792 16730
rect 38752 16516 38804 16522
rect 38752 16458 38804 16464
rect 38660 16176 38712 16182
rect 38660 16118 38712 16124
rect 38568 16040 38620 16046
rect 38568 15982 38620 15988
rect 38660 16040 38712 16046
rect 38660 15982 38712 15988
rect 38396 15830 38608 15858
rect 38476 15496 38528 15502
rect 38476 15438 38528 15444
rect 38200 15360 38252 15366
rect 38200 15302 38252 15308
rect 38384 15360 38436 15366
rect 38384 15302 38436 15308
rect 38108 15088 38160 15094
rect 38108 15030 38160 15036
rect 38212 15026 38240 15302
rect 38200 15020 38252 15026
rect 38200 14962 38252 14968
rect 38028 14878 38332 14906
rect 37924 13864 37976 13870
rect 37924 13806 37976 13812
rect 38108 13864 38160 13870
rect 38108 13806 38160 13812
rect 37936 13530 37964 13806
rect 37924 13524 37976 13530
rect 37924 13466 37976 13472
rect 38120 12782 38148 13806
rect 38108 12776 38160 12782
rect 38028 12736 38108 12764
rect 37752 12406 37872 12434
rect 37648 12232 37700 12238
rect 37648 12174 37700 12180
rect 37738 12200 37794 12209
rect 37660 11762 37688 12174
rect 37738 12135 37794 12144
rect 37752 12102 37780 12135
rect 37740 12096 37792 12102
rect 37740 12038 37792 12044
rect 37752 11830 37780 12038
rect 37740 11824 37792 11830
rect 37740 11766 37792 11772
rect 37648 11756 37700 11762
rect 37648 11698 37700 11704
rect 37556 11552 37608 11558
rect 37556 11494 37608 11500
rect 37740 11552 37792 11558
rect 37740 11494 37792 11500
rect 37372 11008 37424 11014
rect 37372 10950 37424 10956
rect 37372 8356 37424 8362
rect 37372 8298 37424 8304
rect 37384 7886 37412 8298
rect 37568 7886 37596 11494
rect 37648 8968 37700 8974
rect 37648 8910 37700 8916
rect 37660 8430 37688 8910
rect 37648 8424 37700 8430
rect 37648 8366 37700 8372
rect 37372 7880 37424 7886
rect 37372 7822 37424 7828
rect 37464 7880 37516 7886
rect 37464 7822 37516 7828
rect 37556 7880 37608 7886
rect 37556 7822 37608 7828
rect 37384 7410 37412 7822
rect 37476 7546 37504 7822
rect 37464 7540 37516 7546
rect 37464 7482 37516 7488
rect 37372 7404 37424 7410
rect 37372 7346 37424 7352
rect 37292 7262 37688 7290
rect 37280 6860 37332 6866
rect 37280 6802 37332 6808
rect 37096 6656 37148 6662
rect 37096 6598 37148 6604
rect 37108 6390 37136 6598
rect 37096 6384 37148 6390
rect 37096 6326 37148 6332
rect 36728 5228 36780 5234
rect 36728 5170 36780 5176
rect 37188 4684 37240 4690
rect 37292 4672 37320 6802
rect 37464 6316 37516 6322
rect 37464 6258 37516 6264
rect 37240 4644 37320 4672
rect 37188 4626 37240 4632
rect 37096 4616 37148 4622
rect 37096 4558 37148 4564
rect 36636 4480 36688 4486
rect 36634 4448 36636 4457
rect 36688 4448 36690 4457
rect 36634 4383 36690 4392
rect 36544 4208 36596 4214
rect 36544 4150 36596 4156
rect 36556 3738 36584 4150
rect 36728 3936 36780 3942
rect 36728 3878 36780 3884
rect 36544 3732 36596 3738
rect 36544 3674 36596 3680
rect 36360 3528 36412 3534
rect 36360 3470 36412 3476
rect 36266 3224 36322 3233
rect 36266 3159 36322 3168
rect 36176 2984 36228 2990
rect 36176 2926 36228 2932
rect 36004 2746 36124 2774
rect 35716 1148 35768 1154
rect 35716 1090 35768 1096
rect 35176 870 35388 898
rect 35440 944 35492 950
rect 35440 886 35492 892
rect 35176 800 35204 870
rect 35452 800 35480 886
rect 35728 800 35756 1090
rect 36004 800 36032 2746
rect 36084 2372 36136 2378
rect 36084 2314 36136 2320
rect 36096 1018 36124 2314
rect 36188 1222 36216 2926
rect 36740 2446 36768 3878
rect 36728 2440 36780 2446
rect 36728 2382 36780 2388
rect 36268 1284 36320 1290
rect 36268 1226 36320 1232
rect 36176 1216 36228 1222
rect 36176 1158 36228 1164
rect 36084 1012 36136 1018
rect 36084 954 36136 960
rect 36280 800 36308 1226
rect 36820 1216 36872 1222
rect 36820 1158 36872 1164
rect 36544 1012 36596 1018
rect 36544 954 36596 960
rect 36556 800 36584 954
rect 36832 800 36860 1158
rect 37108 800 37136 4558
rect 37188 4480 37240 4486
rect 37188 4422 37240 4428
rect 37200 4282 37228 4422
rect 37292 4282 37320 4644
rect 37188 4276 37240 4282
rect 37188 4218 37240 4224
rect 37280 4276 37332 4282
rect 37280 4218 37332 4224
rect 37200 4185 37228 4218
rect 37186 4176 37242 4185
rect 37186 4111 37242 4120
rect 37476 3738 37504 6258
rect 37556 6248 37608 6254
rect 37556 6190 37608 6196
rect 37568 6118 37596 6190
rect 37556 6112 37608 6118
rect 37556 6054 37608 6060
rect 37568 5234 37596 6054
rect 37556 5228 37608 5234
rect 37556 5170 37608 5176
rect 37556 4548 37608 4554
rect 37556 4490 37608 4496
rect 37464 3732 37516 3738
rect 37464 3674 37516 3680
rect 37372 3596 37424 3602
rect 37372 3538 37424 3544
rect 37280 2984 37332 2990
rect 37280 2926 37332 2932
rect 37292 950 37320 2926
rect 37280 944 37332 950
rect 37280 886 37332 892
rect 37384 800 37412 3538
rect 37568 2446 37596 4490
rect 37660 2774 37688 7262
rect 37752 6769 37780 11494
rect 37844 7886 37872 12406
rect 38028 11694 38056 12736
rect 38108 12718 38160 12724
rect 38108 12436 38160 12442
rect 38304 12434 38332 14878
rect 38396 14822 38424 15302
rect 38384 14816 38436 14822
rect 38384 14758 38436 14764
rect 38488 13870 38516 15438
rect 38476 13864 38528 13870
rect 38476 13806 38528 13812
rect 38580 12646 38608 15830
rect 38672 15638 38700 15982
rect 38660 15632 38712 15638
rect 38660 15574 38712 15580
rect 38568 12640 38620 12646
rect 38568 12582 38620 12588
rect 38304 12406 38516 12434
rect 38108 12378 38160 12384
rect 38016 11688 38068 11694
rect 38016 11630 38068 11636
rect 38120 11286 38148 12378
rect 38200 11688 38252 11694
rect 38200 11630 38252 11636
rect 38108 11280 38160 11286
rect 38108 11222 38160 11228
rect 38106 10704 38162 10713
rect 38212 10674 38240 11630
rect 38292 11144 38344 11150
rect 38292 11086 38344 11092
rect 38106 10639 38162 10648
rect 38200 10668 38252 10674
rect 38016 9920 38068 9926
rect 38016 9862 38068 9868
rect 37924 8900 37976 8906
rect 37924 8842 37976 8848
rect 37936 8673 37964 8842
rect 37922 8664 37978 8673
rect 37922 8599 37978 8608
rect 37832 7880 37884 7886
rect 37832 7822 37884 7828
rect 37936 6866 37964 8599
rect 37924 6860 37976 6866
rect 37924 6802 37976 6808
rect 37738 6760 37794 6769
rect 37738 6695 37794 6704
rect 37832 6112 37884 6118
rect 37832 6054 37884 6060
rect 37844 5166 37872 6054
rect 38028 5574 38056 9862
rect 38120 8022 38148 10639
rect 38200 10610 38252 10616
rect 38304 9586 38332 11086
rect 38384 10464 38436 10470
rect 38384 10406 38436 10412
rect 38396 9994 38424 10406
rect 38384 9988 38436 9994
rect 38384 9930 38436 9936
rect 38292 9580 38344 9586
rect 38292 9522 38344 9528
rect 38396 9466 38424 9930
rect 38304 9438 38424 9466
rect 38108 8016 38160 8022
rect 38108 7958 38160 7964
rect 38200 7404 38252 7410
rect 38200 7346 38252 7352
rect 38212 7002 38240 7346
rect 38200 6996 38252 7002
rect 38200 6938 38252 6944
rect 38304 6934 38332 9438
rect 38382 7440 38438 7449
rect 38382 7375 38438 7384
rect 38396 7274 38424 7375
rect 38384 7268 38436 7274
rect 38384 7210 38436 7216
rect 38292 6928 38344 6934
rect 38292 6870 38344 6876
rect 38108 6860 38160 6866
rect 38108 6802 38160 6808
rect 38016 5568 38068 5574
rect 38016 5510 38068 5516
rect 37832 5160 37884 5166
rect 37832 5102 37884 5108
rect 37844 4758 37872 5102
rect 38120 4826 38148 6802
rect 38200 6180 38252 6186
rect 38200 6122 38252 6128
rect 38212 5642 38240 6122
rect 38200 5636 38252 5642
rect 38200 5578 38252 5584
rect 38292 5636 38344 5642
rect 38292 5578 38344 5584
rect 38108 4820 38160 4826
rect 38108 4762 38160 4768
rect 37832 4752 37884 4758
rect 37738 4720 37794 4729
rect 37832 4694 37884 4700
rect 37738 4655 37794 4664
rect 37752 4622 37780 4655
rect 37740 4616 37792 4622
rect 37740 4558 37792 4564
rect 38212 4146 38240 5578
rect 38200 4140 38252 4146
rect 38200 4082 38252 4088
rect 38212 3942 38240 4082
rect 38200 3936 38252 3942
rect 38200 3878 38252 3884
rect 37924 3732 37976 3738
rect 37924 3674 37976 3680
rect 37660 2746 37780 2774
rect 37752 2530 37780 2746
rect 37752 2502 37872 2530
rect 37556 2440 37608 2446
rect 37556 2382 37608 2388
rect 37844 2378 37872 2502
rect 37740 2372 37792 2378
rect 37740 2314 37792 2320
rect 37832 2372 37884 2378
rect 37832 2314 37884 2320
rect 37752 1086 37780 2314
rect 37740 1080 37792 1086
rect 37740 1022 37792 1028
rect 37648 944 37700 950
rect 37648 886 37700 892
rect 37660 800 37688 886
rect 37936 800 37964 3674
rect 38200 3664 38252 3670
rect 38200 3606 38252 3612
rect 38212 800 38240 3606
rect 38304 3058 38332 5578
rect 38488 3777 38516 12406
rect 38856 11898 38884 18566
rect 38948 14074 38976 20402
rect 39040 17882 39068 20810
rect 39120 20460 39172 20466
rect 39120 20402 39172 20408
rect 39132 20058 39160 20402
rect 39120 20052 39172 20058
rect 39120 19994 39172 20000
rect 39120 18624 39172 18630
rect 39120 18566 39172 18572
rect 39132 18290 39160 18566
rect 39120 18284 39172 18290
rect 39120 18226 39172 18232
rect 39028 17876 39080 17882
rect 39028 17818 39080 17824
rect 39040 17338 39068 17818
rect 39028 17332 39080 17338
rect 39028 17274 39080 17280
rect 38936 14068 38988 14074
rect 38936 14010 38988 14016
rect 39316 12850 39344 22222
rect 39394 22264 39450 22273
rect 39394 22199 39450 22208
rect 39408 21554 39436 22199
rect 39396 21548 39448 21554
rect 39396 21490 39448 21496
rect 39304 12844 39356 12850
rect 39304 12786 39356 12792
rect 39500 12322 39528 25298
rect 40224 24064 40276 24070
rect 40224 24006 40276 24012
rect 40132 23588 40184 23594
rect 40132 23530 40184 23536
rect 40040 23520 40092 23526
rect 40040 23462 40092 23468
rect 40052 23202 40080 23462
rect 39960 23186 40080 23202
rect 39948 23180 40080 23186
rect 40000 23174 40080 23180
rect 39948 23122 40000 23128
rect 39580 23112 39632 23118
rect 39580 23054 39632 23060
rect 40040 23112 40092 23118
rect 40040 23054 40092 23060
rect 39592 22030 39620 23054
rect 40052 22778 40080 23054
rect 40144 23050 40172 23530
rect 40132 23044 40184 23050
rect 40132 22986 40184 22992
rect 39948 22772 40000 22778
rect 39948 22714 40000 22720
rect 40040 22772 40092 22778
rect 40040 22714 40092 22720
rect 39960 22681 39988 22714
rect 39946 22672 40002 22681
rect 39946 22607 40002 22616
rect 39856 22228 39908 22234
rect 39856 22170 39908 22176
rect 39672 22092 39724 22098
rect 39672 22034 39724 22040
rect 39580 22024 39632 22030
rect 39580 21966 39632 21972
rect 39592 20466 39620 21966
rect 39684 21622 39712 22034
rect 39868 22030 39896 22170
rect 40236 22094 40264 24006
rect 40144 22066 40264 22094
rect 39856 22024 39908 22030
rect 39856 21966 39908 21972
rect 39672 21616 39724 21622
rect 39672 21558 39724 21564
rect 39684 20466 39712 21558
rect 39580 20460 39632 20466
rect 39580 20402 39632 20408
rect 39672 20460 39724 20466
rect 39672 20402 39724 20408
rect 39592 20346 39620 20402
rect 39592 20318 39712 20346
rect 39578 20088 39634 20097
rect 39578 20023 39634 20032
rect 39592 18698 39620 20023
rect 39684 19310 39712 20318
rect 40040 19916 40092 19922
rect 40040 19858 40092 19864
rect 40052 19514 40080 19858
rect 40144 19854 40172 22066
rect 40500 22024 40552 22030
rect 40500 21966 40552 21972
rect 40408 21956 40460 21962
rect 40408 21898 40460 21904
rect 40224 21888 40276 21894
rect 40420 21865 40448 21898
rect 40224 21830 40276 21836
rect 40406 21856 40462 21865
rect 40236 20942 40264 21830
rect 40406 21791 40462 21800
rect 40420 21554 40448 21791
rect 40408 21548 40460 21554
rect 40408 21490 40460 21496
rect 40512 21350 40540 21966
rect 40500 21344 40552 21350
rect 40500 21286 40552 21292
rect 40512 21078 40540 21286
rect 40316 21072 40368 21078
rect 40316 21014 40368 21020
rect 40500 21072 40552 21078
rect 40500 21014 40552 21020
rect 40328 20942 40356 21014
rect 40224 20936 40276 20942
rect 40224 20878 40276 20884
rect 40316 20936 40368 20942
rect 40316 20878 40368 20884
rect 40224 20800 40276 20806
rect 40224 20742 40276 20748
rect 40316 20800 40368 20806
rect 40316 20742 40368 20748
rect 40236 20505 40264 20742
rect 40222 20496 40278 20505
rect 40222 20431 40278 20440
rect 40222 19952 40278 19961
rect 40222 19887 40278 19896
rect 40236 19854 40264 19887
rect 40132 19848 40184 19854
rect 40132 19790 40184 19796
rect 40224 19848 40276 19854
rect 40224 19790 40276 19796
rect 40040 19508 40092 19514
rect 40040 19450 40092 19456
rect 40040 19372 40092 19378
rect 40040 19314 40092 19320
rect 40224 19372 40276 19378
rect 40224 19314 40276 19320
rect 39672 19304 39724 19310
rect 39672 19246 39724 19252
rect 39684 18766 39712 19246
rect 39672 18760 39724 18766
rect 39672 18702 39724 18708
rect 39580 18692 39632 18698
rect 39580 18634 39632 18640
rect 39948 18420 40000 18426
rect 40052 18408 40080 19314
rect 40132 18760 40184 18766
rect 40132 18702 40184 18708
rect 40000 18380 40080 18408
rect 39948 18362 40000 18368
rect 40144 18154 40172 18702
rect 40236 18426 40264 19314
rect 40224 18420 40276 18426
rect 40224 18362 40276 18368
rect 40328 18222 40356 20742
rect 40408 20596 40460 20602
rect 40408 20538 40460 20544
rect 40420 18970 40448 20538
rect 40500 20460 40552 20466
rect 40500 20402 40552 20408
rect 40512 19786 40540 20402
rect 40500 19780 40552 19786
rect 40500 19722 40552 19728
rect 40408 18964 40460 18970
rect 40408 18906 40460 18912
rect 40408 18760 40460 18766
rect 40408 18702 40460 18708
rect 40316 18216 40368 18222
rect 40316 18158 40368 18164
rect 40132 18148 40184 18154
rect 40132 18090 40184 18096
rect 40420 17746 40448 18702
rect 40512 17746 40540 19722
rect 40408 17740 40460 17746
rect 40408 17682 40460 17688
rect 40500 17740 40552 17746
rect 40500 17682 40552 17688
rect 40224 17672 40276 17678
rect 40224 17614 40276 17620
rect 39672 17604 39724 17610
rect 39672 17546 39724 17552
rect 39684 17338 39712 17546
rect 40236 17513 40264 17614
rect 40222 17504 40278 17513
rect 40222 17439 40278 17448
rect 39672 17332 39724 17338
rect 39672 17274 39724 17280
rect 40316 17264 40368 17270
rect 40316 17206 40368 17212
rect 39580 16788 39632 16794
rect 39580 16730 39632 16736
rect 39592 12434 39620 16730
rect 40040 16448 40092 16454
rect 40040 16390 40092 16396
rect 40132 16448 40184 16454
rect 40132 16390 40184 16396
rect 40052 16182 40080 16390
rect 40040 16176 40092 16182
rect 40040 16118 40092 16124
rect 39764 16108 39816 16114
rect 39764 16050 39816 16056
rect 39776 15434 39804 16050
rect 39948 16040 40000 16046
rect 40144 16028 40172 16390
rect 39948 15982 40000 15988
rect 40052 16000 40172 16028
rect 39960 15706 39988 15982
rect 40052 15910 40080 16000
rect 40040 15904 40092 15910
rect 40040 15846 40092 15852
rect 39948 15700 40000 15706
rect 39948 15642 40000 15648
rect 39764 15428 39816 15434
rect 39764 15370 39816 15376
rect 40052 15201 40080 15846
rect 40038 15192 40094 15201
rect 40038 15127 40094 15136
rect 39946 14920 40002 14929
rect 39946 14855 40002 14864
rect 39960 14822 39988 14855
rect 39948 14816 40000 14822
rect 39948 14758 40000 14764
rect 40038 12880 40094 12889
rect 40038 12815 40094 12824
rect 40052 12714 40080 12815
rect 40040 12708 40092 12714
rect 40040 12650 40092 12656
rect 39592 12406 39804 12434
rect 39776 12374 39804 12406
rect 39764 12368 39816 12374
rect 39670 12336 39726 12345
rect 39500 12294 39620 12322
rect 38844 11892 38896 11898
rect 38844 11834 38896 11840
rect 39120 11620 39172 11626
rect 39120 11562 39172 11568
rect 39132 11150 39160 11562
rect 39120 11144 39172 11150
rect 39120 11086 39172 11092
rect 39304 11144 39356 11150
rect 39304 11086 39356 11092
rect 39212 11076 39264 11082
rect 39212 11018 39264 11024
rect 39028 10668 39080 10674
rect 39028 10610 39080 10616
rect 39040 10130 39068 10610
rect 39028 10124 39080 10130
rect 39028 10066 39080 10072
rect 38568 10056 38620 10062
rect 38568 9998 38620 10004
rect 38580 9042 38608 9998
rect 39040 9926 39068 10066
rect 39028 9920 39080 9926
rect 39028 9862 39080 9868
rect 39224 9738 39252 11018
rect 39316 10266 39344 11086
rect 39396 11076 39448 11082
rect 39396 11018 39448 11024
rect 39304 10260 39356 10266
rect 39304 10202 39356 10208
rect 39302 9752 39358 9761
rect 39224 9710 39302 9738
rect 39302 9687 39358 9696
rect 38844 9648 38896 9654
rect 38896 9608 38976 9636
rect 38844 9590 38896 9596
rect 38948 9518 38976 9608
rect 39316 9586 39344 9687
rect 39304 9580 39356 9586
rect 39304 9522 39356 9528
rect 38936 9512 38988 9518
rect 38936 9454 38988 9460
rect 39028 9172 39080 9178
rect 39028 9114 39080 9120
rect 38568 9036 38620 9042
rect 38568 8978 38620 8984
rect 38844 7880 38896 7886
rect 38844 7822 38896 7828
rect 38660 4548 38712 4554
rect 38660 4490 38712 4496
rect 38566 4312 38622 4321
rect 38566 4247 38622 4256
rect 38580 4146 38608 4247
rect 38568 4140 38620 4146
rect 38568 4082 38620 4088
rect 38474 3768 38530 3777
rect 38474 3703 38530 3712
rect 38488 3466 38516 3703
rect 38476 3460 38528 3466
rect 38476 3402 38528 3408
rect 38476 3188 38528 3194
rect 38476 3130 38528 3136
rect 38292 3052 38344 3058
rect 38292 2994 38344 3000
rect 38384 3052 38436 3058
rect 38384 2994 38436 3000
rect 38396 2553 38424 2994
rect 38382 2544 38438 2553
rect 38382 2479 38438 2488
rect 38488 800 38516 3130
rect 38672 3058 38700 4490
rect 38752 4072 38804 4078
rect 38752 4014 38804 4020
rect 38660 3052 38712 3058
rect 38660 2994 38712 3000
rect 38660 2372 38712 2378
rect 38660 2314 38712 2320
rect 38672 1154 38700 2314
rect 38764 1222 38792 4014
rect 38856 2922 38884 7822
rect 39040 6322 39068 9114
rect 39120 8492 39172 8498
rect 39120 8434 39172 8440
rect 39028 6316 39080 6322
rect 39028 6258 39080 6264
rect 38936 5636 38988 5642
rect 38936 5578 38988 5584
rect 38948 3738 38976 5578
rect 39132 5234 39160 8434
rect 39408 8090 39436 11018
rect 39592 11014 39620 12294
rect 39764 12310 39816 12316
rect 39670 12271 39726 12280
rect 39488 11008 39540 11014
rect 39488 10950 39540 10956
rect 39580 11008 39632 11014
rect 39580 10950 39632 10956
rect 39500 10742 39528 10950
rect 39488 10736 39540 10742
rect 39488 10678 39540 10684
rect 39580 10464 39632 10470
rect 39580 10406 39632 10412
rect 39592 10198 39620 10406
rect 39580 10192 39632 10198
rect 39580 10134 39632 10140
rect 39396 8084 39448 8090
rect 39396 8026 39448 8032
rect 39488 7336 39540 7342
rect 39684 7290 39712 12271
rect 39762 10840 39818 10849
rect 39762 10775 39818 10784
rect 39488 7278 39540 7284
rect 39304 6724 39356 6730
rect 39304 6666 39356 6672
rect 39316 6322 39344 6666
rect 39500 6458 39528 7278
rect 39592 7262 39712 7290
rect 39488 6452 39540 6458
rect 39488 6394 39540 6400
rect 39592 6338 39620 7262
rect 39672 7200 39724 7206
rect 39672 7142 39724 7148
rect 39684 7002 39712 7142
rect 39672 6996 39724 7002
rect 39672 6938 39724 6944
rect 39304 6316 39356 6322
rect 39304 6258 39356 6264
rect 39500 6310 39620 6338
rect 39304 6180 39356 6186
rect 39304 6122 39356 6128
rect 39120 5228 39172 5234
rect 39120 5170 39172 5176
rect 39118 4448 39174 4457
rect 39118 4383 39174 4392
rect 39132 4214 39160 4383
rect 39212 4276 39264 4282
rect 39212 4218 39264 4224
rect 39120 4208 39172 4214
rect 39120 4150 39172 4156
rect 39028 4140 39080 4146
rect 39028 4082 39080 4088
rect 39040 3913 39068 4082
rect 39120 4072 39172 4078
rect 39120 4014 39172 4020
rect 39026 3904 39082 3913
rect 39026 3839 39082 3848
rect 38936 3732 38988 3738
rect 38936 3674 38988 3680
rect 39132 3466 39160 4014
rect 39224 3534 39252 4218
rect 39212 3528 39264 3534
rect 39212 3470 39264 3476
rect 39120 3460 39172 3466
rect 39120 3402 39172 3408
rect 39132 3126 39160 3402
rect 39120 3120 39172 3126
rect 39120 3062 39172 3068
rect 38844 2916 38896 2922
rect 38844 2858 38896 2864
rect 39224 2582 39252 3470
rect 39212 2576 39264 2582
rect 39212 2518 39264 2524
rect 39316 2446 39344 6122
rect 39396 5228 39448 5234
rect 39396 5170 39448 5176
rect 39408 4826 39436 5170
rect 39396 4820 39448 4826
rect 39396 4762 39448 4768
rect 39396 3528 39448 3534
rect 39396 3470 39448 3476
rect 39408 3058 39436 3470
rect 39396 3052 39448 3058
rect 39396 2994 39448 3000
rect 39304 2440 39356 2446
rect 39304 2382 39356 2388
rect 39500 1834 39528 6310
rect 39580 5704 39632 5710
rect 39580 5646 39632 5652
rect 39488 1828 39540 1834
rect 39488 1770 39540 1776
rect 38752 1216 38804 1222
rect 38752 1158 38804 1164
rect 39028 1216 39080 1222
rect 39028 1158 39080 1164
rect 38660 1148 38712 1154
rect 38660 1090 38712 1096
rect 38752 944 38804 950
rect 38752 886 38804 892
rect 38764 800 38792 886
rect 39040 800 39068 1158
rect 39304 1080 39356 1086
rect 39304 1022 39356 1028
rect 39316 800 39344 1022
rect 39592 800 39620 5646
rect 39672 2984 39724 2990
rect 39672 2926 39724 2932
rect 39684 1290 39712 2926
rect 39776 2650 39804 10775
rect 40224 10464 40276 10470
rect 40224 10406 40276 10412
rect 40236 9654 40264 10406
rect 40224 9648 40276 9654
rect 40224 9590 40276 9596
rect 39856 6792 39908 6798
rect 39856 6734 39908 6740
rect 39948 6792 40000 6798
rect 39948 6734 40000 6740
rect 39868 6458 39896 6734
rect 39856 6452 39908 6458
rect 39856 6394 39908 6400
rect 39960 5914 39988 6734
rect 40224 6656 40276 6662
rect 40224 6598 40276 6604
rect 40040 6316 40092 6322
rect 40040 6258 40092 6264
rect 40052 6118 40080 6258
rect 40040 6112 40092 6118
rect 40040 6054 40092 6060
rect 39948 5908 40000 5914
rect 39948 5850 40000 5856
rect 40236 5778 40264 6598
rect 40328 5914 40356 17206
rect 40500 15020 40552 15026
rect 40500 14962 40552 14968
rect 40512 14618 40540 14962
rect 40500 14612 40552 14618
rect 40500 14554 40552 14560
rect 40604 12434 40632 40462
rect 41432 38282 41460 44338
rect 41708 43790 41736 44406
rect 41696 43784 41748 43790
rect 41696 43726 41748 43732
rect 41420 38276 41472 38282
rect 41420 38218 41472 38224
rect 41144 35556 41196 35562
rect 41144 35498 41196 35504
rect 41156 34746 41184 35498
rect 41144 34740 41196 34746
rect 41144 34682 41196 34688
rect 41432 30802 41460 38218
rect 41696 34536 41748 34542
rect 41696 34478 41748 34484
rect 41420 30796 41472 30802
rect 41420 30738 41472 30744
rect 41708 28490 41736 34478
rect 41880 30048 41932 30054
rect 41880 29990 41932 29996
rect 41696 28484 41748 28490
rect 41696 28426 41748 28432
rect 41236 28416 41288 28422
rect 41236 28358 41288 28364
rect 40684 24812 40736 24818
rect 40684 24754 40736 24760
rect 40512 12406 40632 12434
rect 40696 12434 40724 24754
rect 40776 24608 40828 24614
rect 40776 24550 40828 24556
rect 40788 17270 40816 24550
rect 40868 23724 40920 23730
rect 40868 23666 40920 23672
rect 40880 21622 40908 23666
rect 41144 23044 41196 23050
rect 41144 22986 41196 22992
rect 40960 22704 41012 22710
rect 40960 22646 41012 22652
rect 40972 22080 41000 22646
rect 40972 22052 41092 22080
rect 40868 21616 40920 21622
rect 40868 21558 40920 21564
rect 40868 20596 40920 20602
rect 40868 20538 40920 20544
rect 40880 19854 40908 20538
rect 41064 20466 41092 22052
rect 41052 20460 41104 20466
rect 41052 20402 41104 20408
rect 41156 20346 41184 22986
rect 41248 21876 41276 28358
rect 41788 26036 41840 26042
rect 41788 25978 41840 25984
rect 41800 25906 41828 25978
rect 41788 25900 41840 25906
rect 41788 25842 41840 25848
rect 41328 24404 41380 24410
rect 41328 24346 41380 24352
rect 41340 23594 41368 24346
rect 41696 23724 41748 23730
rect 41696 23666 41748 23672
rect 41328 23588 41380 23594
rect 41328 23530 41380 23536
rect 41420 23180 41472 23186
rect 41340 23140 41420 23168
rect 41340 23050 41368 23140
rect 41420 23122 41472 23128
rect 41708 23089 41736 23666
rect 41892 23118 41920 29990
rect 42168 28558 42196 47398
rect 42352 45354 42380 52430
rect 42536 51406 42564 52430
rect 42708 52352 42760 52358
rect 42708 52294 42760 52300
rect 42524 51400 42576 51406
rect 42524 51342 42576 51348
rect 42536 49842 42564 51342
rect 42524 49836 42576 49842
rect 42524 49778 42576 49784
rect 42536 45554 42564 49778
rect 42616 49768 42668 49774
rect 42614 49736 42616 49745
rect 42668 49736 42670 49745
rect 42614 49671 42670 49680
rect 42536 45526 42656 45554
rect 42340 45348 42392 45354
rect 42340 45290 42392 45296
rect 42628 44470 42656 45526
rect 42616 44464 42668 44470
rect 42616 44406 42668 44412
rect 42248 35080 42300 35086
rect 42248 35022 42300 35028
rect 42260 32910 42288 35022
rect 42432 34672 42484 34678
rect 42432 34614 42484 34620
rect 42248 32904 42300 32910
rect 42248 32846 42300 32852
rect 42156 28552 42208 28558
rect 42156 28494 42208 28500
rect 42064 28484 42116 28490
rect 42064 28426 42116 28432
rect 42076 25974 42104 28426
rect 42064 25968 42116 25974
rect 42064 25910 42116 25916
rect 42156 23860 42208 23866
rect 42156 23802 42208 23808
rect 42168 23730 42196 23802
rect 42156 23724 42208 23730
rect 42156 23666 42208 23672
rect 41880 23112 41932 23118
rect 41694 23080 41750 23089
rect 41328 23044 41380 23050
rect 41694 23015 41750 23024
rect 41800 23060 41880 23066
rect 41972 23112 42024 23118
rect 41800 23054 41932 23060
rect 41970 23080 41972 23089
rect 42064 23112 42116 23118
rect 42024 23080 42026 23089
rect 41800 23038 41920 23054
rect 41328 22986 41380 22992
rect 41512 22976 41564 22982
rect 41512 22918 41564 22924
rect 41328 22568 41380 22574
rect 41328 22510 41380 22516
rect 41340 22030 41368 22510
rect 41420 22500 41472 22506
rect 41420 22442 41472 22448
rect 41328 22024 41380 22030
rect 41328 21966 41380 21972
rect 41432 21962 41460 22442
rect 41420 21956 41472 21962
rect 41420 21898 41472 21904
rect 41248 21848 41368 21876
rect 41236 21616 41288 21622
rect 41236 21558 41288 21564
rect 41248 20874 41276 21558
rect 41236 20868 41288 20874
rect 41236 20810 41288 20816
rect 41340 20754 41368 21848
rect 41432 21418 41460 21898
rect 41420 21412 41472 21418
rect 41420 21354 41472 21360
rect 41524 20942 41552 22918
rect 41604 22772 41656 22778
rect 41604 22714 41656 22720
rect 41616 22642 41644 22714
rect 41604 22636 41656 22642
rect 41604 22578 41656 22584
rect 41604 21888 41656 21894
rect 41604 21830 41656 21836
rect 41616 21690 41644 21830
rect 41604 21684 41656 21690
rect 41604 21626 41656 21632
rect 41512 20936 41564 20942
rect 41512 20878 41564 20884
rect 41064 20318 41184 20346
rect 41248 20726 41368 20754
rect 40868 19848 40920 19854
rect 40866 19816 40868 19825
rect 40920 19816 40922 19825
rect 40866 19751 40922 19760
rect 40960 19780 41012 19786
rect 40960 19722 41012 19728
rect 40972 19514 41000 19722
rect 40960 19508 41012 19514
rect 40960 19450 41012 19456
rect 40868 18896 40920 18902
rect 40868 18838 40920 18844
rect 40880 18086 40908 18838
rect 40868 18080 40920 18086
rect 40868 18022 40920 18028
rect 40868 17536 40920 17542
rect 40868 17478 40920 17484
rect 40880 17270 40908 17478
rect 40776 17264 40828 17270
rect 40776 17206 40828 17212
rect 40868 17264 40920 17270
rect 40868 17206 40920 17212
rect 41064 16590 41092 20318
rect 41144 20256 41196 20262
rect 41144 20198 41196 20204
rect 41156 19922 41184 20198
rect 41144 19916 41196 19922
rect 41144 19858 41196 19864
rect 41144 19508 41196 19514
rect 41144 19450 41196 19456
rect 41156 18766 41184 19450
rect 41248 19378 41276 20726
rect 41696 20460 41748 20466
rect 41696 20402 41748 20408
rect 41512 20324 41564 20330
rect 41512 20266 41564 20272
rect 41420 19848 41472 19854
rect 41420 19790 41472 19796
rect 41328 19712 41380 19718
rect 41328 19654 41380 19660
rect 41236 19372 41288 19378
rect 41236 19314 41288 19320
rect 41340 19174 41368 19654
rect 41328 19168 41380 19174
rect 41328 19110 41380 19116
rect 41144 18760 41196 18766
rect 41144 18702 41196 18708
rect 41432 18426 41460 19790
rect 41524 18834 41552 20266
rect 41708 19718 41736 20402
rect 41696 19712 41748 19718
rect 41696 19654 41748 19660
rect 41604 19168 41656 19174
rect 41604 19110 41656 19116
rect 41512 18828 41564 18834
rect 41512 18770 41564 18776
rect 41420 18420 41472 18426
rect 41420 18362 41472 18368
rect 41616 18290 41644 19110
rect 41696 18828 41748 18834
rect 41696 18770 41748 18776
rect 41604 18284 41656 18290
rect 41604 18226 41656 18232
rect 41708 18154 41736 18770
rect 41696 18148 41748 18154
rect 41696 18090 41748 18096
rect 41328 17740 41380 17746
rect 41328 17682 41380 17688
rect 41236 17536 41288 17542
rect 41236 17478 41288 17484
rect 41248 17202 41276 17478
rect 41236 17196 41288 17202
rect 41236 17138 41288 17144
rect 41144 16652 41196 16658
rect 41144 16594 41196 16600
rect 41052 16584 41104 16590
rect 41052 16526 41104 16532
rect 40776 15496 40828 15502
rect 41156 15450 41184 16594
rect 41236 15904 41288 15910
rect 41236 15846 41288 15852
rect 41248 15502 41276 15846
rect 40828 15444 41184 15450
rect 40776 15438 41184 15444
rect 41236 15496 41288 15502
rect 41236 15438 41288 15444
rect 40788 15422 41184 15438
rect 40960 14816 41012 14822
rect 40960 14758 41012 14764
rect 40972 14482 41000 14758
rect 41156 14482 41184 15422
rect 40960 14476 41012 14482
rect 40960 14418 41012 14424
rect 41144 14476 41196 14482
rect 41144 14418 41196 14424
rect 41156 13258 41184 14418
rect 41144 13252 41196 13258
rect 41144 13194 41196 13200
rect 40696 12406 40816 12434
rect 40512 9568 40540 12406
rect 40592 11688 40644 11694
rect 40592 11630 40644 11636
rect 40604 11218 40632 11630
rect 40592 11212 40644 11218
rect 40592 11154 40644 11160
rect 40512 9540 40632 9568
rect 40500 6792 40552 6798
rect 40500 6734 40552 6740
rect 40512 6458 40540 6734
rect 40500 6452 40552 6458
rect 40500 6394 40552 6400
rect 40500 6316 40552 6322
rect 40500 6258 40552 6264
rect 40316 5908 40368 5914
rect 40316 5850 40368 5856
rect 40512 5817 40540 6258
rect 40498 5808 40554 5817
rect 40224 5772 40276 5778
rect 40498 5743 40554 5752
rect 40224 5714 40276 5720
rect 40040 5568 40092 5574
rect 40040 5510 40092 5516
rect 40052 4146 40080 5510
rect 40512 5370 40540 5743
rect 40224 5364 40276 5370
rect 40224 5306 40276 5312
rect 40500 5364 40552 5370
rect 40500 5306 40552 5312
rect 40132 4752 40184 4758
rect 40132 4694 40184 4700
rect 40144 4486 40172 4694
rect 40236 4690 40264 5306
rect 40512 4706 40540 5306
rect 40224 4684 40276 4690
rect 40224 4626 40276 4632
rect 40328 4678 40540 4706
rect 40328 4486 40356 4678
rect 40408 4616 40460 4622
rect 40408 4558 40460 4564
rect 40132 4480 40184 4486
rect 40132 4422 40184 4428
rect 40316 4480 40368 4486
rect 40316 4422 40368 4428
rect 40132 4276 40184 4282
rect 40132 4218 40184 4224
rect 40040 4140 40092 4146
rect 40040 4082 40092 4088
rect 40040 3936 40092 3942
rect 40040 3878 40092 3884
rect 40052 3466 40080 3878
rect 40040 3460 40092 3466
rect 40040 3402 40092 3408
rect 39764 2644 39816 2650
rect 39764 2586 39816 2592
rect 39672 1284 39724 1290
rect 39672 1226 39724 1232
rect 39856 1148 39908 1154
rect 39856 1090 39908 1096
rect 39868 800 39896 1090
rect 40144 800 40172 4218
rect 40224 3936 40276 3942
rect 40222 3904 40224 3913
rect 40276 3904 40278 3913
rect 40222 3839 40278 3848
rect 40316 2372 40368 2378
rect 40316 2314 40368 2320
rect 40328 1018 40356 2314
rect 40316 1012 40368 1018
rect 40316 954 40368 960
rect 40420 800 40448 4558
rect 40604 2922 40632 9540
rect 40684 8832 40736 8838
rect 40684 8774 40736 8780
rect 40696 8498 40724 8774
rect 40684 8492 40736 8498
rect 40684 8434 40736 8440
rect 40684 6928 40736 6934
rect 40684 6870 40736 6876
rect 40696 4690 40724 6870
rect 40684 4684 40736 4690
rect 40684 4626 40736 4632
rect 40696 4457 40724 4626
rect 40682 4448 40738 4457
rect 40682 4383 40738 4392
rect 40788 4078 40816 12406
rect 41340 12170 41368 17682
rect 41800 16250 41828 23038
rect 42064 23054 42116 23060
rect 41970 23015 42026 23024
rect 41984 20534 42012 23015
rect 42076 21690 42104 23054
rect 42064 21684 42116 21690
rect 42064 21626 42116 21632
rect 42168 20874 42196 23666
rect 42248 23112 42300 23118
rect 42248 23054 42300 23060
rect 42260 22642 42288 23054
rect 42340 22976 42392 22982
rect 42340 22918 42392 22924
rect 42248 22636 42300 22642
rect 42248 22578 42300 22584
rect 42246 22400 42302 22409
rect 42246 22335 42302 22344
rect 42260 21842 42288 22335
rect 42352 22030 42380 22918
rect 42340 22024 42392 22030
rect 42340 21966 42392 21972
rect 42260 21814 42380 21842
rect 42156 20868 42208 20874
rect 42156 20810 42208 20816
rect 41972 20528 42024 20534
rect 41972 20470 42024 20476
rect 41972 20392 42024 20398
rect 41972 20334 42024 20340
rect 41880 20256 41932 20262
rect 41880 20198 41932 20204
rect 41892 19990 41920 20198
rect 41880 19984 41932 19990
rect 41880 19926 41932 19932
rect 41984 19310 42012 20334
rect 42064 20256 42116 20262
rect 42064 20198 42116 20204
rect 42076 19922 42104 20198
rect 42168 19990 42196 20810
rect 42156 19984 42208 19990
rect 42156 19926 42208 19932
rect 42064 19916 42116 19922
rect 42064 19858 42116 19864
rect 41972 19304 42024 19310
rect 41972 19246 42024 19252
rect 41984 18630 42012 19246
rect 42076 18766 42104 19858
rect 42156 19712 42208 19718
rect 42156 19654 42208 19660
rect 42064 18760 42116 18766
rect 42064 18702 42116 18708
rect 41972 18624 42024 18630
rect 41972 18566 42024 18572
rect 42064 18624 42116 18630
rect 42168 18612 42196 19654
rect 42116 18584 42196 18612
rect 42064 18566 42116 18572
rect 41880 18284 41932 18290
rect 41880 18226 41932 18232
rect 41892 17882 41920 18226
rect 41972 18216 42024 18222
rect 41972 18158 42024 18164
rect 41880 17876 41932 17882
rect 41880 17818 41932 17824
rect 41892 17678 41920 17818
rect 41984 17814 42012 18158
rect 41972 17808 42024 17814
rect 41972 17750 42024 17756
rect 41880 17672 41932 17678
rect 41880 17614 41932 17620
rect 41880 17128 41932 17134
rect 41880 17070 41932 17076
rect 41788 16244 41840 16250
rect 41788 16186 41840 16192
rect 41696 16040 41748 16046
rect 41696 15982 41748 15988
rect 41708 15638 41736 15982
rect 41696 15632 41748 15638
rect 41696 15574 41748 15580
rect 41696 12640 41748 12646
rect 41696 12582 41748 12588
rect 41328 12164 41380 12170
rect 41328 12106 41380 12112
rect 41512 12096 41564 12102
rect 41512 12038 41564 12044
rect 41524 11830 41552 12038
rect 41512 11824 41564 11830
rect 41512 11766 41564 11772
rect 41418 9752 41474 9761
rect 41418 9687 41474 9696
rect 40868 9648 40920 9654
rect 40868 9590 40920 9596
rect 40880 4758 40908 9590
rect 41144 8832 41196 8838
rect 41144 8774 41196 8780
rect 41156 8634 41184 8774
rect 41144 8628 41196 8634
rect 41144 8570 41196 8576
rect 41432 7002 41460 9687
rect 41420 6996 41472 7002
rect 41420 6938 41472 6944
rect 41234 5400 41290 5409
rect 41234 5335 41236 5344
rect 41288 5335 41290 5344
rect 41236 5306 41288 5312
rect 41052 5228 41104 5234
rect 41052 5170 41104 5176
rect 41236 5228 41288 5234
rect 41236 5170 41288 5176
rect 40868 4752 40920 4758
rect 40868 4694 40920 4700
rect 40776 4072 40828 4078
rect 40776 4014 40828 4020
rect 40880 3058 40908 4694
rect 41064 4282 41092 5170
rect 41052 4276 41104 4282
rect 41052 4218 41104 4224
rect 41052 4140 41104 4146
rect 41052 4082 41104 4088
rect 41064 3466 41092 4082
rect 41052 3460 41104 3466
rect 41052 3402 41104 3408
rect 40960 3392 41012 3398
rect 40960 3334 41012 3340
rect 40868 3052 40920 3058
rect 40868 2994 40920 3000
rect 40592 2916 40644 2922
rect 40592 2858 40644 2864
rect 40972 2774 41000 3334
rect 40880 2746 41000 2774
rect 40880 2310 40908 2746
rect 40960 2372 41012 2378
rect 40960 2314 41012 2320
rect 40868 2304 40920 2310
rect 40868 2246 40920 2252
rect 40684 944 40736 950
rect 40684 886 40736 892
rect 40696 800 40724 886
rect 40972 800 41000 2314
rect 41248 800 41276 5170
rect 41328 4548 41380 4554
rect 41328 4490 41380 4496
rect 41340 3194 41368 4490
rect 41708 3194 41736 12582
rect 41892 12238 41920 17070
rect 41984 16522 42012 17750
rect 42076 17377 42104 18566
rect 42248 17672 42300 17678
rect 42248 17614 42300 17620
rect 42062 17368 42118 17377
rect 42062 17303 42118 17312
rect 42260 16590 42288 17614
rect 42248 16584 42300 16590
rect 42248 16526 42300 16532
rect 41972 16516 42024 16522
rect 41972 16458 42024 16464
rect 42260 15706 42288 16526
rect 42248 15700 42300 15706
rect 42248 15642 42300 15648
rect 42154 13832 42210 13841
rect 42154 13767 42210 13776
rect 41880 12232 41932 12238
rect 41880 12174 41932 12180
rect 41972 12096 42024 12102
rect 41972 12038 42024 12044
rect 41984 11558 42012 12038
rect 41972 11552 42024 11558
rect 41972 11494 42024 11500
rect 41984 10169 42012 11494
rect 41970 10160 42026 10169
rect 41970 10095 42026 10104
rect 41970 9616 42026 9625
rect 41970 9551 42026 9560
rect 41880 9444 41932 9450
rect 41880 9386 41932 9392
rect 41892 5098 41920 9386
rect 41984 5098 42012 9551
rect 41880 5092 41932 5098
rect 41880 5034 41932 5040
rect 41972 5092 42024 5098
rect 41972 5034 42024 5040
rect 42168 4826 42196 13767
rect 42352 8974 42380 21814
rect 42340 8968 42392 8974
rect 42340 8910 42392 8916
rect 42444 5098 42472 34614
rect 42720 34066 42748 52294
rect 43076 50176 43128 50182
rect 43076 50118 43128 50124
rect 43088 49842 43116 50118
rect 43076 49836 43128 49842
rect 43076 49778 43128 49784
rect 43260 49836 43312 49842
rect 43260 49778 43312 49784
rect 43076 47592 43128 47598
rect 43076 47534 43128 47540
rect 42892 43716 42944 43722
rect 42892 43658 42944 43664
rect 42904 43450 42932 43658
rect 42892 43444 42944 43450
rect 42892 43386 42944 43392
rect 43088 41449 43116 47534
rect 43074 41440 43130 41449
rect 43074 41375 43130 41384
rect 43272 35086 43300 49778
rect 42800 35080 42852 35086
rect 42800 35022 42852 35028
rect 43260 35080 43312 35086
rect 43260 35022 43312 35028
rect 42812 34746 42840 35022
rect 42800 34740 42852 34746
rect 42800 34682 42852 34688
rect 43640 34610 43668 57190
rect 43720 40452 43772 40458
rect 43720 40394 43772 40400
rect 43732 35630 43760 40394
rect 45008 36032 45060 36038
rect 45008 35974 45060 35980
rect 43720 35624 43772 35630
rect 43720 35566 43772 35572
rect 43732 34610 43760 35566
rect 42800 34604 42852 34610
rect 42800 34546 42852 34552
rect 43628 34604 43680 34610
rect 43628 34546 43680 34552
rect 43720 34604 43772 34610
rect 43720 34546 43772 34552
rect 42812 34134 42840 34546
rect 42984 34400 43036 34406
rect 42984 34342 43036 34348
rect 42800 34128 42852 34134
rect 42800 34070 42852 34076
rect 42708 34060 42760 34066
rect 42708 34002 42760 34008
rect 42616 27872 42668 27878
rect 42616 27814 42668 27820
rect 42524 23112 42576 23118
rect 42524 23054 42576 23060
rect 42536 22506 42564 23054
rect 42628 22778 42656 27814
rect 42800 26988 42852 26994
rect 42800 26930 42852 26936
rect 42812 26382 42840 26930
rect 42996 26874 43024 34342
rect 43076 33992 43128 33998
rect 43076 33934 43128 33940
rect 43168 33992 43220 33998
rect 43168 33934 43220 33940
rect 43088 32502 43116 33934
rect 43076 32496 43128 32502
rect 43076 32438 43128 32444
rect 43180 26994 43208 33934
rect 43904 30864 43956 30870
rect 43904 30806 43956 30812
rect 43168 26988 43220 26994
rect 43168 26930 43220 26936
rect 42996 26846 43668 26874
rect 43260 26512 43312 26518
rect 43260 26454 43312 26460
rect 43272 26382 43300 26454
rect 42800 26376 42852 26382
rect 42800 26318 42852 26324
rect 43076 26376 43128 26382
rect 43076 26318 43128 26324
rect 43260 26376 43312 26382
rect 43260 26318 43312 26324
rect 42984 24676 43036 24682
rect 42984 24618 43036 24624
rect 42800 24200 42852 24206
rect 42800 24142 42852 24148
rect 42708 23792 42760 23798
rect 42708 23734 42760 23740
rect 42720 22778 42748 23734
rect 42812 23168 42840 24142
rect 42892 23656 42944 23662
rect 42892 23598 42944 23604
rect 42904 23322 42932 23598
rect 42892 23316 42944 23322
rect 42892 23258 42944 23264
rect 42812 23140 42932 23168
rect 42616 22772 42668 22778
rect 42616 22714 42668 22720
rect 42708 22772 42760 22778
rect 42708 22714 42760 22720
rect 42524 22500 42576 22506
rect 42524 22442 42576 22448
rect 42628 22409 42656 22714
rect 42706 22672 42762 22681
rect 42706 22607 42708 22616
rect 42760 22607 42762 22616
rect 42708 22578 42760 22584
rect 42708 22432 42760 22438
rect 42614 22400 42670 22409
rect 42708 22374 42760 22380
rect 42614 22335 42670 22344
rect 42616 22024 42668 22030
rect 42616 21966 42668 21972
rect 42628 21690 42656 21966
rect 42616 21684 42668 21690
rect 42616 21626 42668 21632
rect 42720 21554 42748 22374
rect 42800 22092 42852 22098
rect 42800 22034 42852 22040
rect 42812 21690 42840 22034
rect 42800 21684 42852 21690
rect 42800 21626 42852 21632
rect 42904 21570 42932 23140
rect 42524 21548 42576 21554
rect 42524 21490 42576 21496
rect 42708 21548 42760 21554
rect 42708 21490 42760 21496
rect 42812 21542 42932 21570
rect 42536 20942 42564 21490
rect 42524 20936 42576 20942
rect 42524 20878 42576 20884
rect 42812 20874 42840 21542
rect 42996 21321 43024 24618
rect 42982 21312 43038 21321
rect 42982 21247 43038 21256
rect 42800 20868 42852 20874
rect 42800 20810 42852 20816
rect 42812 20641 42840 20810
rect 42798 20632 42854 20641
rect 42798 20567 42854 20576
rect 42616 20460 42668 20466
rect 42616 20402 42668 20408
rect 42628 19922 42656 20402
rect 42616 19916 42668 19922
rect 42616 19858 42668 19864
rect 42984 19848 43036 19854
rect 42984 19790 43036 19796
rect 42708 19440 42760 19446
rect 42708 19382 42760 19388
rect 42720 19334 42748 19382
rect 42628 19306 42748 19334
rect 42628 18222 42656 19306
rect 42708 18760 42760 18766
rect 42708 18702 42760 18708
rect 42720 18426 42748 18702
rect 42708 18420 42760 18426
rect 42708 18362 42760 18368
rect 42616 18216 42668 18222
rect 42616 18158 42668 18164
rect 42616 17604 42668 17610
rect 42616 17546 42668 17552
rect 42628 17338 42656 17546
rect 42708 17536 42760 17542
rect 42708 17478 42760 17484
rect 42720 17338 42748 17478
rect 42616 17332 42668 17338
rect 42616 17274 42668 17280
rect 42708 17332 42760 17338
rect 42708 17274 42760 17280
rect 42800 17196 42852 17202
rect 42800 17138 42852 17144
rect 42812 16250 42840 17138
rect 42800 16244 42852 16250
rect 42800 16186 42852 16192
rect 42800 15088 42852 15094
rect 42800 15030 42852 15036
rect 42812 13954 42840 15030
rect 42720 13938 42932 13954
rect 42708 13932 42932 13938
rect 42760 13926 42932 13932
rect 42708 13874 42760 13880
rect 42708 12096 42760 12102
rect 42708 12038 42760 12044
rect 42720 11150 42748 12038
rect 42800 11756 42852 11762
rect 42800 11698 42852 11704
rect 42708 11144 42760 11150
rect 42708 11086 42760 11092
rect 42812 9042 42840 11698
rect 42904 11694 42932 13926
rect 42996 12850 43024 19790
rect 43088 18222 43116 26318
rect 43168 26308 43220 26314
rect 43168 26250 43220 26256
rect 43180 19854 43208 26250
rect 43260 25900 43312 25906
rect 43260 25842 43312 25848
rect 43444 25900 43496 25906
rect 43444 25842 43496 25848
rect 43272 25294 43300 25842
rect 43260 25288 43312 25294
rect 43260 25230 43312 25236
rect 43456 24993 43484 25842
rect 43442 24984 43498 24993
rect 43442 24919 43498 24928
rect 43444 23180 43496 23186
rect 43444 23122 43496 23128
rect 43456 22710 43484 23122
rect 43444 22704 43496 22710
rect 43444 22646 43496 22652
rect 43352 22636 43404 22642
rect 43352 22578 43404 22584
rect 43364 21894 43392 22578
rect 43536 22432 43588 22438
rect 43536 22374 43588 22380
rect 43444 21956 43496 21962
rect 43444 21898 43496 21904
rect 43352 21888 43404 21894
rect 43352 21830 43404 21836
rect 43364 21690 43392 21830
rect 43352 21684 43404 21690
rect 43352 21626 43404 21632
rect 43456 21554 43484 21898
rect 43444 21548 43496 21554
rect 43444 21490 43496 21496
rect 43260 21072 43312 21078
rect 43260 21014 43312 21020
rect 43168 19848 43220 19854
rect 43168 19790 43220 19796
rect 43272 18630 43300 21014
rect 43352 20936 43404 20942
rect 43456 20924 43484 21490
rect 43548 21146 43576 22374
rect 43640 22094 43668 26846
rect 43720 26852 43772 26858
rect 43720 26794 43772 26800
rect 43732 26314 43760 26794
rect 43720 26308 43772 26314
rect 43720 26250 43772 26256
rect 43812 25900 43864 25906
rect 43812 25842 43864 25848
rect 43824 25430 43852 25842
rect 43812 25424 43864 25430
rect 43812 25366 43864 25372
rect 43812 22976 43864 22982
rect 43812 22918 43864 22924
rect 43640 22066 43760 22094
rect 43536 21140 43588 21146
rect 43536 21082 43588 21088
rect 43404 20896 43484 20924
rect 43352 20878 43404 20884
rect 43352 20800 43404 20806
rect 43352 20742 43404 20748
rect 43364 19854 43392 20742
rect 43352 19848 43404 19854
rect 43352 19790 43404 19796
rect 43456 19446 43484 20896
rect 43628 20936 43680 20942
rect 43628 20878 43680 20884
rect 43536 20460 43588 20466
rect 43536 20402 43588 20408
rect 43548 20058 43576 20402
rect 43536 20052 43588 20058
rect 43536 19994 43588 20000
rect 43444 19440 43496 19446
rect 43444 19382 43496 19388
rect 43444 18760 43496 18766
rect 43444 18702 43496 18708
rect 43260 18624 43312 18630
rect 43260 18566 43312 18572
rect 43076 18216 43128 18222
rect 43076 18158 43128 18164
rect 43456 18086 43484 18702
rect 43076 18080 43128 18086
rect 43444 18080 43496 18086
rect 43076 18022 43128 18028
rect 43442 18048 43444 18057
rect 43496 18048 43498 18057
rect 43088 17202 43116 18022
rect 43442 17983 43498 17992
rect 43076 17196 43128 17202
rect 43076 17138 43128 17144
rect 43260 17196 43312 17202
rect 43260 17138 43312 17144
rect 43076 17060 43128 17066
rect 43076 17002 43128 17008
rect 43088 16182 43116 17002
rect 43166 16688 43222 16697
rect 43166 16623 43222 16632
rect 43076 16176 43128 16182
rect 43076 16118 43128 16124
rect 43076 15904 43128 15910
rect 43076 15846 43128 15852
rect 43088 15434 43116 15846
rect 43076 15428 43128 15434
rect 43076 15370 43128 15376
rect 43180 14090 43208 16623
rect 43272 15910 43300 17138
rect 43352 16516 43404 16522
rect 43352 16458 43404 16464
rect 43364 16114 43392 16458
rect 43352 16108 43404 16114
rect 43352 16050 43404 16056
rect 43260 15904 43312 15910
rect 43260 15846 43312 15852
rect 43536 15428 43588 15434
rect 43536 15370 43588 15376
rect 43548 15162 43576 15370
rect 43536 15156 43588 15162
rect 43536 15098 43588 15104
rect 43536 14952 43588 14958
rect 43536 14894 43588 14900
rect 43180 14062 43300 14090
rect 43168 13932 43220 13938
rect 43168 13874 43220 13880
rect 43076 13184 43128 13190
rect 43076 13126 43128 13132
rect 43088 12918 43116 13126
rect 43076 12912 43128 12918
rect 43076 12854 43128 12860
rect 42984 12844 43036 12850
rect 42984 12786 43036 12792
rect 43180 12646 43208 13874
rect 43168 12640 43220 12646
rect 43168 12582 43220 12588
rect 43272 12434 43300 14062
rect 43352 13252 43404 13258
rect 43352 13194 43404 13200
rect 43364 12782 43392 13194
rect 43548 13025 43576 14894
rect 43534 13016 43590 13025
rect 43534 12951 43590 12960
rect 43352 12776 43404 12782
rect 43352 12718 43404 12724
rect 43180 12406 43300 12434
rect 42984 12300 43036 12306
rect 42984 12242 43036 12248
rect 42996 11898 43024 12242
rect 43076 12096 43128 12102
rect 43076 12038 43128 12044
rect 42984 11892 43036 11898
rect 42984 11834 43036 11840
rect 42892 11688 42944 11694
rect 42892 11630 42944 11636
rect 43088 11286 43116 12038
rect 43076 11280 43128 11286
rect 43074 11248 43076 11257
rect 43128 11248 43130 11257
rect 43074 11183 43130 11192
rect 43074 9752 43130 9761
rect 43074 9687 43130 9696
rect 42800 9036 42852 9042
rect 42800 8978 42852 8984
rect 42720 8498 42840 8514
rect 42708 8492 42840 8498
rect 42760 8486 42840 8492
rect 42708 8434 42760 8440
rect 42616 8288 42668 8294
rect 42616 8230 42668 8236
rect 42628 6633 42656 8230
rect 42708 7268 42760 7274
rect 42708 7210 42760 7216
rect 42720 6662 42748 7210
rect 42708 6656 42760 6662
rect 42614 6624 42670 6633
rect 42708 6598 42760 6604
rect 42614 6559 42670 6568
rect 42812 6322 42840 8486
rect 42892 8492 42944 8498
rect 42892 8434 42944 8440
rect 42904 8090 42932 8434
rect 42892 8084 42944 8090
rect 42892 8026 42944 8032
rect 42982 7984 43038 7993
rect 42982 7919 42984 7928
rect 43036 7919 43038 7928
rect 42984 7890 43036 7896
rect 42984 7200 43036 7206
rect 42984 7142 43036 7148
rect 42800 6316 42852 6322
rect 42800 6258 42852 6264
rect 42892 5636 42944 5642
rect 42892 5578 42944 5584
rect 42904 5166 42932 5578
rect 42892 5160 42944 5166
rect 42892 5102 42944 5108
rect 42432 5092 42484 5098
rect 42432 5034 42484 5040
rect 42156 4820 42208 4826
rect 42156 4762 42208 4768
rect 42904 4758 42932 5102
rect 42892 4752 42944 4758
rect 42892 4694 42944 4700
rect 42064 4548 42116 4554
rect 42064 4490 42116 4496
rect 41788 4140 41840 4146
rect 41788 4082 41840 4088
rect 41800 3670 41828 4082
rect 41788 3664 41840 3670
rect 41788 3606 41840 3612
rect 41880 3460 41932 3466
rect 41880 3402 41932 3408
rect 41892 3369 41920 3402
rect 41878 3360 41934 3369
rect 41878 3295 41934 3304
rect 41328 3188 41380 3194
rect 41328 3130 41380 3136
rect 41696 3188 41748 3194
rect 41696 3130 41748 3136
rect 41512 3052 41564 3058
rect 41512 2994 41564 3000
rect 41418 2680 41474 2689
rect 41418 2615 41420 2624
rect 41472 2615 41474 2624
rect 41420 2586 41472 2592
rect 41420 2440 41472 2446
rect 41420 2382 41472 2388
rect 41432 814 41460 2382
rect 41420 808 41472 814
rect 5906 0 5962 800
rect 6182 0 6238 800
rect 6458 0 6514 800
rect 6734 0 6790 800
rect 7010 0 7066 800
rect 7286 0 7342 800
rect 7562 0 7618 800
rect 7838 0 7894 800
rect 8114 0 8170 800
rect 8390 0 8446 800
rect 8666 0 8722 800
rect 8942 0 8998 800
rect 9218 0 9274 800
rect 9494 0 9550 800
rect 9770 0 9826 800
rect 10046 0 10102 800
rect 10322 0 10378 800
rect 10598 0 10654 800
rect 10874 0 10930 800
rect 11150 0 11206 800
rect 11426 0 11482 800
rect 11702 0 11758 800
rect 11978 0 12034 800
rect 12254 0 12310 800
rect 12530 0 12586 800
rect 12806 0 12862 800
rect 13082 0 13138 800
rect 13358 0 13414 800
rect 13634 0 13690 800
rect 13910 0 13966 800
rect 14186 0 14242 800
rect 14462 0 14518 800
rect 14738 0 14794 800
rect 15014 0 15070 800
rect 15290 0 15346 800
rect 15566 0 15622 800
rect 15842 0 15898 800
rect 16118 0 16174 800
rect 16394 0 16450 800
rect 16670 0 16726 800
rect 16946 0 17002 800
rect 17222 0 17278 800
rect 17498 0 17554 800
rect 17774 0 17830 800
rect 18050 0 18106 800
rect 18326 0 18382 800
rect 18602 0 18658 800
rect 18878 0 18934 800
rect 19154 0 19210 800
rect 19430 0 19486 800
rect 19706 0 19762 800
rect 19982 0 20038 800
rect 20258 0 20314 800
rect 20534 0 20590 800
rect 20810 0 20866 800
rect 21086 0 21142 800
rect 21362 0 21418 800
rect 21638 0 21694 800
rect 21914 0 21970 800
rect 22190 0 22246 800
rect 22466 0 22522 800
rect 22742 0 22798 800
rect 23018 0 23074 800
rect 23294 0 23350 800
rect 23570 0 23626 800
rect 23846 0 23902 800
rect 24122 0 24178 800
rect 24398 0 24454 800
rect 24674 0 24730 800
rect 24950 0 25006 800
rect 25226 0 25282 800
rect 25502 0 25558 800
rect 25778 0 25834 800
rect 26054 0 26110 800
rect 26330 0 26386 800
rect 26606 0 26662 800
rect 26882 0 26938 800
rect 27158 0 27214 800
rect 27434 0 27490 800
rect 27710 0 27766 800
rect 27986 0 28042 800
rect 28262 0 28318 800
rect 28538 0 28594 800
rect 28814 0 28870 800
rect 29090 0 29146 800
rect 29366 0 29422 800
rect 29642 0 29698 800
rect 29918 0 29974 800
rect 30194 0 30250 800
rect 30470 0 30526 800
rect 30746 0 30802 800
rect 31022 0 31078 800
rect 31298 0 31354 800
rect 31574 0 31630 800
rect 31850 0 31906 800
rect 32126 0 32182 800
rect 32402 0 32458 800
rect 32678 0 32734 800
rect 32954 0 33010 800
rect 33230 0 33286 800
rect 33506 0 33562 800
rect 33782 0 33838 800
rect 34058 0 34114 800
rect 34334 0 34390 800
rect 34610 0 34666 800
rect 34886 0 34942 800
rect 35162 0 35218 800
rect 35438 0 35494 800
rect 35714 0 35770 800
rect 35990 0 36046 800
rect 36266 0 36322 800
rect 36542 0 36598 800
rect 36818 0 36874 800
rect 37094 0 37150 800
rect 37370 0 37426 800
rect 37646 0 37702 800
rect 37922 0 37978 800
rect 38198 0 38254 800
rect 38474 0 38530 800
rect 38750 0 38806 800
rect 39026 0 39082 800
rect 39302 0 39358 800
rect 39578 0 39634 800
rect 39854 0 39910 800
rect 40130 0 40186 800
rect 40406 0 40462 800
rect 40682 0 40738 800
rect 40958 0 41014 800
rect 41234 0 41290 800
rect 41524 800 41552 2994
rect 41788 2372 41840 2378
rect 41788 2314 41840 2320
rect 41800 800 41828 2314
rect 42076 800 42104 4490
rect 42892 4480 42944 4486
rect 42892 4422 42944 4428
rect 42708 4140 42760 4146
rect 42708 4082 42760 4088
rect 42616 4072 42668 4078
rect 42616 4014 42668 4020
rect 42628 2774 42656 4014
rect 42720 3738 42748 4082
rect 42708 3732 42760 3738
rect 42708 3674 42760 3680
rect 42904 3534 42932 4422
rect 42996 4146 43024 7142
rect 42984 4140 43036 4146
rect 42984 4082 43036 4088
rect 42984 3732 43036 3738
rect 42984 3674 43036 3680
rect 42996 3534 43024 3674
rect 43088 3534 43116 9687
rect 43180 5710 43208 12406
rect 43260 9036 43312 9042
rect 43260 8978 43312 8984
rect 43272 7954 43300 8978
rect 43536 8288 43588 8294
rect 43456 8236 43536 8242
rect 43456 8230 43588 8236
rect 43456 8214 43576 8230
rect 43260 7948 43312 7954
rect 43260 7890 43312 7896
rect 43456 7750 43484 8214
rect 43640 7886 43668 20878
rect 43732 19718 43760 22066
rect 43824 20777 43852 22918
rect 43916 20942 43944 30806
rect 44272 22772 44324 22778
rect 44272 22714 44324 22720
rect 44364 22772 44416 22778
rect 44364 22714 44416 22720
rect 44180 22636 44232 22642
rect 44180 22578 44232 22584
rect 44088 22568 44140 22574
rect 44088 22510 44140 22516
rect 44100 22030 44128 22510
rect 44088 22024 44140 22030
rect 44088 21966 44140 21972
rect 44100 21622 44128 21966
rect 44088 21616 44140 21622
rect 44088 21558 44140 21564
rect 44192 21146 44220 22578
rect 44180 21140 44232 21146
rect 44180 21082 44232 21088
rect 44284 20942 44312 22714
rect 44376 22681 44404 22714
rect 44362 22672 44418 22681
rect 44362 22607 44418 22616
rect 44376 21962 44404 22607
rect 44640 22024 44692 22030
rect 44640 21966 44692 21972
rect 44364 21956 44416 21962
rect 44364 21898 44416 21904
rect 44548 21888 44600 21894
rect 44548 21830 44600 21836
rect 44560 21010 44588 21830
rect 44548 21004 44600 21010
rect 44548 20946 44600 20952
rect 43904 20936 43956 20942
rect 43904 20878 43956 20884
rect 43996 20936 44048 20942
rect 44272 20936 44324 20942
rect 43996 20878 44048 20884
rect 44192 20896 44272 20924
rect 43810 20768 43866 20777
rect 43810 20703 43866 20712
rect 44008 19922 44036 20878
rect 44192 20058 44220 20896
rect 44272 20878 44324 20884
rect 44546 20632 44602 20641
rect 44546 20567 44602 20576
rect 44560 20398 44588 20567
rect 44652 20534 44680 21966
rect 44640 20528 44692 20534
rect 44640 20470 44692 20476
rect 44548 20392 44600 20398
rect 44548 20334 44600 20340
rect 44364 20324 44416 20330
rect 44364 20266 44416 20272
rect 44180 20052 44232 20058
rect 44180 19994 44232 20000
rect 43996 19916 44048 19922
rect 43996 19858 44048 19864
rect 44192 19854 44220 19994
rect 44376 19990 44404 20266
rect 44560 20262 44588 20334
rect 44548 20256 44600 20262
rect 44548 20198 44600 20204
rect 44548 20052 44600 20058
rect 44548 19994 44600 20000
rect 44364 19984 44416 19990
rect 44270 19952 44326 19961
rect 44364 19926 44416 19932
rect 44270 19887 44326 19896
rect 44284 19854 44312 19887
rect 44560 19854 44588 19994
rect 44180 19848 44232 19854
rect 44180 19790 44232 19796
rect 44272 19848 44324 19854
rect 44456 19848 44508 19854
rect 44272 19790 44324 19796
rect 44362 19816 44418 19825
rect 43720 19712 43772 19718
rect 43720 19654 43772 19660
rect 43994 19544 44050 19553
rect 43994 19479 44050 19488
rect 44008 19446 44036 19479
rect 43996 19440 44048 19446
rect 43996 19382 44048 19388
rect 43996 18284 44048 18290
rect 43996 18226 44048 18232
rect 43904 18216 43956 18222
rect 43904 18158 43956 18164
rect 43720 17876 43772 17882
rect 43720 17818 43772 17824
rect 43732 17202 43760 17818
rect 43916 17814 43944 18158
rect 43904 17808 43956 17814
rect 43904 17750 43956 17756
rect 43720 17196 43772 17202
rect 43720 17138 43772 17144
rect 43904 13728 43956 13734
rect 43904 13670 43956 13676
rect 43916 12714 43944 13670
rect 43904 12708 43956 12714
rect 43904 12650 43956 12656
rect 43916 12434 43944 12650
rect 43824 12406 43944 12434
rect 43718 11792 43774 11801
rect 43718 11727 43774 11736
rect 43628 7880 43680 7886
rect 43628 7822 43680 7828
rect 43444 7744 43496 7750
rect 43444 7686 43496 7692
rect 43456 7478 43484 7686
rect 43444 7472 43496 7478
rect 43444 7414 43496 7420
rect 43350 6760 43406 6769
rect 43350 6695 43406 6704
rect 43260 6656 43312 6662
rect 43260 6598 43312 6604
rect 43168 5704 43220 5710
rect 43168 5646 43220 5652
rect 43180 4826 43208 5646
rect 43272 5234 43300 6598
rect 43364 6390 43392 6695
rect 43352 6384 43404 6390
rect 43352 6326 43404 6332
rect 43444 6316 43496 6322
rect 43444 6258 43496 6264
rect 43350 5672 43406 5681
rect 43350 5607 43406 5616
rect 43364 5574 43392 5607
rect 43352 5568 43404 5574
rect 43352 5510 43404 5516
rect 43260 5228 43312 5234
rect 43260 5170 43312 5176
rect 43168 4820 43220 4826
rect 43168 4762 43220 4768
rect 43364 4622 43392 5510
rect 43456 5302 43484 6258
rect 43732 5658 43760 11727
rect 43824 5846 43852 12406
rect 44008 11778 44036 18226
rect 44192 17882 44220 19790
rect 44456 19790 44508 19796
rect 44548 19848 44600 19854
rect 44548 19790 44600 19796
rect 44362 19751 44418 19760
rect 44376 19310 44404 19751
rect 44468 19514 44496 19790
rect 44456 19508 44508 19514
rect 44456 19450 44508 19456
rect 44652 19378 44680 20470
rect 44732 20256 44784 20262
rect 44732 20198 44784 20204
rect 44456 19372 44508 19378
rect 44456 19314 44508 19320
rect 44640 19372 44692 19378
rect 44640 19314 44692 19320
rect 44364 19304 44416 19310
rect 44364 19246 44416 19252
rect 44272 19168 44324 19174
rect 44272 19110 44324 19116
rect 44180 17876 44232 17882
rect 44180 17818 44232 17824
rect 44180 17740 44232 17746
rect 44180 17682 44232 17688
rect 44088 17672 44140 17678
rect 44088 17614 44140 17620
rect 44100 17202 44128 17614
rect 44192 17241 44220 17682
rect 44178 17232 44234 17241
rect 44088 17196 44140 17202
rect 44178 17167 44234 17176
rect 44088 17138 44140 17144
rect 44180 17128 44232 17134
rect 44180 17070 44232 17076
rect 44192 16794 44220 17070
rect 44180 16788 44232 16794
rect 44180 16730 44232 16736
rect 44284 16590 44312 19110
rect 44364 17876 44416 17882
rect 44364 17818 44416 17824
rect 44376 16590 44404 17818
rect 44468 17678 44496 19314
rect 44456 17672 44508 17678
rect 44456 17614 44508 17620
rect 44548 16788 44600 16794
rect 44548 16730 44600 16736
rect 44456 16720 44508 16726
rect 44456 16662 44508 16668
rect 44468 16590 44496 16662
rect 44272 16584 44324 16590
rect 44272 16526 44324 16532
rect 44364 16584 44416 16590
rect 44364 16526 44416 16532
rect 44456 16584 44508 16590
rect 44560 16574 44588 16730
rect 44652 16726 44680 19314
rect 44744 18358 44772 20198
rect 44822 19952 44878 19961
rect 44822 19887 44878 19896
rect 44732 18352 44784 18358
rect 44732 18294 44784 18300
rect 44640 16720 44692 16726
rect 44640 16662 44692 16668
rect 44732 16584 44784 16590
rect 44560 16546 44680 16574
rect 44456 16526 44508 16532
rect 44180 16108 44232 16114
rect 44180 16050 44232 16056
rect 44088 15972 44140 15978
rect 44088 15914 44140 15920
rect 44100 14958 44128 15914
rect 44088 14952 44140 14958
rect 44088 14894 44140 14900
rect 44100 12306 44128 14894
rect 44192 13190 44220 16050
rect 44180 13184 44232 13190
rect 44180 13126 44232 13132
rect 44088 12300 44140 12306
rect 44088 12242 44140 12248
rect 44284 12238 44312 16526
rect 44376 16182 44404 16526
rect 44364 16176 44416 16182
rect 44364 16118 44416 16124
rect 44364 15360 44416 15366
rect 44364 15302 44416 15308
rect 44456 15360 44508 15366
rect 44456 15302 44508 15308
rect 44376 15026 44404 15302
rect 44468 15094 44496 15302
rect 44456 15088 44508 15094
rect 44456 15030 44508 15036
rect 44364 15020 44416 15026
rect 44364 14962 44416 14968
rect 44272 12232 44324 12238
rect 44272 12174 44324 12180
rect 44008 11750 44220 11778
rect 44088 11688 44140 11694
rect 44088 11630 44140 11636
rect 43996 11212 44048 11218
rect 43996 11154 44048 11160
rect 43904 9512 43956 9518
rect 43904 9454 43956 9460
rect 43916 8974 43944 9454
rect 43904 8968 43956 8974
rect 43904 8910 43956 8916
rect 43904 6860 43956 6866
rect 43904 6802 43956 6808
rect 43916 6186 43944 6802
rect 44008 6730 44036 11154
rect 44100 10606 44128 11630
rect 44088 10600 44140 10606
rect 44088 10542 44140 10548
rect 43996 6724 44048 6730
rect 43996 6666 44048 6672
rect 44008 6361 44036 6666
rect 43994 6352 44050 6361
rect 43994 6287 44050 6296
rect 43904 6180 43956 6186
rect 43904 6122 43956 6128
rect 44088 6112 44140 6118
rect 44088 6054 44140 6060
rect 43812 5840 43864 5846
rect 43812 5782 43864 5788
rect 43732 5630 43852 5658
rect 44100 5642 44128 6054
rect 43444 5296 43496 5302
rect 43444 5238 43496 5244
rect 43352 4616 43404 4622
rect 43352 4558 43404 4564
rect 43352 4140 43404 4146
rect 43352 4082 43404 4088
rect 43168 3936 43220 3942
rect 43168 3878 43220 3884
rect 42800 3528 42852 3534
rect 42706 3496 42762 3505
rect 42800 3470 42852 3476
rect 42892 3528 42944 3534
rect 42892 3470 42944 3476
rect 42984 3528 43036 3534
rect 42984 3470 43036 3476
rect 43076 3528 43128 3534
rect 43076 3470 43128 3476
rect 42706 3431 42762 3440
rect 42720 3058 42748 3431
rect 42812 3126 42840 3470
rect 42996 3398 43024 3470
rect 42984 3392 43036 3398
rect 42984 3334 43036 3340
rect 42800 3120 42852 3126
rect 42800 3062 42852 3068
rect 42708 3052 42760 3058
rect 42708 2994 42760 3000
rect 42892 2848 42944 2854
rect 42892 2790 42944 2796
rect 42628 2746 42748 2774
rect 42720 2122 42748 2746
rect 42628 2094 42748 2122
rect 42340 1012 42392 1018
rect 42340 954 42392 960
rect 42352 800 42380 954
rect 42628 800 42656 2094
rect 42904 800 42932 2790
rect 43180 800 43208 3878
rect 43260 3052 43312 3058
rect 43260 2994 43312 3000
rect 43272 1086 43300 2994
rect 43364 1222 43392 4082
rect 43534 4040 43590 4049
rect 43534 3975 43536 3984
rect 43588 3975 43590 3984
rect 43536 3946 43588 3952
rect 43444 3596 43496 3602
rect 43444 3538 43496 3544
rect 43352 1216 43404 1222
rect 43352 1158 43404 1164
rect 43260 1080 43312 1086
rect 43260 1022 43312 1028
rect 43456 800 43484 3538
rect 43720 3528 43772 3534
rect 43720 3470 43772 3476
rect 43628 3392 43680 3398
rect 43628 3334 43680 3340
rect 43640 3233 43668 3334
rect 43626 3224 43682 3233
rect 43626 3159 43682 3168
rect 43732 2922 43760 3470
rect 43720 2916 43772 2922
rect 43720 2858 43772 2864
rect 43824 2650 43852 5630
rect 44088 5636 44140 5642
rect 44088 5578 44140 5584
rect 44192 3738 44220 11750
rect 44456 11008 44508 11014
rect 44456 10950 44508 10956
rect 44364 8968 44416 8974
rect 44364 8910 44416 8916
rect 44272 7404 44324 7410
rect 44272 7346 44324 7352
rect 44284 6798 44312 7346
rect 44272 6792 44324 6798
rect 44272 6734 44324 6740
rect 44284 6458 44312 6734
rect 44272 6452 44324 6458
rect 44272 6394 44324 6400
rect 44376 6322 44404 8910
rect 44468 7342 44496 10950
rect 44548 10600 44600 10606
rect 44548 10542 44600 10548
rect 44560 10062 44588 10542
rect 44548 10056 44600 10062
rect 44548 9998 44600 10004
rect 44652 9654 44680 16546
rect 44732 16526 44784 16532
rect 44744 15910 44772 16526
rect 44732 15904 44784 15910
rect 44732 15846 44784 15852
rect 44744 15094 44772 15846
rect 44836 15162 44864 19887
rect 44916 19712 44968 19718
rect 44916 19654 44968 19660
rect 44928 19446 44956 19654
rect 44916 19440 44968 19446
rect 44916 19382 44968 19388
rect 45020 19334 45048 35974
rect 45388 25974 45416 57190
rect 46308 36038 46336 57190
rect 46296 36032 46348 36038
rect 46296 35974 46348 35980
rect 46020 33924 46072 33930
rect 46020 33866 46072 33872
rect 45560 31136 45612 31142
rect 45560 31078 45612 31084
rect 45572 30122 45600 31078
rect 45560 30116 45612 30122
rect 45560 30058 45612 30064
rect 45468 27600 45520 27606
rect 45468 27542 45520 27548
rect 45480 26790 45508 27542
rect 45468 26784 45520 26790
rect 45468 26726 45520 26732
rect 45376 25968 45428 25974
rect 45376 25910 45428 25916
rect 45100 25424 45152 25430
rect 45100 25366 45152 25372
rect 44928 19306 45048 19334
rect 44928 18290 44956 19306
rect 45008 18896 45060 18902
rect 45008 18838 45060 18844
rect 45020 18426 45048 18838
rect 45008 18420 45060 18426
rect 45008 18362 45060 18368
rect 44916 18284 44968 18290
rect 44916 18226 44968 18232
rect 45112 18222 45140 25366
rect 45928 25288 45980 25294
rect 45926 25256 45928 25265
rect 45980 25256 45982 25265
rect 45926 25191 45982 25200
rect 45192 24268 45244 24274
rect 45192 24210 45244 24216
rect 45100 18216 45152 18222
rect 45100 18158 45152 18164
rect 45204 18034 45232 24210
rect 45744 23316 45796 23322
rect 45744 23258 45796 23264
rect 45560 22432 45612 22438
rect 45560 22374 45612 22380
rect 45284 21956 45336 21962
rect 45284 21898 45336 21904
rect 45296 21146 45324 21898
rect 45284 21140 45336 21146
rect 45284 21082 45336 21088
rect 45572 20942 45600 22374
rect 45652 21412 45704 21418
rect 45652 21354 45704 21360
rect 45664 20942 45692 21354
rect 45560 20936 45612 20942
rect 45560 20878 45612 20884
rect 45652 20936 45704 20942
rect 45652 20878 45704 20884
rect 45376 20392 45428 20398
rect 45376 20334 45428 20340
rect 45388 18426 45416 20334
rect 45572 19854 45600 20878
rect 45560 19848 45612 19854
rect 45756 19825 45784 23258
rect 46032 21486 46060 33866
rect 46400 25294 46428 57190
rect 48884 56681 48912 57190
rect 48870 56672 48926 56681
rect 48870 56607 48926 56616
rect 47860 53440 47912 53446
rect 47860 53382 47912 53388
rect 47674 52728 47730 52737
rect 47674 52663 47676 52672
rect 47728 52663 47730 52672
rect 47676 52634 47728 52640
rect 47872 52494 47900 53382
rect 48136 53032 48188 53038
rect 48136 52974 48188 52980
rect 48504 53032 48556 53038
rect 48504 52974 48556 52980
rect 48044 52896 48096 52902
rect 48044 52838 48096 52844
rect 48056 52601 48084 52838
rect 48042 52592 48098 52601
rect 48042 52527 48098 52536
rect 48148 52494 48176 52974
rect 48516 52494 48544 52974
rect 47860 52488 47912 52494
rect 47860 52430 47912 52436
rect 48136 52488 48188 52494
rect 48136 52430 48188 52436
rect 48504 52488 48556 52494
rect 48504 52430 48556 52436
rect 48148 51950 48176 52430
rect 48516 51950 48544 52430
rect 47768 51944 47820 51950
rect 47768 51886 47820 51892
rect 48136 51944 48188 51950
rect 48136 51886 48188 51892
rect 48504 51944 48556 51950
rect 48504 51886 48556 51892
rect 46848 51808 46900 51814
rect 46848 51750 46900 51756
rect 46860 51406 46888 51750
rect 46848 51400 46900 51406
rect 46848 51342 46900 51348
rect 47032 51332 47084 51338
rect 47032 51274 47084 51280
rect 47492 51332 47544 51338
rect 47492 51274 47544 51280
rect 47044 50998 47072 51274
rect 47032 50992 47084 50998
rect 47032 50934 47084 50940
rect 47044 49910 47072 50934
rect 47308 50856 47360 50862
rect 47308 50798 47360 50804
rect 47032 49904 47084 49910
rect 47032 49846 47084 49852
rect 47216 44872 47268 44878
rect 47216 44814 47268 44820
rect 47228 43722 47256 44814
rect 47216 43716 47268 43722
rect 47216 43658 47268 43664
rect 46480 32564 46532 32570
rect 46480 32506 46532 32512
rect 46204 25288 46256 25294
rect 46204 25230 46256 25236
rect 46388 25288 46440 25294
rect 46388 25230 46440 25236
rect 46020 21480 46072 21486
rect 46018 21448 46020 21457
rect 46072 21448 46074 21457
rect 46018 21383 46074 21392
rect 45836 21072 45888 21078
rect 45836 21014 45888 21020
rect 45560 19790 45612 19796
rect 45742 19816 45798 19825
rect 45376 18420 45428 18426
rect 45376 18362 45428 18368
rect 45468 18216 45520 18222
rect 45468 18158 45520 18164
rect 45112 18006 45232 18034
rect 44824 15156 44876 15162
rect 44824 15098 44876 15104
rect 44916 15156 44968 15162
rect 44916 15098 44968 15104
rect 44732 15088 44784 15094
rect 44732 15030 44784 15036
rect 44928 14618 44956 15098
rect 44916 14612 44968 14618
rect 44916 14554 44968 14560
rect 44916 14000 44968 14006
rect 44916 13942 44968 13948
rect 44928 12434 44956 13942
rect 44744 12406 44956 12434
rect 44640 9648 44692 9654
rect 44640 9590 44692 9596
rect 44638 8392 44694 8401
rect 44638 8327 44694 8336
rect 44456 7336 44508 7342
rect 44456 7278 44508 7284
rect 44456 6792 44508 6798
rect 44456 6734 44508 6740
rect 44364 6316 44416 6322
rect 44364 6258 44416 6264
rect 44468 5302 44496 6734
rect 44548 6656 44600 6662
rect 44548 6598 44600 6604
rect 44560 5710 44588 6598
rect 44548 5704 44600 5710
rect 44548 5646 44600 5652
rect 44456 5296 44508 5302
rect 44456 5238 44508 5244
rect 44548 5228 44600 5234
rect 44548 5170 44600 5176
rect 44364 4208 44416 4214
rect 44364 4150 44416 4156
rect 44270 4040 44326 4049
rect 44270 3975 44272 3984
rect 44324 3975 44326 3984
rect 44272 3946 44324 3952
rect 44088 3732 44140 3738
rect 44088 3674 44140 3680
rect 44180 3732 44232 3738
rect 44180 3674 44232 3680
rect 44100 3618 44128 3674
rect 44100 3590 44220 3618
rect 44192 3534 44220 3590
rect 43904 3528 43956 3534
rect 44180 3528 44232 3534
rect 43956 3488 44128 3516
rect 43904 3470 43956 3476
rect 44100 3398 44128 3488
rect 44180 3470 44232 3476
rect 44088 3392 44140 3398
rect 44088 3334 44140 3340
rect 43904 3188 43956 3194
rect 43904 3130 43956 3136
rect 43916 3097 43944 3130
rect 43902 3088 43958 3097
rect 43902 3023 43958 3032
rect 44088 3052 44140 3058
rect 44088 2994 44140 3000
rect 43812 2644 43864 2650
rect 43812 2586 43864 2592
rect 43812 2372 43864 2378
rect 43812 2314 43864 2320
rect 43720 1080 43772 1086
rect 43720 1022 43772 1028
rect 43732 800 43760 1022
rect 43824 882 43852 2314
rect 44100 1154 44128 2994
rect 44192 2990 44220 3470
rect 44180 2984 44232 2990
rect 44180 2926 44232 2932
rect 44376 2122 44404 4150
rect 44456 3460 44508 3466
rect 44456 3402 44508 3408
rect 44468 3233 44496 3402
rect 44454 3224 44510 3233
rect 44454 3159 44510 3168
rect 44560 2774 44588 5170
rect 44652 4282 44680 8327
rect 44640 4276 44692 4282
rect 44640 4218 44692 4224
rect 44638 3224 44694 3233
rect 44638 3159 44640 3168
rect 44692 3159 44694 3168
rect 44640 3130 44692 3136
rect 44744 2774 44772 12406
rect 44824 10464 44876 10470
rect 44824 10406 44876 10412
rect 44836 9110 44864 10406
rect 44824 9104 44876 9110
rect 44824 9046 44876 9052
rect 45112 8430 45140 18006
rect 45480 17746 45508 18158
rect 45572 17882 45600 19790
rect 45742 19751 45798 19760
rect 45560 17876 45612 17882
rect 45560 17818 45612 17824
rect 45468 17740 45520 17746
rect 45468 17682 45520 17688
rect 45652 17672 45704 17678
rect 45652 17614 45704 17620
rect 45284 17604 45336 17610
rect 45284 17546 45336 17552
rect 45296 17134 45324 17546
rect 45664 17270 45692 17614
rect 45756 17270 45784 19751
rect 45652 17264 45704 17270
rect 45652 17206 45704 17212
rect 45744 17264 45796 17270
rect 45744 17206 45796 17212
rect 45284 17128 45336 17134
rect 45284 17070 45336 17076
rect 45652 17128 45704 17134
rect 45848 17116 45876 21014
rect 45928 20460 45980 20466
rect 45928 20402 45980 20408
rect 45940 18970 45968 20402
rect 46020 19508 46072 19514
rect 46020 19450 46072 19456
rect 46032 19174 46060 19450
rect 46020 19168 46072 19174
rect 46020 19110 46072 19116
rect 45928 18964 45980 18970
rect 45928 18906 45980 18912
rect 46032 18766 46060 19110
rect 46020 18760 46072 18766
rect 46020 18702 46072 18708
rect 46032 18630 46060 18702
rect 46020 18624 46072 18630
rect 46020 18566 46072 18572
rect 46112 17332 46164 17338
rect 46112 17274 46164 17280
rect 45928 17264 45980 17270
rect 45928 17206 45980 17212
rect 45652 17070 45704 17076
rect 45756 17088 45876 17116
rect 45560 17060 45612 17066
rect 45560 17002 45612 17008
rect 45192 16652 45244 16658
rect 45192 16594 45244 16600
rect 45204 16182 45232 16594
rect 45192 16176 45244 16182
rect 45192 16118 45244 16124
rect 45204 15570 45232 16118
rect 45192 15564 45244 15570
rect 45192 15506 45244 15512
rect 45284 14476 45336 14482
rect 45284 14418 45336 14424
rect 45192 11756 45244 11762
rect 45192 11698 45244 11704
rect 45204 11354 45232 11698
rect 45192 11348 45244 11354
rect 45192 11290 45244 11296
rect 45192 9172 45244 9178
rect 45192 9114 45244 9120
rect 45100 8424 45152 8430
rect 45100 8366 45152 8372
rect 44824 7880 44876 7886
rect 44824 7822 44876 7828
rect 44836 7546 44864 7822
rect 44824 7540 44876 7546
rect 44824 7482 44876 7488
rect 45204 7410 45232 9114
rect 45192 7404 45244 7410
rect 45192 7346 45244 7352
rect 44824 7336 44876 7342
rect 44824 7278 44876 7284
rect 45008 7336 45060 7342
rect 45060 7284 45140 7290
rect 45008 7278 45140 7284
rect 44836 5234 44864 7278
rect 45020 7262 45140 7278
rect 44914 6896 44970 6905
rect 44914 6831 44970 6840
rect 44928 6798 44956 6831
rect 44916 6792 44968 6798
rect 44916 6734 44968 6740
rect 45008 6724 45060 6730
rect 45008 6666 45060 6672
rect 45020 5794 45048 6666
rect 45112 6322 45140 7262
rect 45204 6458 45232 7346
rect 45192 6452 45244 6458
rect 45192 6394 45244 6400
rect 45100 6316 45152 6322
rect 45100 6258 45152 6264
rect 45192 6316 45244 6322
rect 45192 6258 45244 6264
rect 45112 5914 45140 6258
rect 45100 5908 45152 5914
rect 45100 5850 45152 5856
rect 45204 5794 45232 6258
rect 45020 5766 45232 5794
rect 45204 5642 45232 5766
rect 45192 5636 45244 5642
rect 45192 5578 45244 5584
rect 44824 5228 44876 5234
rect 45296 5216 45324 14418
rect 45468 11552 45520 11558
rect 45468 11494 45520 11500
rect 45480 11150 45508 11494
rect 45468 11144 45520 11150
rect 45468 11086 45520 11092
rect 45468 9988 45520 9994
rect 45468 9930 45520 9936
rect 45480 9722 45508 9930
rect 45468 9716 45520 9722
rect 45468 9658 45520 9664
rect 45376 6656 45428 6662
rect 45376 6598 45428 6604
rect 45388 6497 45416 6598
rect 45374 6488 45430 6497
rect 45374 6423 45430 6432
rect 45468 6452 45520 6458
rect 45468 6394 45520 6400
rect 45480 6338 45508 6394
rect 45388 6310 45508 6338
rect 45388 5234 45416 6310
rect 45468 6248 45520 6254
rect 45468 6190 45520 6196
rect 44824 5170 44876 5176
rect 45020 5188 45324 5216
rect 45376 5228 45428 5234
rect 45020 4978 45048 5188
rect 45376 5170 45428 5176
rect 45480 5166 45508 6190
rect 45572 5914 45600 17002
rect 45664 6458 45692 17070
rect 45756 11082 45784 17088
rect 45940 15026 45968 17206
rect 46124 16574 46152 17274
rect 46032 16546 46152 16574
rect 45928 15020 45980 15026
rect 45928 14962 45980 14968
rect 45836 12776 45888 12782
rect 45836 12718 45888 12724
rect 45848 11218 45876 12718
rect 46032 12434 46060 16546
rect 46032 12406 46152 12434
rect 45836 11212 45888 11218
rect 45836 11154 45888 11160
rect 45744 11076 45796 11082
rect 45744 11018 45796 11024
rect 45836 10260 45888 10266
rect 45836 10202 45888 10208
rect 45848 9518 45876 10202
rect 45836 9512 45888 9518
rect 45836 9454 45888 9460
rect 46124 8838 46152 12406
rect 46216 9058 46244 25230
rect 46296 25220 46348 25226
rect 46296 25162 46348 25168
rect 46308 24954 46336 25162
rect 46296 24948 46348 24954
rect 46296 24890 46348 24896
rect 46492 21434 46520 32506
rect 46572 30728 46624 30734
rect 46572 30670 46624 30676
rect 46584 22574 46612 30670
rect 47216 26920 47268 26926
rect 47216 26862 47268 26868
rect 47124 25832 47176 25838
rect 47124 25774 47176 25780
rect 46756 25696 46808 25702
rect 46756 25638 46808 25644
rect 46664 22772 46716 22778
rect 46664 22714 46716 22720
rect 46572 22568 46624 22574
rect 46572 22510 46624 22516
rect 46572 21888 46624 21894
rect 46572 21830 46624 21836
rect 46584 21622 46612 21830
rect 46572 21616 46624 21622
rect 46572 21558 46624 21564
rect 46308 21406 46520 21434
rect 46308 11286 46336 21406
rect 46480 18080 46532 18086
rect 46480 18022 46532 18028
rect 46388 15904 46440 15910
rect 46388 15846 46440 15852
rect 46400 15502 46428 15846
rect 46388 15496 46440 15502
rect 46388 15438 46440 15444
rect 46492 12434 46520 18022
rect 46572 16448 46624 16454
rect 46572 16390 46624 16396
rect 46584 16046 46612 16390
rect 46572 16040 46624 16046
rect 46572 15982 46624 15988
rect 46572 15904 46624 15910
rect 46572 15846 46624 15852
rect 46584 15434 46612 15846
rect 46572 15428 46624 15434
rect 46572 15370 46624 15376
rect 46676 14006 46704 22714
rect 46768 21078 46796 25638
rect 47136 25294 47164 25774
rect 47124 25288 47176 25294
rect 46938 25256 46994 25265
rect 47122 25256 47124 25265
rect 47176 25256 47178 25265
rect 46938 25191 46994 25200
rect 47032 25220 47084 25226
rect 46952 24206 46980 25191
rect 47122 25191 47178 25200
rect 47032 25162 47084 25168
rect 46940 24200 46992 24206
rect 46940 24142 46992 24148
rect 46848 22568 46900 22574
rect 46848 22510 46900 22516
rect 46756 21072 46808 21078
rect 46756 21014 46808 21020
rect 46860 20369 46888 22510
rect 46940 21480 46992 21486
rect 46940 21422 46992 21428
rect 46846 20360 46902 20369
rect 46768 20318 46846 20346
rect 46768 18834 46796 20318
rect 46846 20295 46902 20304
rect 46846 19680 46902 19689
rect 46846 19615 46902 19624
rect 46860 19446 46888 19615
rect 46848 19440 46900 19446
rect 46848 19382 46900 19388
rect 46756 18828 46808 18834
rect 46756 18770 46808 18776
rect 46952 18698 46980 21422
rect 46940 18692 46992 18698
rect 46940 18634 46992 18640
rect 46952 18426 46980 18634
rect 46940 18420 46992 18426
rect 46940 18362 46992 18368
rect 46952 18222 46980 18362
rect 46940 18216 46992 18222
rect 46940 18158 46992 18164
rect 46754 16144 46810 16153
rect 46754 16079 46756 16088
rect 46808 16079 46810 16088
rect 46756 16050 46808 16056
rect 46848 16040 46900 16046
rect 46848 15982 46900 15988
rect 46860 15638 46888 15982
rect 46848 15632 46900 15638
rect 46846 15600 46848 15609
rect 46900 15600 46902 15609
rect 46846 15535 46902 15544
rect 46848 15360 46900 15366
rect 46848 15302 46900 15308
rect 46860 14346 46888 15302
rect 46848 14340 46900 14346
rect 46848 14282 46900 14288
rect 46664 14000 46716 14006
rect 46664 13942 46716 13948
rect 46940 12844 46992 12850
rect 46940 12786 46992 12792
rect 46400 12406 46520 12434
rect 46296 11280 46348 11286
rect 46296 11222 46348 11228
rect 46216 9030 46336 9058
rect 46204 8900 46256 8906
rect 46204 8842 46256 8848
rect 46112 8832 46164 8838
rect 46112 8774 46164 8780
rect 46020 7404 46072 7410
rect 46020 7346 46072 7352
rect 46032 6934 46060 7346
rect 46020 6928 46072 6934
rect 45834 6896 45890 6905
rect 46020 6870 46072 6876
rect 45834 6831 45890 6840
rect 45744 6792 45796 6798
rect 45744 6734 45796 6740
rect 45652 6452 45704 6458
rect 45652 6394 45704 6400
rect 45756 6390 45784 6734
rect 45848 6662 45876 6831
rect 45836 6656 45888 6662
rect 45836 6598 45888 6604
rect 45744 6384 45796 6390
rect 45744 6326 45796 6332
rect 45560 5908 45612 5914
rect 45560 5850 45612 5856
rect 46032 5710 46060 6870
rect 46124 6798 46152 8774
rect 46216 8634 46244 8842
rect 46204 8628 46256 8634
rect 46204 8570 46256 8576
rect 46112 6792 46164 6798
rect 46112 6734 46164 6740
rect 46020 5704 46072 5710
rect 46020 5646 46072 5652
rect 46204 5228 46256 5234
rect 46204 5170 46256 5176
rect 45468 5160 45520 5166
rect 45468 5102 45520 5108
rect 45376 5092 45428 5098
rect 45376 5034 45428 5040
rect 44468 2746 44588 2774
rect 44652 2746 44772 2774
rect 44836 4950 45048 4978
rect 44468 2650 44496 2746
rect 44456 2644 44508 2650
rect 44456 2586 44508 2592
rect 44456 2372 44508 2378
rect 44456 2314 44508 2320
rect 44284 2094 44404 2122
rect 44088 1148 44140 1154
rect 44088 1090 44140 1096
rect 43812 876 43864 882
rect 43812 818 43864 824
rect 44008 836 44128 864
rect 44008 800 44036 836
rect 41420 750 41472 756
rect 41510 0 41566 800
rect 41786 0 41842 800
rect 42062 0 42118 800
rect 42338 0 42394 800
rect 42614 0 42670 800
rect 42890 0 42946 800
rect 43166 0 43222 800
rect 43442 0 43498 800
rect 43718 0 43774 800
rect 43994 0 44050 800
rect 44100 134 44128 836
rect 44284 800 44312 2094
rect 44468 950 44496 2314
rect 44652 2038 44680 2746
rect 44836 2514 44864 4950
rect 45192 4276 45244 4282
rect 45192 4218 45244 4224
rect 44916 3120 44968 3126
rect 44916 3062 44968 3068
rect 44824 2508 44876 2514
rect 44824 2450 44876 2456
rect 44640 2032 44692 2038
rect 44640 1974 44692 1980
rect 44928 1578 44956 3062
rect 45204 2122 45232 4218
rect 45388 3058 45416 5034
rect 45652 4548 45704 4554
rect 45652 4490 45704 4496
rect 46020 4548 46072 4554
rect 46020 4490 46072 4496
rect 45468 3460 45520 3466
rect 45468 3402 45520 3408
rect 45284 3052 45336 3058
rect 45284 2994 45336 3000
rect 45376 3052 45428 3058
rect 45376 2994 45428 3000
rect 45296 2854 45324 2994
rect 45284 2848 45336 2854
rect 45284 2790 45336 2796
rect 44560 1550 44956 1578
rect 45112 2094 45232 2122
rect 44456 944 44508 950
rect 44456 886 44508 892
rect 44560 800 44588 1550
rect 44824 944 44876 950
rect 44824 886 44876 892
rect 44836 800 44864 886
rect 45112 800 45140 2094
rect 45480 932 45508 3402
rect 45388 904 45508 932
rect 45388 800 45416 904
rect 45664 800 45692 4490
rect 46032 2774 46060 4490
rect 46112 3188 46164 3194
rect 46112 3130 46164 3136
rect 45940 2746 46060 2774
rect 45940 800 45968 2746
rect 46124 2650 46152 3130
rect 46112 2644 46164 2650
rect 46112 2586 46164 2592
rect 46020 2372 46072 2378
rect 46020 2314 46072 2320
rect 46112 2372 46164 2378
rect 46112 2314 46164 2320
rect 46032 1018 46060 2314
rect 46020 1012 46072 1018
rect 46020 954 46072 960
rect 46124 950 46152 2314
rect 46112 944 46164 950
rect 46112 886 46164 892
rect 46216 800 46244 5170
rect 46308 3194 46336 9030
rect 46400 8945 46428 12406
rect 46480 11824 46532 11830
rect 46480 11766 46532 11772
rect 46492 11150 46520 11766
rect 46664 11756 46716 11762
rect 46664 11698 46716 11704
rect 46480 11144 46532 11150
rect 46480 11086 46532 11092
rect 46386 8936 46442 8945
rect 46386 8871 46442 8880
rect 46480 8424 46532 8430
rect 46480 8366 46532 8372
rect 46388 6656 46440 6662
rect 46388 6598 46440 6604
rect 46400 6458 46428 6598
rect 46388 6452 46440 6458
rect 46388 6394 46440 6400
rect 46388 6112 46440 6118
rect 46388 6054 46440 6060
rect 46400 5846 46428 6054
rect 46388 5840 46440 5846
rect 46388 5782 46440 5788
rect 46492 5098 46520 8366
rect 46572 7404 46624 7410
rect 46572 7346 46624 7352
rect 46584 5914 46612 7346
rect 46676 6798 46704 11698
rect 46756 11212 46808 11218
rect 46756 11154 46808 11160
rect 46768 10674 46796 11154
rect 46848 11144 46900 11150
rect 46848 11086 46900 11092
rect 46756 10668 46808 10674
rect 46756 10610 46808 10616
rect 46768 9518 46796 10610
rect 46756 9512 46808 9518
rect 46756 9454 46808 9460
rect 46664 6792 46716 6798
rect 46664 6734 46716 6740
rect 46664 6656 46716 6662
rect 46662 6624 46664 6633
rect 46716 6624 46718 6633
rect 46662 6559 46718 6568
rect 46676 6186 46704 6559
rect 46754 6488 46810 6497
rect 46754 6423 46810 6432
rect 46664 6180 46716 6186
rect 46664 6122 46716 6128
rect 46768 5914 46796 6423
rect 46572 5908 46624 5914
rect 46572 5850 46624 5856
rect 46756 5908 46808 5914
rect 46756 5850 46808 5856
rect 46664 5704 46716 5710
rect 46664 5646 46716 5652
rect 46676 5166 46704 5646
rect 46664 5160 46716 5166
rect 46664 5102 46716 5108
rect 46480 5092 46532 5098
rect 46480 5034 46532 5040
rect 46388 4684 46440 4690
rect 46388 4626 46440 4632
rect 46296 3188 46348 3194
rect 46296 3130 46348 3136
rect 46400 3126 46428 4626
rect 46480 4616 46532 4622
rect 46480 4558 46532 4564
rect 46388 3120 46440 3126
rect 46388 3062 46440 3068
rect 46296 3052 46348 3058
rect 46296 2994 46348 3000
rect 46308 1086 46336 2994
rect 46296 1080 46348 1086
rect 46296 1022 46348 1028
rect 46492 800 46520 4558
rect 46676 3942 46704 5102
rect 46860 4826 46888 11086
rect 46952 7886 46980 12786
rect 46940 7880 46992 7886
rect 46940 7822 46992 7828
rect 46952 7546 46980 7822
rect 46940 7540 46992 7546
rect 46940 7482 46992 7488
rect 46952 7002 46980 7482
rect 46940 6996 46992 7002
rect 46940 6938 46992 6944
rect 46848 4820 46900 4826
rect 46848 4762 46900 4768
rect 46664 3936 46716 3942
rect 46664 3878 46716 3884
rect 47044 2582 47072 25162
rect 47124 19236 47176 19242
rect 47124 19178 47176 19184
rect 47136 18970 47164 19178
rect 47124 18964 47176 18970
rect 47124 18906 47176 18912
rect 47124 16516 47176 16522
rect 47124 16458 47176 16464
rect 47136 16250 47164 16458
rect 47124 16244 47176 16250
rect 47124 16186 47176 16192
rect 47124 12232 47176 12238
rect 47124 12174 47176 12180
rect 47136 7342 47164 12174
rect 47228 8430 47256 26862
rect 47216 8424 47268 8430
rect 47216 8366 47268 8372
rect 47124 7336 47176 7342
rect 47124 7278 47176 7284
rect 47216 6996 47268 7002
rect 47216 6938 47268 6944
rect 47228 6662 47256 6938
rect 47216 6656 47268 6662
rect 47216 6598 47268 6604
rect 47228 5574 47256 6598
rect 47216 5568 47268 5574
rect 47216 5510 47268 5516
rect 47124 4072 47176 4078
rect 47124 4014 47176 4020
rect 47136 2650 47164 4014
rect 47320 3670 47348 50798
rect 47400 25288 47452 25294
rect 47400 25230 47452 25236
rect 47412 24954 47440 25230
rect 47400 24948 47452 24954
rect 47400 24890 47452 24896
rect 47400 24132 47452 24138
rect 47400 24074 47452 24080
rect 47412 4706 47440 24074
rect 47504 15638 47532 51274
rect 47780 51105 47808 51886
rect 48148 51542 48176 51886
rect 47952 51536 48004 51542
rect 47952 51478 48004 51484
rect 48136 51536 48188 51542
rect 48136 51478 48188 51484
rect 47766 51096 47822 51105
rect 47766 51031 47822 51040
rect 47964 34066 47992 51478
rect 48148 50998 48176 51478
rect 48228 51400 48280 51406
rect 48516 51354 48544 51886
rect 48596 51468 48648 51474
rect 48596 51410 48648 51416
rect 48280 51348 48544 51354
rect 48228 51342 48544 51348
rect 48240 51326 48544 51342
rect 48136 50992 48188 50998
rect 48136 50934 48188 50940
rect 48516 50862 48544 51326
rect 48504 50856 48556 50862
rect 48504 50798 48556 50804
rect 48516 50522 48544 50798
rect 48504 50516 48556 50522
rect 48504 50458 48556 50464
rect 48516 49774 48544 50458
rect 48608 50454 48636 51410
rect 48872 51400 48924 51406
rect 48872 51342 48924 51348
rect 48688 50992 48740 50998
rect 48688 50934 48740 50940
rect 48596 50448 48648 50454
rect 48596 50390 48648 50396
rect 48504 49768 48556 49774
rect 48504 49710 48556 49716
rect 48700 45830 48728 50934
rect 48884 50930 48912 51342
rect 48872 50924 48924 50930
rect 48872 50866 48924 50872
rect 48780 50244 48832 50250
rect 48780 50186 48832 50192
rect 48688 45824 48740 45830
rect 48688 45766 48740 45772
rect 48688 44736 48740 44742
rect 48688 44678 48740 44684
rect 48700 44305 48728 44678
rect 48686 44296 48742 44305
rect 48686 44231 48742 44240
rect 47952 34060 48004 34066
rect 47952 34002 48004 34008
rect 47676 33992 47728 33998
rect 47676 33934 47728 33940
rect 47584 30728 47636 30734
rect 47584 30670 47636 30676
rect 47596 30258 47624 30670
rect 47584 30252 47636 30258
rect 47584 30194 47636 30200
rect 47584 24948 47636 24954
rect 47584 24890 47636 24896
rect 47596 24206 47624 24890
rect 47688 24410 47716 33934
rect 47860 33856 47912 33862
rect 47860 33798 47912 33804
rect 47768 32020 47820 32026
rect 47768 31962 47820 31968
rect 47780 30734 47808 31962
rect 47768 30728 47820 30734
rect 47768 30670 47820 30676
rect 47872 25498 47900 33798
rect 48792 31754 48820 50186
rect 48608 31726 48820 31754
rect 48136 31340 48188 31346
rect 48136 31282 48188 31288
rect 48320 31340 48372 31346
rect 48320 31282 48372 31288
rect 48148 30938 48176 31282
rect 48136 30932 48188 30938
rect 48136 30874 48188 30880
rect 48228 30320 48280 30326
rect 48228 30262 48280 30268
rect 47952 26512 48004 26518
rect 47952 26454 48004 26460
rect 47860 25492 47912 25498
rect 47860 25434 47912 25440
rect 47768 25152 47820 25158
rect 47768 25094 47820 25100
rect 47860 25152 47912 25158
rect 47860 25094 47912 25100
rect 47780 24886 47808 25094
rect 47768 24880 47820 24886
rect 47768 24822 47820 24828
rect 47676 24404 47728 24410
rect 47676 24346 47728 24352
rect 47584 24200 47636 24206
rect 47584 24142 47636 24148
rect 47676 22092 47728 22098
rect 47676 22034 47728 22040
rect 47688 21486 47716 22034
rect 47872 22001 47900 25094
rect 47964 24818 47992 26454
rect 48240 26382 48268 30262
rect 48332 28150 48360 31282
rect 48320 28144 48372 28150
rect 48320 28086 48372 28092
rect 48228 26376 48280 26382
rect 48228 26318 48280 26324
rect 48228 26240 48280 26246
rect 48228 26182 48280 26188
rect 48412 26240 48464 26246
rect 48412 26182 48464 26188
rect 48240 24886 48268 26182
rect 48424 25294 48452 26182
rect 48412 25288 48464 25294
rect 48412 25230 48464 25236
rect 48228 24880 48280 24886
rect 48228 24822 48280 24828
rect 47952 24812 48004 24818
rect 47952 24754 48004 24760
rect 48044 24608 48096 24614
rect 48044 24550 48096 24556
rect 48056 22778 48084 24550
rect 48226 23216 48282 23225
rect 48226 23151 48282 23160
rect 48240 23118 48268 23151
rect 48228 23112 48280 23118
rect 48228 23054 48280 23060
rect 48320 23044 48372 23050
rect 48320 22986 48372 22992
rect 48504 23044 48556 23050
rect 48504 22986 48556 22992
rect 48044 22772 48096 22778
rect 48044 22714 48096 22720
rect 47858 21992 47914 22001
rect 47858 21927 47860 21936
rect 47912 21927 47914 21936
rect 47860 21898 47912 21904
rect 47676 21480 47728 21486
rect 47676 21422 47728 21428
rect 48136 20800 48188 20806
rect 48136 20742 48188 20748
rect 47768 20596 47820 20602
rect 47768 20538 47820 20544
rect 47780 19854 47808 20538
rect 47952 20460 48004 20466
rect 47952 20402 48004 20408
rect 47768 19848 47820 19854
rect 47768 19790 47820 19796
rect 47860 19848 47912 19854
rect 47860 19790 47912 19796
rect 47676 18420 47728 18426
rect 47676 18362 47728 18368
rect 47584 17672 47636 17678
rect 47584 17614 47636 17620
rect 47492 15632 47544 15638
rect 47492 15574 47544 15580
rect 47492 15496 47544 15502
rect 47492 15438 47544 15444
rect 47504 15026 47532 15438
rect 47492 15020 47544 15026
rect 47492 14962 47544 14968
rect 47492 13184 47544 13190
rect 47492 13126 47544 13132
rect 47504 10062 47532 13126
rect 47492 10056 47544 10062
rect 47492 9998 47544 10004
rect 47504 7954 47532 9998
rect 47492 7948 47544 7954
rect 47492 7890 47544 7896
rect 47492 7336 47544 7342
rect 47492 7278 47544 7284
rect 47504 5846 47532 7278
rect 47492 5840 47544 5846
rect 47492 5782 47544 5788
rect 47412 4678 47532 4706
rect 47398 4584 47454 4593
rect 47398 4519 47454 4528
rect 47412 4486 47440 4519
rect 47400 4480 47452 4486
rect 47400 4422 47452 4428
rect 47504 4146 47532 4678
rect 47492 4140 47544 4146
rect 47492 4082 47544 4088
rect 47398 3768 47454 3777
rect 47596 3738 47624 17614
rect 47688 16574 47716 18362
rect 47780 17882 47808 19790
rect 47872 18086 47900 19790
rect 47964 18698 47992 20402
rect 48148 19854 48176 20742
rect 48332 20210 48360 22986
rect 48516 22778 48544 22986
rect 48504 22772 48556 22778
rect 48504 22714 48556 22720
rect 48412 22568 48464 22574
rect 48412 22510 48464 22516
rect 48424 20942 48452 22510
rect 48608 22094 48636 31726
rect 48688 30592 48740 30598
rect 48688 30534 48740 30540
rect 48700 28490 48728 30534
rect 48688 28484 48740 28490
rect 48688 28426 48740 28432
rect 48700 27402 48728 28426
rect 48884 28422 48912 50866
rect 49068 34066 49096 57190
rect 50294 56604 50602 56613
rect 50294 56602 50300 56604
rect 50356 56602 50380 56604
rect 50436 56602 50460 56604
rect 50516 56602 50540 56604
rect 50596 56602 50602 56604
rect 50356 56550 50358 56602
rect 50538 56550 50540 56602
rect 50294 56548 50300 56550
rect 50356 56548 50380 56550
rect 50436 56548 50460 56550
rect 50516 56548 50540 56550
rect 50596 56548 50602 56550
rect 50294 56539 50602 56548
rect 50294 55516 50602 55525
rect 50294 55514 50300 55516
rect 50356 55514 50380 55516
rect 50436 55514 50460 55516
rect 50516 55514 50540 55516
rect 50596 55514 50602 55516
rect 50356 55462 50358 55514
rect 50538 55462 50540 55514
rect 50294 55460 50300 55462
rect 50356 55460 50380 55462
rect 50436 55460 50460 55462
rect 50516 55460 50540 55462
rect 50596 55460 50602 55462
rect 50294 55451 50602 55460
rect 50294 54428 50602 54437
rect 50294 54426 50300 54428
rect 50356 54426 50380 54428
rect 50436 54426 50460 54428
rect 50516 54426 50540 54428
rect 50596 54426 50602 54428
rect 50356 54374 50358 54426
rect 50538 54374 50540 54426
rect 50294 54372 50300 54374
rect 50356 54372 50380 54374
rect 50436 54372 50460 54374
rect 50516 54372 50540 54374
rect 50596 54372 50602 54374
rect 50294 54363 50602 54372
rect 50294 53340 50602 53349
rect 50294 53338 50300 53340
rect 50356 53338 50380 53340
rect 50436 53338 50460 53340
rect 50516 53338 50540 53340
rect 50596 53338 50602 53340
rect 50356 53286 50358 53338
rect 50538 53286 50540 53338
rect 50294 53284 50300 53286
rect 50356 53284 50380 53286
rect 50436 53284 50460 53286
rect 50516 53284 50540 53286
rect 50596 53284 50602 53286
rect 50294 53275 50602 53284
rect 50294 52252 50602 52261
rect 50294 52250 50300 52252
rect 50356 52250 50380 52252
rect 50436 52250 50460 52252
rect 50516 52250 50540 52252
rect 50596 52250 50602 52252
rect 50356 52198 50358 52250
rect 50538 52198 50540 52250
rect 50294 52196 50300 52198
rect 50356 52196 50380 52198
rect 50436 52196 50460 52198
rect 50516 52196 50540 52198
rect 50596 52196 50602 52198
rect 50294 52187 50602 52196
rect 50294 51164 50602 51173
rect 50294 51162 50300 51164
rect 50356 51162 50380 51164
rect 50436 51162 50460 51164
rect 50516 51162 50540 51164
rect 50596 51162 50602 51164
rect 50356 51110 50358 51162
rect 50538 51110 50540 51162
rect 50294 51108 50300 51110
rect 50356 51108 50380 51110
rect 50436 51108 50460 51110
rect 50516 51108 50540 51110
rect 50596 51108 50602 51110
rect 50294 51099 50602 51108
rect 49240 50788 49292 50794
rect 49240 50730 49292 50736
rect 49148 50720 49200 50726
rect 49148 50662 49200 50668
rect 49160 50386 49188 50662
rect 49252 50454 49280 50730
rect 49424 50516 49476 50522
rect 49424 50458 49476 50464
rect 49240 50448 49292 50454
rect 49240 50390 49292 50396
rect 49148 50380 49200 50386
rect 49148 50322 49200 50328
rect 49252 45554 49280 50390
rect 49436 50386 49464 50458
rect 49424 50380 49476 50386
rect 49424 50322 49476 50328
rect 49608 50244 49660 50250
rect 49608 50186 49660 50192
rect 49160 45526 49280 45554
rect 49160 40458 49188 45526
rect 49332 44940 49384 44946
rect 49332 44882 49384 44888
rect 49344 44402 49372 44882
rect 49332 44396 49384 44402
rect 49332 44338 49384 44344
rect 49148 40452 49200 40458
rect 49148 40394 49200 40400
rect 49056 34060 49108 34066
rect 49056 34002 49108 34008
rect 49240 28552 49292 28558
rect 49240 28494 49292 28500
rect 48872 28416 48924 28422
rect 48872 28358 48924 28364
rect 48688 27396 48740 27402
rect 48688 27338 48740 27344
rect 48700 26314 48728 27338
rect 48780 26444 48832 26450
rect 48780 26386 48832 26392
rect 48688 26308 48740 26314
rect 48688 26250 48740 26256
rect 48792 25650 48820 26386
rect 48884 25838 48912 28358
rect 48964 27532 49016 27538
rect 48964 27474 49016 27480
rect 48976 26382 49004 27474
rect 49252 26450 49280 28494
rect 49424 27464 49476 27470
rect 49424 27406 49476 27412
rect 49436 26926 49464 27406
rect 49424 26920 49476 26926
rect 49424 26862 49476 26868
rect 49240 26444 49292 26450
rect 49240 26386 49292 26392
rect 48964 26376 49016 26382
rect 48964 26318 49016 26324
rect 49252 26330 49280 26386
rect 49424 26376 49476 26382
rect 49252 26324 49424 26330
rect 49252 26318 49476 26324
rect 49252 26302 49464 26318
rect 48872 25832 48924 25838
rect 48872 25774 48924 25780
rect 48792 25622 48912 25650
rect 48688 22976 48740 22982
rect 48688 22918 48740 22924
rect 48516 22066 48636 22094
rect 48516 21457 48544 22066
rect 48700 22030 48728 22918
rect 48780 22636 48832 22642
rect 48780 22578 48832 22584
rect 48792 22234 48820 22578
rect 48780 22228 48832 22234
rect 48780 22170 48832 22176
rect 48596 22024 48648 22030
rect 48596 21966 48648 21972
rect 48688 22024 48740 22030
rect 48688 21966 48740 21972
rect 48502 21448 48558 21457
rect 48502 21383 48558 21392
rect 48502 21312 48558 21321
rect 48502 21247 48558 21256
rect 48412 20936 48464 20942
rect 48412 20878 48464 20884
rect 48424 20534 48452 20878
rect 48412 20528 48464 20534
rect 48412 20470 48464 20476
rect 48240 20182 48360 20210
rect 48136 19848 48188 19854
rect 48136 19790 48188 19796
rect 48240 19530 48268 20182
rect 48320 20052 48372 20058
rect 48320 19994 48372 20000
rect 48056 19502 48268 19530
rect 48056 19446 48084 19502
rect 48044 19440 48096 19446
rect 48044 19382 48096 19388
rect 48056 19258 48084 19382
rect 48136 19372 48188 19378
rect 48332 19360 48360 19994
rect 48424 19378 48452 20470
rect 48188 19332 48360 19360
rect 48412 19372 48464 19378
rect 48136 19314 48188 19320
rect 48412 19314 48464 19320
rect 48056 19230 48360 19258
rect 47952 18692 48004 18698
rect 47952 18634 48004 18640
rect 47860 18080 47912 18086
rect 47860 18022 47912 18028
rect 47768 17876 47820 17882
rect 47768 17818 47820 17824
rect 47964 16574 47992 18634
rect 48332 18086 48360 19230
rect 48516 18834 48544 21247
rect 48608 19854 48636 21966
rect 48780 21548 48832 21554
rect 48780 21490 48832 21496
rect 48688 21344 48740 21350
rect 48688 21286 48740 21292
rect 48700 20942 48728 21286
rect 48688 20936 48740 20942
rect 48688 20878 48740 20884
rect 48792 20602 48820 21490
rect 48780 20596 48832 20602
rect 48780 20538 48832 20544
rect 48688 20460 48740 20466
rect 48688 20402 48740 20408
rect 48700 20369 48728 20402
rect 48686 20360 48742 20369
rect 48686 20295 48742 20304
rect 48596 19848 48648 19854
rect 48596 19790 48648 19796
rect 48884 19666 48912 25622
rect 49056 25220 49108 25226
rect 49056 25162 49108 25168
rect 48964 19780 49016 19786
rect 48964 19722 49016 19728
rect 48608 19638 48912 19666
rect 48504 18828 48556 18834
rect 48504 18770 48556 18776
rect 48516 18222 48544 18770
rect 48504 18216 48556 18222
rect 48504 18158 48556 18164
rect 48320 18080 48372 18086
rect 48320 18022 48372 18028
rect 48410 17912 48466 17921
rect 48410 17847 48466 17856
rect 48424 17678 48452 17847
rect 48412 17672 48464 17678
rect 48412 17614 48464 17620
rect 48516 17338 48544 18158
rect 48504 17332 48556 17338
rect 48504 17274 48556 17280
rect 48320 17196 48372 17202
rect 48320 17138 48372 17144
rect 48504 17196 48556 17202
rect 48504 17138 48556 17144
rect 48228 17128 48280 17134
rect 48226 17096 48228 17105
rect 48280 17096 48282 17105
rect 48226 17031 48282 17040
rect 48332 16640 48360 17138
rect 48412 17128 48464 17134
rect 48410 17096 48412 17105
rect 48464 17096 48466 17105
rect 48410 17031 48466 17040
rect 48412 16992 48464 16998
rect 48412 16934 48464 16940
rect 47688 16546 47808 16574
rect 47676 16448 47728 16454
rect 47676 16390 47728 16396
rect 47688 15502 47716 16390
rect 47780 16250 47808 16546
rect 47872 16546 47992 16574
rect 48240 16612 48360 16640
rect 48240 16561 48268 16612
rect 48226 16552 48282 16561
rect 47768 16244 47820 16250
rect 47768 16186 47820 16192
rect 47768 15632 47820 15638
rect 47768 15574 47820 15580
rect 47676 15496 47728 15502
rect 47676 15438 47728 15444
rect 47780 11898 47808 15574
rect 47768 11892 47820 11898
rect 47768 11834 47820 11840
rect 47872 8616 47900 16546
rect 48424 16522 48452 16934
rect 48226 16487 48282 16496
rect 48412 16516 48464 16522
rect 48412 16458 48464 16464
rect 48136 16244 48188 16250
rect 48136 16186 48188 16192
rect 48044 16108 48096 16114
rect 48044 16050 48096 16056
rect 47952 15428 48004 15434
rect 47952 15370 48004 15376
rect 47964 12850 47992 15370
rect 48056 15162 48084 16050
rect 48148 15502 48176 16186
rect 48320 16176 48372 16182
rect 48320 16118 48372 16124
rect 48136 15496 48188 15502
rect 48136 15438 48188 15444
rect 48044 15156 48096 15162
rect 48044 15098 48096 15104
rect 48332 13530 48360 16118
rect 48424 14482 48452 16458
rect 48412 14476 48464 14482
rect 48412 14418 48464 14424
rect 48320 13524 48372 13530
rect 48320 13466 48372 13472
rect 47952 12844 48004 12850
rect 47952 12786 48004 12792
rect 48332 12434 48360 13466
rect 48332 12406 48452 12434
rect 48320 11552 48372 11558
rect 48320 11494 48372 11500
rect 48332 9994 48360 11494
rect 48320 9988 48372 9994
rect 48320 9930 48372 9936
rect 48424 8906 48452 12406
rect 48412 8900 48464 8906
rect 48412 8842 48464 8848
rect 47780 8588 47900 8616
rect 47676 8560 47728 8566
rect 47676 8502 47728 8508
rect 47688 7206 47716 8502
rect 47676 7200 47728 7206
rect 47676 7142 47728 7148
rect 47676 6724 47728 6730
rect 47676 6666 47728 6672
rect 47688 6322 47716 6666
rect 47676 6316 47728 6322
rect 47676 6258 47728 6264
rect 47780 4434 47808 8588
rect 47872 8498 48360 8514
rect 47860 8492 48372 8498
rect 47912 8486 48320 8492
rect 47860 8434 47912 8440
rect 48320 8434 48372 8440
rect 48136 8356 48188 8362
rect 48136 8298 48188 8304
rect 48148 7993 48176 8298
rect 48134 7984 48190 7993
rect 48134 7919 48190 7928
rect 48136 7812 48188 7818
rect 48136 7754 48188 7760
rect 47952 7744 48004 7750
rect 47952 7686 48004 7692
rect 47964 7410 47992 7686
rect 48148 7546 48176 7754
rect 48136 7540 48188 7546
rect 48136 7482 48188 7488
rect 47952 7404 48004 7410
rect 47952 7346 48004 7352
rect 48136 7200 48188 7206
rect 48136 7142 48188 7148
rect 47860 6792 47912 6798
rect 47860 6734 47912 6740
rect 47872 6118 47900 6734
rect 47860 6112 47912 6118
rect 47860 6054 47912 6060
rect 48042 5536 48098 5545
rect 48042 5471 48098 5480
rect 47952 5296 48004 5302
rect 47952 5238 48004 5244
rect 47688 4406 47808 4434
rect 47398 3703 47454 3712
rect 47584 3732 47636 3738
rect 47308 3664 47360 3670
rect 47308 3606 47360 3612
rect 47412 3534 47440 3703
rect 47584 3674 47636 3680
rect 47688 3641 47716 4406
rect 47766 4312 47822 4321
rect 47766 4247 47822 4256
rect 47780 4146 47808 4247
rect 47768 4140 47820 4146
rect 47768 4082 47820 4088
rect 47858 4040 47914 4049
rect 47858 3975 47914 3984
rect 47674 3632 47730 3641
rect 47674 3567 47730 3576
rect 47400 3528 47452 3534
rect 47400 3470 47452 3476
rect 47216 3460 47268 3466
rect 47216 3402 47268 3408
rect 47308 3460 47360 3466
rect 47308 3402 47360 3408
rect 47228 2990 47256 3402
rect 47320 3126 47348 3402
rect 47308 3120 47360 3126
rect 47308 3062 47360 3068
rect 47872 3058 47900 3975
rect 47964 3534 47992 5238
rect 48056 4622 48084 5471
rect 48148 4842 48176 7142
rect 48226 6760 48282 6769
rect 48226 6695 48282 6704
rect 48240 6662 48268 6695
rect 48228 6656 48280 6662
rect 48228 6598 48280 6604
rect 48424 6458 48452 8842
rect 48412 6452 48464 6458
rect 48412 6394 48464 6400
rect 48148 4814 48360 4842
rect 48228 4752 48280 4758
rect 48228 4694 48280 4700
rect 48044 4616 48096 4622
rect 48044 4558 48096 4564
rect 48044 4276 48096 4282
rect 48096 4236 48176 4264
rect 48044 4218 48096 4224
rect 47952 3528 48004 3534
rect 47952 3470 48004 3476
rect 47860 3052 47912 3058
rect 47860 2994 47912 3000
rect 48044 3052 48096 3058
rect 48044 2994 48096 3000
rect 47216 2984 47268 2990
rect 47216 2926 47268 2932
rect 47768 2984 47820 2990
rect 47768 2926 47820 2932
rect 47124 2644 47176 2650
rect 47124 2586 47176 2592
rect 47032 2576 47084 2582
rect 47032 2518 47084 2524
rect 47780 2378 47808 2926
rect 47950 2680 48006 2689
rect 47950 2615 48006 2624
rect 47964 2446 47992 2615
rect 48056 2582 48084 2994
rect 48044 2576 48096 2582
rect 48044 2518 48096 2524
rect 48148 2530 48176 4236
rect 48240 3058 48268 4694
rect 48332 4622 48360 4814
rect 48412 4752 48464 4758
rect 48412 4694 48464 4700
rect 48320 4616 48372 4622
rect 48320 4558 48372 4564
rect 48320 4140 48372 4146
rect 48424 4128 48452 4694
rect 48372 4100 48452 4128
rect 48320 4082 48372 4088
rect 48320 4004 48372 4010
rect 48320 3946 48372 3952
rect 48228 3052 48280 3058
rect 48228 2994 48280 3000
rect 48148 2502 48268 2530
rect 47952 2440 48004 2446
rect 47952 2382 48004 2388
rect 48136 2440 48188 2446
rect 48136 2382 48188 2388
rect 47768 2372 47820 2378
rect 47768 2314 47820 2320
rect 48148 2106 48176 2382
rect 48136 2100 48188 2106
rect 48136 2042 48188 2048
rect 48240 1986 48268 2502
rect 48332 2446 48360 3946
rect 48424 3194 48452 4100
rect 48516 3194 48544 17138
rect 48608 11150 48636 19638
rect 48780 18760 48832 18766
rect 48780 18702 48832 18708
rect 48688 18284 48740 18290
rect 48688 18226 48740 18232
rect 48596 11144 48648 11150
rect 48596 11086 48648 11092
rect 48596 9036 48648 9042
rect 48596 8978 48648 8984
rect 48608 6798 48636 8978
rect 48596 6792 48648 6798
rect 48596 6734 48648 6740
rect 48608 6186 48636 6734
rect 48596 6180 48648 6186
rect 48596 6122 48648 6128
rect 48700 4826 48728 18226
rect 48792 16674 48820 18702
rect 48976 18426 49004 19722
rect 49068 18834 49096 25162
rect 49240 23112 49292 23118
rect 49240 23054 49292 23060
rect 49252 22642 49280 23054
rect 49240 22636 49292 22642
rect 49240 22578 49292 22584
rect 49148 22432 49200 22438
rect 49148 22374 49200 22380
rect 49160 22234 49188 22374
rect 49148 22228 49200 22234
rect 49148 22170 49200 22176
rect 49252 22094 49280 22578
rect 49160 22066 49280 22094
rect 49160 20602 49188 22066
rect 49148 20596 49200 20602
rect 49148 20538 49200 20544
rect 49160 20058 49188 20538
rect 49148 20052 49200 20058
rect 49148 19994 49200 20000
rect 49148 19848 49200 19854
rect 49148 19790 49200 19796
rect 49160 19514 49188 19790
rect 49240 19780 49292 19786
rect 49240 19722 49292 19728
rect 49516 19780 49568 19786
rect 49516 19722 49568 19728
rect 49148 19508 49200 19514
rect 49148 19450 49200 19456
rect 49252 19258 49280 19722
rect 49332 19712 49384 19718
rect 49332 19654 49384 19660
rect 49344 19446 49372 19654
rect 49528 19514 49556 19722
rect 49516 19508 49568 19514
rect 49516 19450 49568 19456
rect 49332 19440 49384 19446
rect 49332 19382 49384 19388
rect 49252 19230 49372 19258
rect 49056 18828 49108 18834
rect 49056 18770 49108 18776
rect 48964 18420 49016 18426
rect 48964 18362 49016 18368
rect 48872 18284 48924 18290
rect 48872 18226 48924 18232
rect 48884 17678 48912 18226
rect 48976 17746 49004 18362
rect 49068 18290 49096 18770
rect 49056 18284 49108 18290
rect 49056 18226 49108 18232
rect 48964 17740 49016 17746
rect 48964 17682 49016 17688
rect 48872 17672 48924 17678
rect 48872 17614 48924 17620
rect 49056 17672 49108 17678
rect 49056 17614 49108 17620
rect 49240 17672 49292 17678
rect 49240 17614 49292 17620
rect 48884 17116 48912 17614
rect 48964 17128 49016 17134
rect 48884 17088 48964 17116
rect 48964 17070 49016 17076
rect 49068 16794 49096 17614
rect 49056 16788 49108 16794
rect 49056 16730 49108 16736
rect 48792 16646 49188 16674
rect 48872 15360 48924 15366
rect 48872 15302 48924 15308
rect 48884 12434 48912 15302
rect 48884 12406 49004 12434
rect 48780 11756 48832 11762
rect 48780 11698 48832 11704
rect 48792 11354 48820 11698
rect 48872 11620 48924 11626
rect 48872 11562 48924 11568
rect 48780 11348 48832 11354
rect 48780 11290 48832 11296
rect 48780 8832 48832 8838
rect 48780 8774 48832 8780
rect 48792 8362 48820 8774
rect 48780 8356 48832 8362
rect 48780 8298 48832 8304
rect 48688 4820 48740 4826
rect 48688 4762 48740 4768
rect 48780 4548 48832 4554
rect 48780 4490 48832 4496
rect 48596 4140 48648 4146
rect 48596 4082 48648 4088
rect 48608 4049 48636 4082
rect 48594 4040 48650 4049
rect 48594 3975 48650 3984
rect 48792 3534 48820 4490
rect 48884 4146 48912 11562
rect 48976 9042 49004 12406
rect 49056 11892 49108 11898
rect 49056 11834 49108 11840
rect 49068 11694 49096 11834
rect 49056 11688 49108 11694
rect 49056 11630 49108 11636
rect 48964 9036 49016 9042
rect 48964 8978 49016 8984
rect 48964 8900 49016 8906
rect 48964 8842 49016 8848
rect 48976 8498 49004 8842
rect 48964 8492 49016 8498
rect 48964 8434 49016 8440
rect 49056 8424 49108 8430
rect 49056 8366 49108 8372
rect 48964 8288 49016 8294
rect 48964 8230 49016 8236
rect 48976 7478 49004 8230
rect 48964 7472 49016 7478
rect 48964 7414 49016 7420
rect 48872 4140 48924 4146
rect 48872 4082 48924 4088
rect 48596 3528 48648 3534
rect 48596 3470 48648 3476
rect 48780 3528 48832 3534
rect 48780 3470 48832 3476
rect 48608 3194 48636 3470
rect 48412 3188 48464 3194
rect 48412 3130 48464 3136
rect 48504 3188 48556 3194
rect 48504 3130 48556 3136
rect 48596 3188 48648 3194
rect 48596 3130 48648 3136
rect 48424 3097 48452 3130
rect 48410 3088 48466 3097
rect 48594 3088 48650 3097
rect 48410 3023 48412 3032
rect 48464 3023 48466 3032
rect 48504 3052 48556 3058
rect 48412 2994 48464 3000
rect 48594 3023 48650 3032
rect 48504 2994 48556 3000
rect 48516 2774 48544 2994
rect 48424 2746 48544 2774
rect 48320 2440 48372 2446
rect 48320 2382 48372 2388
rect 48148 1958 48268 1986
rect 47032 1216 47084 1222
rect 47032 1158 47084 1164
rect 46676 870 46796 898
rect 46676 814 46704 870
rect 46664 808 46716 814
rect 44088 128 44140 134
rect 44088 70 44140 76
rect 44270 0 44326 800
rect 44546 0 44602 800
rect 44822 0 44878 800
rect 45098 0 45154 800
rect 45374 0 45430 800
rect 45650 0 45706 800
rect 45926 0 45982 800
rect 46202 0 46258 800
rect 46478 0 46534 800
rect 46768 800 46796 870
rect 47044 800 47072 1158
rect 47584 1148 47636 1154
rect 47584 1090 47636 1096
rect 47308 1080 47360 1086
rect 47308 1022 47360 1028
rect 47320 800 47348 1022
rect 47596 800 47624 1090
rect 47860 944 47912 950
rect 47860 886 47912 892
rect 47872 800 47900 886
rect 48148 800 48176 1958
rect 48424 800 48452 2746
rect 48608 2446 48636 3023
rect 48792 2990 48820 3470
rect 48780 2984 48832 2990
rect 48780 2926 48832 2932
rect 48884 2514 48912 4082
rect 49068 2990 49096 8366
rect 49056 2984 49108 2990
rect 49056 2926 49108 2932
rect 49160 2650 49188 16646
rect 49252 16590 49280 17614
rect 49240 16584 49292 16590
rect 49344 16561 49372 19230
rect 49516 18624 49568 18630
rect 49516 18566 49568 18572
rect 49424 18284 49476 18290
rect 49424 18226 49476 18232
rect 49240 16526 49292 16532
rect 49330 16552 49386 16561
rect 49252 15366 49280 16526
rect 49330 16487 49386 16496
rect 49240 15360 49292 15366
rect 49240 15302 49292 15308
rect 49344 12238 49372 16487
rect 49436 13258 49464 18226
rect 49528 16250 49556 18566
rect 49516 16244 49568 16250
rect 49516 16186 49568 16192
rect 49424 13252 49476 13258
rect 49424 13194 49476 13200
rect 49436 12918 49464 13194
rect 49424 12912 49476 12918
rect 49424 12854 49476 12860
rect 49332 12232 49384 12238
rect 49332 12174 49384 12180
rect 49332 11280 49384 11286
rect 49332 11222 49384 11228
rect 49240 11008 49292 11014
rect 49240 10950 49292 10956
rect 49252 4622 49280 10950
rect 49240 4616 49292 4622
rect 49240 4558 49292 4564
rect 49252 3534 49280 4558
rect 49240 3528 49292 3534
rect 49240 3470 49292 3476
rect 49238 2952 49294 2961
rect 49238 2887 49294 2896
rect 49252 2854 49280 2887
rect 49240 2848 49292 2854
rect 49240 2790 49292 2796
rect 49344 2650 49372 11222
rect 49620 5302 49648 50186
rect 50294 50076 50602 50085
rect 50294 50074 50300 50076
rect 50356 50074 50380 50076
rect 50436 50074 50460 50076
rect 50516 50074 50540 50076
rect 50596 50074 50602 50076
rect 50356 50022 50358 50074
rect 50538 50022 50540 50074
rect 50294 50020 50300 50022
rect 50356 50020 50380 50022
rect 50436 50020 50460 50022
rect 50516 50020 50540 50022
rect 50596 50020 50602 50022
rect 50294 50011 50602 50020
rect 50294 48988 50602 48997
rect 50294 48986 50300 48988
rect 50356 48986 50380 48988
rect 50436 48986 50460 48988
rect 50516 48986 50540 48988
rect 50596 48986 50602 48988
rect 50356 48934 50358 48986
rect 50538 48934 50540 48986
rect 50294 48932 50300 48934
rect 50356 48932 50380 48934
rect 50436 48932 50460 48934
rect 50516 48932 50540 48934
rect 50596 48932 50602 48934
rect 50294 48923 50602 48932
rect 50294 47900 50602 47909
rect 50294 47898 50300 47900
rect 50356 47898 50380 47900
rect 50436 47898 50460 47900
rect 50516 47898 50540 47900
rect 50596 47898 50602 47900
rect 50356 47846 50358 47898
rect 50538 47846 50540 47898
rect 50294 47844 50300 47846
rect 50356 47844 50380 47846
rect 50436 47844 50460 47846
rect 50516 47844 50540 47846
rect 50596 47844 50602 47846
rect 50294 47835 50602 47844
rect 50294 46812 50602 46821
rect 50294 46810 50300 46812
rect 50356 46810 50380 46812
rect 50436 46810 50460 46812
rect 50516 46810 50540 46812
rect 50596 46810 50602 46812
rect 50356 46758 50358 46810
rect 50538 46758 50540 46810
rect 50294 46756 50300 46758
rect 50356 46756 50380 46758
rect 50436 46756 50460 46758
rect 50516 46756 50540 46758
rect 50596 46756 50602 46758
rect 50294 46747 50602 46756
rect 50712 46504 50764 46510
rect 50712 46446 50764 46452
rect 50294 45724 50602 45733
rect 50294 45722 50300 45724
rect 50356 45722 50380 45724
rect 50436 45722 50460 45724
rect 50516 45722 50540 45724
rect 50596 45722 50602 45724
rect 50356 45670 50358 45722
rect 50538 45670 50540 45722
rect 50294 45668 50300 45670
rect 50356 45668 50380 45670
rect 50436 45668 50460 45670
rect 50516 45668 50540 45670
rect 50596 45668 50602 45670
rect 50294 45659 50602 45668
rect 50294 44636 50602 44645
rect 50294 44634 50300 44636
rect 50356 44634 50380 44636
rect 50436 44634 50460 44636
rect 50516 44634 50540 44636
rect 50596 44634 50602 44636
rect 50356 44582 50358 44634
rect 50538 44582 50540 44634
rect 50294 44580 50300 44582
rect 50356 44580 50380 44582
rect 50436 44580 50460 44582
rect 50516 44580 50540 44582
rect 50596 44580 50602 44582
rect 50294 44571 50602 44580
rect 50294 43548 50602 43557
rect 50294 43546 50300 43548
rect 50356 43546 50380 43548
rect 50436 43546 50460 43548
rect 50516 43546 50540 43548
rect 50596 43546 50602 43548
rect 50356 43494 50358 43546
rect 50538 43494 50540 43546
rect 50294 43492 50300 43494
rect 50356 43492 50380 43494
rect 50436 43492 50460 43494
rect 50516 43492 50540 43494
rect 50596 43492 50602 43494
rect 50294 43483 50602 43492
rect 50294 42460 50602 42469
rect 50294 42458 50300 42460
rect 50356 42458 50380 42460
rect 50436 42458 50460 42460
rect 50516 42458 50540 42460
rect 50596 42458 50602 42460
rect 50356 42406 50358 42458
rect 50538 42406 50540 42458
rect 50294 42404 50300 42406
rect 50356 42404 50380 42406
rect 50436 42404 50460 42406
rect 50516 42404 50540 42406
rect 50596 42404 50602 42406
rect 50294 42395 50602 42404
rect 50294 41372 50602 41381
rect 50294 41370 50300 41372
rect 50356 41370 50380 41372
rect 50436 41370 50460 41372
rect 50516 41370 50540 41372
rect 50596 41370 50602 41372
rect 50356 41318 50358 41370
rect 50538 41318 50540 41370
rect 50294 41316 50300 41318
rect 50356 41316 50380 41318
rect 50436 41316 50460 41318
rect 50516 41316 50540 41318
rect 50596 41316 50602 41318
rect 50294 41307 50602 41316
rect 50294 40284 50602 40293
rect 50294 40282 50300 40284
rect 50356 40282 50380 40284
rect 50436 40282 50460 40284
rect 50516 40282 50540 40284
rect 50596 40282 50602 40284
rect 50356 40230 50358 40282
rect 50538 40230 50540 40282
rect 50294 40228 50300 40230
rect 50356 40228 50380 40230
rect 50436 40228 50460 40230
rect 50516 40228 50540 40230
rect 50596 40228 50602 40230
rect 50294 40219 50602 40228
rect 50294 39196 50602 39205
rect 50294 39194 50300 39196
rect 50356 39194 50380 39196
rect 50436 39194 50460 39196
rect 50516 39194 50540 39196
rect 50596 39194 50602 39196
rect 50356 39142 50358 39194
rect 50538 39142 50540 39194
rect 50294 39140 50300 39142
rect 50356 39140 50380 39142
rect 50436 39140 50460 39142
rect 50516 39140 50540 39142
rect 50596 39140 50602 39142
rect 50294 39131 50602 39140
rect 50294 38108 50602 38117
rect 50294 38106 50300 38108
rect 50356 38106 50380 38108
rect 50436 38106 50460 38108
rect 50516 38106 50540 38108
rect 50596 38106 50602 38108
rect 50356 38054 50358 38106
rect 50538 38054 50540 38106
rect 50294 38052 50300 38054
rect 50356 38052 50380 38054
rect 50436 38052 50460 38054
rect 50516 38052 50540 38054
rect 50596 38052 50602 38054
rect 50294 38043 50602 38052
rect 50294 37020 50602 37029
rect 50294 37018 50300 37020
rect 50356 37018 50380 37020
rect 50436 37018 50460 37020
rect 50516 37018 50540 37020
rect 50596 37018 50602 37020
rect 50356 36966 50358 37018
rect 50538 36966 50540 37018
rect 50294 36964 50300 36966
rect 50356 36964 50380 36966
rect 50436 36964 50460 36966
rect 50516 36964 50540 36966
rect 50596 36964 50602 36966
rect 50294 36955 50602 36964
rect 50294 35932 50602 35941
rect 50294 35930 50300 35932
rect 50356 35930 50380 35932
rect 50436 35930 50460 35932
rect 50516 35930 50540 35932
rect 50596 35930 50602 35932
rect 50356 35878 50358 35930
rect 50538 35878 50540 35930
rect 50294 35876 50300 35878
rect 50356 35876 50380 35878
rect 50436 35876 50460 35878
rect 50516 35876 50540 35878
rect 50596 35876 50602 35878
rect 50294 35867 50602 35876
rect 50294 34844 50602 34853
rect 50294 34842 50300 34844
rect 50356 34842 50380 34844
rect 50436 34842 50460 34844
rect 50516 34842 50540 34844
rect 50596 34842 50602 34844
rect 50356 34790 50358 34842
rect 50538 34790 50540 34842
rect 50294 34788 50300 34790
rect 50356 34788 50380 34790
rect 50436 34788 50460 34790
rect 50516 34788 50540 34790
rect 50596 34788 50602 34790
rect 50294 34779 50602 34788
rect 50294 33756 50602 33765
rect 50294 33754 50300 33756
rect 50356 33754 50380 33756
rect 50436 33754 50460 33756
rect 50516 33754 50540 33756
rect 50596 33754 50602 33756
rect 50356 33702 50358 33754
rect 50538 33702 50540 33754
rect 50294 33700 50300 33702
rect 50356 33700 50380 33702
rect 50436 33700 50460 33702
rect 50516 33700 50540 33702
rect 50596 33700 50602 33702
rect 50294 33691 50602 33700
rect 49884 32904 49936 32910
rect 49884 32846 49936 32852
rect 49700 29708 49752 29714
rect 49700 29650 49752 29656
rect 49608 5296 49660 5302
rect 49608 5238 49660 5244
rect 49516 3936 49568 3942
rect 49516 3878 49568 3884
rect 49424 3052 49476 3058
rect 49424 2994 49476 3000
rect 49148 2644 49200 2650
rect 49148 2586 49200 2592
rect 49332 2644 49384 2650
rect 49332 2586 49384 2592
rect 48872 2508 48924 2514
rect 48872 2450 48924 2456
rect 48596 2440 48648 2446
rect 48596 2382 48648 2388
rect 48504 2372 48556 2378
rect 48504 2314 48556 2320
rect 48516 950 48544 2314
rect 48964 1012 49016 1018
rect 48964 954 49016 960
rect 48504 944 48556 950
rect 48504 886 48556 892
rect 48700 882 48820 898
rect 48700 876 48832 882
rect 48700 870 48780 876
rect 48700 800 48728 870
rect 48780 818 48832 824
rect 48976 800 49004 954
rect 49240 944 49292 950
rect 49240 886 49292 892
rect 49252 800 49280 886
rect 46664 750 46716 756
rect 46754 0 46810 800
rect 47030 0 47086 800
rect 47306 0 47362 800
rect 47582 0 47638 800
rect 47858 0 47914 800
rect 48134 0 48190 800
rect 48410 0 48466 800
rect 48686 0 48742 800
rect 48962 0 49018 800
rect 49238 0 49294 800
rect 49436 134 49464 2994
rect 49528 800 49556 3878
rect 49712 2650 49740 29650
rect 49792 22772 49844 22778
rect 49792 22714 49844 22720
rect 49804 22438 49832 22714
rect 49792 22432 49844 22438
rect 49792 22374 49844 22380
rect 49792 21548 49844 21554
rect 49792 21490 49844 21496
rect 49804 19446 49832 21490
rect 49896 21146 49924 32846
rect 50294 32668 50602 32677
rect 50294 32666 50300 32668
rect 50356 32666 50380 32668
rect 50436 32666 50460 32668
rect 50516 32666 50540 32668
rect 50596 32666 50602 32668
rect 50356 32614 50358 32666
rect 50538 32614 50540 32666
rect 50294 32612 50300 32614
rect 50356 32612 50380 32614
rect 50436 32612 50460 32614
rect 50516 32612 50540 32614
rect 50596 32612 50602 32614
rect 50294 32603 50602 32612
rect 50294 31580 50602 31589
rect 50294 31578 50300 31580
rect 50356 31578 50380 31580
rect 50436 31578 50460 31580
rect 50516 31578 50540 31580
rect 50596 31578 50602 31580
rect 50356 31526 50358 31578
rect 50538 31526 50540 31578
rect 50294 31524 50300 31526
rect 50356 31524 50380 31526
rect 50436 31524 50460 31526
rect 50516 31524 50540 31526
rect 50596 31524 50602 31526
rect 50294 31515 50602 31524
rect 50294 30492 50602 30501
rect 50294 30490 50300 30492
rect 50356 30490 50380 30492
rect 50436 30490 50460 30492
rect 50516 30490 50540 30492
rect 50596 30490 50602 30492
rect 50356 30438 50358 30490
rect 50538 30438 50540 30490
rect 50294 30436 50300 30438
rect 50356 30436 50380 30438
rect 50436 30436 50460 30438
rect 50516 30436 50540 30438
rect 50596 30436 50602 30438
rect 50294 30427 50602 30436
rect 50294 29404 50602 29413
rect 50294 29402 50300 29404
rect 50356 29402 50380 29404
rect 50436 29402 50460 29404
rect 50516 29402 50540 29404
rect 50596 29402 50602 29404
rect 50356 29350 50358 29402
rect 50538 29350 50540 29402
rect 50294 29348 50300 29350
rect 50356 29348 50380 29350
rect 50436 29348 50460 29350
rect 50516 29348 50540 29350
rect 50596 29348 50602 29350
rect 50294 29339 50602 29348
rect 50724 28490 50752 46446
rect 50896 42288 50948 42294
rect 50896 42230 50948 42236
rect 50804 33108 50856 33114
rect 50804 33050 50856 33056
rect 50712 28484 50764 28490
rect 50712 28426 50764 28432
rect 50294 28316 50602 28325
rect 50294 28314 50300 28316
rect 50356 28314 50380 28316
rect 50436 28314 50460 28316
rect 50516 28314 50540 28316
rect 50596 28314 50602 28316
rect 50356 28262 50358 28314
rect 50538 28262 50540 28314
rect 50294 28260 50300 28262
rect 50356 28260 50380 28262
rect 50436 28260 50460 28262
rect 50516 28260 50540 28262
rect 50596 28260 50602 28262
rect 50294 28251 50602 28260
rect 50294 27228 50602 27237
rect 50294 27226 50300 27228
rect 50356 27226 50380 27228
rect 50436 27226 50460 27228
rect 50516 27226 50540 27228
rect 50596 27226 50602 27228
rect 50356 27174 50358 27226
rect 50538 27174 50540 27226
rect 50294 27172 50300 27174
rect 50356 27172 50380 27174
rect 50436 27172 50460 27174
rect 50516 27172 50540 27174
rect 50596 27172 50602 27174
rect 50294 27163 50602 27172
rect 50294 26140 50602 26149
rect 50294 26138 50300 26140
rect 50356 26138 50380 26140
rect 50436 26138 50460 26140
rect 50516 26138 50540 26140
rect 50596 26138 50602 26140
rect 50356 26086 50358 26138
rect 50538 26086 50540 26138
rect 50294 26084 50300 26086
rect 50356 26084 50380 26086
rect 50436 26084 50460 26086
rect 50516 26084 50540 26086
rect 50596 26084 50602 26086
rect 50294 26075 50602 26084
rect 50068 25764 50120 25770
rect 50068 25706 50120 25712
rect 49884 21140 49936 21146
rect 49884 21082 49936 21088
rect 49896 20466 49924 21082
rect 49884 20460 49936 20466
rect 49884 20402 49936 20408
rect 50080 20346 50108 25706
rect 50294 25052 50602 25061
rect 50294 25050 50300 25052
rect 50356 25050 50380 25052
rect 50436 25050 50460 25052
rect 50516 25050 50540 25052
rect 50596 25050 50602 25052
rect 50356 24998 50358 25050
rect 50538 24998 50540 25050
rect 50294 24996 50300 24998
rect 50356 24996 50380 24998
rect 50436 24996 50460 24998
rect 50516 24996 50540 24998
rect 50596 24996 50602 24998
rect 50294 24987 50602 24996
rect 50294 23964 50602 23973
rect 50294 23962 50300 23964
rect 50356 23962 50380 23964
rect 50436 23962 50460 23964
rect 50516 23962 50540 23964
rect 50596 23962 50602 23964
rect 50356 23910 50358 23962
rect 50538 23910 50540 23962
rect 50294 23908 50300 23910
rect 50356 23908 50380 23910
rect 50436 23908 50460 23910
rect 50516 23908 50540 23910
rect 50596 23908 50602 23910
rect 50294 23899 50602 23908
rect 50294 22876 50602 22885
rect 50294 22874 50300 22876
rect 50356 22874 50380 22876
rect 50436 22874 50460 22876
rect 50516 22874 50540 22876
rect 50596 22874 50602 22876
rect 50356 22822 50358 22874
rect 50538 22822 50540 22874
rect 50294 22820 50300 22822
rect 50356 22820 50380 22822
rect 50436 22820 50460 22822
rect 50516 22820 50540 22822
rect 50596 22820 50602 22822
rect 50294 22811 50602 22820
rect 50294 21788 50602 21797
rect 50294 21786 50300 21788
rect 50356 21786 50380 21788
rect 50436 21786 50460 21788
rect 50516 21786 50540 21788
rect 50596 21786 50602 21788
rect 50356 21734 50358 21786
rect 50538 21734 50540 21786
rect 50294 21732 50300 21734
rect 50356 21732 50380 21734
rect 50436 21732 50460 21734
rect 50516 21732 50540 21734
rect 50596 21732 50602 21734
rect 50294 21723 50602 21732
rect 50294 20700 50602 20709
rect 50294 20698 50300 20700
rect 50356 20698 50380 20700
rect 50436 20698 50460 20700
rect 50516 20698 50540 20700
rect 50596 20698 50602 20700
rect 50356 20646 50358 20698
rect 50538 20646 50540 20698
rect 50294 20644 50300 20646
rect 50356 20644 50380 20646
rect 50436 20644 50460 20646
rect 50516 20644 50540 20646
rect 50596 20644 50602 20646
rect 50294 20635 50602 20644
rect 50528 20596 50580 20602
rect 50528 20538 50580 20544
rect 50160 20460 50212 20466
rect 50160 20402 50212 20408
rect 49896 20318 50108 20346
rect 49792 19440 49844 19446
rect 49792 19382 49844 19388
rect 49896 16574 49924 20318
rect 50172 19802 50200 20402
rect 50436 20052 50488 20058
rect 50436 19994 50488 20000
rect 50080 19774 50200 19802
rect 50080 19514 50108 19774
rect 50448 19718 50476 19994
rect 50540 19854 50568 20538
rect 50528 19848 50580 19854
rect 50528 19790 50580 19796
rect 50160 19712 50212 19718
rect 50160 19654 50212 19660
rect 50436 19712 50488 19718
rect 50436 19654 50488 19660
rect 50068 19508 50120 19514
rect 50068 19450 50120 19456
rect 50172 19378 50200 19654
rect 50294 19612 50602 19621
rect 50294 19610 50300 19612
rect 50356 19610 50380 19612
rect 50436 19610 50460 19612
rect 50516 19610 50540 19612
rect 50596 19610 50602 19612
rect 50356 19558 50358 19610
rect 50538 19558 50540 19610
rect 50294 19556 50300 19558
rect 50356 19556 50380 19558
rect 50436 19556 50460 19558
rect 50516 19556 50540 19558
rect 50596 19556 50602 19558
rect 50294 19547 50602 19556
rect 50160 19372 50212 19378
rect 50160 19314 50212 19320
rect 50294 18524 50602 18533
rect 50294 18522 50300 18524
rect 50356 18522 50380 18524
rect 50436 18522 50460 18524
rect 50516 18522 50540 18524
rect 50596 18522 50602 18524
rect 50356 18470 50358 18522
rect 50538 18470 50540 18522
rect 50294 18468 50300 18470
rect 50356 18468 50380 18470
rect 50436 18468 50460 18470
rect 50516 18468 50540 18470
rect 50596 18468 50602 18470
rect 50294 18459 50602 18468
rect 50294 17436 50602 17445
rect 50294 17434 50300 17436
rect 50356 17434 50380 17436
rect 50436 17434 50460 17436
rect 50516 17434 50540 17436
rect 50596 17434 50602 17436
rect 50356 17382 50358 17434
rect 50538 17382 50540 17434
rect 50294 17380 50300 17382
rect 50356 17380 50380 17382
rect 50436 17380 50460 17382
rect 50516 17380 50540 17382
rect 50596 17380 50602 17382
rect 50294 17371 50602 17380
rect 49896 16546 50016 16574
rect 49884 15088 49936 15094
rect 49884 15030 49936 15036
rect 49792 14884 49844 14890
rect 49792 14826 49844 14832
rect 49804 14414 49832 14826
rect 49792 14408 49844 14414
rect 49792 14350 49844 14356
rect 49896 14006 49924 15030
rect 49884 14000 49936 14006
rect 49884 13942 49936 13948
rect 49884 13456 49936 13462
rect 49884 13398 49936 13404
rect 49792 13388 49844 13394
rect 49792 13330 49844 13336
rect 49804 13258 49832 13330
rect 49792 13252 49844 13258
rect 49792 13194 49844 13200
rect 49896 12238 49924 13398
rect 49884 12232 49936 12238
rect 49884 12174 49936 12180
rect 49988 3738 50016 16546
rect 50294 16348 50602 16357
rect 50294 16346 50300 16348
rect 50356 16346 50380 16348
rect 50436 16346 50460 16348
rect 50516 16346 50540 16348
rect 50596 16346 50602 16348
rect 50356 16294 50358 16346
rect 50538 16294 50540 16346
rect 50294 16292 50300 16294
rect 50356 16292 50380 16294
rect 50436 16292 50460 16294
rect 50516 16292 50540 16294
rect 50596 16292 50602 16294
rect 50294 16283 50602 16292
rect 50160 16108 50212 16114
rect 50160 16050 50212 16056
rect 50620 16108 50672 16114
rect 50620 16050 50672 16056
rect 50068 15360 50120 15366
rect 50068 15302 50120 15308
rect 50080 15026 50108 15302
rect 50068 15020 50120 15026
rect 50068 14962 50120 14968
rect 50172 14414 50200 16050
rect 50294 15260 50602 15269
rect 50294 15258 50300 15260
rect 50356 15258 50380 15260
rect 50436 15258 50460 15260
rect 50516 15258 50540 15260
rect 50596 15258 50602 15260
rect 50356 15206 50358 15258
rect 50538 15206 50540 15258
rect 50294 15204 50300 15206
rect 50356 15204 50380 15206
rect 50436 15204 50460 15206
rect 50516 15204 50540 15206
rect 50596 15204 50602 15206
rect 50294 15195 50602 15204
rect 50632 15162 50660 16050
rect 50620 15156 50672 15162
rect 50620 15098 50672 15104
rect 50160 14408 50212 14414
rect 50160 14350 50212 14356
rect 50068 14272 50120 14278
rect 50068 14214 50120 14220
rect 50080 13870 50108 14214
rect 50068 13864 50120 13870
rect 50068 13806 50120 13812
rect 50172 13190 50200 14350
rect 50294 14172 50602 14181
rect 50294 14170 50300 14172
rect 50356 14170 50380 14172
rect 50436 14170 50460 14172
rect 50516 14170 50540 14172
rect 50596 14170 50602 14172
rect 50356 14118 50358 14170
rect 50538 14118 50540 14170
rect 50294 14116 50300 14118
rect 50356 14116 50380 14118
rect 50436 14116 50460 14118
rect 50516 14116 50540 14118
rect 50596 14116 50602 14118
rect 50294 14107 50602 14116
rect 50620 13864 50672 13870
rect 50620 13806 50672 13812
rect 50632 13326 50660 13806
rect 50620 13320 50672 13326
rect 50620 13262 50672 13268
rect 50160 13184 50212 13190
rect 50160 13126 50212 13132
rect 50172 12306 50200 13126
rect 50294 13084 50602 13093
rect 50294 13082 50300 13084
rect 50356 13082 50380 13084
rect 50436 13082 50460 13084
rect 50516 13082 50540 13084
rect 50596 13082 50602 13084
rect 50356 13030 50358 13082
rect 50538 13030 50540 13082
rect 50294 13028 50300 13030
rect 50356 13028 50380 13030
rect 50436 13028 50460 13030
rect 50516 13028 50540 13030
rect 50596 13028 50602 13030
rect 50294 13019 50602 13028
rect 50160 12300 50212 12306
rect 50160 12242 50212 12248
rect 50294 11996 50602 12005
rect 50294 11994 50300 11996
rect 50356 11994 50380 11996
rect 50436 11994 50460 11996
rect 50516 11994 50540 11996
rect 50596 11994 50602 11996
rect 50356 11942 50358 11994
rect 50538 11942 50540 11994
rect 50294 11940 50300 11942
rect 50356 11940 50380 11942
rect 50436 11940 50460 11942
rect 50516 11940 50540 11942
rect 50596 11940 50602 11942
rect 50294 11931 50602 11940
rect 50816 11082 50844 33050
rect 50908 27402 50936 42230
rect 51460 33318 51488 57190
rect 50988 33312 51040 33318
rect 50988 33254 51040 33260
rect 51448 33312 51500 33318
rect 51448 33254 51500 33260
rect 50896 27396 50948 27402
rect 50896 27338 50948 27344
rect 51000 18358 51028 33254
rect 51540 29776 51592 29782
rect 51540 29718 51592 29724
rect 51356 27532 51408 27538
rect 51356 27474 51408 27480
rect 51080 22636 51132 22642
rect 51080 22578 51132 22584
rect 51092 22098 51120 22578
rect 51080 22092 51132 22098
rect 51080 22034 51132 22040
rect 51080 20528 51132 20534
rect 51080 20470 51132 20476
rect 51092 19786 51120 20470
rect 51264 20256 51316 20262
rect 51264 20198 51316 20204
rect 51172 20052 51224 20058
rect 51172 19994 51224 20000
rect 51080 19780 51132 19786
rect 51080 19722 51132 19728
rect 51092 18426 51120 19722
rect 51080 18420 51132 18426
rect 51080 18362 51132 18368
rect 50988 18352 51040 18358
rect 50988 18294 51040 18300
rect 51080 17740 51132 17746
rect 51080 17682 51132 17688
rect 51092 17270 51120 17682
rect 51184 17270 51212 19994
rect 51276 19854 51304 20198
rect 51264 19848 51316 19854
rect 51264 19790 51316 19796
rect 51080 17264 51132 17270
rect 51080 17206 51132 17212
rect 51172 17264 51224 17270
rect 51172 17206 51224 17212
rect 51184 16794 51212 17206
rect 51172 16788 51224 16794
rect 51172 16730 51224 16736
rect 50988 16516 51040 16522
rect 50988 16458 51040 16464
rect 51000 15094 51028 16458
rect 51080 16448 51132 16454
rect 51080 16390 51132 16396
rect 51092 16114 51120 16390
rect 51080 16108 51132 16114
rect 51080 16050 51132 16056
rect 51080 15496 51132 15502
rect 51080 15438 51132 15444
rect 50988 15088 51040 15094
rect 50988 15030 51040 15036
rect 50896 15020 50948 15026
rect 50896 14962 50948 14968
rect 50908 14074 50936 14962
rect 50896 14068 50948 14074
rect 50896 14010 50948 14016
rect 50908 13258 50936 14010
rect 51092 13870 51120 15438
rect 51184 15434 51212 16730
rect 51172 15428 51224 15434
rect 51172 15370 51224 15376
rect 51080 13864 51132 13870
rect 51080 13806 51132 13812
rect 50896 13252 50948 13258
rect 50896 13194 50948 13200
rect 50908 12782 50936 13194
rect 50896 12776 50948 12782
rect 50896 12718 50948 12724
rect 50804 11076 50856 11082
rect 50804 11018 50856 11024
rect 50294 10908 50602 10917
rect 50294 10906 50300 10908
rect 50356 10906 50380 10908
rect 50436 10906 50460 10908
rect 50516 10906 50540 10908
rect 50596 10906 50602 10908
rect 50356 10854 50358 10906
rect 50538 10854 50540 10906
rect 50294 10852 50300 10854
rect 50356 10852 50380 10854
rect 50436 10852 50460 10854
rect 50516 10852 50540 10854
rect 50596 10852 50602 10854
rect 50294 10843 50602 10852
rect 50294 9820 50602 9829
rect 50294 9818 50300 9820
rect 50356 9818 50380 9820
rect 50436 9818 50460 9820
rect 50516 9818 50540 9820
rect 50596 9818 50602 9820
rect 50356 9766 50358 9818
rect 50538 9766 50540 9818
rect 50294 9764 50300 9766
rect 50356 9764 50380 9766
rect 50436 9764 50460 9766
rect 50516 9764 50540 9766
rect 50596 9764 50602 9766
rect 50294 9755 50602 9764
rect 50294 8732 50602 8741
rect 50294 8730 50300 8732
rect 50356 8730 50380 8732
rect 50436 8730 50460 8732
rect 50516 8730 50540 8732
rect 50596 8730 50602 8732
rect 50356 8678 50358 8730
rect 50538 8678 50540 8730
rect 50294 8676 50300 8678
rect 50356 8676 50380 8678
rect 50436 8676 50460 8678
rect 50516 8676 50540 8678
rect 50596 8676 50602 8678
rect 50294 8667 50602 8676
rect 50294 7644 50602 7653
rect 50294 7642 50300 7644
rect 50356 7642 50380 7644
rect 50436 7642 50460 7644
rect 50516 7642 50540 7644
rect 50596 7642 50602 7644
rect 50356 7590 50358 7642
rect 50538 7590 50540 7642
rect 50294 7588 50300 7590
rect 50356 7588 50380 7590
rect 50436 7588 50460 7590
rect 50516 7588 50540 7590
rect 50596 7588 50602 7590
rect 50294 7579 50602 7588
rect 50294 6556 50602 6565
rect 50294 6554 50300 6556
rect 50356 6554 50380 6556
rect 50436 6554 50460 6556
rect 50516 6554 50540 6556
rect 50596 6554 50602 6556
rect 50356 6502 50358 6554
rect 50538 6502 50540 6554
rect 50294 6500 50300 6502
rect 50356 6500 50380 6502
rect 50436 6500 50460 6502
rect 50516 6500 50540 6502
rect 50596 6500 50602 6502
rect 50294 6491 50602 6500
rect 50294 5468 50602 5477
rect 50294 5466 50300 5468
rect 50356 5466 50380 5468
rect 50436 5466 50460 5468
rect 50516 5466 50540 5468
rect 50596 5466 50602 5468
rect 50356 5414 50358 5466
rect 50538 5414 50540 5466
rect 50294 5412 50300 5414
rect 50356 5412 50380 5414
rect 50436 5412 50460 5414
rect 50516 5412 50540 5414
rect 50596 5412 50602 5414
rect 50294 5403 50602 5412
rect 50294 4380 50602 4389
rect 50294 4378 50300 4380
rect 50356 4378 50380 4380
rect 50436 4378 50460 4380
rect 50516 4378 50540 4380
rect 50596 4378 50602 4380
rect 50356 4326 50358 4378
rect 50538 4326 50540 4378
rect 50294 4324 50300 4326
rect 50356 4324 50380 4326
rect 50436 4324 50460 4326
rect 50516 4324 50540 4326
rect 50596 4324 50602 4326
rect 50294 4315 50602 4324
rect 51172 4276 51224 4282
rect 51172 4218 51224 4224
rect 50528 4208 50580 4214
rect 50528 4150 50580 4156
rect 50712 4208 50764 4214
rect 50712 4150 50764 4156
rect 50540 3942 50568 4150
rect 50528 3936 50580 3942
rect 50528 3878 50580 3884
rect 50620 3936 50672 3942
rect 50620 3878 50672 3884
rect 49976 3732 50028 3738
rect 49976 3674 50028 3680
rect 50632 3670 50660 3878
rect 50620 3664 50672 3670
rect 50620 3606 50672 3612
rect 49976 3528 50028 3534
rect 50436 3528 50488 3534
rect 49976 3470 50028 3476
rect 50434 3496 50436 3505
rect 50488 3496 50490 3505
rect 49792 3460 49844 3466
rect 49792 3402 49844 3408
rect 49700 2644 49752 2650
rect 49700 2586 49752 2592
rect 49804 800 49832 3402
rect 49882 3360 49938 3369
rect 49882 3295 49938 3304
rect 49896 2854 49924 3295
rect 49884 2848 49936 2854
rect 49884 2790 49936 2796
rect 49884 2372 49936 2378
rect 49884 2314 49936 2320
rect 49896 950 49924 2314
rect 49988 1154 50016 3470
rect 50434 3431 50490 3440
rect 50068 3392 50120 3398
rect 50068 3334 50120 3340
rect 49976 1148 50028 1154
rect 49976 1090 50028 1096
rect 49884 944 49936 950
rect 49884 886 49936 892
rect 50080 800 50108 3334
rect 50294 3292 50602 3301
rect 50294 3290 50300 3292
rect 50356 3290 50380 3292
rect 50436 3290 50460 3292
rect 50516 3290 50540 3292
rect 50596 3290 50602 3292
rect 50356 3238 50358 3290
rect 50538 3238 50540 3290
rect 50294 3236 50300 3238
rect 50356 3236 50380 3238
rect 50436 3236 50460 3238
rect 50516 3236 50540 3238
rect 50596 3236 50602 3238
rect 50294 3227 50602 3236
rect 50294 2204 50602 2213
rect 50294 2202 50300 2204
rect 50356 2202 50380 2204
rect 50436 2202 50460 2204
rect 50516 2202 50540 2204
rect 50596 2202 50602 2204
rect 50356 2150 50358 2202
rect 50538 2150 50540 2202
rect 50294 2148 50300 2150
rect 50356 2148 50380 2150
rect 50436 2148 50460 2150
rect 50516 2148 50540 2150
rect 50596 2148 50602 2150
rect 50294 2139 50602 2148
rect 50724 2122 50752 4150
rect 50804 3052 50856 3058
rect 50804 2994 50856 3000
rect 50632 2094 50752 2122
rect 50344 1284 50396 1290
rect 50344 1226 50396 1232
rect 50356 800 50384 1226
rect 50632 800 50660 2094
rect 50816 814 50844 2994
rect 51080 2440 51132 2446
rect 51080 2382 51132 2388
rect 50896 944 50948 950
rect 50896 886 50948 892
rect 50804 808 50856 814
rect 49424 128 49476 134
rect 49424 70 49476 76
rect 49514 0 49570 800
rect 49790 0 49846 800
rect 50066 0 50122 800
rect 50342 0 50398 800
rect 50618 0 50674 800
rect 50908 800 50936 886
rect 51092 882 51120 2382
rect 51080 876 51132 882
rect 51080 818 51132 824
rect 51184 800 51212 4218
rect 51368 4146 51396 27474
rect 51448 24880 51500 24886
rect 51448 24822 51500 24828
rect 51356 4140 51408 4146
rect 51356 4082 51408 4088
rect 51460 3942 51488 24822
rect 51552 22094 51580 29718
rect 51736 25362 51764 57190
rect 52460 56772 52512 56778
rect 52460 56714 52512 56720
rect 52472 55894 52500 56714
rect 52552 56160 52604 56166
rect 52552 56102 52604 56108
rect 52460 55888 52512 55894
rect 52460 55830 52512 55836
rect 52564 55706 52592 56102
rect 52472 55678 52592 55706
rect 52472 53106 52500 55678
rect 52460 53100 52512 53106
rect 52460 53042 52512 53048
rect 52656 51338 52684 57258
rect 53932 57248 53984 57254
rect 53932 57190 53984 57196
rect 54116 57248 54168 57254
rect 54116 57190 54168 57196
rect 53564 56976 53616 56982
rect 53564 56918 53616 56924
rect 53196 55888 53248 55894
rect 53196 55830 53248 55836
rect 52644 51332 52696 51338
rect 52644 51274 52696 51280
rect 52828 32428 52880 32434
rect 52828 32370 52880 32376
rect 52736 30252 52788 30258
rect 52736 30194 52788 30200
rect 52184 28620 52236 28626
rect 52184 28562 52236 28568
rect 51724 25356 51776 25362
rect 51724 25298 51776 25304
rect 51908 23180 51960 23186
rect 51908 23122 51960 23128
rect 51632 23112 51684 23118
rect 51632 23054 51684 23060
rect 51644 22778 51672 23054
rect 51632 22772 51684 22778
rect 51632 22714 51684 22720
rect 51724 22636 51776 22642
rect 51724 22578 51776 22584
rect 51736 22166 51764 22578
rect 51920 22574 51948 23122
rect 52000 22976 52052 22982
rect 52000 22918 52052 22924
rect 51908 22568 51960 22574
rect 51908 22510 51960 22516
rect 51724 22160 51776 22166
rect 51724 22102 51776 22108
rect 51552 22066 51672 22094
rect 51540 16992 51592 16998
rect 51540 16934 51592 16940
rect 51552 16726 51580 16934
rect 51540 16720 51592 16726
rect 51540 16662 51592 16668
rect 51540 15904 51592 15910
rect 51540 15846 51592 15852
rect 51552 15570 51580 15846
rect 51540 15564 51592 15570
rect 51540 15506 51592 15512
rect 51540 13388 51592 13394
rect 51540 13330 51592 13336
rect 51552 12714 51580 13330
rect 51540 12708 51592 12714
rect 51540 12650 51592 12656
rect 51448 3936 51500 3942
rect 51448 3878 51500 3884
rect 51448 3528 51500 3534
rect 51448 3470 51500 3476
rect 51264 2372 51316 2378
rect 51264 2314 51316 2320
rect 51276 1086 51304 2314
rect 51264 1080 51316 1086
rect 51264 1022 51316 1028
rect 51460 800 51488 3470
rect 51540 3052 51592 3058
rect 51540 2994 51592 3000
rect 51552 1222 51580 2994
rect 51644 2650 51672 22066
rect 52012 21962 52040 22918
rect 52000 21956 52052 21962
rect 52000 21898 52052 21904
rect 52000 20256 52052 20262
rect 52000 20198 52052 20204
rect 51908 19848 51960 19854
rect 51908 19790 51960 19796
rect 51920 19446 51948 19790
rect 51908 19440 51960 19446
rect 51908 19382 51960 19388
rect 51724 17672 51776 17678
rect 51724 17614 51776 17620
rect 51736 17338 51764 17614
rect 51724 17332 51776 17338
rect 51724 17274 51776 17280
rect 51920 16998 51948 19382
rect 52012 19378 52040 20198
rect 52092 19780 52144 19786
rect 52092 19722 52144 19728
rect 52104 19514 52132 19722
rect 52092 19508 52144 19514
rect 52092 19450 52144 19456
rect 52000 19372 52052 19378
rect 52000 19314 52052 19320
rect 52092 19372 52144 19378
rect 52092 19314 52144 19320
rect 52104 19258 52132 19314
rect 52012 19230 52132 19258
rect 52012 17678 52040 19230
rect 52000 17672 52052 17678
rect 52000 17614 52052 17620
rect 51908 16992 51960 16998
rect 51908 16934 51960 16940
rect 51816 16584 51868 16590
rect 51816 16526 51868 16532
rect 51828 16046 51856 16526
rect 51816 16040 51868 16046
rect 51816 15982 51868 15988
rect 51724 14272 51776 14278
rect 51724 14214 51776 14220
rect 51736 13938 51764 14214
rect 51724 13932 51776 13938
rect 51724 13874 51776 13880
rect 51724 13252 51776 13258
rect 51724 13194 51776 13200
rect 51736 12102 51764 13194
rect 51828 12918 51856 15982
rect 51920 15706 51948 16934
rect 51908 15700 51960 15706
rect 51908 15642 51960 15648
rect 51920 15434 51948 15642
rect 51908 15428 51960 15434
rect 51908 15370 51960 15376
rect 52012 14890 52040 17614
rect 52092 17536 52144 17542
rect 52092 17478 52144 17484
rect 52104 16590 52132 17478
rect 52092 16584 52144 16590
rect 52092 16526 52144 16532
rect 52092 15496 52144 15502
rect 52092 15438 52144 15444
rect 52000 14884 52052 14890
rect 52000 14826 52052 14832
rect 51816 12912 51868 12918
rect 51816 12854 51868 12860
rect 51724 12096 51776 12102
rect 51724 12038 51776 12044
rect 51736 11150 51764 12038
rect 51724 11144 51776 11150
rect 51724 11086 51776 11092
rect 52104 9450 52132 15438
rect 52092 9444 52144 9450
rect 52092 9386 52144 9392
rect 52196 3670 52224 28562
rect 52368 22024 52420 22030
rect 52368 21966 52420 21972
rect 52380 21486 52408 21966
rect 52368 21480 52420 21486
rect 52368 21422 52420 21428
rect 52276 20460 52328 20466
rect 52276 20402 52328 20408
rect 52288 19310 52316 20402
rect 52380 19786 52408 21422
rect 52368 19780 52420 19786
rect 52368 19722 52420 19728
rect 52380 19446 52408 19722
rect 52368 19440 52420 19446
rect 52368 19382 52420 19388
rect 52276 19304 52328 19310
rect 52276 19246 52328 19252
rect 52288 18358 52316 19246
rect 52460 18896 52512 18902
rect 52460 18838 52512 18844
rect 52472 18737 52500 18838
rect 52458 18728 52514 18737
rect 52458 18663 52514 18672
rect 52276 18352 52328 18358
rect 52276 18294 52328 18300
rect 52288 18034 52316 18294
rect 52288 18006 52408 18034
rect 52274 17096 52330 17105
rect 52274 17031 52276 17040
rect 52328 17031 52330 17040
rect 52276 17002 52328 17008
rect 52380 16402 52408 18006
rect 52380 16374 52500 16402
rect 52472 16182 52500 16374
rect 52460 16176 52512 16182
rect 52460 16118 52512 16124
rect 52276 4140 52328 4146
rect 52276 4082 52328 4088
rect 52184 3664 52236 3670
rect 52184 3606 52236 3612
rect 52000 3460 52052 3466
rect 52000 3402 52052 3408
rect 51632 2644 51684 2650
rect 51632 2586 51684 2592
rect 51540 1216 51592 1222
rect 51540 1158 51592 1164
rect 51724 1080 51776 1086
rect 51724 1022 51776 1028
rect 51736 800 51764 1022
rect 52012 800 52040 3402
rect 52288 800 52316 4082
rect 52644 3052 52696 3058
rect 52644 2994 52696 3000
rect 52460 2848 52512 2854
rect 52460 2790 52512 2796
rect 52472 2553 52500 2790
rect 52458 2544 52514 2553
rect 52458 2479 52514 2488
rect 52552 1148 52604 1154
rect 52552 1090 52604 1096
rect 52564 800 52592 1090
rect 52656 1018 52684 2994
rect 52748 2650 52776 30194
rect 52840 3194 52868 32370
rect 53208 30326 53236 55830
rect 53576 52018 53604 56918
rect 53840 56228 53892 56234
rect 53840 56170 53892 56176
rect 53564 52012 53616 52018
rect 53564 51954 53616 51960
rect 53852 51270 53880 56170
rect 53840 51264 53892 51270
rect 53840 51206 53892 51212
rect 53288 37936 53340 37942
rect 53288 37878 53340 37884
rect 53196 30320 53248 30326
rect 53196 30262 53248 30268
rect 53300 26874 53328 37878
rect 53944 31754 53972 57190
rect 54128 50998 54156 57190
rect 56232 56704 56284 56710
rect 56232 56646 56284 56652
rect 55220 56296 55272 56302
rect 55220 56238 55272 56244
rect 55232 51066 55260 56238
rect 56048 56160 56100 56166
rect 56048 56102 56100 56108
rect 55956 52624 56008 52630
rect 55956 52566 56008 52572
rect 55220 51060 55272 51066
rect 55220 51002 55272 51008
rect 54116 50992 54168 50998
rect 54116 50934 54168 50940
rect 55864 50856 55916 50862
rect 55864 50798 55916 50804
rect 55876 39030 55904 50798
rect 55968 42090 55996 52566
rect 56060 50454 56088 56102
rect 56048 50448 56100 50454
rect 56048 50390 56100 50396
rect 56140 50176 56192 50182
rect 56140 50118 56192 50124
rect 56048 48544 56100 48550
rect 56048 48486 56100 48492
rect 56060 42158 56088 48486
rect 56152 43790 56180 50118
rect 56140 43784 56192 43790
rect 56140 43726 56192 43732
rect 56048 42152 56100 42158
rect 56048 42094 56100 42100
rect 55956 42084 56008 42090
rect 55956 42026 56008 42032
rect 55864 39024 55916 39030
rect 55864 38966 55916 38972
rect 55956 36168 56008 36174
rect 55956 36110 56008 36116
rect 54576 32496 54628 32502
rect 54576 32438 54628 32444
rect 54484 31952 54536 31958
rect 54484 31894 54536 31900
rect 53944 31726 54064 31754
rect 53208 26846 53328 26874
rect 52920 26444 52972 26450
rect 52920 26386 52972 26392
rect 52932 4078 52960 26386
rect 53104 26376 53156 26382
rect 53104 26318 53156 26324
rect 53116 22658 53144 26318
rect 53024 22642 53144 22658
rect 53012 22636 53144 22642
rect 53064 22630 53144 22636
rect 53012 22578 53064 22584
rect 53012 22500 53064 22506
rect 53012 22442 53064 22448
rect 53024 22098 53052 22442
rect 53116 22234 53144 22630
rect 53104 22228 53156 22234
rect 53104 22170 53156 22176
rect 53012 22092 53064 22098
rect 53012 22034 53064 22040
rect 53104 20596 53156 20602
rect 53104 20538 53156 20544
rect 53116 20330 53144 20538
rect 53012 20324 53064 20330
rect 53012 20266 53064 20272
rect 53104 20324 53156 20330
rect 53104 20266 53156 20272
rect 53024 19378 53052 20266
rect 53012 19372 53064 19378
rect 53012 19314 53064 19320
rect 53012 17332 53064 17338
rect 53012 17274 53064 17280
rect 53024 16726 53052 17274
rect 53012 16720 53064 16726
rect 53012 16662 53064 16668
rect 53208 8566 53236 26846
rect 53380 24064 53432 24070
rect 53380 24006 53432 24012
rect 53288 22432 53340 22438
rect 53288 22374 53340 22380
rect 53300 21622 53328 22374
rect 53288 21616 53340 21622
rect 53288 21558 53340 21564
rect 53196 8560 53248 8566
rect 53196 8502 53248 8508
rect 53392 8362 53420 24006
rect 53748 23044 53800 23050
rect 53748 22986 53800 22992
rect 53840 23044 53892 23050
rect 53840 22986 53892 22992
rect 53760 22778 53788 22986
rect 53748 22772 53800 22778
rect 53748 22714 53800 22720
rect 53748 22092 53800 22098
rect 53748 22034 53800 22040
rect 53564 22024 53616 22030
rect 53564 21966 53616 21972
rect 53576 21690 53604 21966
rect 53760 21962 53788 22034
rect 53748 21956 53800 21962
rect 53748 21898 53800 21904
rect 53564 21684 53616 21690
rect 53564 21626 53616 21632
rect 53852 20482 53880 22986
rect 54036 22098 54064 31726
rect 54300 24268 54352 24274
rect 54300 24210 54352 24216
rect 54116 22636 54168 22642
rect 54116 22578 54168 22584
rect 54128 22234 54156 22578
rect 54116 22228 54168 22234
rect 54116 22170 54168 22176
rect 54024 22092 54076 22098
rect 54024 22034 54076 22040
rect 53932 22024 53984 22030
rect 53932 21966 53984 21972
rect 54208 22024 54260 22030
rect 54208 21966 54260 21972
rect 53944 21298 53972 21966
rect 54024 21956 54076 21962
rect 54024 21898 54076 21904
rect 54036 21690 54064 21898
rect 54024 21684 54076 21690
rect 54024 21626 54076 21632
rect 53944 21270 54064 21298
rect 53484 20454 53696 20482
rect 53852 20466 53972 20482
rect 53484 20398 53512 20454
rect 53472 20392 53524 20398
rect 53472 20334 53524 20340
rect 53564 20392 53616 20398
rect 53564 20334 53616 20340
rect 53472 20256 53524 20262
rect 53472 20198 53524 20204
rect 53484 20058 53512 20198
rect 53472 20052 53524 20058
rect 53472 19994 53524 20000
rect 53576 19922 53604 20334
rect 53668 20058 53696 20454
rect 53840 20460 53972 20466
rect 53892 20454 53972 20460
rect 53840 20402 53892 20408
rect 53656 20052 53708 20058
rect 53656 19994 53708 20000
rect 53944 19990 53972 20454
rect 53932 19984 53984 19990
rect 53932 19926 53984 19932
rect 53564 19916 53616 19922
rect 53564 19858 53616 19864
rect 53576 19514 53604 19858
rect 54036 19718 54064 21270
rect 54116 19848 54168 19854
rect 54116 19790 54168 19796
rect 54024 19712 54076 19718
rect 54024 19654 54076 19660
rect 54128 19514 54156 19790
rect 53564 19508 53616 19514
rect 53564 19450 53616 19456
rect 54116 19508 54168 19514
rect 54116 19450 54168 19456
rect 54220 18766 54248 21966
rect 54208 18760 54260 18766
rect 54208 18702 54260 18708
rect 53472 17196 53524 17202
rect 53472 17138 53524 17144
rect 53484 16794 53512 17138
rect 53472 16788 53524 16794
rect 53472 16730 53524 16736
rect 53656 16448 53708 16454
rect 53656 16390 53708 16396
rect 53668 16250 53696 16390
rect 53656 16244 53708 16250
rect 53656 16186 53708 16192
rect 53564 16176 53616 16182
rect 53564 16118 53616 16124
rect 53576 15994 53604 16118
rect 53484 15966 53604 15994
rect 53484 15910 53512 15966
rect 53472 15904 53524 15910
rect 53472 15846 53524 15852
rect 54208 11756 54260 11762
rect 54208 11698 54260 11704
rect 53380 8356 53432 8362
rect 53380 8298 53432 8304
rect 53656 5772 53708 5778
rect 53656 5714 53708 5720
rect 53472 4480 53524 4486
rect 53472 4422 53524 4428
rect 52920 4072 52972 4078
rect 52920 4014 52972 4020
rect 53484 3738 53512 4422
rect 53472 3732 53524 3738
rect 53472 3674 53524 3680
rect 53668 3670 53696 5714
rect 53746 4176 53802 4185
rect 53746 4111 53802 4120
rect 53760 4078 53788 4111
rect 53748 4072 53800 4078
rect 53748 4014 53800 4020
rect 54220 3738 54248 11698
rect 54208 3732 54260 3738
rect 54208 3674 54260 3680
rect 53656 3664 53708 3670
rect 53656 3606 53708 3612
rect 53104 3528 53156 3534
rect 53104 3470 53156 3476
rect 52828 3188 52880 3194
rect 52828 3130 52880 3136
rect 53012 3052 53064 3058
rect 53012 2994 53064 3000
rect 52736 2644 52788 2650
rect 52736 2586 52788 2592
rect 52644 1012 52696 1018
rect 52644 954 52696 960
rect 52828 1012 52880 1018
rect 52828 954 52880 960
rect 52840 800 52868 954
rect 53024 950 53052 2994
rect 53012 944 53064 950
rect 53012 886 53064 892
rect 53116 800 53144 3470
rect 54312 2514 54340 24210
rect 54392 19848 54444 19854
rect 54392 19790 54444 19796
rect 54404 18154 54432 19790
rect 54392 18148 54444 18154
rect 54392 18090 54444 18096
rect 54496 15502 54524 31894
rect 54484 15496 54536 15502
rect 54484 15438 54536 15444
rect 54496 15026 54524 15438
rect 54484 15020 54536 15026
rect 54484 14962 54536 14968
rect 54588 3194 54616 32438
rect 55220 24200 55272 24206
rect 55220 24142 55272 24148
rect 55232 22506 55260 24142
rect 55404 23112 55456 23118
rect 55404 23054 55456 23060
rect 55416 22574 55444 23054
rect 55404 22568 55456 22574
rect 55404 22510 55456 22516
rect 55220 22500 55272 22506
rect 55220 22442 55272 22448
rect 55416 21554 55444 22510
rect 55772 22024 55824 22030
rect 55772 21966 55824 21972
rect 55680 21956 55732 21962
rect 55680 21898 55732 21904
rect 55692 21690 55720 21898
rect 55680 21684 55732 21690
rect 55680 21626 55732 21632
rect 55404 21548 55456 21554
rect 55404 21490 55456 21496
rect 55496 21548 55548 21554
rect 55496 21490 55548 21496
rect 55218 21040 55274 21049
rect 55218 20975 55274 20984
rect 55232 20534 55260 20975
rect 55220 20528 55272 20534
rect 55220 20470 55272 20476
rect 55416 19922 55444 21490
rect 55508 21146 55536 21490
rect 55496 21140 55548 21146
rect 55496 21082 55548 21088
rect 55784 21010 55812 21966
rect 55864 21888 55916 21894
rect 55864 21830 55916 21836
rect 55876 21690 55904 21830
rect 55864 21684 55916 21690
rect 55864 21626 55916 21632
rect 55772 21004 55824 21010
rect 55772 20946 55824 20952
rect 55680 20460 55732 20466
rect 55680 20402 55732 20408
rect 55404 19916 55456 19922
rect 55404 19858 55456 19864
rect 55692 18970 55720 20402
rect 55784 19378 55812 20946
rect 55876 20942 55904 21626
rect 55864 20936 55916 20942
rect 55864 20878 55916 20884
rect 55876 20466 55904 20878
rect 55864 20460 55916 20466
rect 55864 20402 55916 20408
rect 55772 19372 55824 19378
rect 55772 19314 55824 19320
rect 55864 19372 55916 19378
rect 55864 19314 55916 19320
rect 55680 18964 55732 18970
rect 55680 18906 55732 18912
rect 55680 18828 55732 18834
rect 55680 18770 55732 18776
rect 55692 18290 55720 18770
rect 55680 18284 55732 18290
rect 55680 18226 55732 18232
rect 55404 18148 55456 18154
rect 55404 18090 55456 18096
rect 54944 18080 54996 18086
rect 54944 18022 54996 18028
rect 54668 17128 54720 17134
rect 54668 17070 54720 17076
rect 54680 16590 54708 17070
rect 54668 16584 54720 16590
rect 54668 16526 54720 16532
rect 54680 15094 54708 16526
rect 54956 15094 54984 18022
rect 54668 15088 54720 15094
rect 54668 15030 54720 15036
rect 54944 15088 54996 15094
rect 54944 15030 54996 15036
rect 54956 12238 54984 15030
rect 54944 12232 54996 12238
rect 54944 12174 54996 12180
rect 55312 8356 55364 8362
rect 55312 8298 55364 8304
rect 54668 6384 54720 6390
rect 54668 6326 54720 6332
rect 54680 5846 54708 6326
rect 54760 6112 54812 6118
rect 54760 6054 54812 6060
rect 54668 5840 54720 5846
rect 54668 5782 54720 5788
rect 54772 3924 54800 6054
rect 55220 4208 55272 4214
rect 55220 4150 55272 4156
rect 54852 3936 54904 3942
rect 54772 3896 54852 3924
rect 54772 3534 54800 3896
rect 54852 3878 54904 3884
rect 54760 3528 54812 3534
rect 54760 3470 54812 3476
rect 55232 3233 55260 4150
rect 55218 3224 55274 3233
rect 54576 3188 54628 3194
rect 55324 3194 55352 8298
rect 55416 6730 55444 18090
rect 55784 17814 55812 19314
rect 55876 18426 55904 19314
rect 55864 18420 55916 18426
rect 55864 18362 55916 18368
rect 55772 17808 55824 17814
rect 55772 17750 55824 17756
rect 55968 16658 55996 36110
rect 56244 26246 56272 56646
rect 56704 56438 56732 57258
rect 56796 56846 56824 57938
rect 57244 57248 57296 57254
rect 57244 57190 57296 57196
rect 56784 56840 56836 56846
rect 56784 56782 56836 56788
rect 56692 56432 56744 56438
rect 56692 56374 56744 56380
rect 56600 54528 56652 54534
rect 56600 54470 56652 54476
rect 56612 49842 56640 54470
rect 56600 49836 56652 49842
rect 56600 49778 56652 49784
rect 56692 33992 56744 33998
rect 56692 33934 56744 33940
rect 56704 31754 56732 33934
rect 57256 33114 57284 57190
rect 57428 57044 57480 57050
rect 57428 56986 57480 56992
rect 57440 55758 57468 56986
rect 57624 56846 57652 59200
rect 58990 58712 59046 58721
rect 58990 58647 59046 58656
rect 58714 58304 58770 58313
rect 58714 58239 58770 58248
rect 58256 57248 58308 57254
rect 58256 57190 58308 57196
rect 58268 56982 58296 57190
rect 58256 56976 58308 56982
rect 58256 56918 58308 56924
rect 57612 56840 57664 56846
rect 57612 56782 57664 56788
rect 58728 56506 58756 58239
rect 59004 58002 59032 58647
rect 58992 57996 59044 58002
rect 58992 57938 59044 57944
rect 58990 57896 59046 57905
rect 58990 57831 59046 57840
rect 59004 57526 59032 57831
rect 58992 57520 59044 57526
rect 58806 57488 58862 57497
rect 58992 57462 59044 57468
rect 58806 57423 58862 57432
rect 58900 57452 58952 57458
rect 58820 57322 58848 57423
rect 58900 57394 58952 57400
rect 58808 57316 58860 57322
rect 58808 57258 58860 57264
rect 58716 56500 58768 56506
rect 58716 56442 58768 56448
rect 58164 56364 58216 56370
rect 58164 56306 58216 56312
rect 57428 55752 57480 55758
rect 57428 55694 57480 55700
rect 57520 55616 57572 55622
rect 57520 55558 57572 55564
rect 57532 52494 57560 55558
rect 58176 55457 58204 56306
rect 58912 56273 58940 57394
rect 58990 57080 59046 57089
rect 58990 57015 58992 57024
rect 59044 57015 59046 57024
rect 58992 56986 59044 56992
rect 58992 56908 59044 56914
rect 58992 56850 59044 56856
rect 59004 56681 59032 56850
rect 59452 56772 59504 56778
rect 59452 56714 59504 56720
rect 58990 56672 59046 56681
rect 58990 56607 59046 56616
rect 58992 56432 59044 56438
rect 58992 56374 59044 56380
rect 58898 56264 58954 56273
rect 58898 56199 58954 56208
rect 59004 55865 59032 56374
rect 58990 55856 59046 55865
rect 58990 55791 59046 55800
rect 58992 55752 59044 55758
rect 58992 55694 59044 55700
rect 58162 55448 58218 55457
rect 58162 55383 58218 55392
rect 58808 55276 58860 55282
rect 58808 55218 58860 55224
rect 58256 54528 58308 54534
rect 58256 54470 58308 54476
rect 58164 53508 58216 53514
rect 58164 53450 58216 53456
rect 58176 53009 58204 53450
rect 58162 53000 58218 53009
rect 58162 52935 58218 52944
rect 58072 52896 58124 52902
rect 58072 52838 58124 52844
rect 57520 52488 57572 52494
rect 57520 52430 57572 52436
rect 57980 51808 58032 51814
rect 57980 51750 58032 51756
rect 57520 51264 57572 51270
rect 57520 51206 57572 51212
rect 57336 48000 57388 48006
rect 57336 47942 57388 47948
rect 57348 45014 57376 47942
rect 57428 47456 57480 47462
rect 57428 47398 57480 47404
rect 57336 45008 57388 45014
rect 57336 44950 57388 44956
rect 57336 44736 57388 44742
rect 57336 44678 57388 44684
rect 57348 43654 57376 44678
rect 57336 43648 57388 43654
rect 57336 43590 57388 43596
rect 57440 35222 57468 47398
rect 57532 37874 57560 51206
rect 57992 49314 58020 51750
rect 58084 50862 58112 52838
rect 58164 52624 58216 52630
rect 58164 52566 58216 52572
rect 58176 52426 58204 52566
rect 58268 52562 58296 54470
rect 58820 54233 58848 55218
rect 59004 55049 59032 55694
rect 59084 55412 59136 55418
rect 59084 55354 59136 55360
rect 58990 55040 59046 55049
rect 58990 54975 59046 54984
rect 58992 54664 59044 54670
rect 58990 54632 58992 54641
rect 59044 54632 59046 54641
rect 58900 54596 58952 54602
rect 58990 54567 59046 54576
rect 58900 54538 58952 54544
rect 58806 54224 58862 54233
rect 58806 54159 58862 54168
rect 58532 53984 58584 53990
rect 58532 53926 58584 53932
rect 58440 53508 58492 53514
rect 58440 53450 58492 53456
rect 58256 52556 58308 52562
rect 58256 52498 58308 52504
rect 58164 52420 58216 52426
rect 58164 52362 58216 52368
rect 58256 50924 58308 50930
rect 58256 50866 58308 50872
rect 58072 50856 58124 50862
rect 58072 50798 58124 50804
rect 58072 50720 58124 50726
rect 58072 50662 58124 50668
rect 57900 49286 58020 49314
rect 57900 48822 57928 49286
rect 58084 49178 58112 50662
rect 58164 50244 58216 50250
rect 58164 50186 58216 50192
rect 58176 49745 58204 50186
rect 58268 50153 58296 50866
rect 58348 50380 58400 50386
rect 58348 50322 58400 50328
rect 58254 50144 58310 50153
rect 58254 50079 58310 50088
rect 58162 49736 58218 49745
rect 58162 49671 58218 49680
rect 57980 49156 58032 49162
rect 58084 49150 58204 49178
rect 57980 49098 58032 49104
rect 57992 48929 58020 49098
rect 58072 49088 58124 49094
rect 58072 49030 58124 49036
rect 57978 48920 58034 48929
rect 57978 48855 58034 48864
rect 57888 48816 57940 48822
rect 57888 48758 57940 48764
rect 57888 48340 57940 48346
rect 57888 48282 57940 48288
rect 57900 48142 57928 48282
rect 57888 48136 57940 48142
rect 57888 48078 57940 48084
rect 58084 47274 58112 49030
rect 58176 48278 58204 49150
rect 58164 48272 58216 48278
rect 58164 48214 58216 48220
rect 57992 47246 58112 47274
rect 57992 44010 58020 47246
rect 58164 46572 58216 46578
rect 58164 46514 58216 46520
rect 58072 45892 58124 45898
rect 58072 45834 58124 45840
rect 57900 43982 58020 44010
rect 57900 43450 57928 43982
rect 58084 43874 58112 45834
rect 58176 45665 58204 46514
rect 58256 46368 58308 46374
rect 58256 46310 58308 46316
rect 58162 45656 58218 45665
rect 58162 45591 58218 45600
rect 58164 45484 58216 45490
rect 58164 45426 58216 45432
rect 58176 44441 58204 45426
rect 58268 45370 58296 46310
rect 58360 45490 58388 50322
rect 58452 47734 58480 53450
rect 58440 47728 58492 47734
rect 58440 47670 58492 47676
rect 58440 47456 58492 47462
rect 58440 47398 58492 47404
rect 58348 45484 58400 45490
rect 58348 45426 58400 45432
rect 58268 45342 58388 45370
rect 58256 45280 58308 45286
rect 58256 45222 58308 45228
rect 58162 44432 58218 44441
rect 58162 44367 58218 44376
rect 58268 44282 58296 45222
rect 58360 45082 58388 45342
rect 58348 45076 58400 45082
rect 58348 45018 58400 45024
rect 57992 43846 58112 43874
rect 58176 44254 58296 44282
rect 57888 43444 57940 43450
rect 57888 43386 57940 43392
rect 57520 37868 57572 37874
rect 57520 37810 57572 37816
rect 57520 37256 57572 37262
rect 57520 37198 57572 37204
rect 57428 35216 57480 35222
rect 57428 35158 57480 35164
rect 57244 33108 57296 33114
rect 57244 33050 57296 33056
rect 57060 31816 57112 31822
rect 57060 31758 57112 31764
rect 56704 31726 56824 31754
rect 56324 30592 56376 30598
rect 56324 30534 56376 30540
rect 56232 26240 56284 26246
rect 56232 26182 56284 26188
rect 56336 22642 56364 30534
rect 56600 28552 56652 28558
rect 56600 28494 56652 28500
rect 56416 22976 56468 22982
rect 56416 22918 56468 22924
rect 56428 22658 56456 22918
rect 56324 22636 56376 22642
rect 56428 22630 56548 22658
rect 56324 22578 56376 22584
rect 56416 22568 56468 22574
rect 56416 22510 56468 22516
rect 56324 21956 56376 21962
rect 56324 21898 56376 21904
rect 56232 21548 56284 21554
rect 56232 21490 56284 21496
rect 56140 21480 56192 21486
rect 56140 21422 56192 21428
rect 56152 21010 56180 21422
rect 56140 21004 56192 21010
rect 56140 20946 56192 20952
rect 56046 20904 56102 20913
rect 56046 20839 56048 20848
rect 56100 20839 56102 20848
rect 56048 20810 56100 20816
rect 56048 20256 56100 20262
rect 56048 20198 56100 20204
rect 56060 19854 56088 20198
rect 56244 20058 56272 21490
rect 56336 20874 56364 21898
rect 56324 20868 56376 20874
rect 56324 20810 56376 20816
rect 56336 20466 56364 20810
rect 56428 20806 56456 22510
rect 56416 20800 56468 20806
rect 56416 20742 56468 20748
rect 56324 20460 56376 20466
rect 56324 20402 56376 20408
rect 56336 20262 56364 20402
rect 56428 20369 56456 20742
rect 56414 20360 56470 20369
rect 56414 20295 56416 20304
rect 56468 20295 56470 20304
rect 56416 20266 56468 20272
rect 56324 20256 56376 20262
rect 56324 20198 56376 20204
rect 56232 20052 56284 20058
rect 56232 19994 56284 20000
rect 56048 19848 56100 19854
rect 56048 19790 56100 19796
rect 56140 18896 56192 18902
rect 56140 18838 56192 18844
rect 56048 18760 56100 18766
rect 56048 18702 56100 18708
rect 56060 18426 56088 18702
rect 56048 18420 56100 18426
rect 56048 18362 56100 18368
rect 56060 17134 56088 18362
rect 56152 17202 56180 18838
rect 56336 18766 56364 20198
rect 56428 19394 56456 20266
rect 56520 19514 56548 22630
rect 56612 21622 56640 28494
rect 56796 21894 56824 31726
rect 56876 27464 56928 27470
rect 56876 27406 56928 27412
rect 56784 21888 56836 21894
rect 56784 21830 56836 21836
rect 56600 21616 56652 21622
rect 56600 21558 56652 21564
rect 56796 20942 56824 21830
rect 56784 20936 56836 20942
rect 56784 20878 56836 20884
rect 56508 19508 56560 19514
rect 56508 19450 56560 19456
rect 56600 19508 56652 19514
rect 56600 19450 56652 19456
rect 56428 19366 56548 19394
rect 56324 18760 56376 18766
rect 56324 18702 56376 18708
rect 56416 18352 56468 18358
rect 56416 18294 56468 18300
rect 56428 18154 56456 18294
rect 56416 18148 56468 18154
rect 56416 18090 56468 18096
rect 56428 17678 56456 18090
rect 56416 17672 56468 17678
rect 56416 17614 56468 17620
rect 56140 17196 56192 17202
rect 56140 17138 56192 17144
rect 56048 17128 56100 17134
rect 56048 17070 56100 17076
rect 56046 16688 56102 16697
rect 55956 16652 56008 16658
rect 56046 16623 56048 16632
rect 55956 16594 56008 16600
rect 56100 16623 56102 16632
rect 56048 16594 56100 16600
rect 55968 16250 55996 16594
rect 55956 16244 56008 16250
rect 55956 16186 56008 16192
rect 56152 15638 56180 17138
rect 56232 16992 56284 16998
rect 56232 16934 56284 16940
rect 56244 16590 56272 16934
rect 56232 16584 56284 16590
rect 56232 16526 56284 16532
rect 55864 15632 55916 15638
rect 55864 15574 55916 15580
rect 56140 15632 56192 15638
rect 56140 15574 56192 15580
rect 55876 13326 55904 15574
rect 56048 14884 56100 14890
rect 56048 14826 56100 14832
rect 55864 13320 55916 13326
rect 55864 13262 55916 13268
rect 55772 12912 55824 12918
rect 55586 12880 55642 12889
rect 55876 12900 55904 13262
rect 55956 13252 56008 13258
rect 55956 13194 56008 13200
rect 55824 12872 55904 12900
rect 55772 12854 55824 12860
rect 55586 12815 55588 12824
rect 55640 12815 55642 12824
rect 55588 12786 55640 12792
rect 55784 12306 55812 12854
rect 55864 12708 55916 12714
rect 55864 12650 55916 12656
rect 55772 12300 55824 12306
rect 55772 12242 55824 12248
rect 55496 7404 55548 7410
rect 55496 7346 55548 7352
rect 55772 7404 55824 7410
rect 55772 7346 55824 7352
rect 55404 6724 55456 6730
rect 55404 6666 55456 6672
rect 55416 4622 55444 6666
rect 55404 4616 55456 4622
rect 55404 4558 55456 4564
rect 55508 4554 55536 7346
rect 55680 6316 55732 6322
rect 55680 6258 55732 6264
rect 55692 5574 55720 6258
rect 55784 5914 55812 7346
rect 55772 5908 55824 5914
rect 55772 5850 55824 5856
rect 55680 5568 55732 5574
rect 55680 5510 55732 5516
rect 55692 5234 55720 5510
rect 55680 5228 55732 5234
rect 55680 5170 55732 5176
rect 55496 4548 55548 4554
rect 55496 4490 55548 4496
rect 55508 3534 55536 4490
rect 55496 3528 55548 3534
rect 55496 3470 55548 3476
rect 55218 3159 55274 3168
rect 55312 3188 55364 3194
rect 54576 3130 54628 3136
rect 55312 3130 55364 3136
rect 54392 3052 54444 3058
rect 54392 2994 54444 3000
rect 55220 3052 55272 3058
rect 55220 2994 55272 3000
rect 54300 2508 54352 2514
rect 54300 2450 54352 2456
rect 53932 2440 53984 2446
rect 53932 2382 53984 2388
rect 53656 1216 53708 1222
rect 53656 1158 53708 1164
rect 53380 944 53432 950
rect 53380 886 53432 892
rect 53392 800 53420 886
rect 53668 800 53696 1158
rect 53944 800 53972 2382
rect 54404 1290 54432 2994
rect 54392 1284 54444 1290
rect 54392 1226 54444 1232
rect 55232 1086 55260 2994
rect 55588 2372 55640 2378
rect 55588 2314 55640 2320
rect 55220 1080 55272 1086
rect 55220 1022 55272 1028
rect 55600 950 55628 2314
rect 55876 1193 55904 12650
rect 55968 11830 55996 13194
rect 55956 11824 56008 11830
rect 55956 11766 56008 11772
rect 56060 10674 56088 14826
rect 56416 13932 56468 13938
rect 56416 13874 56468 13880
rect 56232 13864 56284 13870
rect 56232 13806 56284 13812
rect 56140 13252 56192 13258
rect 56140 13194 56192 13200
rect 56152 12850 56180 13194
rect 56140 12844 56192 12850
rect 56140 12786 56192 12792
rect 56244 12434 56272 13806
rect 56428 13530 56456 13874
rect 56416 13524 56468 13530
rect 56416 13466 56468 13472
rect 56520 12850 56548 19366
rect 56612 18698 56640 19450
rect 56784 18760 56836 18766
rect 56690 18728 56746 18737
rect 56600 18692 56652 18698
rect 56784 18702 56836 18708
rect 56690 18663 56746 18672
rect 56600 18634 56652 18640
rect 56704 18358 56732 18663
rect 56692 18352 56744 18358
rect 56692 18294 56744 18300
rect 56692 18080 56744 18086
rect 56692 18022 56744 18028
rect 56704 17542 56732 18022
rect 56692 17536 56744 17542
rect 56692 17478 56744 17484
rect 56796 16794 56824 18702
rect 56888 18340 56916 27406
rect 56968 23248 57020 23254
rect 56968 23190 57020 23196
rect 56980 20942 57008 23190
rect 57072 22098 57100 31758
rect 57152 22228 57204 22234
rect 57152 22170 57204 22176
rect 57060 22092 57112 22098
rect 57060 22034 57112 22040
rect 57164 22030 57192 22170
rect 57152 22024 57204 22030
rect 57152 21966 57204 21972
rect 57428 21956 57480 21962
rect 57428 21898 57480 21904
rect 57440 21690 57468 21898
rect 57428 21684 57480 21690
rect 57428 21626 57480 21632
rect 57428 21548 57480 21554
rect 57428 21490 57480 21496
rect 56968 20936 57020 20942
rect 56968 20878 57020 20884
rect 57440 20602 57468 21490
rect 57532 21350 57560 37198
rect 57992 35766 58020 43846
rect 58072 43784 58124 43790
rect 58072 43726 58124 43732
rect 58084 43625 58112 43726
rect 58070 43616 58126 43625
rect 58070 43551 58126 43560
rect 58072 43444 58124 43450
rect 58072 43386 58124 43392
rect 58084 37942 58112 43386
rect 58176 38486 58204 44254
rect 58256 44192 58308 44198
rect 58256 44134 58308 44140
rect 58164 38480 58216 38486
rect 58164 38422 58216 38428
rect 58072 37936 58124 37942
rect 58072 37878 58124 37884
rect 58070 37088 58126 37097
rect 58070 37023 58126 37032
rect 58084 36786 58112 37023
rect 58072 36780 58124 36786
rect 58072 36722 58124 36728
rect 58162 36272 58218 36281
rect 58162 36207 58164 36216
rect 58216 36207 58218 36216
rect 58164 36178 58216 36184
rect 58162 35864 58218 35873
rect 58162 35799 58218 35808
rect 58176 35766 58204 35799
rect 57980 35760 58032 35766
rect 57980 35702 58032 35708
rect 58164 35760 58216 35766
rect 58164 35702 58216 35708
rect 57612 35080 57664 35086
rect 57612 35022 57664 35028
rect 58162 35048 58218 35057
rect 57624 21434 57652 35022
rect 58162 34983 58164 34992
rect 58216 34983 58218 34992
rect 58164 34954 58216 34960
rect 58070 34640 58126 34649
rect 58070 34575 58072 34584
rect 58124 34575 58126 34584
rect 58072 34546 58124 34552
rect 58164 33924 58216 33930
rect 58164 33866 58216 33872
rect 58176 33833 58204 33866
rect 58162 33824 58218 33833
rect 58162 33759 58218 33768
rect 58072 33516 58124 33522
rect 58072 33458 58124 33464
rect 58084 33425 58112 33458
rect 58070 33416 58126 33425
rect 58070 33351 58126 33360
rect 58164 32836 58216 32842
rect 58164 32778 58216 32784
rect 58176 32609 58204 32778
rect 58162 32600 58218 32609
rect 58162 32535 58218 32544
rect 58072 32428 58124 32434
rect 58072 32370 58124 32376
rect 57980 32224 58032 32230
rect 58084 32201 58112 32370
rect 57980 32166 58032 32172
rect 58070 32192 58126 32201
rect 57704 29640 57756 29646
rect 57704 29582 57756 29588
rect 57716 21554 57744 29582
rect 57888 25288 57940 25294
rect 57888 25230 57940 25236
rect 57796 22092 57848 22098
rect 57796 22034 57848 22040
rect 57704 21548 57756 21554
rect 57704 21490 57756 21496
rect 57624 21406 57744 21434
rect 57520 21344 57572 21350
rect 57520 21286 57572 21292
rect 57612 21344 57664 21350
rect 57612 21286 57664 21292
rect 57428 20596 57480 20602
rect 57428 20538 57480 20544
rect 57532 20466 57560 21286
rect 57520 20460 57572 20466
rect 57520 20402 57572 20408
rect 57624 20097 57652 21286
rect 57610 20088 57666 20097
rect 57610 20023 57666 20032
rect 56968 18352 57020 18358
rect 56888 18312 56968 18340
rect 56888 17882 56916 18312
rect 56968 18294 57020 18300
rect 56876 17876 56928 17882
rect 56876 17818 56928 17824
rect 56784 16788 56836 16794
rect 56784 16730 56836 16736
rect 56876 16652 56928 16658
rect 56876 16594 56928 16600
rect 56888 16114 56916 16594
rect 56876 16108 56928 16114
rect 56876 16050 56928 16056
rect 56600 13728 56652 13734
rect 56600 13670 56652 13676
rect 56612 13326 56640 13670
rect 56784 13388 56836 13394
rect 56888 13376 56916 16050
rect 57060 13932 57112 13938
rect 57060 13874 57112 13880
rect 56836 13348 56916 13376
rect 56784 13330 56836 13336
rect 56600 13320 56652 13326
rect 56600 13262 56652 13268
rect 56416 12844 56468 12850
rect 56416 12786 56468 12792
rect 56508 12844 56560 12850
rect 56508 12786 56560 12792
rect 56152 12406 56272 12434
rect 56152 12170 56180 12406
rect 56140 12164 56192 12170
rect 56140 12106 56192 12112
rect 56152 11694 56180 12106
rect 56140 11688 56192 11694
rect 56140 11630 56192 11636
rect 56048 10668 56100 10674
rect 56048 10610 56100 10616
rect 56060 9994 56088 10610
rect 56048 9988 56100 9994
rect 56048 9930 56100 9936
rect 56060 7478 56088 9930
rect 56048 7472 56100 7478
rect 56048 7414 56100 7420
rect 56048 7200 56100 7206
rect 56048 7142 56100 7148
rect 56060 6322 56088 7142
rect 56048 6316 56100 6322
rect 56048 6258 56100 6264
rect 56152 3058 56180 11630
rect 56428 10606 56456 12786
rect 56508 12640 56560 12646
rect 56508 12582 56560 12588
rect 56520 11762 56548 12582
rect 56600 12436 56652 12442
rect 56600 12378 56652 12384
rect 56508 11756 56560 11762
rect 56508 11698 56560 11704
rect 56612 10674 56640 12378
rect 56796 12306 56824 13330
rect 57072 12918 57100 13874
rect 57716 13530 57744 21406
rect 57808 21146 57836 22034
rect 57796 21140 57848 21146
rect 57796 21082 57848 21088
rect 57900 19514 57928 25230
rect 57992 22710 58020 32166
rect 58070 32127 58126 32136
rect 58268 31754 58296 44134
rect 58346 42392 58402 42401
rect 58346 42327 58402 42336
rect 58360 42226 58388 42327
rect 58348 42220 58400 42226
rect 58348 42162 58400 42168
rect 58346 39944 58402 39953
rect 58346 39879 58348 39888
rect 58400 39879 58402 39888
rect 58348 39850 58400 39856
rect 58348 38752 58400 38758
rect 58346 38720 58348 38729
rect 58400 38720 58402 38729
rect 58346 38655 58402 38664
rect 58452 38570 58480 47398
rect 58544 46510 58572 53926
rect 58912 53825 58940 54538
rect 58992 54188 59044 54194
rect 58992 54130 59044 54136
rect 58898 53816 58954 53825
rect 58898 53751 58954 53760
rect 59004 53417 59032 54130
rect 58990 53408 59046 53417
rect 58990 53343 59046 53352
rect 58900 53100 58952 53106
rect 58900 53042 58952 53048
rect 58912 52193 58940 53042
rect 58990 52592 59046 52601
rect 58990 52527 59046 52536
rect 59004 52494 59032 52527
rect 58992 52488 59044 52494
rect 58992 52430 59044 52436
rect 58898 52184 58954 52193
rect 58898 52119 58954 52128
rect 58992 52080 59044 52086
rect 58992 52022 59044 52028
rect 58808 52012 58860 52018
rect 58808 51954 58860 51960
rect 58716 51264 58768 51270
rect 58716 51206 58768 51212
rect 58624 49768 58676 49774
rect 58624 49710 58676 49716
rect 58532 46504 58584 46510
rect 58532 46446 58584 46452
rect 58532 45484 58584 45490
rect 58532 45426 58584 45432
rect 58544 42294 58572 45426
rect 58532 42288 58584 42294
rect 58532 42230 58584 42236
rect 58532 40928 58584 40934
rect 58532 40870 58584 40876
rect 58360 38542 58480 38570
rect 58360 35154 58388 38542
rect 58440 38480 58492 38486
rect 58440 38422 58492 38428
rect 58348 35148 58400 35154
rect 58348 35090 58400 35096
rect 58268 31726 58388 31754
rect 58072 31340 58124 31346
rect 58072 31282 58124 31288
rect 58084 30977 58112 31282
rect 58256 31136 58308 31142
rect 58256 31078 58308 31084
rect 58070 30968 58126 30977
rect 58268 30938 58296 31078
rect 58070 30903 58126 30912
rect 58256 30932 58308 30938
rect 58256 30874 58308 30880
rect 58164 30660 58216 30666
rect 58164 30602 58216 30608
rect 58176 30569 58204 30602
rect 58162 30560 58218 30569
rect 58162 30495 58218 30504
rect 58072 30252 58124 30258
rect 58072 30194 58124 30200
rect 58084 29753 58112 30194
rect 58162 30152 58218 30161
rect 58162 30087 58218 30096
rect 58070 29744 58126 29753
rect 58176 29714 58204 30087
rect 58070 29679 58126 29688
rect 58164 29708 58216 29714
rect 58164 29650 58216 29656
rect 58070 29336 58126 29345
rect 58070 29271 58126 29280
rect 58084 29170 58112 29271
rect 58360 29238 58388 31726
rect 58452 31414 58480 38422
rect 58544 34202 58572 40870
rect 58532 34196 58584 34202
rect 58532 34138 58584 34144
rect 58440 31408 58492 31414
rect 58440 31350 58492 31356
rect 58636 30734 58664 49710
rect 58728 44742 58756 51206
rect 58820 50969 58848 51954
rect 59004 51785 59032 52022
rect 58990 51776 59046 51785
rect 58990 51711 59046 51720
rect 58992 51400 59044 51406
rect 58990 51368 58992 51377
rect 59044 51368 59046 51377
rect 58900 51332 58952 51338
rect 58990 51303 59046 51312
rect 58900 51274 58952 51280
rect 58806 50960 58862 50969
rect 58806 50895 58862 50904
rect 58912 50561 58940 51274
rect 58898 50552 58954 50561
rect 58898 50487 58954 50496
rect 59096 50386 59124 55354
rect 59084 50380 59136 50386
rect 59084 50322 59136 50328
rect 58992 49836 59044 49842
rect 58992 49778 59044 49784
rect 59004 49337 59032 49778
rect 58990 49328 59046 49337
rect 58990 49263 59046 49272
rect 58808 48748 58860 48754
rect 58808 48690 58860 48696
rect 58820 47705 58848 48690
rect 58990 48512 59046 48521
rect 58990 48447 59046 48456
rect 59004 48346 59032 48447
rect 58992 48340 59044 48346
rect 58992 48282 59044 48288
rect 58992 48136 59044 48142
rect 58990 48104 58992 48113
rect 59044 48104 59046 48113
rect 58990 48039 59046 48048
rect 59084 48068 59136 48074
rect 59084 48010 59136 48016
rect 58806 47696 58862 47705
rect 58806 47631 58862 47640
rect 58900 47660 58952 47666
rect 58900 47602 58952 47608
rect 58808 47184 58860 47190
rect 58808 47126 58860 47132
rect 58716 44736 58768 44742
rect 58716 44678 58768 44684
rect 58716 43648 58768 43654
rect 58716 43590 58768 43596
rect 58624 30728 58676 30734
rect 58624 30670 58676 30676
rect 58348 29232 58400 29238
rect 58348 29174 58400 29180
rect 58072 29164 58124 29170
rect 58072 29106 58124 29112
rect 58440 29028 58492 29034
rect 58440 28970 58492 28976
rect 58162 28928 58218 28937
rect 58162 28863 58218 28872
rect 58176 28626 58204 28863
rect 58164 28620 58216 28626
rect 58164 28562 58216 28568
rect 58070 28520 58126 28529
rect 58070 28455 58126 28464
rect 58084 28082 58112 28455
rect 58072 28076 58124 28082
rect 58072 28018 58124 28024
rect 58162 27296 58218 27305
rect 58162 27231 58218 27240
rect 58176 27062 58204 27231
rect 58164 27056 58216 27062
rect 58164 26998 58216 27004
rect 58162 26480 58218 26489
rect 58162 26415 58164 26424
rect 58216 26415 58218 26424
rect 58164 26386 58216 26392
rect 58162 26072 58218 26081
rect 58162 26007 58218 26016
rect 58176 25974 58204 26007
rect 58164 25968 58216 25974
rect 58164 25910 58216 25916
rect 58162 25256 58218 25265
rect 58162 25191 58164 25200
rect 58216 25191 58218 25200
rect 58164 25162 58216 25168
rect 58070 24848 58126 24857
rect 58070 24783 58072 24792
rect 58124 24783 58126 24792
rect 58072 24754 58124 24760
rect 58164 24132 58216 24138
rect 58164 24074 58216 24080
rect 58176 24041 58204 24074
rect 58162 24032 58218 24041
rect 58162 23967 58218 23976
rect 58072 23724 58124 23730
rect 58072 23666 58124 23672
rect 58084 23633 58112 23666
rect 58070 23624 58126 23633
rect 58070 23559 58126 23568
rect 58256 23180 58308 23186
rect 58256 23122 58308 23128
rect 58164 23044 58216 23050
rect 58164 22986 58216 22992
rect 58176 22817 58204 22986
rect 58162 22808 58218 22817
rect 58162 22743 58218 22752
rect 57980 22704 58032 22710
rect 57980 22646 58032 22652
rect 58072 22636 58124 22642
rect 58072 22578 58124 22584
rect 58084 22409 58112 22578
rect 58070 22400 58126 22409
rect 58070 22335 58126 22344
rect 58268 22234 58296 23122
rect 58256 22228 58308 22234
rect 58256 22170 58308 22176
rect 58072 21548 58124 21554
rect 58072 21490 58124 21496
rect 58084 21185 58112 21490
rect 58070 21176 58126 21185
rect 58070 21111 58126 21120
rect 58164 20460 58216 20466
rect 58164 20402 58216 20408
rect 57980 20256 58032 20262
rect 57980 20198 58032 20204
rect 57992 19961 58020 20198
rect 58176 19961 58204 20402
rect 58254 20360 58310 20369
rect 58254 20295 58310 20304
rect 57978 19952 58034 19961
rect 57978 19887 58034 19896
rect 58162 19952 58218 19961
rect 58268 19922 58296 20295
rect 58162 19887 58218 19896
rect 58256 19916 58308 19922
rect 58256 19858 58308 19864
rect 57888 19508 57940 19514
rect 57888 19450 57940 19456
rect 58162 19136 58218 19145
rect 58162 19071 58218 19080
rect 58176 18834 58204 19071
rect 58164 18828 58216 18834
rect 58164 18770 58216 18776
rect 58162 17504 58218 17513
rect 58162 17439 58218 17448
rect 58176 17270 58204 17439
rect 58164 17264 58216 17270
rect 58164 17206 58216 17212
rect 58256 17196 58308 17202
rect 58256 17138 58308 17144
rect 58268 16794 58296 17138
rect 58256 16788 58308 16794
rect 58256 16730 58308 16736
rect 58162 16280 58218 16289
rect 58162 16215 58218 16224
rect 58176 16182 58204 16215
rect 58164 16176 58216 16182
rect 58164 16118 58216 16124
rect 58162 15464 58218 15473
rect 58162 15399 58164 15408
rect 58216 15399 58218 15408
rect 58164 15370 58216 15376
rect 58070 15056 58126 15065
rect 58070 14991 58072 15000
rect 58124 14991 58126 15000
rect 58072 14962 58124 14968
rect 58256 14816 58308 14822
rect 58256 14758 58308 14764
rect 58164 14340 58216 14346
rect 58164 14282 58216 14288
rect 58176 14249 58204 14282
rect 58162 14240 58218 14249
rect 58162 14175 58218 14184
rect 58268 14006 58296 14758
rect 58256 14000 58308 14006
rect 58162 13968 58218 13977
rect 58072 13932 58124 13938
rect 58256 13942 58308 13948
rect 58162 13903 58218 13912
rect 58072 13874 58124 13880
rect 58084 13841 58112 13874
rect 58070 13832 58126 13841
rect 58176 13802 58204 13903
rect 58070 13767 58126 13776
rect 58164 13796 58216 13802
rect 58164 13738 58216 13744
rect 57704 13524 57756 13530
rect 57704 13466 57756 13472
rect 57716 13258 57744 13466
rect 57704 13252 57756 13258
rect 57704 13194 57756 13200
rect 57152 13184 57204 13190
rect 57152 13126 57204 13132
rect 57164 12918 57192 13126
rect 57060 12912 57112 12918
rect 57060 12854 57112 12860
rect 57152 12912 57204 12918
rect 57152 12854 57204 12860
rect 57072 12442 57100 12854
rect 58072 12844 58124 12850
rect 58072 12786 58124 12792
rect 58084 12617 58112 12786
rect 58070 12608 58126 12617
rect 58070 12543 58126 12552
rect 57060 12436 57112 12442
rect 57060 12378 57112 12384
rect 56784 12300 56836 12306
rect 56784 12242 56836 12248
rect 56692 12164 56744 12170
rect 56692 12106 56744 12112
rect 56704 11898 56732 12106
rect 56692 11892 56744 11898
rect 56692 11834 56744 11840
rect 56508 10668 56560 10674
rect 56508 10610 56560 10616
rect 56600 10668 56652 10674
rect 56600 10610 56652 10616
rect 56416 10600 56468 10606
rect 56416 10542 56468 10548
rect 56324 10056 56376 10062
rect 56324 9998 56376 10004
rect 56232 9920 56284 9926
rect 56232 9862 56284 9868
rect 56244 9722 56272 9862
rect 56232 9716 56284 9722
rect 56232 9658 56284 9664
rect 56336 9382 56364 9998
rect 56428 9586 56456 10542
rect 56520 10538 56548 10610
rect 56508 10532 56560 10538
rect 56508 10474 56560 10480
rect 56692 10192 56744 10198
rect 56692 10134 56744 10140
rect 56416 9580 56468 9586
rect 56416 9522 56468 9528
rect 56324 9376 56376 9382
rect 56324 9318 56376 9324
rect 56428 7886 56456 9522
rect 56704 8974 56732 10134
rect 56796 10130 56824 12242
rect 58162 11792 58218 11801
rect 58072 11756 58124 11762
rect 58162 11727 58218 11736
rect 58072 11698 58124 11704
rect 58084 11393 58112 11698
rect 58070 11384 58126 11393
rect 58070 11319 58126 11328
rect 58176 11218 58204 11727
rect 58164 11212 58216 11218
rect 58164 11154 58216 11160
rect 57060 10668 57112 10674
rect 57060 10610 57112 10616
rect 58256 10668 58308 10674
rect 58256 10610 58308 10616
rect 56876 10464 56928 10470
rect 56876 10406 56928 10412
rect 56784 10124 56836 10130
rect 56784 10066 56836 10072
rect 56796 9042 56824 10066
rect 56888 10062 56916 10406
rect 57072 10266 57100 10610
rect 57888 10600 57940 10606
rect 57940 10548 58020 10554
rect 57888 10542 58020 10548
rect 57900 10526 58020 10542
rect 57992 10470 58020 10526
rect 57980 10464 58032 10470
rect 57980 10406 58032 10412
rect 58268 10266 58296 10610
rect 57060 10260 57112 10266
rect 57060 10202 57112 10208
rect 58256 10260 58308 10266
rect 58256 10202 58308 10208
rect 56876 10056 56928 10062
rect 56876 9998 56928 10004
rect 57060 9580 57112 9586
rect 57060 9522 57112 9528
rect 57072 9178 57100 9522
rect 57060 9172 57112 9178
rect 57060 9114 57112 9120
rect 56784 9036 56836 9042
rect 56784 8978 56836 8984
rect 56692 8968 56744 8974
rect 56692 8910 56744 8916
rect 56600 8288 56652 8294
rect 56600 8230 56652 8236
rect 56416 7880 56468 7886
rect 56416 7822 56468 7828
rect 56324 7472 56376 7478
rect 56324 7414 56376 7420
rect 56336 6322 56364 7414
rect 56324 6316 56376 6322
rect 56324 6258 56376 6264
rect 56428 6118 56456 7822
rect 56508 7744 56560 7750
rect 56508 7686 56560 7692
rect 56520 7546 56548 7686
rect 56508 7540 56560 7546
rect 56508 7482 56560 7488
rect 56612 7410 56640 8230
rect 56600 7404 56652 7410
rect 56600 7346 56652 7352
rect 56796 6798 56824 8978
rect 58070 8936 58126 8945
rect 58070 8871 58126 8880
rect 58084 8498 58112 8871
rect 58072 8492 58124 8498
rect 58072 8434 58124 8440
rect 58162 8120 58218 8129
rect 58162 8055 58218 8064
rect 58176 7954 58204 8055
rect 57980 7948 58032 7954
rect 57980 7890 58032 7896
rect 58164 7948 58216 7954
rect 58164 7890 58216 7896
rect 57992 7410 58020 7890
rect 58070 7712 58126 7721
rect 58070 7647 58126 7656
rect 58084 7410 58112 7647
rect 57980 7404 58032 7410
rect 57980 7346 58032 7352
rect 58072 7404 58124 7410
rect 58072 7346 58124 7352
rect 56968 7200 57020 7206
rect 56968 7142 57020 7148
rect 56980 6798 57008 7142
rect 57992 7002 58020 7346
rect 58254 7304 58310 7313
rect 58254 7239 58256 7248
rect 58308 7239 58310 7248
rect 58256 7210 58308 7216
rect 57980 6996 58032 7002
rect 57980 6938 58032 6944
rect 56784 6792 56836 6798
rect 56784 6734 56836 6740
rect 56968 6792 57020 6798
rect 56968 6734 57020 6740
rect 56796 6390 56824 6734
rect 56784 6384 56836 6390
rect 56784 6326 56836 6332
rect 56416 6112 56468 6118
rect 56416 6054 56468 6060
rect 56428 5778 56456 6054
rect 56796 5778 56824 6326
rect 57152 6248 57204 6254
rect 57152 6190 57204 6196
rect 57060 6112 57112 6118
rect 57060 6054 57112 6060
rect 56416 5772 56468 5778
rect 56416 5714 56468 5720
rect 56784 5772 56836 5778
rect 56784 5714 56836 5720
rect 56796 4690 56824 5714
rect 56876 5704 56928 5710
rect 57072 5658 57100 6054
rect 56928 5652 57100 5658
rect 56876 5646 57100 5652
rect 56888 5630 57100 5646
rect 57164 5642 57192 6190
rect 58072 6112 58124 6118
rect 58072 6054 58124 6060
rect 58084 5710 58112 6054
rect 58452 5914 58480 28970
rect 58728 28150 58756 43590
rect 58820 40934 58848 47126
rect 58912 46889 58940 47602
rect 58992 47592 59044 47598
rect 58992 47534 59044 47540
rect 59004 47297 59032 47534
rect 58990 47288 59046 47297
rect 58990 47223 59046 47232
rect 58992 47048 59044 47054
rect 58992 46990 59044 46996
rect 58898 46880 58954 46889
rect 58898 46815 58954 46824
rect 59004 46481 59032 46990
rect 58990 46472 59046 46481
rect 58990 46407 59046 46416
rect 58990 46064 59046 46073
rect 58990 45999 59046 46008
rect 59004 45966 59032 45999
rect 58992 45960 59044 45966
rect 58992 45902 59044 45908
rect 58990 45248 59046 45257
rect 58990 45183 59046 45192
rect 58900 44940 58952 44946
rect 58900 44882 58952 44888
rect 58912 44849 58940 44882
rect 59004 44878 59032 45183
rect 58992 44872 59044 44878
rect 58898 44840 58954 44849
rect 58992 44814 59044 44820
rect 58898 44775 58954 44784
rect 58992 44396 59044 44402
rect 58992 44338 59044 44344
rect 59004 44033 59032 44338
rect 58990 44024 59046 44033
rect 58990 43959 59046 43968
rect 58992 43308 59044 43314
rect 58992 43250 59044 43256
rect 58898 43208 58954 43217
rect 58898 43143 58954 43152
rect 58912 42702 58940 43143
rect 59004 42809 59032 43250
rect 58990 42800 59046 42809
rect 58990 42735 59046 42744
rect 58900 42696 58952 42702
rect 58900 42638 58952 42644
rect 58900 42560 58952 42566
rect 58900 42502 58952 42508
rect 58808 40928 58860 40934
rect 58808 40870 58860 40876
rect 58808 40724 58860 40730
rect 58808 40666 58860 40672
rect 58716 28144 58768 28150
rect 58716 28086 58768 28092
rect 58820 12434 58848 40666
rect 58912 35894 58940 42502
rect 58992 41608 59044 41614
rect 58992 41550 59044 41556
rect 59004 41177 59032 41550
rect 58990 41168 59046 41177
rect 58990 41103 59046 41112
rect 59096 40730 59124 48010
rect 59268 44804 59320 44810
rect 59268 44746 59320 44752
rect 59176 43104 59228 43110
rect 59176 43046 59228 43052
rect 59084 40724 59136 40730
rect 59084 40666 59136 40672
rect 59188 39522 59216 43046
rect 59096 39494 59216 39522
rect 58990 37496 59046 37505
rect 58990 37431 59046 37440
rect 59004 37262 59032 37431
rect 58992 37256 59044 37262
rect 58992 37198 59044 37204
rect 58912 35866 59032 35894
rect 59004 34898 59032 35866
rect 59096 35018 59124 39494
rect 59084 35012 59136 35018
rect 59084 34954 59136 34960
rect 59004 34870 59216 34898
rect 59084 34740 59136 34746
rect 59084 34682 59136 34688
rect 58900 31884 58952 31890
rect 58900 31826 58952 31832
rect 58912 31385 58940 31826
rect 58992 31816 59044 31822
rect 58990 31784 58992 31793
rect 59044 31784 59046 31793
rect 58990 31719 59046 31728
rect 58898 31376 58954 31385
rect 58898 31311 58954 31320
rect 58990 27704 59046 27713
rect 58990 27639 59046 27648
rect 59004 27538 59032 27639
rect 58992 27532 59044 27538
rect 58992 27474 59044 27480
rect 59096 26874 59124 34682
rect 59188 27130 59216 34870
rect 59280 32774 59308 44746
rect 59360 35012 59412 35018
rect 59360 34954 59412 34960
rect 59268 32768 59320 32774
rect 59268 32710 59320 32716
rect 59176 27124 59228 27130
rect 59176 27066 59228 27072
rect 58728 12406 58848 12434
rect 58912 26846 59124 26874
rect 58728 8537 58756 12406
rect 58912 11234 58940 26846
rect 59372 26586 59400 34954
rect 59360 26580 59412 26586
rect 59360 26522 59412 26528
rect 58992 22976 59044 22982
rect 58992 22918 59044 22924
rect 59004 21593 59032 22918
rect 58990 21584 59046 21593
rect 58990 21519 59046 21528
rect 58992 19372 59044 19378
rect 58992 19314 59044 19320
rect 59004 18737 59032 19314
rect 58990 18728 59046 18737
rect 58990 18663 59046 18672
rect 58992 18624 59044 18630
rect 58992 18566 59044 18572
rect 59004 17921 59032 18566
rect 58990 17912 59046 17921
rect 58990 17847 59046 17856
rect 59464 17678 59492 56714
rect 59544 36576 59596 36582
rect 59544 36518 59596 36524
rect 59452 17672 59504 17678
rect 59452 17614 59504 17620
rect 58992 17128 59044 17134
rect 58992 17070 59044 17076
rect 59004 16697 59032 17070
rect 58990 16688 59046 16697
rect 58990 16623 59046 16632
rect 59084 16176 59136 16182
rect 59082 16144 59084 16153
rect 59136 16144 59138 16153
rect 59082 16079 59138 16088
rect 59556 14618 59584 36518
rect 59728 35556 59780 35562
rect 59728 35498 59780 35504
rect 59636 33312 59688 33318
rect 59636 33254 59688 33260
rect 59544 14612 59596 14618
rect 59544 14554 59596 14560
rect 58992 13864 59044 13870
rect 58992 13806 59044 13812
rect 59004 13025 59032 13806
rect 58990 13016 59046 13025
rect 58990 12951 59046 12960
rect 58820 11206 58940 11234
rect 58820 9654 58848 11206
rect 58900 11076 58952 11082
rect 58900 11018 58952 11024
rect 58912 10169 58940 11018
rect 59648 10810 59676 33254
rect 59740 16182 59768 35498
rect 59728 16176 59780 16182
rect 59728 16118 59780 16124
rect 59636 10804 59688 10810
rect 59636 10746 59688 10752
rect 58990 10568 59046 10577
rect 58990 10503 59046 10512
rect 59004 10470 59032 10503
rect 58992 10464 59044 10470
rect 58992 10406 59044 10412
rect 58898 10160 58954 10169
rect 58898 10095 58954 10104
rect 58808 9648 58860 9654
rect 58808 9590 58860 9596
rect 58992 9512 59044 9518
rect 58992 9454 59044 9460
rect 59004 9353 59032 9454
rect 58990 9344 59046 9353
rect 58990 9279 59046 9288
rect 58714 8528 58770 8537
rect 58714 8463 58770 8472
rect 58992 7336 59044 7342
rect 58992 7278 59044 7284
rect 59004 6905 59032 7278
rect 58990 6896 59046 6905
rect 58990 6831 59046 6840
rect 58992 6724 59044 6730
rect 58992 6666 59044 6672
rect 59004 6497 59032 6666
rect 58990 6488 59046 6497
rect 58990 6423 59046 6432
rect 58440 5908 58492 5914
rect 58440 5850 58492 5856
rect 58072 5704 58124 5710
rect 58072 5646 58124 5652
rect 58990 5672 59046 5681
rect 57072 5234 57100 5630
rect 57152 5636 57204 5642
rect 57152 5578 57204 5584
rect 57336 5636 57388 5642
rect 58990 5607 58992 5616
rect 57336 5578 57388 5584
rect 59044 5607 59046 5616
rect 58992 5578 59044 5584
rect 57348 5302 57376 5578
rect 57336 5296 57388 5302
rect 57336 5238 57388 5244
rect 58070 5264 58126 5273
rect 57060 5228 57112 5234
rect 58070 5199 58072 5208
rect 57060 5170 57112 5176
rect 58124 5199 58126 5208
rect 58072 5170 58124 5176
rect 58992 5160 59044 5166
rect 58992 5102 59044 5108
rect 57336 5092 57388 5098
rect 57336 5034 57388 5040
rect 56416 4684 56468 4690
rect 56416 4626 56468 4632
rect 56784 4684 56836 4690
rect 56784 4626 56836 4632
rect 56324 4616 56376 4622
rect 56324 4558 56376 4564
rect 56336 4078 56364 4558
rect 56324 4072 56376 4078
rect 56324 4014 56376 4020
rect 56428 3534 56456 4626
rect 56968 4548 57020 4554
rect 56968 4490 57020 4496
rect 56876 4140 56928 4146
rect 56876 4082 56928 4088
rect 56416 3528 56468 3534
rect 56416 3470 56468 3476
rect 56888 3466 56916 4082
rect 56876 3460 56928 3466
rect 56876 3402 56928 3408
rect 56784 3392 56836 3398
rect 56784 3334 56836 3340
rect 56796 3058 56824 3334
rect 55956 3052 56008 3058
rect 55956 2994 56008 3000
rect 56140 3052 56192 3058
rect 56140 2994 56192 3000
rect 56784 3052 56836 3058
rect 56784 2994 56836 3000
rect 55862 1184 55918 1193
rect 55968 1154 55996 2994
rect 56048 2848 56100 2854
rect 56048 2790 56100 2796
rect 56060 2106 56088 2790
rect 56888 2582 56916 3402
rect 56980 3194 57008 4490
rect 57348 4146 57376 5034
rect 58900 5024 58952 5030
rect 58900 4966 58952 4972
rect 58256 4480 58308 4486
rect 58256 4422 58308 4428
rect 57336 4140 57388 4146
rect 57336 4082 57388 4088
rect 58072 4140 58124 4146
rect 58072 4082 58124 4088
rect 57348 3602 57376 4082
rect 58084 4049 58112 4082
rect 58070 4040 58126 4049
rect 58070 3975 58126 3984
rect 57336 3596 57388 3602
rect 57336 3538 57388 3544
rect 56968 3188 57020 3194
rect 56968 3130 57020 3136
rect 56968 3052 57020 3058
rect 56968 2994 57020 3000
rect 56876 2576 56928 2582
rect 56876 2518 56928 2524
rect 56048 2100 56100 2106
rect 56048 2042 56100 2048
rect 56980 1222 57008 2994
rect 58268 2582 58296 4422
rect 58808 4208 58860 4214
rect 58808 4150 58860 4156
rect 58348 3120 58400 3126
rect 58348 3062 58400 3068
rect 58360 2582 58388 3062
rect 58256 2576 58308 2582
rect 58256 2518 58308 2524
rect 58348 2576 58400 2582
rect 58348 2518 58400 2524
rect 57336 2372 57388 2378
rect 57336 2314 57388 2320
rect 56968 1216 57020 1222
rect 56968 1158 57020 1164
rect 55862 1119 55918 1128
rect 55956 1148 56008 1154
rect 55956 1090 56008 1096
rect 57348 1018 57376 2314
rect 58820 1601 58848 4150
rect 58912 2825 58940 4966
rect 59004 4457 59032 5102
rect 58990 4448 59046 4457
rect 58990 4383 59046 4392
rect 58898 2816 58954 2825
rect 58898 2751 58954 2760
rect 58900 2508 58952 2514
rect 58900 2450 58952 2456
rect 58912 2009 58940 2450
rect 58992 2440 59044 2446
rect 58990 2408 58992 2417
rect 59044 2408 59046 2417
rect 58990 2343 59046 2352
rect 58898 2000 58954 2009
rect 58898 1935 58954 1944
rect 58806 1592 58862 1601
rect 58806 1527 58862 1536
rect 57336 1012 57388 1018
rect 57336 954 57388 960
rect 55588 944 55640 950
rect 55588 886 55640 892
rect 50804 750 50856 756
rect 50894 0 50950 800
rect 51170 0 51226 800
rect 51446 0 51502 800
rect 51722 0 51778 800
rect 51998 0 52054 800
rect 52274 0 52330 800
rect 52550 0 52606 800
rect 52826 0 52882 800
rect 53102 0 53158 800
rect 53378 0 53434 800
rect 53654 0 53710 800
rect 53930 0 53986 800
<< via2 >>
rect 19580 57690 19636 57692
rect 19660 57690 19716 57692
rect 19740 57690 19796 57692
rect 19820 57690 19876 57692
rect 19580 57638 19626 57690
rect 19626 57638 19636 57690
rect 19660 57638 19690 57690
rect 19690 57638 19702 57690
rect 19702 57638 19716 57690
rect 19740 57638 19754 57690
rect 19754 57638 19766 57690
rect 19766 57638 19796 57690
rect 19820 57638 19830 57690
rect 19830 57638 19876 57690
rect 19580 57636 19636 57638
rect 19660 57636 19716 57638
rect 19740 57636 19796 57638
rect 19820 57636 19876 57638
rect 50300 57690 50356 57692
rect 50380 57690 50436 57692
rect 50460 57690 50516 57692
rect 50540 57690 50596 57692
rect 50300 57638 50346 57690
rect 50346 57638 50356 57690
rect 50380 57638 50410 57690
rect 50410 57638 50422 57690
rect 50422 57638 50436 57690
rect 50460 57638 50474 57690
rect 50474 57638 50486 57690
rect 50486 57638 50516 57690
rect 50540 57638 50550 57690
rect 50550 57638 50596 57690
rect 50300 57636 50356 57638
rect 50380 57636 50436 57638
rect 50460 57636 50516 57638
rect 50540 57636 50596 57638
rect 938 55800 994 55856
rect 938 55256 994 55312
rect 1030 54712 1086 54768
rect 938 54168 994 54224
rect 1030 53624 1086 53680
rect 938 53080 994 53136
rect 1030 52536 1086 52592
rect 938 51992 994 52048
rect 1030 51448 1086 51504
rect 938 50904 994 50960
rect 1030 50360 1086 50416
rect 938 49816 994 49872
rect 1030 49272 1086 49328
rect 938 48728 994 48784
rect 1030 48184 1086 48240
rect 938 47640 994 47696
rect 1030 47096 1086 47152
rect 938 46552 994 46608
rect 1030 46008 1086 46064
rect 938 45464 994 45520
rect 1030 44920 1086 44976
rect 938 44376 994 44432
rect 1030 43832 1086 43888
rect 938 43288 994 43344
rect 1030 42744 1086 42800
rect 938 42200 994 42256
rect 1030 41656 1086 41712
rect 938 41112 994 41168
rect 1030 40568 1086 40624
rect 938 40024 994 40080
rect 1030 39480 1086 39536
rect 938 38936 994 38992
rect 1030 38392 1086 38448
rect 938 37848 994 37904
rect 1030 37304 1086 37360
rect 938 36760 994 36816
rect 1030 36216 1086 36272
rect 938 35672 994 35728
rect 1030 35128 1086 35184
rect 938 34584 994 34640
rect 1030 34040 1086 34096
rect 938 33496 994 33552
rect 1030 32952 1086 33008
rect 938 32408 994 32464
rect 938 31864 994 31920
rect 1030 31320 1086 31376
rect 938 30776 994 30832
rect 938 30268 940 30288
rect 940 30268 992 30288
rect 992 30268 994 30288
rect 938 30232 994 30268
rect 938 29688 994 29744
rect 1030 29144 1086 29200
rect 938 28600 994 28656
rect 938 28092 940 28112
rect 940 28092 992 28112
rect 992 28092 994 28112
rect 938 28056 994 28092
rect 938 27512 994 27568
rect 938 27004 940 27024
rect 940 27004 992 27024
rect 992 27004 994 27024
rect 938 26968 994 27004
rect 1030 26424 1086 26480
rect 938 25880 994 25936
rect 938 25336 994 25392
rect 938 24792 994 24848
rect 938 24248 994 24304
rect 938 23704 994 23760
rect 938 23160 994 23216
rect 938 22616 994 22672
rect 938 22092 994 22128
rect 938 22072 940 22092
rect 940 22072 992 22092
rect 992 22072 994 22092
rect 938 21528 994 21584
rect 938 21004 994 21040
rect 938 20984 940 21004
rect 940 20984 992 21004
rect 992 20984 994 21004
rect 938 20440 994 20496
rect 938 19916 994 19952
rect 938 19896 940 19916
rect 940 19896 992 19916
rect 992 19896 994 19916
rect 938 19352 994 19408
rect 1030 18808 1086 18864
rect 938 18264 994 18320
rect 938 17720 994 17776
rect 4220 57146 4276 57148
rect 4300 57146 4356 57148
rect 4380 57146 4436 57148
rect 4460 57146 4516 57148
rect 4220 57094 4266 57146
rect 4266 57094 4276 57146
rect 4300 57094 4330 57146
rect 4330 57094 4342 57146
rect 4342 57094 4356 57146
rect 4380 57094 4394 57146
rect 4394 57094 4406 57146
rect 4406 57094 4436 57146
rect 4460 57094 4470 57146
rect 4470 57094 4516 57146
rect 4220 57092 4276 57094
rect 4300 57092 4356 57094
rect 4380 57092 4436 57094
rect 4460 57092 4516 57094
rect 4220 56058 4276 56060
rect 4300 56058 4356 56060
rect 4380 56058 4436 56060
rect 4460 56058 4516 56060
rect 4220 56006 4266 56058
rect 4266 56006 4276 56058
rect 4300 56006 4330 56058
rect 4330 56006 4342 56058
rect 4342 56006 4356 56058
rect 4380 56006 4394 56058
rect 4394 56006 4406 56058
rect 4406 56006 4436 56058
rect 4460 56006 4470 56058
rect 4470 56006 4516 56058
rect 4220 56004 4276 56006
rect 4300 56004 4356 56006
rect 4380 56004 4436 56006
rect 4460 56004 4516 56006
rect 4220 54970 4276 54972
rect 4300 54970 4356 54972
rect 4380 54970 4436 54972
rect 4460 54970 4516 54972
rect 4220 54918 4266 54970
rect 4266 54918 4276 54970
rect 4300 54918 4330 54970
rect 4330 54918 4342 54970
rect 4342 54918 4356 54970
rect 4380 54918 4394 54970
rect 4394 54918 4406 54970
rect 4406 54918 4436 54970
rect 4460 54918 4470 54970
rect 4470 54918 4516 54970
rect 4220 54916 4276 54918
rect 4300 54916 4356 54918
rect 4380 54916 4436 54918
rect 4460 54916 4516 54918
rect 4220 53882 4276 53884
rect 4300 53882 4356 53884
rect 4380 53882 4436 53884
rect 4460 53882 4516 53884
rect 4220 53830 4266 53882
rect 4266 53830 4276 53882
rect 4300 53830 4330 53882
rect 4330 53830 4342 53882
rect 4342 53830 4356 53882
rect 4380 53830 4394 53882
rect 4394 53830 4406 53882
rect 4406 53830 4436 53882
rect 4460 53830 4470 53882
rect 4470 53830 4516 53882
rect 4220 53828 4276 53830
rect 4300 53828 4356 53830
rect 4380 53828 4436 53830
rect 4460 53828 4516 53830
rect 4220 52794 4276 52796
rect 4300 52794 4356 52796
rect 4380 52794 4436 52796
rect 4460 52794 4516 52796
rect 4220 52742 4266 52794
rect 4266 52742 4276 52794
rect 4300 52742 4330 52794
rect 4330 52742 4342 52794
rect 4342 52742 4356 52794
rect 4380 52742 4394 52794
rect 4394 52742 4406 52794
rect 4406 52742 4436 52794
rect 4460 52742 4470 52794
rect 4470 52742 4516 52794
rect 4220 52740 4276 52742
rect 4300 52740 4356 52742
rect 4380 52740 4436 52742
rect 4460 52740 4516 52742
rect 4220 51706 4276 51708
rect 4300 51706 4356 51708
rect 4380 51706 4436 51708
rect 4460 51706 4516 51708
rect 4220 51654 4266 51706
rect 4266 51654 4276 51706
rect 4300 51654 4330 51706
rect 4330 51654 4342 51706
rect 4342 51654 4356 51706
rect 4380 51654 4394 51706
rect 4394 51654 4406 51706
rect 4406 51654 4436 51706
rect 4460 51654 4470 51706
rect 4470 51654 4516 51706
rect 4220 51652 4276 51654
rect 4300 51652 4356 51654
rect 4380 51652 4436 51654
rect 4460 51652 4516 51654
rect 4220 50618 4276 50620
rect 4300 50618 4356 50620
rect 4380 50618 4436 50620
rect 4460 50618 4516 50620
rect 4220 50566 4266 50618
rect 4266 50566 4276 50618
rect 4300 50566 4330 50618
rect 4330 50566 4342 50618
rect 4342 50566 4356 50618
rect 4380 50566 4394 50618
rect 4394 50566 4406 50618
rect 4406 50566 4436 50618
rect 4460 50566 4470 50618
rect 4470 50566 4516 50618
rect 4220 50564 4276 50566
rect 4300 50564 4356 50566
rect 4380 50564 4436 50566
rect 4460 50564 4516 50566
rect 4220 49530 4276 49532
rect 4300 49530 4356 49532
rect 4380 49530 4436 49532
rect 4460 49530 4516 49532
rect 4220 49478 4266 49530
rect 4266 49478 4276 49530
rect 4300 49478 4330 49530
rect 4330 49478 4342 49530
rect 4342 49478 4356 49530
rect 4380 49478 4394 49530
rect 4394 49478 4406 49530
rect 4406 49478 4436 49530
rect 4460 49478 4470 49530
rect 4470 49478 4516 49530
rect 4220 49476 4276 49478
rect 4300 49476 4356 49478
rect 4380 49476 4436 49478
rect 4460 49476 4516 49478
rect 4220 48442 4276 48444
rect 4300 48442 4356 48444
rect 4380 48442 4436 48444
rect 4460 48442 4516 48444
rect 4220 48390 4266 48442
rect 4266 48390 4276 48442
rect 4300 48390 4330 48442
rect 4330 48390 4342 48442
rect 4342 48390 4356 48442
rect 4380 48390 4394 48442
rect 4394 48390 4406 48442
rect 4406 48390 4436 48442
rect 4460 48390 4470 48442
rect 4470 48390 4516 48442
rect 4220 48388 4276 48390
rect 4300 48388 4356 48390
rect 4380 48388 4436 48390
rect 4460 48388 4516 48390
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 938 17176 994 17232
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 938 16632 994 16688
rect 938 16088 994 16144
rect 938 15544 994 15600
rect 938 15000 994 15056
rect 938 14456 994 14512
rect 938 13912 994 13968
rect 938 13368 994 13424
rect 938 12824 994 12880
rect 938 12280 994 12336
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 938 11736 994 11792
rect 938 11192 994 11248
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 938 10648 994 10704
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 938 10104 994 10160
rect 938 9560 994 9616
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 938 9016 994 9072
rect 938 8472 994 8528
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 938 7928 994 7984
rect 938 7384 994 7440
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 938 6840 994 6896
rect 938 6296 994 6352
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 938 5752 994 5808
rect 938 5208 994 5264
rect 938 4664 994 4720
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 938 4120 994 4176
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 9494 5752 9550 5808
rect 12438 13232 12494 13288
rect 10046 4020 10048 4040
rect 10048 4020 10100 4040
rect 10100 4020 10102 4040
rect 10046 3984 10102 4020
rect 12622 10124 12678 10160
rect 12622 10104 12624 10124
rect 12624 10104 12676 10124
rect 12676 10104 12678 10124
rect 11702 7384 11758 7440
rect 14554 11212 14610 11248
rect 14554 11192 14556 11212
rect 14556 11192 14608 11212
rect 14608 11192 14610 11212
rect 19580 56602 19636 56604
rect 19660 56602 19716 56604
rect 19740 56602 19796 56604
rect 19820 56602 19876 56604
rect 19580 56550 19626 56602
rect 19626 56550 19636 56602
rect 19660 56550 19690 56602
rect 19690 56550 19702 56602
rect 19702 56550 19716 56602
rect 19740 56550 19754 56602
rect 19754 56550 19766 56602
rect 19766 56550 19796 56602
rect 19820 56550 19830 56602
rect 19830 56550 19876 56602
rect 19580 56548 19636 56550
rect 19660 56548 19716 56550
rect 19740 56548 19796 56550
rect 19820 56548 19876 56550
rect 15842 15564 15898 15600
rect 15842 15544 15844 15564
rect 15844 15544 15896 15564
rect 15896 15544 15898 15564
rect 16762 3460 16818 3496
rect 16762 3440 16764 3460
rect 16764 3440 16816 3460
rect 16816 3440 16818 3460
rect 17958 3068 17960 3088
rect 17960 3068 18012 3088
rect 18012 3068 18014 3088
rect 17958 3032 18014 3068
rect 19580 55514 19636 55516
rect 19660 55514 19716 55516
rect 19740 55514 19796 55516
rect 19820 55514 19876 55516
rect 19580 55462 19626 55514
rect 19626 55462 19636 55514
rect 19660 55462 19690 55514
rect 19690 55462 19702 55514
rect 19702 55462 19716 55514
rect 19740 55462 19754 55514
rect 19754 55462 19766 55514
rect 19766 55462 19796 55514
rect 19820 55462 19830 55514
rect 19830 55462 19876 55514
rect 19580 55460 19636 55462
rect 19660 55460 19716 55462
rect 19740 55460 19796 55462
rect 19820 55460 19876 55462
rect 19580 54426 19636 54428
rect 19660 54426 19716 54428
rect 19740 54426 19796 54428
rect 19820 54426 19876 54428
rect 19580 54374 19626 54426
rect 19626 54374 19636 54426
rect 19660 54374 19690 54426
rect 19690 54374 19702 54426
rect 19702 54374 19716 54426
rect 19740 54374 19754 54426
rect 19754 54374 19766 54426
rect 19766 54374 19796 54426
rect 19820 54374 19830 54426
rect 19830 54374 19876 54426
rect 19580 54372 19636 54374
rect 19660 54372 19716 54374
rect 19740 54372 19796 54374
rect 19820 54372 19876 54374
rect 19580 53338 19636 53340
rect 19660 53338 19716 53340
rect 19740 53338 19796 53340
rect 19820 53338 19876 53340
rect 19580 53286 19626 53338
rect 19626 53286 19636 53338
rect 19660 53286 19690 53338
rect 19690 53286 19702 53338
rect 19702 53286 19716 53338
rect 19740 53286 19754 53338
rect 19754 53286 19766 53338
rect 19766 53286 19796 53338
rect 19820 53286 19830 53338
rect 19830 53286 19876 53338
rect 19580 53284 19636 53286
rect 19660 53284 19716 53286
rect 19740 53284 19796 53286
rect 19820 53284 19876 53286
rect 19580 52250 19636 52252
rect 19660 52250 19716 52252
rect 19740 52250 19796 52252
rect 19820 52250 19876 52252
rect 19580 52198 19626 52250
rect 19626 52198 19636 52250
rect 19660 52198 19690 52250
rect 19690 52198 19702 52250
rect 19702 52198 19716 52250
rect 19740 52198 19754 52250
rect 19754 52198 19766 52250
rect 19766 52198 19796 52250
rect 19820 52198 19830 52250
rect 19830 52198 19876 52250
rect 19580 52196 19636 52198
rect 19660 52196 19716 52198
rect 19740 52196 19796 52198
rect 19820 52196 19876 52198
rect 19580 51162 19636 51164
rect 19660 51162 19716 51164
rect 19740 51162 19796 51164
rect 19820 51162 19876 51164
rect 19580 51110 19626 51162
rect 19626 51110 19636 51162
rect 19660 51110 19690 51162
rect 19690 51110 19702 51162
rect 19702 51110 19716 51162
rect 19740 51110 19754 51162
rect 19754 51110 19766 51162
rect 19766 51110 19796 51162
rect 19820 51110 19830 51162
rect 19830 51110 19876 51162
rect 19580 51108 19636 51110
rect 19660 51108 19716 51110
rect 19740 51108 19796 51110
rect 19820 51108 19876 51110
rect 19580 50074 19636 50076
rect 19660 50074 19716 50076
rect 19740 50074 19796 50076
rect 19820 50074 19876 50076
rect 19580 50022 19626 50074
rect 19626 50022 19636 50074
rect 19660 50022 19690 50074
rect 19690 50022 19702 50074
rect 19702 50022 19716 50074
rect 19740 50022 19754 50074
rect 19754 50022 19766 50074
rect 19766 50022 19796 50074
rect 19820 50022 19830 50074
rect 19830 50022 19876 50074
rect 19580 50020 19636 50022
rect 19660 50020 19716 50022
rect 19740 50020 19796 50022
rect 19820 50020 19876 50022
rect 19580 48986 19636 48988
rect 19660 48986 19716 48988
rect 19740 48986 19796 48988
rect 19820 48986 19876 48988
rect 19580 48934 19626 48986
rect 19626 48934 19636 48986
rect 19660 48934 19690 48986
rect 19690 48934 19702 48986
rect 19702 48934 19716 48986
rect 19740 48934 19754 48986
rect 19754 48934 19766 48986
rect 19766 48934 19796 48986
rect 19820 48934 19830 48986
rect 19830 48934 19876 48986
rect 19580 48932 19636 48934
rect 19660 48932 19716 48934
rect 19740 48932 19796 48934
rect 19820 48932 19876 48934
rect 19580 47898 19636 47900
rect 19660 47898 19716 47900
rect 19740 47898 19796 47900
rect 19820 47898 19876 47900
rect 19580 47846 19626 47898
rect 19626 47846 19636 47898
rect 19660 47846 19690 47898
rect 19690 47846 19702 47898
rect 19702 47846 19716 47898
rect 19740 47846 19754 47898
rect 19754 47846 19766 47898
rect 19766 47846 19796 47898
rect 19820 47846 19830 47898
rect 19830 47846 19876 47898
rect 19580 47844 19636 47846
rect 19660 47844 19716 47846
rect 19740 47844 19796 47846
rect 19820 47844 19876 47846
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 22282 29996 22284 30016
rect 22284 29996 22336 30016
rect 22336 29996 22338 30016
rect 22282 29960 22338 29996
rect 22282 29300 22338 29336
rect 22282 29280 22284 29300
rect 22284 29280 22336 29300
rect 22336 29280 22338 29300
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 23570 29280 23626 29336
rect 23202 29008 23258 29064
rect 23662 29008 23718 29064
rect 23018 26988 23074 27024
rect 23018 26968 23020 26988
rect 23020 26968 23072 26988
rect 23072 26968 23074 26988
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19798 5228 19854 5264
rect 19798 5208 19800 5228
rect 19800 5208 19852 5228
rect 19852 5208 19854 5228
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19890 4120 19946 4176
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 20166 15816 20222 15872
rect 20718 12144 20774 12200
rect 23294 21936 23350 21992
rect 21914 17312 21970 17368
rect 20994 6432 21050 6488
rect 20718 3984 20774 4040
rect 20902 4428 20904 4448
rect 20904 4428 20956 4448
rect 20956 4428 20958 4448
rect 20902 4392 20958 4428
rect 21822 13096 21878 13152
rect 22742 11600 22798 11656
rect 22098 10648 22154 10704
rect 22006 10512 22062 10568
rect 22098 9424 22154 9480
rect 23202 15700 23258 15736
rect 23202 15680 23204 15700
rect 23204 15680 23256 15700
rect 23256 15680 23258 15700
rect 23202 14456 23258 14512
rect 23018 9016 23074 9072
rect 23662 20984 23718 21040
rect 26054 27124 26110 27160
rect 26054 27104 26056 27124
rect 26056 27104 26108 27124
rect 26108 27104 26110 27124
rect 26422 26968 26478 27024
rect 23386 14864 23442 14920
rect 23294 12280 23350 12336
rect 23478 12008 23534 12064
rect 22006 4700 22008 4720
rect 22008 4700 22060 4720
rect 22060 4700 22062 4720
rect 22006 4664 22062 4700
rect 22558 4428 22560 4448
rect 22560 4428 22612 4448
rect 22612 4428 22614 4448
rect 22558 4392 22614 4428
rect 22558 4140 22614 4176
rect 22558 4120 22560 4140
rect 22560 4120 22612 4140
rect 22612 4120 22614 4140
rect 22558 3032 22614 3088
rect 22650 2896 22706 2952
rect 22834 3168 22890 3224
rect 23110 3304 23166 3360
rect 24490 17176 24546 17232
rect 24674 15136 24730 15192
rect 24214 8880 24270 8936
rect 23570 2896 23626 2952
rect 24950 14456 25006 14512
rect 26330 9424 26386 9480
rect 26974 27412 26976 27432
rect 26976 27412 27028 27432
rect 27028 27412 27030 27432
rect 26974 27376 27030 27412
rect 27618 32408 27674 32464
rect 27802 32272 27858 32328
rect 26882 18128 26938 18184
rect 25226 6332 25228 6352
rect 25228 6332 25280 6352
rect 25280 6332 25282 6352
rect 25226 6296 25282 6332
rect 25686 6196 25688 6216
rect 25688 6196 25740 6216
rect 25740 6196 25742 6216
rect 25686 6160 25742 6196
rect 25594 4700 25596 4720
rect 25596 4700 25648 4720
rect 25648 4700 25650 4720
rect 25594 4664 25650 4700
rect 24950 3576 25006 3632
rect 26790 11600 26846 11656
rect 25686 3304 25742 3360
rect 25226 2388 25228 2408
rect 25228 2388 25280 2408
rect 25280 2388 25282 2408
rect 25226 2352 25282 2388
rect 26974 9152 27030 9208
rect 27158 12280 27214 12336
rect 27250 9424 27306 9480
rect 28078 32136 28134 32192
rect 28446 32272 28502 32328
rect 28446 29960 28502 30016
rect 28630 32172 28632 32192
rect 28632 32172 28684 32192
rect 28684 32172 28686 32192
rect 28630 32136 28686 32172
rect 28722 29688 28778 29744
rect 28446 27412 28448 27432
rect 28448 27412 28500 27432
rect 28500 27412 28502 27432
rect 28446 27376 28502 27412
rect 27802 19760 27858 19816
rect 27710 10376 27766 10432
rect 28630 27104 28686 27160
rect 29090 24132 29146 24168
rect 29090 24112 29092 24132
rect 29092 24112 29144 24132
rect 29144 24112 29146 24132
rect 28538 19624 28594 19680
rect 28814 19780 28870 19816
rect 28814 19760 28816 19780
rect 28816 19760 28868 19780
rect 28868 19760 28870 19780
rect 27802 9424 27858 9480
rect 27618 8336 27674 8392
rect 28906 19624 28962 19680
rect 28722 15680 28778 15736
rect 29550 32000 29606 32056
rect 29642 28056 29698 28112
rect 30470 35980 30472 36000
rect 30472 35980 30524 36000
rect 30524 35980 30526 36000
rect 30470 35944 30526 35980
rect 30746 34584 30802 34640
rect 29918 28056 29974 28112
rect 28814 13912 28870 13968
rect 28630 11056 28686 11112
rect 28354 9832 28410 9888
rect 28630 10376 28686 10432
rect 28538 9444 28594 9480
rect 28538 9424 28540 9444
rect 28540 9424 28592 9444
rect 28592 9424 28594 9444
rect 28538 8472 28594 8528
rect 27802 6196 27804 6216
rect 27804 6196 27856 6216
rect 27856 6196 27858 6216
rect 27802 6160 27858 6196
rect 27618 5616 27674 5672
rect 27894 5208 27950 5264
rect 27526 3848 27582 3904
rect 28354 7248 28410 7304
rect 29090 13776 29146 13832
rect 29090 12960 29146 13016
rect 28998 11328 29054 11384
rect 28814 8472 28870 8528
rect 29090 6704 29146 6760
rect 28998 6180 29054 6216
rect 28998 6160 29000 6180
rect 29000 6160 29052 6180
rect 29052 6160 29054 6180
rect 28262 4528 28318 4584
rect 28906 3476 28908 3496
rect 28908 3476 28960 3496
rect 28960 3476 28962 3496
rect 28906 3440 28962 3476
rect 29734 21548 29790 21584
rect 29734 21528 29736 21548
rect 29736 21528 29788 21548
rect 29788 21528 29790 21548
rect 30562 27004 30564 27024
rect 30564 27004 30616 27024
rect 30616 27004 30618 27024
rect 30562 26968 30618 27004
rect 32678 45484 32734 45520
rect 32678 45464 32680 45484
rect 32680 45464 32732 45484
rect 32732 45464 32734 45484
rect 31114 28056 31170 28112
rect 30286 24148 30288 24168
rect 30288 24148 30340 24168
rect 30340 24148 30342 24168
rect 30286 24112 30342 24148
rect 30286 21392 30342 21448
rect 30470 21800 30526 21856
rect 29550 14764 29552 14784
rect 29552 14764 29604 14784
rect 29604 14764 29606 14784
rect 29550 14728 29606 14764
rect 30102 13368 30158 13424
rect 30378 15000 30434 15056
rect 29826 10920 29882 10976
rect 29826 8608 29882 8664
rect 29918 8472 29974 8528
rect 30470 9288 30526 9344
rect 30286 6568 30342 6624
rect 31390 21528 31446 21584
rect 30930 12008 30986 12064
rect 30746 11328 30802 11384
rect 30746 9632 30802 9688
rect 30930 9424 30986 9480
rect 30838 9288 30894 9344
rect 30930 7520 30986 7576
rect 31666 26444 31722 26480
rect 31666 26424 31668 26444
rect 31668 26424 31720 26444
rect 31720 26424 31722 26444
rect 31758 17040 31814 17096
rect 34940 57146 34996 57148
rect 35020 57146 35076 57148
rect 35100 57146 35156 57148
rect 35180 57146 35236 57148
rect 34940 57094 34986 57146
rect 34986 57094 34996 57146
rect 35020 57094 35050 57146
rect 35050 57094 35062 57146
rect 35062 57094 35076 57146
rect 35100 57094 35114 57146
rect 35114 57094 35126 57146
rect 35126 57094 35156 57146
rect 35180 57094 35190 57146
rect 35190 57094 35236 57146
rect 34940 57092 34996 57094
rect 35020 57092 35076 57094
rect 35100 57092 35156 57094
rect 35180 57092 35236 57094
rect 34940 56058 34996 56060
rect 35020 56058 35076 56060
rect 35100 56058 35156 56060
rect 35180 56058 35236 56060
rect 34940 56006 34986 56058
rect 34986 56006 34996 56058
rect 35020 56006 35050 56058
rect 35050 56006 35062 56058
rect 35062 56006 35076 56058
rect 35100 56006 35114 56058
rect 35114 56006 35126 56058
rect 35126 56006 35156 56058
rect 35180 56006 35190 56058
rect 35190 56006 35236 56058
rect 34940 56004 34996 56006
rect 35020 56004 35076 56006
rect 35100 56004 35156 56006
rect 35180 56004 35236 56006
rect 34940 54970 34996 54972
rect 35020 54970 35076 54972
rect 35100 54970 35156 54972
rect 35180 54970 35236 54972
rect 34940 54918 34986 54970
rect 34986 54918 34996 54970
rect 35020 54918 35050 54970
rect 35050 54918 35062 54970
rect 35062 54918 35076 54970
rect 35100 54918 35114 54970
rect 35114 54918 35126 54970
rect 35126 54918 35156 54970
rect 35180 54918 35190 54970
rect 35190 54918 35236 54970
rect 34940 54916 34996 54918
rect 35020 54916 35076 54918
rect 35100 54916 35156 54918
rect 35180 54916 35236 54918
rect 34940 53882 34996 53884
rect 35020 53882 35076 53884
rect 35100 53882 35156 53884
rect 35180 53882 35236 53884
rect 34940 53830 34986 53882
rect 34986 53830 34996 53882
rect 35020 53830 35050 53882
rect 35050 53830 35062 53882
rect 35062 53830 35076 53882
rect 35100 53830 35114 53882
rect 35114 53830 35126 53882
rect 35126 53830 35156 53882
rect 35180 53830 35190 53882
rect 35190 53830 35236 53882
rect 34940 53828 34996 53830
rect 35020 53828 35076 53830
rect 35100 53828 35156 53830
rect 35180 53828 35236 53830
rect 34940 52794 34996 52796
rect 35020 52794 35076 52796
rect 35100 52794 35156 52796
rect 35180 52794 35236 52796
rect 34940 52742 34986 52794
rect 34986 52742 34996 52794
rect 35020 52742 35050 52794
rect 35050 52742 35062 52794
rect 35062 52742 35076 52794
rect 35100 52742 35114 52794
rect 35114 52742 35126 52794
rect 35126 52742 35156 52794
rect 35180 52742 35190 52794
rect 35190 52742 35236 52794
rect 34940 52740 34996 52742
rect 35020 52740 35076 52742
rect 35100 52740 35156 52742
rect 35180 52740 35236 52742
rect 34940 51706 34996 51708
rect 35020 51706 35076 51708
rect 35100 51706 35156 51708
rect 35180 51706 35236 51708
rect 34940 51654 34986 51706
rect 34986 51654 34996 51706
rect 35020 51654 35050 51706
rect 35050 51654 35062 51706
rect 35062 51654 35076 51706
rect 35100 51654 35114 51706
rect 35114 51654 35126 51706
rect 35126 51654 35156 51706
rect 35180 51654 35190 51706
rect 35190 51654 35236 51706
rect 34940 51652 34996 51654
rect 35020 51652 35076 51654
rect 35100 51652 35156 51654
rect 35180 51652 35236 51654
rect 34940 50618 34996 50620
rect 35020 50618 35076 50620
rect 35100 50618 35156 50620
rect 35180 50618 35236 50620
rect 34940 50566 34986 50618
rect 34986 50566 34996 50618
rect 35020 50566 35050 50618
rect 35050 50566 35062 50618
rect 35062 50566 35076 50618
rect 35100 50566 35114 50618
rect 35114 50566 35126 50618
rect 35126 50566 35156 50618
rect 35180 50566 35190 50618
rect 35190 50566 35236 50618
rect 34940 50564 34996 50566
rect 35020 50564 35076 50566
rect 35100 50564 35156 50566
rect 35180 50564 35236 50566
rect 34940 49530 34996 49532
rect 35020 49530 35076 49532
rect 35100 49530 35156 49532
rect 35180 49530 35236 49532
rect 34940 49478 34986 49530
rect 34986 49478 34996 49530
rect 35020 49478 35050 49530
rect 35050 49478 35062 49530
rect 35062 49478 35076 49530
rect 35100 49478 35114 49530
rect 35114 49478 35126 49530
rect 35126 49478 35156 49530
rect 35180 49478 35190 49530
rect 35190 49478 35236 49530
rect 34940 49476 34996 49478
rect 35020 49476 35076 49478
rect 35100 49476 35156 49478
rect 35180 49476 35236 49478
rect 34940 48442 34996 48444
rect 35020 48442 35076 48444
rect 35100 48442 35156 48444
rect 35180 48442 35236 48444
rect 34940 48390 34986 48442
rect 34986 48390 34996 48442
rect 35020 48390 35050 48442
rect 35050 48390 35062 48442
rect 35062 48390 35076 48442
rect 35100 48390 35114 48442
rect 35114 48390 35126 48442
rect 35126 48390 35156 48442
rect 35180 48390 35190 48442
rect 35190 48390 35236 48442
rect 34940 48388 34996 48390
rect 35020 48388 35076 48390
rect 35100 48388 35156 48390
rect 35180 48388 35236 48390
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 31850 13640 31906 13696
rect 31298 9560 31354 9616
rect 32034 27004 32036 27024
rect 32036 27004 32088 27024
rect 32088 27004 32090 27024
rect 32034 26968 32090 27004
rect 33138 26424 33194 26480
rect 32310 24112 32366 24168
rect 31298 8744 31354 8800
rect 30930 7112 30986 7168
rect 31574 9288 31630 9344
rect 31482 9172 31538 9208
rect 31482 9152 31484 9172
rect 31484 9152 31536 9172
rect 31536 9152 31538 9172
rect 31482 8744 31538 8800
rect 31942 7928 31998 7984
rect 31298 3984 31354 4040
rect 32218 17040 32274 17096
rect 31022 3032 31078 3088
rect 32862 14728 32918 14784
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 35346 36488 35402 36544
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 33322 13368 33378 13424
rect 33230 13096 33286 13152
rect 32402 8472 32458 8528
rect 32954 10920 33010 10976
rect 33138 10920 33194 10976
rect 33322 9560 33378 9616
rect 33046 9016 33102 9072
rect 33230 6296 33286 6352
rect 32862 3460 32918 3496
rect 32862 3440 32864 3460
rect 32864 3440 32916 3460
rect 32916 3440 32918 3460
rect 33782 26288 33838 26344
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 36818 31764 36820 31784
rect 36820 31764 36872 31784
rect 36872 31764 36874 31784
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 36818 31728 36874 31764
rect 36542 29008 36598 29064
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 33690 10920 33746 10976
rect 33874 11056 33930 11112
rect 33690 8508 33692 8528
rect 33692 8508 33744 8528
rect 33744 8508 33746 8528
rect 33690 8472 33746 8508
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34426 20596 34482 20632
rect 34426 20576 34428 20596
rect 34428 20576 34480 20596
rect 34480 20576 34482 20596
rect 35254 20460 35310 20496
rect 35254 20440 35256 20460
rect 35256 20440 35308 20460
rect 35308 20440 35310 20460
rect 34702 19896 34758 19952
rect 34426 19624 34482 19680
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34242 15816 34298 15872
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34058 13368 34114 13424
rect 34426 13776 34482 13832
rect 34242 11600 34298 11656
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 35530 17040 35586 17096
rect 36082 19760 36138 19816
rect 35806 17584 35862 17640
rect 36082 17448 36138 17504
rect 35898 17076 35900 17096
rect 35900 17076 35952 17096
rect 35952 17076 35954 17096
rect 35898 17040 35954 17076
rect 37002 21392 37058 21448
rect 36818 19488 36874 19544
rect 36450 17448 36506 17504
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34702 9832 34758 9888
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 35898 13368 35954 13424
rect 36082 13232 36138 13288
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34794 7112 34850 7168
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 35990 7948 36046 7984
rect 35990 7928 35992 7948
rect 35992 7928 36044 7948
rect 36044 7928 36046 7948
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 35162 4664 35218 4720
rect 35714 6568 35770 6624
rect 35898 6160 35954 6216
rect 36542 15952 36598 16008
rect 36174 8744 36230 8800
rect 36266 7520 36322 7576
rect 36450 8356 36506 8392
rect 36450 8336 36452 8356
rect 36452 8336 36504 8356
rect 36504 8336 36506 8356
rect 36174 6432 36230 6488
rect 36266 5636 36322 5672
rect 36266 5616 36268 5636
rect 36268 5616 36320 5636
rect 36320 5616 36322 5636
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 35990 4392 36046 4448
rect 35898 4256 35954 4312
rect 36634 9424 36690 9480
rect 37922 24112 37978 24168
rect 38106 21800 38162 21856
rect 39118 23160 39174 23216
rect 38750 22208 38806 22264
rect 38658 21800 38714 21856
rect 39210 23060 39212 23080
rect 39212 23060 39264 23080
rect 39264 23060 39266 23080
rect 39210 23024 39266 23060
rect 41326 42880 41382 42936
rect 38106 17584 38162 17640
rect 38198 15952 38254 16008
rect 38934 20712 38990 20768
rect 37738 12144 37794 12200
rect 36634 4428 36636 4448
rect 36636 4428 36688 4448
rect 36688 4428 36690 4448
rect 36634 4392 36690 4428
rect 36266 3168 36322 3224
rect 37186 4120 37242 4176
rect 38106 10648 38162 10704
rect 37922 8608 37978 8664
rect 37738 6704 37794 6760
rect 38382 7384 38438 7440
rect 37738 4664 37794 4720
rect 39394 22208 39450 22264
rect 39946 22616 40002 22672
rect 39578 20032 39634 20088
rect 40406 21800 40462 21856
rect 40222 20440 40278 20496
rect 40222 19896 40278 19952
rect 40222 17448 40278 17504
rect 40038 15136 40094 15192
rect 39946 14864 40002 14920
rect 40038 12824 40094 12880
rect 39302 9696 39358 9752
rect 38566 4256 38622 4312
rect 38474 3712 38530 3768
rect 38382 2488 38438 2544
rect 39670 12280 39726 12336
rect 39762 10784 39818 10840
rect 39118 4392 39174 4448
rect 39026 3848 39082 3904
rect 42614 49716 42616 49736
rect 42616 49716 42668 49736
rect 42668 49716 42670 49736
rect 42614 49680 42670 49716
rect 41694 23024 41750 23080
rect 41970 23060 41972 23080
rect 41972 23060 42024 23080
rect 42024 23060 42026 23080
rect 40866 19796 40868 19816
rect 40868 19796 40920 19816
rect 40920 19796 40922 19816
rect 40866 19760 40922 19796
rect 40498 5752 40554 5808
rect 40222 3884 40224 3904
rect 40224 3884 40276 3904
rect 40276 3884 40278 3904
rect 40222 3848 40278 3884
rect 40682 4392 40738 4448
rect 41970 23024 42026 23060
rect 42246 22344 42302 22400
rect 41418 9696 41474 9752
rect 41234 5364 41290 5400
rect 41234 5344 41236 5364
rect 41236 5344 41288 5364
rect 41288 5344 41290 5364
rect 42062 17312 42118 17368
rect 42154 13776 42210 13832
rect 41970 10104 42026 10160
rect 41970 9560 42026 9616
rect 43074 41384 43130 41440
rect 42706 22636 42762 22672
rect 42706 22616 42708 22636
rect 42708 22616 42760 22636
rect 42760 22616 42762 22636
rect 42614 22344 42670 22400
rect 42982 21256 43038 21312
rect 42798 20576 42854 20632
rect 43442 24928 43498 24984
rect 43442 18028 43444 18048
rect 43444 18028 43496 18048
rect 43496 18028 43498 18048
rect 43442 17992 43498 18028
rect 43166 16632 43222 16688
rect 43534 12960 43590 13016
rect 43074 11228 43076 11248
rect 43076 11228 43128 11248
rect 43128 11228 43130 11248
rect 43074 11192 43130 11228
rect 43074 9696 43130 9752
rect 42614 6568 42670 6624
rect 42982 7948 43038 7984
rect 42982 7928 42984 7948
rect 42984 7928 43036 7948
rect 43036 7928 43038 7948
rect 41878 3304 41934 3360
rect 41418 2644 41474 2680
rect 41418 2624 41420 2644
rect 41420 2624 41472 2644
rect 41472 2624 41474 2644
rect 44362 22616 44418 22672
rect 43810 20712 43866 20768
rect 44546 20576 44602 20632
rect 44270 19896 44326 19952
rect 43994 19488 44050 19544
rect 43718 11736 43774 11792
rect 43350 6704 43406 6760
rect 43350 5616 43406 5672
rect 44362 19760 44418 19816
rect 44178 17176 44234 17232
rect 44822 19896 44878 19952
rect 43994 6296 44050 6352
rect 42706 3440 42762 3496
rect 43534 4004 43590 4040
rect 43534 3984 43536 4004
rect 43536 3984 43588 4004
rect 43588 3984 43590 4004
rect 43626 3168 43682 3224
rect 45926 25236 45928 25256
rect 45928 25236 45980 25256
rect 45980 25236 45982 25256
rect 45926 25200 45982 25236
rect 48870 56616 48926 56672
rect 47674 52692 47730 52728
rect 47674 52672 47676 52692
rect 47676 52672 47728 52692
rect 47728 52672 47730 52692
rect 48042 52536 48098 52592
rect 46018 21428 46020 21448
rect 46020 21428 46072 21448
rect 46072 21428 46074 21448
rect 46018 21392 46074 21428
rect 44638 8336 44694 8392
rect 44270 4004 44326 4040
rect 44270 3984 44272 4004
rect 44272 3984 44324 4004
rect 44324 3984 44326 4004
rect 43902 3032 43958 3088
rect 44454 3168 44510 3224
rect 44638 3188 44694 3224
rect 44638 3168 44640 3188
rect 44640 3168 44692 3188
rect 44692 3168 44694 3188
rect 45742 19760 45798 19816
rect 44914 6840 44970 6896
rect 45374 6432 45430 6488
rect 46938 25200 46994 25256
rect 47122 25236 47124 25256
rect 47124 25236 47176 25256
rect 47176 25236 47178 25256
rect 47122 25200 47178 25236
rect 46846 20304 46902 20360
rect 46846 19624 46902 19680
rect 46754 16108 46810 16144
rect 46754 16088 46756 16108
rect 46756 16088 46808 16108
rect 46808 16088 46810 16108
rect 46846 15580 46848 15600
rect 46848 15580 46900 15600
rect 46900 15580 46902 15600
rect 46846 15544 46902 15580
rect 45834 6840 45890 6896
rect 46386 8880 46442 8936
rect 46662 6604 46664 6624
rect 46664 6604 46716 6624
rect 46716 6604 46718 6624
rect 46662 6568 46718 6604
rect 46754 6432 46810 6488
rect 47766 51040 47822 51096
rect 48686 44240 48742 44296
rect 48226 23160 48282 23216
rect 47858 21956 47914 21992
rect 47858 21936 47860 21956
rect 47860 21936 47912 21956
rect 47912 21936 47914 21956
rect 47398 4528 47454 4584
rect 47398 3712 47454 3768
rect 50300 56602 50356 56604
rect 50380 56602 50436 56604
rect 50460 56602 50516 56604
rect 50540 56602 50596 56604
rect 50300 56550 50346 56602
rect 50346 56550 50356 56602
rect 50380 56550 50410 56602
rect 50410 56550 50422 56602
rect 50422 56550 50436 56602
rect 50460 56550 50474 56602
rect 50474 56550 50486 56602
rect 50486 56550 50516 56602
rect 50540 56550 50550 56602
rect 50550 56550 50596 56602
rect 50300 56548 50356 56550
rect 50380 56548 50436 56550
rect 50460 56548 50516 56550
rect 50540 56548 50596 56550
rect 50300 55514 50356 55516
rect 50380 55514 50436 55516
rect 50460 55514 50516 55516
rect 50540 55514 50596 55516
rect 50300 55462 50346 55514
rect 50346 55462 50356 55514
rect 50380 55462 50410 55514
rect 50410 55462 50422 55514
rect 50422 55462 50436 55514
rect 50460 55462 50474 55514
rect 50474 55462 50486 55514
rect 50486 55462 50516 55514
rect 50540 55462 50550 55514
rect 50550 55462 50596 55514
rect 50300 55460 50356 55462
rect 50380 55460 50436 55462
rect 50460 55460 50516 55462
rect 50540 55460 50596 55462
rect 50300 54426 50356 54428
rect 50380 54426 50436 54428
rect 50460 54426 50516 54428
rect 50540 54426 50596 54428
rect 50300 54374 50346 54426
rect 50346 54374 50356 54426
rect 50380 54374 50410 54426
rect 50410 54374 50422 54426
rect 50422 54374 50436 54426
rect 50460 54374 50474 54426
rect 50474 54374 50486 54426
rect 50486 54374 50516 54426
rect 50540 54374 50550 54426
rect 50550 54374 50596 54426
rect 50300 54372 50356 54374
rect 50380 54372 50436 54374
rect 50460 54372 50516 54374
rect 50540 54372 50596 54374
rect 50300 53338 50356 53340
rect 50380 53338 50436 53340
rect 50460 53338 50516 53340
rect 50540 53338 50596 53340
rect 50300 53286 50346 53338
rect 50346 53286 50356 53338
rect 50380 53286 50410 53338
rect 50410 53286 50422 53338
rect 50422 53286 50436 53338
rect 50460 53286 50474 53338
rect 50474 53286 50486 53338
rect 50486 53286 50516 53338
rect 50540 53286 50550 53338
rect 50550 53286 50596 53338
rect 50300 53284 50356 53286
rect 50380 53284 50436 53286
rect 50460 53284 50516 53286
rect 50540 53284 50596 53286
rect 50300 52250 50356 52252
rect 50380 52250 50436 52252
rect 50460 52250 50516 52252
rect 50540 52250 50596 52252
rect 50300 52198 50346 52250
rect 50346 52198 50356 52250
rect 50380 52198 50410 52250
rect 50410 52198 50422 52250
rect 50422 52198 50436 52250
rect 50460 52198 50474 52250
rect 50474 52198 50486 52250
rect 50486 52198 50516 52250
rect 50540 52198 50550 52250
rect 50550 52198 50596 52250
rect 50300 52196 50356 52198
rect 50380 52196 50436 52198
rect 50460 52196 50516 52198
rect 50540 52196 50596 52198
rect 50300 51162 50356 51164
rect 50380 51162 50436 51164
rect 50460 51162 50516 51164
rect 50540 51162 50596 51164
rect 50300 51110 50346 51162
rect 50346 51110 50356 51162
rect 50380 51110 50410 51162
rect 50410 51110 50422 51162
rect 50422 51110 50436 51162
rect 50460 51110 50474 51162
rect 50474 51110 50486 51162
rect 50486 51110 50516 51162
rect 50540 51110 50550 51162
rect 50550 51110 50596 51162
rect 50300 51108 50356 51110
rect 50380 51108 50436 51110
rect 50460 51108 50516 51110
rect 50540 51108 50596 51110
rect 48502 21392 48558 21448
rect 48502 21256 48558 21312
rect 48686 20304 48742 20360
rect 48410 17856 48466 17912
rect 48226 17076 48228 17096
rect 48228 17076 48280 17096
rect 48280 17076 48282 17096
rect 48226 17040 48282 17076
rect 48410 17076 48412 17096
rect 48412 17076 48464 17096
rect 48464 17076 48466 17096
rect 48410 17040 48466 17076
rect 48226 16496 48282 16552
rect 48134 7928 48190 7984
rect 48042 5480 48098 5536
rect 47766 4256 47822 4312
rect 47858 3984 47914 4040
rect 47674 3576 47730 3632
rect 48226 6704 48282 6760
rect 47950 2624 48006 2680
rect 48594 3984 48650 4040
rect 48410 3052 48466 3088
rect 48410 3032 48412 3052
rect 48412 3032 48464 3052
rect 48464 3032 48466 3052
rect 48594 3032 48650 3088
rect 49330 16496 49386 16552
rect 49238 2896 49294 2952
rect 50300 50074 50356 50076
rect 50380 50074 50436 50076
rect 50460 50074 50516 50076
rect 50540 50074 50596 50076
rect 50300 50022 50346 50074
rect 50346 50022 50356 50074
rect 50380 50022 50410 50074
rect 50410 50022 50422 50074
rect 50422 50022 50436 50074
rect 50460 50022 50474 50074
rect 50474 50022 50486 50074
rect 50486 50022 50516 50074
rect 50540 50022 50550 50074
rect 50550 50022 50596 50074
rect 50300 50020 50356 50022
rect 50380 50020 50436 50022
rect 50460 50020 50516 50022
rect 50540 50020 50596 50022
rect 50300 48986 50356 48988
rect 50380 48986 50436 48988
rect 50460 48986 50516 48988
rect 50540 48986 50596 48988
rect 50300 48934 50346 48986
rect 50346 48934 50356 48986
rect 50380 48934 50410 48986
rect 50410 48934 50422 48986
rect 50422 48934 50436 48986
rect 50460 48934 50474 48986
rect 50474 48934 50486 48986
rect 50486 48934 50516 48986
rect 50540 48934 50550 48986
rect 50550 48934 50596 48986
rect 50300 48932 50356 48934
rect 50380 48932 50436 48934
rect 50460 48932 50516 48934
rect 50540 48932 50596 48934
rect 50300 47898 50356 47900
rect 50380 47898 50436 47900
rect 50460 47898 50516 47900
rect 50540 47898 50596 47900
rect 50300 47846 50346 47898
rect 50346 47846 50356 47898
rect 50380 47846 50410 47898
rect 50410 47846 50422 47898
rect 50422 47846 50436 47898
rect 50460 47846 50474 47898
rect 50474 47846 50486 47898
rect 50486 47846 50516 47898
rect 50540 47846 50550 47898
rect 50550 47846 50596 47898
rect 50300 47844 50356 47846
rect 50380 47844 50436 47846
rect 50460 47844 50516 47846
rect 50540 47844 50596 47846
rect 50300 46810 50356 46812
rect 50380 46810 50436 46812
rect 50460 46810 50516 46812
rect 50540 46810 50596 46812
rect 50300 46758 50346 46810
rect 50346 46758 50356 46810
rect 50380 46758 50410 46810
rect 50410 46758 50422 46810
rect 50422 46758 50436 46810
rect 50460 46758 50474 46810
rect 50474 46758 50486 46810
rect 50486 46758 50516 46810
rect 50540 46758 50550 46810
rect 50550 46758 50596 46810
rect 50300 46756 50356 46758
rect 50380 46756 50436 46758
rect 50460 46756 50516 46758
rect 50540 46756 50596 46758
rect 50300 45722 50356 45724
rect 50380 45722 50436 45724
rect 50460 45722 50516 45724
rect 50540 45722 50596 45724
rect 50300 45670 50346 45722
rect 50346 45670 50356 45722
rect 50380 45670 50410 45722
rect 50410 45670 50422 45722
rect 50422 45670 50436 45722
rect 50460 45670 50474 45722
rect 50474 45670 50486 45722
rect 50486 45670 50516 45722
rect 50540 45670 50550 45722
rect 50550 45670 50596 45722
rect 50300 45668 50356 45670
rect 50380 45668 50436 45670
rect 50460 45668 50516 45670
rect 50540 45668 50596 45670
rect 50300 44634 50356 44636
rect 50380 44634 50436 44636
rect 50460 44634 50516 44636
rect 50540 44634 50596 44636
rect 50300 44582 50346 44634
rect 50346 44582 50356 44634
rect 50380 44582 50410 44634
rect 50410 44582 50422 44634
rect 50422 44582 50436 44634
rect 50460 44582 50474 44634
rect 50474 44582 50486 44634
rect 50486 44582 50516 44634
rect 50540 44582 50550 44634
rect 50550 44582 50596 44634
rect 50300 44580 50356 44582
rect 50380 44580 50436 44582
rect 50460 44580 50516 44582
rect 50540 44580 50596 44582
rect 50300 43546 50356 43548
rect 50380 43546 50436 43548
rect 50460 43546 50516 43548
rect 50540 43546 50596 43548
rect 50300 43494 50346 43546
rect 50346 43494 50356 43546
rect 50380 43494 50410 43546
rect 50410 43494 50422 43546
rect 50422 43494 50436 43546
rect 50460 43494 50474 43546
rect 50474 43494 50486 43546
rect 50486 43494 50516 43546
rect 50540 43494 50550 43546
rect 50550 43494 50596 43546
rect 50300 43492 50356 43494
rect 50380 43492 50436 43494
rect 50460 43492 50516 43494
rect 50540 43492 50596 43494
rect 50300 42458 50356 42460
rect 50380 42458 50436 42460
rect 50460 42458 50516 42460
rect 50540 42458 50596 42460
rect 50300 42406 50346 42458
rect 50346 42406 50356 42458
rect 50380 42406 50410 42458
rect 50410 42406 50422 42458
rect 50422 42406 50436 42458
rect 50460 42406 50474 42458
rect 50474 42406 50486 42458
rect 50486 42406 50516 42458
rect 50540 42406 50550 42458
rect 50550 42406 50596 42458
rect 50300 42404 50356 42406
rect 50380 42404 50436 42406
rect 50460 42404 50516 42406
rect 50540 42404 50596 42406
rect 50300 41370 50356 41372
rect 50380 41370 50436 41372
rect 50460 41370 50516 41372
rect 50540 41370 50596 41372
rect 50300 41318 50346 41370
rect 50346 41318 50356 41370
rect 50380 41318 50410 41370
rect 50410 41318 50422 41370
rect 50422 41318 50436 41370
rect 50460 41318 50474 41370
rect 50474 41318 50486 41370
rect 50486 41318 50516 41370
rect 50540 41318 50550 41370
rect 50550 41318 50596 41370
rect 50300 41316 50356 41318
rect 50380 41316 50436 41318
rect 50460 41316 50516 41318
rect 50540 41316 50596 41318
rect 50300 40282 50356 40284
rect 50380 40282 50436 40284
rect 50460 40282 50516 40284
rect 50540 40282 50596 40284
rect 50300 40230 50346 40282
rect 50346 40230 50356 40282
rect 50380 40230 50410 40282
rect 50410 40230 50422 40282
rect 50422 40230 50436 40282
rect 50460 40230 50474 40282
rect 50474 40230 50486 40282
rect 50486 40230 50516 40282
rect 50540 40230 50550 40282
rect 50550 40230 50596 40282
rect 50300 40228 50356 40230
rect 50380 40228 50436 40230
rect 50460 40228 50516 40230
rect 50540 40228 50596 40230
rect 50300 39194 50356 39196
rect 50380 39194 50436 39196
rect 50460 39194 50516 39196
rect 50540 39194 50596 39196
rect 50300 39142 50346 39194
rect 50346 39142 50356 39194
rect 50380 39142 50410 39194
rect 50410 39142 50422 39194
rect 50422 39142 50436 39194
rect 50460 39142 50474 39194
rect 50474 39142 50486 39194
rect 50486 39142 50516 39194
rect 50540 39142 50550 39194
rect 50550 39142 50596 39194
rect 50300 39140 50356 39142
rect 50380 39140 50436 39142
rect 50460 39140 50516 39142
rect 50540 39140 50596 39142
rect 50300 38106 50356 38108
rect 50380 38106 50436 38108
rect 50460 38106 50516 38108
rect 50540 38106 50596 38108
rect 50300 38054 50346 38106
rect 50346 38054 50356 38106
rect 50380 38054 50410 38106
rect 50410 38054 50422 38106
rect 50422 38054 50436 38106
rect 50460 38054 50474 38106
rect 50474 38054 50486 38106
rect 50486 38054 50516 38106
rect 50540 38054 50550 38106
rect 50550 38054 50596 38106
rect 50300 38052 50356 38054
rect 50380 38052 50436 38054
rect 50460 38052 50516 38054
rect 50540 38052 50596 38054
rect 50300 37018 50356 37020
rect 50380 37018 50436 37020
rect 50460 37018 50516 37020
rect 50540 37018 50596 37020
rect 50300 36966 50346 37018
rect 50346 36966 50356 37018
rect 50380 36966 50410 37018
rect 50410 36966 50422 37018
rect 50422 36966 50436 37018
rect 50460 36966 50474 37018
rect 50474 36966 50486 37018
rect 50486 36966 50516 37018
rect 50540 36966 50550 37018
rect 50550 36966 50596 37018
rect 50300 36964 50356 36966
rect 50380 36964 50436 36966
rect 50460 36964 50516 36966
rect 50540 36964 50596 36966
rect 50300 35930 50356 35932
rect 50380 35930 50436 35932
rect 50460 35930 50516 35932
rect 50540 35930 50596 35932
rect 50300 35878 50346 35930
rect 50346 35878 50356 35930
rect 50380 35878 50410 35930
rect 50410 35878 50422 35930
rect 50422 35878 50436 35930
rect 50460 35878 50474 35930
rect 50474 35878 50486 35930
rect 50486 35878 50516 35930
rect 50540 35878 50550 35930
rect 50550 35878 50596 35930
rect 50300 35876 50356 35878
rect 50380 35876 50436 35878
rect 50460 35876 50516 35878
rect 50540 35876 50596 35878
rect 50300 34842 50356 34844
rect 50380 34842 50436 34844
rect 50460 34842 50516 34844
rect 50540 34842 50596 34844
rect 50300 34790 50346 34842
rect 50346 34790 50356 34842
rect 50380 34790 50410 34842
rect 50410 34790 50422 34842
rect 50422 34790 50436 34842
rect 50460 34790 50474 34842
rect 50474 34790 50486 34842
rect 50486 34790 50516 34842
rect 50540 34790 50550 34842
rect 50550 34790 50596 34842
rect 50300 34788 50356 34790
rect 50380 34788 50436 34790
rect 50460 34788 50516 34790
rect 50540 34788 50596 34790
rect 50300 33754 50356 33756
rect 50380 33754 50436 33756
rect 50460 33754 50516 33756
rect 50540 33754 50596 33756
rect 50300 33702 50346 33754
rect 50346 33702 50356 33754
rect 50380 33702 50410 33754
rect 50410 33702 50422 33754
rect 50422 33702 50436 33754
rect 50460 33702 50474 33754
rect 50474 33702 50486 33754
rect 50486 33702 50516 33754
rect 50540 33702 50550 33754
rect 50550 33702 50596 33754
rect 50300 33700 50356 33702
rect 50380 33700 50436 33702
rect 50460 33700 50516 33702
rect 50540 33700 50596 33702
rect 50300 32666 50356 32668
rect 50380 32666 50436 32668
rect 50460 32666 50516 32668
rect 50540 32666 50596 32668
rect 50300 32614 50346 32666
rect 50346 32614 50356 32666
rect 50380 32614 50410 32666
rect 50410 32614 50422 32666
rect 50422 32614 50436 32666
rect 50460 32614 50474 32666
rect 50474 32614 50486 32666
rect 50486 32614 50516 32666
rect 50540 32614 50550 32666
rect 50550 32614 50596 32666
rect 50300 32612 50356 32614
rect 50380 32612 50436 32614
rect 50460 32612 50516 32614
rect 50540 32612 50596 32614
rect 50300 31578 50356 31580
rect 50380 31578 50436 31580
rect 50460 31578 50516 31580
rect 50540 31578 50596 31580
rect 50300 31526 50346 31578
rect 50346 31526 50356 31578
rect 50380 31526 50410 31578
rect 50410 31526 50422 31578
rect 50422 31526 50436 31578
rect 50460 31526 50474 31578
rect 50474 31526 50486 31578
rect 50486 31526 50516 31578
rect 50540 31526 50550 31578
rect 50550 31526 50596 31578
rect 50300 31524 50356 31526
rect 50380 31524 50436 31526
rect 50460 31524 50516 31526
rect 50540 31524 50596 31526
rect 50300 30490 50356 30492
rect 50380 30490 50436 30492
rect 50460 30490 50516 30492
rect 50540 30490 50596 30492
rect 50300 30438 50346 30490
rect 50346 30438 50356 30490
rect 50380 30438 50410 30490
rect 50410 30438 50422 30490
rect 50422 30438 50436 30490
rect 50460 30438 50474 30490
rect 50474 30438 50486 30490
rect 50486 30438 50516 30490
rect 50540 30438 50550 30490
rect 50550 30438 50596 30490
rect 50300 30436 50356 30438
rect 50380 30436 50436 30438
rect 50460 30436 50516 30438
rect 50540 30436 50596 30438
rect 50300 29402 50356 29404
rect 50380 29402 50436 29404
rect 50460 29402 50516 29404
rect 50540 29402 50596 29404
rect 50300 29350 50346 29402
rect 50346 29350 50356 29402
rect 50380 29350 50410 29402
rect 50410 29350 50422 29402
rect 50422 29350 50436 29402
rect 50460 29350 50474 29402
rect 50474 29350 50486 29402
rect 50486 29350 50516 29402
rect 50540 29350 50550 29402
rect 50550 29350 50596 29402
rect 50300 29348 50356 29350
rect 50380 29348 50436 29350
rect 50460 29348 50516 29350
rect 50540 29348 50596 29350
rect 50300 28314 50356 28316
rect 50380 28314 50436 28316
rect 50460 28314 50516 28316
rect 50540 28314 50596 28316
rect 50300 28262 50346 28314
rect 50346 28262 50356 28314
rect 50380 28262 50410 28314
rect 50410 28262 50422 28314
rect 50422 28262 50436 28314
rect 50460 28262 50474 28314
rect 50474 28262 50486 28314
rect 50486 28262 50516 28314
rect 50540 28262 50550 28314
rect 50550 28262 50596 28314
rect 50300 28260 50356 28262
rect 50380 28260 50436 28262
rect 50460 28260 50516 28262
rect 50540 28260 50596 28262
rect 50300 27226 50356 27228
rect 50380 27226 50436 27228
rect 50460 27226 50516 27228
rect 50540 27226 50596 27228
rect 50300 27174 50346 27226
rect 50346 27174 50356 27226
rect 50380 27174 50410 27226
rect 50410 27174 50422 27226
rect 50422 27174 50436 27226
rect 50460 27174 50474 27226
rect 50474 27174 50486 27226
rect 50486 27174 50516 27226
rect 50540 27174 50550 27226
rect 50550 27174 50596 27226
rect 50300 27172 50356 27174
rect 50380 27172 50436 27174
rect 50460 27172 50516 27174
rect 50540 27172 50596 27174
rect 50300 26138 50356 26140
rect 50380 26138 50436 26140
rect 50460 26138 50516 26140
rect 50540 26138 50596 26140
rect 50300 26086 50346 26138
rect 50346 26086 50356 26138
rect 50380 26086 50410 26138
rect 50410 26086 50422 26138
rect 50422 26086 50436 26138
rect 50460 26086 50474 26138
rect 50474 26086 50486 26138
rect 50486 26086 50516 26138
rect 50540 26086 50550 26138
rect 50550 26086 50596 26138
rect 50300 26084 50356 26086
rect 50380 26084 50436 26086
rect 50460 26084 50516 26086
rect 50540 26084 50596 26086
rect 50300 25050 50356 25052
rect 50380 25050 50436 25052
rect 50460 25050 50516 25052
rect 50540 25050 50596 25052
rect 50300 24998 50346 25050
rect 50346 24998 50356 25050
rect 50380 24998 50410 25050
rect 50410 24998 50422 25050
rect 50422 24998 50436 25050
rect 50460 24998 50474 25050
rect 50474 24998 50486 25050
rect 50486 24998 50516 25050
rect 50540 24998 50550 25050
rect 50550 24998 50596 25050
rect 50300 24996 50356 24998
rect 50380 24996 50436 24998
rect 50460 24996 50516 24998
rect 50540 24996 50596 24998
rect 50300 23962 50356 23964
rect 50380 23962 50436 23964
rect 50460 23962 50516 23964
rect 50540 23962 50596 23964
rect 50300 23910 50346 23962
rect 50346 23910 50356 23962
rect 50380 23910 50410 23962
rect 50410 23910 50422 23962
rect 50422 23910 50436 23962
rect 50460 23910 50474 23962
rect 50474 23910 50486 23962
rect 50486 23910 50516 23962
rect 50540 23910 50550 23962
rect 50550 23910 50596 23962
rect 50300 23908 50356 23910
rect 50380 23908 50436 23910
rect 50460 23908 50516 23910
rect 50540 23908 50596 23910
rect 50300 22874 50356 22876
rect 50380 22874 50436 22876
rect 50460 22874 50516 22876
rect 50540 22874 50596 22876
rect 50300 22822 50346 22874
rect 50346 22822 50356 22874
rect 50380 22822 50410 22874
rect 50410 22822 50422 22874
rect 50422 22822 50436 22874
rect 50460 22822 50474 22874
rect 50474 22822 50486 22874
rect 50486 22822 50516 22874
rect 50540 22822 50550 22874
rect 50550 22822 50596 22874
rect 50300 22820 50356 22822
rect 50380 22820 50436 22822
rect 50460 22820 50516 22822
rect 50540 22820 50596 22822
rect 50300 21786 50356 21788
rect 50380 21786 50436 21788
rect 50460 21786 50516 21788
rect 50540 21786 50596 21788
rect 50300 21734 50346 21786
rect 50346 21734 50356 21786
rect 50380 21734 50410 21786
rect 50410 21734 50422 21786
rect 50422 21734 50436 21786
rect 50460 21734 50474 21786
rect 50474 21734 50486 21786
rect 50486 21734 50516 21786
rect 50540 21734 50550 21786
rect 50550 21734 50596 21786
rect 50300 21732 50356 21734
rect 50380 21732 50436 21734
rect 50460 21732 50516 21734
rect 50540 21732 50596 21734
rect 50300 20698 50356 20700
rect 50380 20698 50436 20700
rect 50460 20698 50516 20700
rect 50540 20698 50596 20700
rect 50300 20646 50346 20698
rect 50346 20646 50356 20698
rect 50380 20646 50410 20698
rect 50410 20646 50422 20698
rect 50422 20646 50436 20698
rect 50460 20646 50474 20698
rect 50474 20646 50486 20698
rect 50486 20646 50516 20698
rect 50540 20646 50550 20698
rect 50550 20646 50596 20698
rect 50300 20644 50356 20646
rect 50380 20644 50436 20646
rect 50460 20644 50516 20646
rect 50540 20644 50596 20646
rect 50300 19610 50356 19612
rect 50380 19610 50436 19612
rect 50460 19610 50516 19612
rect 50540 19610 50596 19612
rect 50300 19558 50346 19610
rect 50346 19558 50356 19610
rect 50380 19558 50410 19610
rect 50410 19558 50422 19610
rect 50422 19558 50436 19610
rect 50460 19558 50474 19610
rect 50474 19558 50486 19610
rect 50486 19558 50516 19610
rect 50540 19558 50550 19610
rect 50550 19558 50596 19610
rect 50300 19556 50356 19558
rect 50380 19556 50436 19558
rect 50460 19556 50516 19558
rect 50540 19556 50596 19558
rect 50300 18522 50356 18524
rect 50380 18522 50436 18524
rect 50460 18522 50516 18524
rect 50540 18522 50596 18524
rect 50300 18470 50346 18522
rect 50346 18470 50356 18522
rect 50380 18470 50410 18522
rect 50410 18470 50422 18522
rect 50422 18470 50436 18522
rect 50460 18470 50474 18522
rect 50474 18470 50486 18522
rect 50486 18470 50516 18522
rect 50540 18470 50550 18522
rect 50550 18470 50596 18522
rect 50300 18468 50356 18470
rect 50380 18468 50436 18470
rect 50460 18468 50516 18470
rect 50540 18468 50596 18470
rect 50300 17434 50356 17436
rect 50380 17434 50436 17436
rect 50460 17434 50516 17436
rect 50540 17434 50596 17436
rect 50300 17382 50346 17434
rect 50346 17382 50356 17434
rect 50380 17382 50410 17434
rect 50410 17382 50422 17434
rect 50422 17382 50436 17434
rect 50460 17382 50474 17434
rect 50474 17382 50486 17434
rect 50486 17382 50516 17434
rect 50540 17382 50550 17434
rect 50550 17382 50596 17434
rect 50300 17380 50356 17382
rect 50380 17380 50436 17382
rect 50460 17380 50516 17382
rect 50540 17380 50596 17382
rect 50300 16346 50356 16348
rect 50380 16346 50436 16348
rect 50460 16346 50516 16348
rect 50540 16346 50596 16348
rect 50300 16294 50346 16346
rect 50346 16294 50356 16346
rect 50380 16294 50410 16346
rect 50410 16294 50422 16346
rect 50422 16294 50436 16346
rect 50460 16294 50474 16346
rect 50474 16294 50486 16346
rect 50486 16294 50516 16346
rect 50540 16294 50550 16346
rect 50550 16294 50596 16346
rect 50300 16292 50356 16294
rect 50380 16292 50436 16294
rect 50460 16292 50516 16294
rect 50540 16292 50596 16294
rect 50300 15258 50356 15260
rect 50380 15258 50436 15260
rect 50460 15258 50516 15260
rect 50540 15258 50596 15260
rect 50300 15206 50346 15258
rect 50346 15206 50356 15258
rect 50380 15206 50410 15258
rect 50410 15206 50422 15258
rect 50422 15206 50436 15258
rect 50460 15206 50474 15258
rect 50474 15206 50486 15258
rect 50486 15206 50516 15258
rect 50540 15206 50550 15258
rect 50550 15206 50596 15258
rect 50300 15204 50356 15206
rect 50380 15204 50436 15206
rect 50460 15204 50516 15206
rect 50540 15204 50596 15206
rect 50300 14170 50356 14172
rect 50380 14170 50436 14172
rect 50460 14170 50516 14172
rect 50540 14170 50596 14172
rect 50300 14118 50346 14170
rect 50346 14118 50356 14170
rect 50380 14118 50410 14170
rect 50410 14118 50422 14170
rect 50422 14118 50436 14170
rect 50460 14118 50474 14170
rect 50474 14118 50486 14170
rect 50486 14118 50516 14170
rect 50540 14118 50550 14170
rect 50550 14118 50596 14170
rect 50300 14116 50356 14118
rect 50380 14116 50436 14118
rect 50460 14116 50516 14118
rect 50540 14116 50596 14118
rect 50300 13082 50356 13084
rect 50380 13082 50436 13084
rect 50460 13082 50516 13084
rect 50540 13082 50596 13084
rect 50300 13030 50346 13082
rect 50346 13030 50356 13082
rect 50380 13030 50410 13082
rect 50410 13030 50422 13082
rect 50422 13030 50436 13082
rect 50460 13030 50474 13082
rect 50474 13030 50486 13082
rect 50486 13030 50516 13082
rect 50540 13030 50550 13082
rect 50550 13030 50596 13082
rect 50300 13028 50356 13030
rect 50380 13028 50436 13030
rect 50460 13028 50516 13030
rect 50540 13028 50596 13030
rect 50300 11994 50356 11996
rect 50380 11994 50436 11996
rect 50460 11994 50516 11996
rect 50540 11994 50596 11996
rect 50300 11942 50346 11994
rect 50346 11942 50356 11994
rect 50380 11942 50410 11994
rect 50410 11942 50422 11994
rect 50422 11942 50436 11994
rect 50460 11942 50474 11994
rect 50474 11942 50486 11994
rect 50486 11942 50516 11994
rect 50540 11942 50550 11994
rect 50550 11942 50596 11994
rect 50300 11940 50356 11942
rect 50380 11940 50436 11942
rect 50460 11940 50516 11942
rect 50540 11940 50596 11942
rect 50300 10906 50356 10908
rect 50380 10906 50436 10908
rect 50460 10906 50516 10908
rect 50540 10906 50596 10908
rect 50300 10854 50346 10906
rect 50346 10854 50356 10906
rect 50380 10854 50410 10906
rect 50410 10854 50422 10906
rect 50422 10854 50436 10906
rect 50460 10854 50474 10906
rect 50474 10854 50486 10906
rect 50486 10854 50516 10906
rect 50540 10854 50550 10906
rect 50550 10854 50596 10906
rect 50300 10852 50356 10854
rect 50380 10852 50436 10854
rect 50460 10852 50516 10854
rect 50540 10852 50596 10854
rect 50300 9818 50356 9820
rect 50380 9818 50436 9820
rect 50460 9818 50516 9820
rect 50540 9818 50596 9820
rect 50300 9766 50346 9818
rect 50346 9766 50356 9818
rect 50380 9766 50410 9818
rect 50410 9766 50422 9818
rect 50422 9766 50436 9818
rect 50460 9766 50474 9818
rect 50474 9766 50486 9818
rect 50486 9766 50516 9818
rect 50540 9766 50550 9818
rect 50550 9766 50596 9818
rect 50300 9764 50356 9766
rect 50380 9764 50436 9766
rect 50460 9764 50516 9766
rect 50540 9764 50596 9766
rect 50300 8730 50356 8732
rect 50380 8730 50436 8732
rect 50460 8730 50516 8732
rect 50540 8730 50596 8732
rect 50300 8678 50346 8730
rect 50346 8678 50356 8730
rect 50380 8678 50410 8730
rect 50410 8678 50422 8730
rect 50422 8678 50436 8730
rect 50460 8678 50474 8730
rect 50474 8678 50486 8730
rect 50486 8678 50516 8730
rect 50540 8678 50550 8730
rect 50550 8678 50596 8730
rect 50300 8676 50356 8678
rect 50380 8676 50436 8678
rect 50460 8676 50516 8678
rect 50540 8676 50596 8678
rect 50300 7642 50356 7644
rect 50380 7642 50436 7644
rect 50460 7642 50516 7644
rect 50540 7642 50596 7644
rect 50300 7590 50346 7642
rect 50346 7590 50356 7642
rect 50380 7590 50410 7642
rect 50410 7590 50422 7642
rect 50422 7590 50436 7642
rect 50460 7590 50474 7642
rect 50474 7590 50486 7642
rect 50486 7590 50516 7642
rect 50540 7590 50550 7642
rect 50550 7590 50596 7642
rect 50300 7588 50356 7590
rect 50380 7588 50436 7590
rect 50460 7588 50516 7590
rect 50540 7588 50596 7590
rect 50300 6554 50356 6556
rect 50380 6554 50436 6556
rect 50460 6554 50516 6556
rect 50540 6554 50596 6556
rect 50300 6502 50346 6554
rect 50346 6502 50356 6554
rect 50380 6502 50410 6554
rect 50410 6502 50422 6554
rect 50422 6502 50436 6554
rect 50460 6502 50474 6554
rect 50474 6502 50486 6554
rect 50486 6502 50516 6554
rect 50540 6502 50550 6554
rect 50550 6502 50596 6554
rect 50300 6500 50356 6502
rect 50380 6500 50436 6502
rect 50460 6500 50516 6502
rect 50540 6500 50596 6502
rect 50300 5466 50356 5468
rect 50380 5466 50436 5468
rect 50460 5466 50516 5468
rect 50540 5466 50596 5468
rect 50300 5414 50346 5466
rect 50346 5414 50356 5466
rect 50380 5414 50410 5466
rect 50410 5414 50422 5466
rect 50422 5414 50436 5466
rect 50460 5414 50474 5466
rect 50474 5414 50486 5466
rect 50486 5414 50516 5466
rect 50540 5414 50550 5466
rect 50550 5414 50596 5466
rect 50300 5412 50356 5414
rect 50380 5412 50436 5414
rect 50460 5412 50516 5414
rect 50540 5412 50596 5414
rect 50300 4378 50356 4380
rect 50380 4378 50436 4380
rect 50460 4378 50516 4380
rect 50540 4378 50596 4380
rect 50300 4326 50346 4378
rect 50346 4326 50356 4378
rect 50380 4326 50410 4378
rect 50410 4326 50422 4378
rect 50422 4326 50436 4378
rect 50460 4326 50474 4378
rect 50474 4326 50486 4378
rect 50486 4326 50516 4378
rect 50540 4326 50550 4378
rect 50550 4326 50596 4378
rect 50300 4324 50356 4326
rect 50380 4324 50436 4326
rect 50460 4324 50516 4326
rect 50540 4324 50596 4326
rect 50434 3476 50436 3496
rect 50436 3476 50488 3496
rect 50488 3476 50490 3496
rect 49882 3304 49938 3360
rect 50434 3440 50490 3476
rect 50300 3290 50356 3292
rect 50380 3290 50436 3292
rect 50460 3290 50516 3292
rect 50540 3290 50596 3292
rect 50300 3238 50346 3290
rect 50346 3238 50356 3290
rect 50380 3238 50410 3290
rect 50410 3238 50422 3290
rect 50422 3238 50436 3290
rect 50460 3238 50474 3290
rect 50474 3238 50486 3290
rect 50486 3238 50516 3290
rect 50540 3238 50550 3290
rect 50550 3238 50596 3290
rect 50300 3236 50356 3238
rect 50380 3236 50436 3238
rect 50460 3236 50516 3238
rect 50540 3236 50596 3238
rect 50300 2202 50356 2204
rect 50380 2202 50436 2204
rect 50460 2202 50516 2204
rect 50540 2202 50596 2204
rect 50300 2150 50346 2202
rect 50346 2150 50356 2202
rect 50380 2150 50410 2202
rect 50410 2150 50422 2202
rect 50422 2150 50436 2202
rect 50460 2150 50474 2202
rect 50474 2150 50486 2202
rect 50486 2150 50516 2202
rect 50540 2150 50550 2202
rect 50550 2150 50596 2202
rect 50300 2148 50356 2150
rect 50380 2148 50436 2150
rect 50460 2148 50516 2150
rect 50540 2148 50596 2150
rect 52458 18672 52514 18728
rect 52274 17060 52330 17096
rect 52274 17040 52276 17060
rect 52276 17040 52328 17060
rect 52328 17040 52330 17060
rect 52458 2488 52514 2544
rect 53746 4120 53802 4176
rect 55218 20984 55274 21040
rect 55218 3168 55274 3224
rect 58990 58656 59046 58712
rect 58714 58248 58770 58304
rect 58990 57840 59046 57896
rect 58806 57432 58862 57488
rect 58990 57044 59046 57080
rect 58990 57024 58992 57044
rect 58992 57024 59044 57044
rect 59044 57024 59046 57044
rect 58990 56616 59046 56672
rect 58898 56208 58954 56264
rect 58990 55800 59046 55856
rect 58162 55392 58218 55448
rect 58162 52944 58218 53000
rect 58990 54984 59046 55040
rect 58990 54612 58992 54632
rect 58992 54612 59044 54632
rect 59044 54612 59046 54632
rect 58990 54576 59046 54612
rect 58806 54168 58862 54224
rect 58254 50088 58310 50144
rect 58162 49680 58218 49736
rect 57978 48864 58034 48920
rect 58162 45600 58218 45656
rect 58162 44376 58218 44432
rect 56046 20868 56102 20904
rect 56046 20848 56048 20868
rect 56048 20848 56100 20868
rect 56100 20848 56102 20868
rect 56414 20324 56470 20360
rect 56414 20304 56416 20324
rect 56416 20304 56468 20324
rect 56468 20304 56470 20324
rect 56046 16652 56102 16688
rect 56046 16632 56048 16652
rect 56048 16632 56100 16652
rect 56100 16632 56102 16652
rect 55586 12844 55642 12880
rect 55586 12824 55588 12844
rect 55588 12824 55640 12844
rect 55640 12824 55642 12844
rect 56690 18672 56746 18728
rect 58070 43560 58126 43616
rect 58070 37032 58126 37088
rect 58162 36236 58218 36272
rect 58162 36216 58164 36236
rect 58164 36216 58216 36236
rect 58216 36216 58218 36236
rect 58162 35808 58218 35864
rect 58162 35012 58218 35048
rect 58162 34992 58164 35012
rect 58164 34992 58216 35012
rect 58216 34992 58218 35012
rect 58070 34604 58126 34640
rect 58070 34584 58072 34604
rect 58072 34584 58124 34604
rect 58124 34584 58126 34604
rect 58162 33768 58218 33824
rect 58070 33360 58126 33416
rect 58162 32544 58218 32600
rect 57610 20032 57666 20088
rect 58070 32136 58126 32192
rect 58346 42336 58402 42392
rect 58346 39908 58402 39944
rect 58346 39888 58348 39908
rect 58348 39888 58400 39908
rect 58400 39888 58402 39908
rect 58346 38700 58348 38720
rect 58348 38700 58400 38720
rect 58400 38700 58402 38720
rect 58346 38664 58402 38700
rect 58898 53760 58954 53816
rect 58990 53352 59046 53408
rect 58990 52536 59046 52592
rect 58898 52128 58954 52184
rect 58070 30912 58126 30968
rect 58162 30504 58218 30560
rect 58162 30096 58218 30152
rect 58070 29688 58126 29744
rect 58070 29280 58126 29336
rect 58990 51720 59046 51776
rect 58990 51348 58992 51368
rect 58992 51348 59044 51368
rect 59044 51348 59046 51368
rect 58990 51312 59046 51348
rect 58806 50904 58862 50960
rect 58898 50496 58954 50552
rect 58990 49272 59046 49328
rect 58990 48456 59046 48512
rect 58990 48084 58992 48104
rect 58992 48084 59044 48104
rect 59044 48084 59046 48104
rect 58990 48048 59046 48084
rect 58806 47640 58862 47696
rect 58162 28872 58218 28928
rect 58070 28464 58126 28520
rect 58162 27240 58218 27296
rect 58162 26444 58218 26480
rect 58162 26424 58164 26444
rect 58164 26424 58216 26444
rect 58216 26424 58218 26444
rect 58162 26016 58218 26072
rect 58162 25220 58218 25256
rect 58162 25200 58164 25220
rect 58164 25200 58216 25220
rect 58216 25200 58218 25220
rect 58070 24812 58126 24848
rect 58070 24792 58072 24812
rect 58072 24792 58124 24812
rect 58124 24792 58126 24812
rect 58162 23976 58218 24032
rect 58070 23568 58126 23624
rect 58162 22752 58218 22808
rect 58070 22344 58126 22400
rect 58070 21120 58126 21176
rect 58254 20304 58310 20360
rect 57978 19896 58034 19952
rect 58162 19896 58218 19952
rect 58162 19080 58218 19136
rect 58162 17448 58218 17504
rect 58162 16224 58218 16280
rect 58162 15428 58218 15464
rect 58162 15408 58164 15428
rect 58164 15408 58216 15428
rect 58216 15408 58218 15428
rect 58070 15020 58126 15056
rect 58070 15000 58072 15020
rect 58072 15000 58124 15020
rect 58124 15000 58126 15020
rect 58162 14184 58218 14240
rect 58162 13912 58218 13968
rect 58070 13776 58126 13832
rect 58070 12552 58126 12608
rect 58162 11736 58218 11792
rect 58070 11328 58126 11384
rect 58070 8880 58126 8936
rect 58162 8064 58218 8120
rect 58070 7656 58126 7712
rect 58254 7268 58310 7304
rect 58254 7248 58256 7268
rect 58256 7248 58308 7268
rect 58308 7248 58310 7268
rect 58990 47232 59046 47288
rect 58898 46824 58954 46880
rect 58990 46416 59046 46472
rect 58990 46008 59046 46064
rect 58990 45192 59046 45248
rect 58898 44784 58954 44840
rect 58990 43968 59046 44024
rect 58898 43152 58954 43208
rect 58990 42744 59046 42800
rect 58990 41112 59046 41168
rect 58990 37440 59046 37496
rect 58990 31764 58992 31784
rect 58992 31764 59044 31784
rect 59044 31764 59046 31784
rect 58990 31728 59046 31764
rect 58898 31320 58954 31376
rect 58990 27648 59046 27704
rect 58990 21528 59046 21584
rect 58990 18672 59046 18728
rect 58990 17856 59046 17912
rect 58990 16632 59046 16688
rect 59082 16124 59084 16144
rect 59084 16124 59136 16144
rect 59136 16124 59138 16144
rect 59082 16088 59138 16124
rect 58990 12960 59046 13016
rect 58990 10512 59046 10568
rect 58898 10104 58954 10160
rect 58990 9288 59046 9344
rect 58714 8472 58770 8528
rect 58990 6840 59046 6896
rect 58990 6432 59046 6488
rect 58990 5636 59046 5672
rect 58990 5616 58992 5636
rect 58992 5616 59044 5636
rect 59044 5616 59046 5636
rect 58070 5228 58126 5264
rect 58070 5208 58072 5228
rect 58072 5208 58124 5228
rect 58124 5208 58126 5228
rect 55862 1128 55918 1184
rect 58070 3984 58126 4040
rect 58990 4392 59046 4448
rect 58898 2760 58954 2816
rect 58990 2388 58992 2408
rect 58992 2388 59044 2408
rect 59044 2388 59046 2408
rect 58990 2352 59046 2388
rect 58898 1944 58954 2000
rect 58806 1536 58862 1592
<< metal3 >>
rect 58985 58714 59051 58717
rect 59200 58714 60000 58744
rect 58985 58712 60000 58714
rect 58985 58656 58990 58712
rect 59046 58656 60000 58712
rect 58985 58654 60000 58656
rect 58985 58651 59051 58654
rect 59200 58624 60000 58654
rect 58709 58306 58775 58309
rect 59200 58306 60000 58336
rect 58709 58304 60000 58306
rect 58709 58248 58714 58304
rect 58770 58248 60000 58304
rect 58709 58246 60000 58248
rect 58709 58243 58775 58246
rect 59200 58216 60000 58246
rect 58985 57898 59051 57901
rect 59200 57898 60000 57928
rect 58985 57896 60000 57898
rect 58985 57840 58990 57896
rect 59046 57840 60000 57896
rect 58985 57838 60000 57840
rect 58985 57835 59051 57838
rect 59200 57808 60000 57838
rect 19570 57696 19886 57697
rect 19570 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19886 57696
rect 19570 57631 19886 57632
rect 50290 57696 50606 57697
rect 50290 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50606 57696
rect 50290 57631 50606 57632
rect 58801 57490 58867 57493
rect 59200 57490 60000 57520
rect 58801 57488 60000 57490
rect 58801 57432 58806 57488
rect 58862 57432 60000 57488
rect 58801 57430 60000 57432
rect 58801 57427 58867 57430
rect 59200 57400 60000 57430
rect 4210 57152 4526 57153
rect 4210 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4526 57152
rect 4210 57087 4526 57088
rect 34930 57152 35246 57153
rect 34930 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35246 57152
rect 34930 57087 35246 57088
rect 58985 57082 59051 57085
rect 59200 57082 60000 57112
rect 58985 57080 60000 57082
rect 58985 57024 58990 57080
rect 59046 57024 60000 57080
rect 58985 57022 60000 57024
rect 58985 57019 59051 57022
rect 59200 56992 60000 57022
rect 48446 56612 48452 56676
rect 48516 56674 48522 56676
rect 48865 56674 48931 56677
rect 48516 56672 48931 56674
rect 48516 56616 48870 56672
rect 48926 56616 48931 56672
rect 48516 56614 48931 56616
rect 48516 56612 48522 56614
rect 48865 56611 48931 56614
rect 58985 56674 59051 56677
rect 59200 56674 60000 56704
rect 58985 56672 60000 56674
rect 58985 56616 58990 56672
rect 59046 56616 60000 56672
rect 58985 56614 60000 56616
rect 58985 56611 59051 56614
rect 19570 56608 19886 56609
rect 19570 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19886 56608
rect 19570 56543 19886 56544
rect 50290 56608 50606 56609
rect 50290 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50606 56608
rect 59200 56584 60000 56614
rect 50290 56543 50606 56544
rect 58893 56266 58959 56269
rect 59200 56266 60000 56296
rect 58893 56264 60000 56266
rect 58893 56208 58898 56264
rect 58954 56208 60000 56264
rect 58893 56206 60000 56208
rect 58893 56203 58959 56206
rect 59200 56176 60000 56206
rect 4210 56064 4526 56065
rect 4210 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4526 56064
rect 4210 55999 4526 56000
rect 34930 56064 35246 56065
rect 34930 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35246 56064
rect 34930 55999 35246 56000
rect 0 55858 800 55888
rect 933 55858 999 55861
rect 0 55856 999 55858
rect 0 55800 938 55856
rect 994 55800 999 55856
rect 0 55798 999 55800
rect 0 55768 800 55798
rect 933 55795 999 55798
rect 58985 55858 59051 55861
rect 59200 55858 60000 55888
rect 58985 55856 60000 55858
rect 58985 55800 58990 55856
rect 59046 55800 60000 55856
rect 58985 55798 60000 55800
rect 58985 55795 59051 55798
rect 59200 55768 60000 55798
rect 19570 55520 19886 55521
rect 19570 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19886 55520
rect 19570 55455 19886 55456
rect 50290 55520 50606 55521
rect 50290 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50606 55520
rect 50290 55455 50606 55456
rect 58157 55450 58223 55453
rect 59200 55450 60000 55480
rect 58157 55448 60000 55450
rect 58157 55392 58162 55448
rect 58218 55392 60000 55448
rect 58157 55390 60000 55392
rect 58157 55387 58223 55390
rect 59200 55360 60000 55390
rect 0 55314 800 55344
rect 933 55314 999 55317
rect 0 55312 999 55314
rect 0 55256 938 55312
rect 994 55256 999 55312
rect 0 55254 999 55256
rect 0 55224 800 55254
rect 933 55251 999 55254
rect 58985 55042 59051 55045
rect 59200 55042 60000 55072
rect 58985 55040 60000 55042
rect 58985 54984 58990 55040
rect 59046 54984 60000 55040
rect 58985 54982 60000 54984
rect 58985 54979 59051 54982
rect 4210 54976 4526 54977
rect 4210 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4526 54976
rect 4210 54911 4526 54912
rect 34930 54976 35246 54977
rect 34930 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35246 54976
rect 59200 54952 60000 54982
rect 34930 54911 35246 54912
rect 0 54770 800 54800
rect 1025 54770 1091 54773
rect 0 54768 1091 54770
rect 0 54712 1030 54768
rect 1086 54712 1091 54768
rect 0 54710 1091 54712
rect 0 54680 800 54710
rect 1025 54707 1091 54710
rect 58985 54634 59051 54637
rect 59200 54634 60000 54664
rect 58985 54632 60000 54634
rect 58985 54576 58990 54632
rect 59046 54576 60000 54632
rect 58985 54574 60000 54576
rect 58985 54571 59051 54574
rect 59200 54544 60000 54574
rect 19570 54432 19886 54433
rect 19570 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19886 54432
rect 19570 54367 19886 54368
rect 50290 54432 50606 54433
rect 50290 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50606 54432
rect 50290 54367 50606 54368
rect 0 54226 800 54256
rect 933 54226 999 54229
rect 0 54224 999 54226
rect 0 54168 938 54224
rect 994 54168 999 54224
rect 0 54166 999 54168
rect 0 54136 800 54166
rect 933 54163 999 54166
rect 58801 54226 58867 54229
rect 59200 54226 60000 54256
rect 58801 54224 60000 54226
rect 58801 54168 58806 54224
rect 58862 54168 60000 54224
rect 58801 54166 60000 54168
rect 58801 54163 58867 54166
rect 59200 54136 60000 54166
rect 4210 53888 4526 53889
rect 4210 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4526 53888
rect 4210 53823 4526 53824
rect 34930 53888 35246 53889
rect 34930 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35246 53888
rect 34930 53823 35246 53824
rect 58893 53818 58959 53821
rect 59200 53818 60000 53848
rect 58893 53816 60000 53818
rect 58893 53760 58898 53816
rect 58954 53760 60000 53816
rect 58893 53758 60000 53760
rect 58893 53755 58959 53758
rect 59200 53728 60000 53758
rect 0 53682 800 53712
rect 1025 53682 1091 53685
rect 0 53680 1091 53682
rect 0 53624 1030 53680
rect 1086 53624 1091 53680
rect 0 53622 1091 53624
rect 0 53592 800 53622
rect 1025 53619 1091 53622
rect 58985 53410 59051 53413
rect 59200 53410 60000 53440
rect 58985 53408 60000 53410
rect 58985 53352 58990 53408
rect 59046 53352 60000 53408
rect 58985 53350 60000 53352
rect 58985 53347 59051 53350
rect 19570 53344 19886 53345
rect 19570 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19886 53344
rect 19570 53279 19886 53280
rect 50290 53344 50606 53345
rect 50290 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50606 53344
rect 59200 53320 60000 53350
rect 50290 53279 50606 53280
rect 0 53138 800 53168
rect 933 53138 999 53141
rect 0 53136 999 53138
rect 0 53080 938 53136
rect 994 53080 999 53136
rect 0 53078 999 53080
rect 0 53048 800 53078
rect 933 53075 999 53078
rect 58157 53002 58223 53005
rect 59200 53002 60000 53032
rect 58157 53000 60000 53002
rect 58157 52944 58162 53000
rect 58218 52944 60000 53000
rect 58157 52942 60000 52944
rect 58157 52939 58223 52942
rect 59200 52912 60000 52942
rect 4210 52800 4526 52801
rect 4210 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4526 52800
rect 4210 52735 4526 52736
rect 34930 52800 35246 52801
rect 34930 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35246 52800
rect 34930 52735 35246 52736
rect 47669 52730 47735 52733
rect 48078 52730 48084 52732
rect 47669 52728 48084 52730
rect 47669 52672 47674 52728
rect 47730 52672 48084 52728
rect 47669 52670 48084 52672
rect 47669 52667 47735 52670
rect 48078 52668 48084 52670
rect 48148 52668 48154 52732
rect 0 52594 800 52624
rect 1025 52594 1091 52597
rect 0 52592 1091 52594
rect 0 52536 1030 52592
rect 1086 52536 1091 52592
rect 0 52534 1091 52536
rect 0 52504 800 52534
rect 1025 52531 1091 52534
rect 47894 52532 47900 52596
rect 47964 52594 47970 52596
rect 48037 52594 48103 52597
rect 47964 52592 48103 52594
rect 47964 52536 48042 52592
rect 48098 52536 48103 52592
rect 47964 52534 48103 52536
rect 47964 52532 47970 52534
rect 48037 52531 48103 52534
rect 58985 52594 59051 52597
rect 59200 52594 60000 52624
rect 58985 52592 60000 52594
rect 58985 52536 58990 52592
rect 59046 52536 60000 52592
rect 58985 52534 60000 52536
rect 58985 52531 59051 52534
rect 59200 52504 60000 52534
rect 19570 52256 19886 52257
rect 19570 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19886 52256
rect 19570 52191 19886 52192
rect 50290 52256 50606 52257
rect 50290 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50606 52256
rect 50290 52191 50606 52192
rect 58893 52186 58959 52189
rect 59200 52186 60000 52216
rect 58893 52184 60000 52186
rect 58893 52128 58898 52184
rect 58954 52128 60000 52184
rect 58893 52126 60000 52128
rect 58893 52123 58959 52126
rect 59200 52096 60000 52126
rect 0 52050 800 52080
rect 933 52050 999 52053
rect 0 52048 999 52050
rect 0 51992 938 52048
rect 994 51992 999 52048
rect 0 51990 999 51992
rect 0 51960 800 51990
rect 933 51987 999 51990
rect 58985 51778 59051 51781
rect 59200 51778 60000 51808
rect 58985 51776 60000 51778
rect 58985 51720 58990 51776
rect 59046 51720 60000 51776
rect 58985 51718 60000 51720
rect 58985 51715 59051 51718
rect 4210 51712 4526 51713
rect 4210 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4526 51712
rect 4210 51647 4526 51648
rect 34930 51712 35246 51713
rect 34930 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35246 51712
rect 59200 51688 60000 51718
rect 34930 51647 35246 51648
rect 0 51506 800 51536
rect 1025 51506 1091 51509
rect 0 51504 1091 51506
rect 0 51448 1030 51504
rect 1086 51448 1091 51504
rect 0 51446 1091 51448
rect 0 51416 800 51446
rect 1025 51443 1091 51446
rect 58985 51370 59051 51373
rect 59200 51370 60000 51400
rect 58985 51368 60000 51370
rect 58985 51312 58990 51368
rect 59046 51312 60000 51368
rect 58985 51310 60000 51312
rect 58985 51307 59051 51310
rect 59200 51280 60000 51310
rect 19570 51168 19886 51169
rect 19570 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19886 51168
rect 19570 51103 19886 51104
rect 50290 51168 50606 51169
rect 50290 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50606 51168
rect 50290 51103 50606 51104
rect 47761 51100 47827 51101
rect 47710 51098 47716 51100
rect 47670 51038 47716 51098
rect 47780 51096 47827 51100
rect 47822 51040 47827 51096
rect 47710 51036 47716 51038
rect 47780 51036 47827 51040
rect 47761 51035 47827 51036
rect 0 50962 800 50992
rect 933 50962 999 50965
rect 0 50960 999 50962
rect 0 50904 938 50960
rect 994 50904 999 50960
rect 0 50902 999 50904
rect 0 50872 800 50902
rect 933 50899 999 50902
rect 58801 50962 58867 50965
rect 59200 50962 60000 50992
rect 58801 50960 60000 50962
rect 58801 50904 58806 50960
rect 58862 50904 60000 50960
rect 58801 50902 60000 50904
rect 58801 50899 58867 50902
rect 59200 50872 60000 50902
rect 4210 50624 4526 50625
rect 4210 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4526 50624
rect 4210 50559 4526 50560
rect 34930 50624 35246 50625
rect 34930 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35246 50624
rect 34930 50559 35246 50560
rect 58893 50554 58959 50557
rect 59200 50554 60000 50584
rect 58893 50552 60000 50554
rect 58893 50496 58898 50552
rect 58954 50496 60000 50552
rect 58893 50494 60000 50496
rect 58893 50491 58959 50494
rect 59200 50464 60000 50494
rect 0 50418 800 50448
rect 1025 50418 1091 50421
rect 0 50416 1091 50418
rect 0 50360 1030 50416
rect 1086 50360 1091 50416
rect 0 50358 1091 50360
rect 0 50328 800 50358
rect 1025 50355 1091 50358
rect 58249 50146 58315 50149
rect 59200 50146 60000 50176
rect 58249 50144 60000 50146
rect 58249 50088 58254 50144
rect 58310 50088 60000 50144
rect 58249 50086 60000 50088
rect 58249 50083 58315 50086
rect 19570 50080 19886 50081
rect 19570 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19886 50080
rect 19570 50015 19886 50016
rect 50290 50080 50606 50081
rect 50290 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50606 50080
rect 59200 50056 60000 50086
rect 50290 50015 50606 50016
rect 0 49874 800 49904
rect 933 49874 999 49877
rect 0 49872 999 49874
rect 0 49816 938 49872
rect 994 49816 999 49872
rect 0 49814 999 49816
rect 0 49784 800 49814
rect 933 49811 999 49814
rect 42609 49740 42675 49741
rect 42558 49738 42564 49740
rect 42518 49678 42564 49738
rect 42628 49736 42675 49740
rect 42670 49680 42675 49736
rect 42558 49676 42564 49678
rect 42628 49676 42675 49680
rect 42609 49675 42675 49676
rect 58157 49738 58223 49741
rect 59200 49738 60000 49768
rect 58157 49736 60000 49738
rect 58157 49680 58162 49736
rect 58218 49680 60000 49736
rect 58157 49678 60000 49680
rect 58157 49675 58223 49678
rect 59200 49648 60000 49678
rect 4210 49536 4526 49537
rect 4210 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4526 49536
rect 4210 49471 4526 49472
rect 34930 49536 35246 49537
rect 34930 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35246 49536
rect 34930 49471 35246 49472
rect 0 49330 800 49360
rect 1025 49330 1091 49333
rect 0 49328 1091 49330
rect 0 49272 1030 49328
rect 1086 49272 1091 49328
rect 0 49270 1091 49272
rect 0 49240 800 49270
rect 1025 49267 1091 49270
rect 58985 49330 59051 49333
rect 59200 49330 60000 49360
rect 58985 49328 60000 49330
rect 58985 49272 58990 49328
rect 59046 49272 60000 49328
rect 58985 49270 60000 49272
rect 58985 49267 59051 49270
rect 59200 49240 60000 49270
rect 19570 48992 19886 48993
rect 19570 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19886 48992
rect 19570 48927 19886 48928
rect 50290 48992 50606 48993
rect 50290 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50606 48992
rect 50290 48927 50606 48928
rect 57973 48922 58039 48925
rect 59200 48922 60000 48952
rect 57973 48920 60000 48922
rect 57973 48864 57978 48920
rect 58034 48864 60000 48920
rect 57973 48862 60000 48864
rect 57973 48859 58039 48862
rect 59200 48832 60000 48862
rect 0 48786 800 48816
rect 933 48786 999 48789
rect 0 48784 999 48786
rect 0 48728 938 48784
rect 994 48728 999 48784
rect 0 48726 999 48728
rect 0 48696 800 48726
rect 933 48723 999 48726
rect 58985 48514 59051 48517
rect 59200 48514 60000 48544
rect 58985 48512 60000 48514
rect 58985 48456 58990 48512
rect 59046 48456 60000 48512
rect 58985 48454 60000 48456
rect 58985 48451 59051 48454
rect 4210 48448 4526 48449
rect 4210 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4526 48448
rect 4210 48383 4526 48384
rect 34930 48448 35246 48449
rect 34930 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35246 48448
rect 59200 48424 60000 48454
rect 34930 48383 35246 48384
rect 0 48242 800 48272
rect 1025 48242 1091 48245
rect 0 48240 1091 48242
rect 0 48184 1030 48240
rect 1086 48184 1091 48240
rect 0 48182 1091 48184
rect 0 48152 800 48182
rect 1025 48179 1091 48182
rect 58985 48106 59051 48109
rect 59200 48106 60000 48136
rect 58985 48104 60000 48106
rect 58985 48048 58990 48104
rect 59046 48048 60000 48104
rect 58985 48046 60000 48048
rect 58985 48043 59051 48046
rect 59200 48016 60000 48046
rect 19570 47904 19886 47905
rect 19570 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19886 47904
rect 19570 47839 19886 47840
rect 50290 47904 50606 47905
rect 50290 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50606 47904
rect 50290 47839 50606 47840
rect 0 47698 800 47728
rect 933 47698 999 47701
rect 0 47696 999 47698
rect 0 47640 938 47696
rect 994 47640 999 47696
rect 0 47638 999 47640
rect 0 47608 800 47638
rect 933 47635 999 47638
rect 58801 47698 58867 47701
rect 59200 47698 60000 47728
rect 58801 47696 60000 47698
rect 58801 47640 58806 47696
rect 58862 47640 60000 47696
rect 58801 47638 60000 47640
rect 58801 47635 58867 47638
rect 59200 47608 60000 47638
rect 4210 47360 4526 47361
rect 4210 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4526 47360
rect 4210 47295 4526 47296
rect 34930 47360 35246 47361
rect 34930 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35246 47360
rect 34930 47295 35246 47296
rect 58985 47290 59051 47293
rect 59200 47290 60000 47320
rect 58985 47288 60000 47290
rect 58985 47232 58990 47288
rect 59046 47232 60000 47288
rect 58985 47230 60000 47232
rect 58985 47227 59051 47230
rect 59200 47200 60000 47230
rect 0 47154 800 47184
rect 1025 47154 1091 47157
rect 0 47152 1091 47154
rect 0 47096 1030 47152
rect 1086 47096 1091 47152
rect 0 47094 1091 47096
rect 0 47064 800 47094
rect 1025 47091 1091 47094
rect 58893 46882 58959 46885
rect 59200 46882 60000 46912
rect 58893 46880 60000 46882
rect 58893 46824 58898 46880
rect 58954 46824 60000 46880
rect 58893 46822 60000 46824
rect 58893 46819 58959 46822
rect 19570 46816 19886 46817
rect 19570 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19886 46816
rect 19570 46751 19886 46752
rect 50290 46816 50606 46817
rect 50290 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50606 46816
rect 59200 46792 60000 46822
rect 50290 46751 50606 46752
rect 0 46610 800 46640
rect 933 46610 999 46613
rect 0 46608 999 46610
rect 0 46552 938 46608
rect 994 46552 999 46608
rect 0 46550 999 46552
rect 0 46520 800 46550
rect 933 46547 999 46550
rect 58985 46474 59051 46477
rect 59200 46474 60000 46504
rect 58985 46472 60000 46474
rect 58985 46416 58990 46472
rect 59046 46416 60000 46472
rect 58985 46414 60000 46416
rect 58985 46411 59051 46414
rect 59200 46384 60000 46414
rect 4210 46272 4526 46273
rect 4210 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4526 46272
rect 4210 46207 4526 46208
rect 34930 46272 35246 46273
rect 34930 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35246 46272
rect 34930 46207 35246 46208
rect 0 46066 800 46096
rect 1025 46066 1091 46069
rect 0 46064 1091 46066
rect 0 46008 1030 46064
rect 1086 46008 1091 46064
rect 0 46006 1091 46008
rect 0 45976 800 46006
rect 1025 46003 1091 46006
rect 58985 46066 59051 46069
rect 59200 46066 60000 46096
rect 58985 46064 60000 46066
rect 58985 46008 58990 46064
rect 59046 46008 60000 46064
rect 58985 46006 60000 46008
rect 58985 46003 59051 46006
rect 59200 45976 60000 46006
rect 19570 45728 19886 45729
rect 19570 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19886 45728
rect 19570 45663 19886 45664
rect 50290 45728 50606 45729
rect 50290 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50606 45728
rect 50290 45663 50606 45664
rect 58157 45658 58223 45661
rect 59200 45658 60000 45688
rect 58157 45656 60000 45658
rect 58157 45600 58162 45656
rect 58218 45600 60000 45656
rect 58157 45598 60000 45600
rect 58157 45595 58223 45598
rect 59200 45568 60000 45598
rect 0 45522 800 45552
rect 933 45522 999 45525
rect 0 45520 999 45522
rect 0 45464 938 45520
rect 994 45464 999 45520
rect 0 45462 999 45464
rect 0 45432 800 45462
rect 933 45459 999 45462
rect 32673 45522 32739 45525
rect 40534 45522 40540 45524
rect 32673 45520 40540 45522
rect 32673 45464 32678 45520
rect 32734 45464 40540 45520
rect 32673 45462 40540 45464
rect 32673 45459 32739 45462
rect 40534 45460 40540 45462
rect 40604 45460 40610 45524
rect 58985 45250 59051 45253
rect 59200 45250 60000 45280
rect 58985 45248 60000 45250
rect 58985 45192 58990 45248
rect 59046 45192 60000 45248
rect 58985 45190 60000 45192
rect 58985 45187 59051 45190
rect 4210 45184 4526 45185
rect 4210 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4526 45184
rect 4210 45119 4526 45120
rect 34930 45184 35246 45185
rect 34930 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35246 45184
rect 59200 45160 60000 45190
rect 34930 45119 35246 45120
rect 0 44978 800 45008
rect 1025 44978 1091 44981
rect 0 44976 1091 44978
rect 0 44920 1030 44976
rect 1086 44920 1091 44976
rect 0 44918 1091 44920
rect 0 44888 800 44918
rect 1025 44915 1091 44918
rect 58893 44842 58959 44845
rect 59200 44842 60000 44872
rect 58893 44840 60000 44842
rect 58893 44784 58898 44840
rect 58954 44784 60000 44840
rect 58893 44782 60000 44784
rect 58893 44779 58959 44782
rect 59200 44752 60000 44782
rect 19570 44640 19886 44641
rect 19570 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19886 44640
rect 19570 44575 19886 44576
rect 50290 44640 50606 44641
rect 50290 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50606 44640
rect 50290 44575 50606 44576
rect 0 44434 800 44464
rect 933 44434 999 44437
rect 0 44432 999 44434
rect 0 44376 938 44432
rect 994 44376 999 44432
rect 0 44374 999 44376
rect 0 44344 800 44374
rect 933 44371 999 44374
rect 58157 44434 58223 44437
rect 59200 44434 60000 44464
rect 58157 44432 60000 44434
rect 58157 44376 58162 44432
rect 58218 44376 60000 44432
rect 58157 44374 60000 44376
rect 58157 44371 58223 44374
rect 59200 44344 60000 44374
rect 48681 44300 48747 44301
rect 48630 44298 48636 44300
rect 48590 44238 48636 44298
rect 48700 44296 48747 44300
rect 48742 44240 48747 44296
rect 48630 44236 48636 44238
rect 48700 44236 48747 44240
rect 48681 44235 48747 44236
rect 4210 44096 4526 44097
rect 4210 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4526 44096
rect 4210 44031 4526 44032
rect 34930 44096 35246 44097
rect 34930 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35246 44096
rect 34930 44031 35246 44032
rect 58985 44026 59051 44029
rect 59200 44026 60000 44056
rect 58985 44024 60000 44026
rect 58985 43968 58990 44024
rect 59046 43968 60000 44024
rect 58985 43966 60000 43968
rect 58985 43963 59051 43966
rect 59200 43936 60000 43966
rect 0 43890 800 43920
rect 1025 43890 1091 43893
rect 0 43888 1091 43890
rect 0 43832 1030 43888
rect 1086 43832 1091 43888
rect 0 43830 1091 43832
rect 0 43800 800 43830
rect 1025 43827 1091 43830
rect 58065 43618 58131 43621
rect 59200 43618 60000 43648
rect 58065 43616 60000 43618
rect 58065 43560 58070 43616
rect 58126 43560 60000 43616
rect 58065 43558 60000 43560
rect 58065 43555 58131 43558
rect 19570 43552 19886 43553
rect 19570 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19886 43552
rect 19570 43487 19886 43488
rect 50290 43552 50606 43553
rect 50290 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50606 43552
rect 59200 43528 60000 43558
rect 50290 43487 50606 43488
rect 0 43346 800 43376
rect 933 43346 999 43349
rect 0 43344 999 43346
rect 0 43288 938 43344
rect 994 43288 999 43344
rect 0 43286 999 43288
rect 0 43256 800 43286
rect 933 43283 999 43286
rect 58893 43210 58959 43213
rect 59200 43210 60000 43240
rect 58893 43208 60000 43210
rect 58893 43152 58898 43208
rect 58954 43152 60000 43208
rect 58893 43150 60000 43152
rect 58893 43147 58959 43150
rect 59200 43120 60000 43150
rect 4210 43008 4526 43009
rect 4210 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4526 43008
rect 4210 42943 4526 42944
rect 34930 43008 35246 43009
rect 34930 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35246 43008
rect 34930 42943 35246 42944
rect 41321 42940 41387 42941
rect 41270 42938 41276 42940
rect 41230 42878 41276 42938
rect 41340 42936 41387 42940
rect 41382 42880 41387 42936
rect 41270 42876 41276 42878
rect 41340 42876 41387 42880
rect 41321 42875 41387 42876
rect 0 42802 800 42832
rect 1025 42802 1091 42805
rect 0 42800 1091 42802
rect 0 42744 1030 42800
rect 1086 42744 1091 42800
rect 0 42742 1091 42744
rect 0 42712 800 42742
rect 1025 42739 1091 42742
rect 58985 42802 59051 42805
rect 59200 42802 60000 42832
rect 58985 42800 60000 42802
rect 58985 42744 58990 42800
rect 59046 42744 60000 42800
rect 58985 42742 60000 42744
rect 58985 42739 59051 42742
rect 59200 42712 60000 42742
rect 19570 42464 19886 42465
rect 19570 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19886 42464
rect 19570 42399 19886 42400
rect 50290 42464 50606 42465
rect 50290 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50606 42464
rect 50290 42399 50606 42400
rect 58341 42394 58407 42397
rect 59200 42394 60000 42424
rect 58341 42392 60000 42394
rect 58341 42336 58346 42392
rect 58402 42336 60000 42392
rect 58341 42334 60000 42336
rect 58341 42331 58407 42334
rect 59200 42304 60000 42334
rect 0 42258 800 42288
rect 933 42258 999 42261
rect 0 42256 999 42258
rect 0 42200 938 42256
rect 994 42200 999 42256
rect 0 42198 999 42200
rect 0 42168 800 42198
rect 933 42195 999 42198
rect 4210 41920 4526 41921
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 34930 41920 35246 41921
rect 34930 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35246 41920
rect 59200 41896 60000 42016
rect 34930 41855 35246 41856
rect 0 41714 800 41744
rect 1025 41714 1091 41717
rect 0 41712 1091 41714
rect 0 41656 1030 41712
rect 1086 41656 1091 41712
rect 0 41654 1091 41656
rect 0 41624 800 41654
rect 1025 41651 1091 41654
rect 59200 41488 60000 41608
rect 43069 41442 43135 41445
rect 44398 41442 44404 41444
rect 43069 41440 44404 41442
rect 43069 41384 43074 41440
rect 43130 41384 44404 41440
rect 43069 41382 44404 41384
rect 43069 41379 43135 41382
rect 44398 41380 44404 41382
rect 44468 41380 44474 41444
rect 19570 41376 19886 41377
rect 19570 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19886 41376
rect 19570 41311 19886 41312
rect 50290 41376 50606 41377
rect 50290 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50606 41376
rect 50290 41311 50606 41312
rect 0 41170 800 41200
rect 933 41170 999 41173
rect 0 41168 999 41170
rect 0 41112 938 41168
rect 994 41112 999 41168
rect 0 41110 999 41112
rect 0 41080 800 41110
rect 933 41107 999 41110
rect 58985 41170 59051 41173
rect 59200 41170 60000 41200
rect 58985 41168 60000 41170
rect 58985 41112 58990 41168
rect 59046 41112 60000 41168
rect 58985 41110 60000 41112
rect 58985 41107 59051 41110
rect 59200 41080 60000 41110
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 34930 40832 35246 40833
rect 34930 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35246 40832
rect 34930 40767 35246 40768
rect 59200 40672 60000 40792
rect 0 40626 800 40656
rect 1025 40626 1091 40629
rect 0 40624 1091 40626
rect 0 40568 1030 40624
rect 1086 40568 1091 40624
rect 0 40566 1091 40568
rect 0 40536 800 40566
rect 1025 40563 1091 40566
rect 19570 40288 19886 40289
rect 19570 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19886 40288
rect 19570 40223 19886 40224
rect 50290 40288 50606 40289
rect 50290 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50606 40288
rect 59200 40264 60000 40384
rect 50290 40223 50606 40224
rect 0 40082 800 40112
rect 933 40082 999 40085
rect 0 40080 999 40082
rect 0 40024 938 40080
rect 994 40024 999 40080
rect 0 40022 999 40024
rect 0 39992 800 40022
rect 933 40019 999 40022
rect 58341 39946 58407 39949
rect 59200 39946 60000 39976
rect 58341 39944 60000 39946
rect 58341 39888 58346 39944
rect 58402 39888 60000 39944
rect 58341 39886 60000 39888
rect 58341 39883 58407 39886
rect 59200 39856 60000 39886
rect 4210 39744 4526 39745
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 34930 39744 35246 39745
rect 34930 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35246 39744
rect 34930 39679 35246 39680
rect 0 39538 800 39568
rect 1025 39538 1091 39541
rect 0 39536 1091 39538
rect 0 39480 1030 39536
rect 1086 39480 1091 39536
rect 0 39478 1091 39480
rect 0 39448 800 39478
rect 1025 39475 1091 39478
rect 59200 39448 60000 39568
rect 19570 39200 19886 39201
rect 19570 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19886 39200
rect 19570 39135 19886 39136
rect 50290 39200 50606 39201
rect 50290 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50606 39200
rect 50290 39135 50606 39136
rect 59200 39040 60000 39160
rect 0 38994 800 39024
rect 933 38994 999 38997
rect 0 38992 999 38994
rect 0 38936 938 38992
rect 994 38936 999 38992
rect 0 38934 999 38936
rect 0 38904 800 38934
rect 933 38931 999 38934
rect 58341 38722 58407 38725
rect 59200 38722 60000 38752
rect 58341 38720 60000 38722
rect 58341 38664 58346 38720
rect 58402 38664 60000 38720
rect 58341 38662 60000 38664
rect 58341 38659 58407 38662
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 59200 38632 60000 38662
rect 34930 38591 35246 38592
rect 0 38450 800 38480
rect 1025 38450 1091 38453
rect 0 38448 1091 38450
rect 0 38392 1030 38448
rect 1086 38392 1091 38448
rect 0 38390 1091 38392
rect 0 38360 800 38390
rect 1025 38387 1091 38390
rect 59200 38224 60000 38344
rect 19570 38112 19886 38113
rect 19570 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19886 38112
rect 19570 38047 19886 38048
rect 50290 38112 50606 38113
rect 50290 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50606 38112
rect 50290 38047 50606 38048
rect 0 37906 800 37936
rect 933 37906 999 37909
rect 0 37904 999 37906
rect 0 37848 938 37904
rect 994 37848 999 37904
rect 0 37846 999 37848
rect 0 37816 800 37846
rect 933 37843 999 37846
rect 59200 37816 60000 37936
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 58985 37498 59051 37501
rect 59200 37498 60000 37528
rect 58985 37496 60000 37498
rect 58985 37440 58990 37496
rect 59046 37440 60000 37496
rect 58985 37438 60000 37440
rect 58985 37435 59051 37438
rect 59200 37408 60000 37438
rect 0 37362 800 37392
rect 1025 37362 1091 37365
rect 0 37360 1091 37362
rect 0 37304 1030 37360
rect 1086 37304 1091 37360
rect 0 37302 1091 37304
rect 0 37272 800 37302
rect 1025 37299 1091 37302
rect 58065 37090 58131 37093
rect 59200 37090 60000 37120
rect 58065 37088 60000 37090
rect 58065 37032 58070 37088
rect 58126 37032 60000 37088
rect 58065 37030 60000 37032
rect 58065 37027 58131 37030
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 50290 37024 50606 37025
rect 50290 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50606 37024
rect 59200 37000 60000 37030
rect 50290 36959 50606 36960
rect 0 36818 800 36848
rect 933 36818 999 36821
rect 0 36816 999 36818
rect 0 36760 938 36816
rect 994 36760 999 36816
rect 0 36758 999 36760
rect 0 36728 800 36758
rect 933 36755 999 36758
rect 59200 36592 60000 36712
rect 35341 36546 35407 36549
rect 41454 36546 41460 36548
rect 35341 36544 41460 36546
rect 35341 36488 35346 36544
rect 35402 36488 41460 36544
rect 35341 36486 41460 36488
rect 35341 36483 35407 36486
rect 41454 36484 41460 36486
rect 41524 36484 41530 36548
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 0 36274 800 36304
rect 1025 36274 1091 36277
rect 0 36272 1091 36274
rect 0 36216 1030 36272
rect 1086 36216 1091 36272
rect 0 36214 1091 36216
rect 0 36184 800 36214
rect 1025 36211 1091 36214
rect 58157 36274 58223 36277
rect 59200 36274 60000 36304
rect 58157 36272 60000 36274
rect 58157 36216 58162 36272
rect 58218 36216 60000 36272
rect 58157 36214 60000 36216
rect 58157 36211 58223 36214
rect 59200 36184 60000 36214
rect 30465 36004 30531 36005
rect 30414 36002 30420 36004
rect 30374 35942 30420 36002
rect 30484 36000 30531 36004
rect 30526 35944 30531 36000
rect 30414 35940 30420 35942
rect 30484 35940 30531 35944
rect 30465 35939 30531 35940
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 50290 35936 50606 35937
rect 50290 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50606 35936
rect 50290 35871 50606 35872
rect 58157 35866 58223 35869
rect 59200 35866 60000 35896
rect 58157 35864 60000 35866
rect 58157 35808 58162 35864
rect 58218 35808 60000 35864
rect 58157 35806 60000 35808
rect 58157 35803 58223 35806
rect 59200 35776 60000 35806
rect 0 35730 800 35760
rect 933 35730 999 35733
rect 0 35728 999 35730
rect 0 35672 938 35728
rect 994 35672 999 35728
rect 0 35670 999 35672
rect 0 35640 800 35670
rect 933 35667 999 35670
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 59200 35368 60000 35488
rect 34930 35327 35246 35328
rect 0 35186 800 35216
rect 1025 35186 1091 35189
rect 0 35184 1091 35186
rect 0 35128 1030 35184
rect 1086 35128 1091 35184
rect 0 35126 1091 35128
rect 0 35096 800 35126
rect 1025 35123 1091 35126
rect 58157 35050 58223 35053
rect 59200 35050 60000 35080
rect 58157 35048 60000 35050
rect 58157 34992 58162 35048
rect 58218 34992 60000 35048
rect 58157 34990 60000 34992
rect 58157 34987 58223 34990
rect 59200 34960 60000 34990
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 50290 34848 50606 34849
rect 50290 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50606 34848
rect 50290 34783 50606 34784
rect 0 34642 800 34672
rect 933 34642 999 34645
rect 0 34640 999 34642
rect 0 34584 938 34640
rect 994 34584 999 34640
rect 0 34582 999 34584
rect 0 34552 800 34582
rect 933 34579 999 34582
rect 30741 34644 30807 34645
rect 30741 34640 30788 34644
rect 30852 34642 30858 34644
rect 58065 34642 58131 34645
rect 59200 34642 60000 34672
rect 30741 34584 30746 34640
rect 30741 34580 30788 34584
rect 30852 34582 30898 34642
rect 58065 34640 60000 34642
rect 58065 34584 58070 34640
rect 58126 34584 60000 34640
rect 58065 34582 60000 34584
rect 30852 34580 30858 34582
rect 30741 34579 30807 34580
rect 58065 34579 58131 34582
rect 59200 34552 60000 34582
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 59200 34144 60000 34264
rect 0 34098 800 34128
rect 1025 34098 1091 34101
rect 0 34096 1091 34098
rect 0 34040 1030 34096
rect 1086 34040 1091 34096
rect 0 34038 1091 34040
rect 0 34008 800 34038
rect 1025 34035 1091 34038
rect 58157 33826 58223 33829
rect 59200 33826 60000 33856
rect 58157 33824 60000 33826
rect 58157 33768 58162 33824
rect 58218 33768 60000 33824
rect 58157 33766 60000 33768
rect 58157 33763 58223 33766
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 50290 33760 50606 33761
rect 50290 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50606 33760
rect 59200 33736 60000 33766
rect 50290 33695 50606 33696
rect 0 33554 800 33584
rect 933 33554 999 33557
rect 0 33552 999 33554
rect 0 33496 938 33552
rect 994 33496 999 33552
rect 0 33494 999 33496
rect 0 33464 800 33494
rect 933 33491 999 33494
rect 58065 33418 58131 33421
rect 59200 33418 60000 33448
rect 58065 33416 60000 33418
rect 58065 33360 58070 33416
rect 58126 33360 60000 33416
rect 58065 33358 60000 33360
rect 58065 33355 58131 33358
rect 59200 33328 60000 33358
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 0 33010 800 33040
rect 1025 33010 1091 33013
rect 0 33008 1091 33010
rect 0 32952 1030 33008
rect 1086 32952 1091 33008
rect 0 32950 1091 32952
rect 0 32920 800 32950
rect 1025 32947 1091 32950
rect 59200 32920 60000 33040
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 50290 32672 50606 32673
rect 50290 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50606 32672
rect 50290 32607 50606 32608
rect 58157 32602 58223 32605
rect 59200 32602 60000 32632
rect 58157 32600 60000 32602
rect 58157 32544 58162 32600
rect 58218 32544 60000 32600
rect 58157 32542 60000 32544
rect 58157 32539 58223 32542
rect 59200 32512 60000 32542
rect 0 32466 800 32496
rect 933 32466 999 32469
rect 0 32464 999 32466
rect 0 32408 938 32464
rect 994 32408 999 32464
rect 0 32406 999 32408
rect 0 32376 800 32406
rect 933 32403 999 32406
rect 27613 32466 27679 32469
rect 39246 32466 39252 32468
rect 27613 32464 39252 32466
rect 27613 32408 27618 32464
rect 27674 32408 39252 32464
rect 27613 32406 39252 32408
rect 27613 32403 27679 32406
rect 39246 32404 39252 32406
rect 39316 32404 39322 32468
rect 27797 32330 27863 32333
rect 28441 32330 28507 32333
rect 27797 32328 28507 32330
rect 27797 32272 27802 32328
rect 27858 32272 28446 32328
rect 28502 32272 28507 32328
rect 27797 32270 28507 32272
rect 27797 32267 27863 32270
rect 28441 32267 28507 32270
rect 28073 32194 28139 32197
rect 28625 32194 28691 32197
rect 28073 32192 28691 32194
rect 28073 32136 28078 32192
rect 28134 32136 28630 32192
rect 28686 32136 28691 32192
rect 28073 32134 28691 32136
rect 28073 32131 28139 32134
rect 28625 32131 28691 32134
rect 58065 32194 58131 32197
rect 59200 32194 60000 32224
rect 58065 32192 60000 32194
rect 58065 32136 58070 32192
rect 58126 32136 60000 32192
rect 58065 32134 60000 32136
rect 58065 32131 58131 32134
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 59200 32104 60000 32134
rect 34930 32063 35246 32064
rect 29545 32060 29611 32061
rect 29494 32058 29500 32060
rect 29454 31998 29500 32058
rect 29564 32056 29611 32060
rect 29606 32000 29611 32056
rect 29494 31996 29500 31998
rect 29564 31996 29611 32000
rect 29545 31995 29611 31996
rect 0 31922 800 31952
rect 933 31922 999 31925
rect 0 31920 999 31922
rect 0 31864 938 31920
rect 994 31864 999 31920
rect 0 31862 999 31864
rect 0 31832 800 31862
rect 933 31859 999 31862
rect 36813 31786 36879 31789
rect 37774 31786 37780 31788
rect 36813 31784 37780 31786
rect 36813 31728 36818 31784
rect 36874 31728 37780 31784
rect 36813 31726 37780 31728
rect 36813 31723 36879 31726
rect 37774 31724 37780 31726
rect 37844 31724 37850 31788
rect 58985 31786 59051 31789
rect 59200 31786 60000 31816
rect 58985 31784 60000 31786
rect 58985 31728 58990 31784
rect 59046 31728 60000 31784
rect 58985 31726 60000 31728
rect 58985 31723 59051 31726
rect 59200 31696 60000 31726
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 50290 31584 50606 31585
rect 50290 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50606 31584
rect 50290 31519 50606 31520
rect 0 31378 800 31408
rect 1025 31378 1091 31381
rect 0 31376 1091 31378
rect 0 31320 1030 31376
rect 1086 31320 1091 31376
rect 0 31318 1091 31320
rect 0 31288 800 31318
rect 1025 31315 1091 31318
rect 58893 31378 58959 31381
rect 59200 31378 60000 31408
rect 58893 31376 60000 31378
rect 58893 31320 58898 31376
rect 58954 31320 60000 31376
rect 58893 31318 60000 31320
rect 58893 31315 58959 31318
rect 59200 31288 60000 31318
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 58065 30970 58131 30973
rect 59200 30970 60000 31000
rect 58065 30968 60000 30970
rect 58065 30912 58070 30968
rect 58126 30912 60000 30968
rect 58065 30910 60000 30912
rect 58065 30907 58131 30910
rect 59200 30880 60000 30910
rect 0 30834 800 30864
rect 933 30834 999 30837
rect 0 30832 999 30834
rect 0 30776 938 30832
rect 994 30776 999 30832
rect 0 30774 999 30776
rect 0 30744 800 30774
rect 933 30771 999 30774
rect 58157 30562 58223 30565
rect 59200 30562 60000 30592
rect 58157 30560 60000 30562
rect 58157 30504 58162 30560
rect 58218 30504 60000 30560
rect 58157 30502 60000 30504
rect 58157 30499 58223 30502
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 50290 30496 50606 30497
rect 50290 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50606 30496
rect 59200 30472 60000 30502
rect 50290 30431 50606 30432
rect 0 30290 800 30320
rect 933 30290 999 30293
rect 0 30288 999 30290
rect 0 30232 938 30288
rect 994 30232 999 30288
rect 0 30230 999 30232
rect 0 30200 800 30230
rect 933 30227 999 30230
rect 58157 30154 58223 30157
rect 59200 30154 60000 30184
rect 58157 30152 60000 30154
rect 58157 30096 58162 30152
rect 58218 30096 60000 30152
rect 58157 30094 60000 30096
rect 58157 30091 58223 30094
rect 59200 30064 60000 30094
rect 22277 30018 22343 30021
rect 28441 30018 28507 30021
rect 22277 30016 28507 30018
rect 22277 29960 22282 30016
rect 22338 29960 28446 30016
rect 28502 29960 28507 30016
rect 22277 29958 28507 29960
rect 22277 29955 22343 29958
rect 28441 29955 28507 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 0 29746 800 29776
rect 933 29746 999 29749
rect 0 29744 999 29746
rect 0 29688 938 29744
rect 994 29688 999 29744
rect 0 29686 999 29688
rect 0 29656 800 29686
rect 933 29683 999 29686
rect 28717 29746 28783 29749
rect 46238 29746 46244 29748
rect 28717 29744 46244 29746
rect 28717 29688 28722 29744
rect 28778 29688 46244 29744
rect 28717 29686 46244 29688
rect 28717 29683 28783 29686
rect 46238 29684 46244 29686
rect 46308 29684 46314 29748
rect 58065 29746 58131 29749
rect 59200 29746 60000 29776
rect 58065 29744 60000 29746
rect 58065 29688 58070 29744
rect 58126 29688 60000 29744
rect 58065 29686 60000 29688
rect 58065 29683 58131 29686
rect 59200 29656 60000 29686
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 50290 29408 50606 29409
rect 50290 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50606 29408
rect 50290 29343 50606 29344
rect 22277 29338 22343 29341
rect 23565 29338 23631 29341
rect 22277 29336 23631 29338
rect 22277 29280 22282 29336
rect 22338 29280 23570 29336
rect 23626 29280 23631 29336
rect 22277 29278 23631 29280
rect 22277 29275 22343 29278
rect 23565 29275 23631 29278
rect 58065 29338 58131 29341
rect 59200 29338 60000 29368
rect 58065 29336 60000 29338
rect 58065 29280 58070 29336
rect 58126 29280 60000 29336
rect 58065 29278 60000 29280
rect 58065 29275 58131 29278
rect 59200 29248 60000 29278
rect 0 29202 800 29232
rect 1025 29202 1091 29205
rect 0 29200 1091 29202
rect 0 29144 1030 29200
rect 1086 29144 1091 29200
rect 0 29142 1091 29144
rect 0 29112 800 29142
rect 1025 29139 1091 29142
rect 23197 29066 23263 29069
rect 23657 29066 23723 29069
rect 23197 29064 23723 29066
rect 23197 29008 23202 29064
rect 23258 29008 23662 29064
rect 23718 29008 23723 29064
rect 23197 29006 23723 29008
rect 23197 29003 23263 29006
rect 23657 29003 23723 29006
rect 36537 29066 36603 29069
rect 44766 29066 44772 29068
rect 36537 29064 44772 29066
rect 36537 29008 36542 29064
rect 36598 29008 44772 29064
rect 36537 29006 44772 29008
rect 36537 29003 36603 29006
rect 44766 29004 44772 29006
rect 44836 29004 44842 29068
rect 58157 28930 58223 28933
rect 59200 28930 60000 28960
rect 58157 28928 60000 28930
rect 58157 28872 58162 28928
rect 58218 28872 60000 28928
rect 58157 28870 60000 28872
rect 58157 28867 58223 28870
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 59200 28840 60000 28870
rect 34930 28799 35246 28800
rect 0 28658 800 28688
rect 933 28658 999 28661
rect 0 28656 999 28658
rect 0 28600 938 28656
rect 994 28600 999 28656
rect 0 28598 999 28600
rect 0 28568 800 28598
rect 933 28595 999 28598
rect 58065 28522 58131 28525
rect 59200 28522 60000 28552
rect 58065 28520 60000 28522
rect 58065 28464 58070 28520
rect 58126 28464 60000 28520
rect 58065 28462 60000 28464
rect 58065 28459 58131 28462
rect 59200 28432 60000 28462
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 50290 28320 50606 28321
rect 50290 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50606 28320
rect 50290 28255 50606 28256
rect 0 28114 800 28144
rect 933 28114 999 28117
rect 0 28112 999 28114
rect 0 28056 938 28112
rect 994 28056 999 28112
rect 0 28054 999 28056
rect 0 28024 800 28054
rect 933 28051 999 28054
rect 29637 28114 29703 28117
rect 29913 28114 29979 28117
rect 31109 28114 31175 28117
rect 29637 28112 31175 28114
rect 29637 28056 29642 28112
rect 29698 28056 29918 28112
rect 29974 28056 31114 28112
rect 31170 28056 31175 28112
rect 29637 28054 31175 28056
rect 29637 28051 29703 28054
rect 29913 28051 29979 28054
rect 31109 28051 31175 28054
rect 59200 28024 60000 28144
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 58985 27706 59051 27709
rect 59200 27706 60000 27736
rect 58985 27704 60000 27706
rect 58985 27648 58990 27704
rect 59046 27648 60000 27704
rect 58985 27646 60000 27648
rect 58985 27643 59051 27646
rect 59200 27616 60000 27646
rect 0 27570 800 27600
rect 933 27570 999 27573
rect 0 27568 999 27570
rect 0 27512 938 27568
rect 994 27512 999 27568
rect 0 27510 999 27512
rect 0 27480 800 27510
rect 933 27507 999 27510
rect 26969 27434 27035 27437
rect 28441 27434 28507 27437
rect 26969 27432 28507 27434
rect 26969 27376 26974 27432
rect 27030 27376 28446 27432
rect 28502 27376 28507 27432
rect 26969 27374 28507 27376
rect 26969 27371 27035 27374
rect 28441 27371 28507 27374
rect 58157 27298 58223 27301
rect 59200 27298 60000 27328
rect 58157 27296 60000 27298
rect 58157 27240 58162 27296
rect 58218 27240 60000 27296
rect 58157 27238 60000 27240
rect 58157 27235 58223 27238
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 50290 27232 50606 27233
rect 50290 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50606 27232
rect 59200 27208 60000 27238
rect 50290 27167 50606 27168
rect 26049 27162 26115 27165
rect 28625 27162 28691 27165
rect 26049 27160 28691 27162
rect 26049 27104 26054 27160
rect 26110 27104 28630 27160
rect 28686 27104 28691 27160
rect 26049 27102 28691 27104
rect 26049 27099 26115 27102
rect 28625 27099 28691 27102
rect 0 27026 800 27056
rect 933 27026 999 27029
rect 0 27024 999 27026
rect 0 26968 938 27024
rect 994 26968 999 27024
rect 0 26966 999 26968
rect 0 26936 800 26966
rect 933 26963 999 26966
rect 23013 27026 23079 27029
rect 26417 27026 26483 27029
rect 23013 27024 26483 27026
rect 23013 26968 23018 27024
rect 23074 26968 26422 27024
rect 26478 26968 26483 27024
rect 23013 26966 26483 26968
rect 23013 26963 23079 26966
rect 26417 26963 26483 26966
rect 30557 27026 30623 27029
rect 32029 27026 32095 27029
rect 30557 27024 32095 27026
rect 30557 26968 30562 27024
rect 30618 26968 32034 27024
rect 32090 26968 32095 27024
rect 30557 26966 32095 26968
rect 30557 26963 30623 26966
rect 32029 26963 32095 26966
rect 59200 26800 60000 26920
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 0 26482 800 26512
rect 1025 26482 1091 26485
rect 0 26480 1091 26482
rect 0 26424 1030 26480
rect 1086 26424 1091 26480
rect 0 26422 1091 26424
rect 0 26392 800 26422
rect 1025 26419 1091 26422
rect 31661 26482 31727 26485
rect 33133 26482 33199 26485
rect 31661 26480 33199 26482
rect 31661 26424 31666 26480
rect 31722 26424 33138 26480
rect 33194 26424 33199 26480
rect 31661 26422 33199 26424
rect 31661 26419 31727 26422
rect 33133 26419 33199 26422
rect 58157 26482 58223 26485
rect 59200 26482 60000 26512
rect 58157 26480 60000 26482
rect 58157 26424 58162 26480
rect 58218 26424 60000 26480
rect 58157 26422 60000 26424
rect 58157 26419 58223 26422
rect 59200 26392 60000 26422
rect 33777 26348 33843 26349
rect 33726 26346 33732 26348
rect 33686 26286 33732 26346
rect 33796 26344 33843 26348
rect 33838 26288 33843 26344
rect 33726 26284 33732 26286
rect 33796 26284 33843 26288
rect 33777 26283 33843 26284
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 50290 26144 50606 26145
rect 50290 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50606 26144
rect 50290 26079 50606 26080
rect 58157 26074 58223 26077
rect 59200 26074 60000 26104
rect 58157 26072 60000 26074
rect 58157 26016 58162 26072
rect 58218 26016 60000 26072
rect 58157 26014 60000 26016
rect 58157 26011 58223 26014
rect 59200 25984 60000 26014
rect 0 25938 800 25968
rect 933 25938 999 25941
rect 0 25936 999 25938
rect 0 25880 938 25936
rect 994 25880 999 25936
rect 0 25878 999 25880
rect 0 25848 800 25878
rect 933 25875 999 25878
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 59200 25576 60000 25696
rect 34930 25535 35246 25536
rect 0 25394 800 25424
rect 933 25394 999 25397
rect 0 25392 999 25394
rect 0 25336 938 25392
rect 994 25336 999 25392
rect 0 25334 999 25336
rect 0 25304 800 25334
rect 933 25331 999 25334
rect 45921 25258 45987 25261
rect 46933 25258 46999 25261
rect 47117 25258 47183 25261
rect 45921 25256 47183 25258
rect 45921 25200 45926 25256
rect 45982 25200 46938 25256
rect 46994 25200 47122 25256
rect 47178 25200 47183 25256
rect 45921 25198 47183 25200
rect 45921 25195 45987 25198
rect 46933 25195 46999 25198
rect 47117 25195 47183 25198
rect 58157 25258 58223 25261
rect 59200 25258 60000 25288
rect 58157 25256 60000 25258
rect 58157 25200 58162 25256
rect 58218 25200 60000 25256
rect 58157 25198 60000 25200
rect 58157 25195 58223 25198
rect 59200 25168 60000 25198
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 50290 25056 50606 25057
rect 50290 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50606 25056
rect 50290 24991 50606 24992
rect 43437 24988 43503 24989
rect 43437 24984 43484 24988
rect 43548 24986 43554 24988
rect 43437 24928 43442 24984
rect 43437 24924 43484 24928
rect 43548 24926 43594 24986
rect 43548 24924 43554 24926
rect 43437 24923 43503 24924
rect 0 24850 800 24880
rect 933 24850 999 24853
rect 0 24848 999 24850
rect 0 24792 938 24848
rect 994 24792 999 24848
rect 0 24790 999 24792
rect 0 24760 800 24790
rect 933 24787 999 24790
rect 58065 24850 58131 24853
rect 59200 24850 60000 24880
rect 58065 24848 60000 24850
rect 58065 24792 58070 24848
rect 58126 24792 60000 24848
rect 58065 24790 60000 24792
rect 58065 24787 58131 24790
rect 59200 24760 60000 24790
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 59200 24352 60000 24472
rect 0 24306 800 24336
rect 933 24306 999 24309
rect 0 24304 999 24306
rect 0 24248 938 24304
rect 994 24248 999 24304
rect 0 24246 999 24248
rect 0 24216 800 24246
rect 933 24243 999 24246
rect 29085 24170 29151 24173
rect 30281 24170 30347 24173
rect 32305 24170 32371 24173
rect 37917 24170 37983 24173
rect 29085 24168 37983 24170
rect 29085 24112 29090 24168
rect 29146 24112 30286 24168
rect 30342 24112 32310 24168
rect 32366 24112 37922 24168
rect 37978 24112 37983 24168
rect 29085 24110 37983 24112
rect 29085 24107 29151 24110
rect 30281 24107 30347 24110
rect 32305 24107 32371 24110
rect 37917 24107 37983 24110
rect 58157 24034 58223 24037
rect 59200 24034 60000 24064
rect 58157 24032 60000 24034
rect 58157 23976 58162 24032
rect 58218 23976 60000 24032
rect 58157 23974 60000 23976
rect 58157 23971 58223 23974
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 50290 23968 50606 23969
rect 50290 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50606 23968
rect 59200 23944 60000 23974
rect 50290 23903 50606 23904
rect 0 23762 800 23792
rect 933 23762 999 23765
rect 0 23760 999 23762
rect 0 23704 938 23760
rect 994 23704 999 23760
rect 0 23702 999 23704
rect 0 23672 800 23702
rect 933 23699 999 23702
rect 58065 23626 58131 23629
rect 59200 23626 60000 23656
rect 58065 23624 60000 23626
rect 58065 23568 58070 23624
rect 58126 23568 60000 23624
rect 58065 23566 60000 23568
rect 58065 23563 58131 23566
rect 59200 23536 60000 23566
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 0 23218 800 23248
rect 933 23218 999 23221
rect 0 23216 999 23218
rect 0 23160 938 23216
rect 994 23160 999 23216
rect 0 23158 999 23160
rect 0 23128 800 23158
rect 933 23155 999 23158
rect 39113 23218 39179 23221
rect 48221 23218 48287 23221
rect 39113 23216 48287 23218
rect 39113 23160 39118 23216
rect 39174 23160 48226 23216
rect 48282 23160 48287 23216
rect 39113 23158 48287 23160
rect 39113 23155 39179 23158
rect 48221 23155 48287 23158
rect 59200 23128 60000 23248
rect 39205 23082 39271 23085
rect 41689 23082 41755 23085
rect 41965 23082 42031 23085
rect 39205 23080 42031 23082
rect 39205 23024 39210 23080
rect 39266 23024 41694 23080
rect 41750 23024 41970 23080
rect 42026 23024 42031 23080
rect 39205 23022 42031 23024
rect 39205 23019 39271 23022
rect 41689 23019 41755 23022
rect 41965 23019 42031 23022
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 50290 22880 50606 22881
rect 50290 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50606 22880
rect 50290 22815 50606 22816
rect 58157 22810 58223 22813
rect 59200 22810 60000 22840
rect 58157 22808 60000 22810
rect 58157 22752 58162 22808
rect 58218 22752 60000 22808
rect 58157 22750 60000 22752
rect 58157 22747 58223 22750
rect 59200 22720 60000 22750
rect 0 22674 800 22704
rect 933 22674 999 22677
rect 0 22672 999 22674
rect 0 22616 938 22672
rect 994 22616 999 22672
rect 0 22614 999 22616
rect 0 22584 800 22614
rect 933 22611 999 22614
rect 39941 22674 40007 22677
rect 42701 22674 42767 22677
rect 44357 22674 44423 22677
rect 39941 22672 44423 22674
rect 39941 22616 39946 22672
rect 40002 22616 42706 22672
rect 42762 22616 44362 22672
rect 44418 22616 44423 22672
rect 39941 22614 44423 22616
rect 39941 22611 40007 22614
rect 42701 22611 42767 22614
rect 44357 22611 44423 22614
rect 42241 22402 42307 22405
rect 42609 22402 42675 22405
rect 42241 22400 42675 22402
rect 42241 22344 42246 22400
rect 42302 22344 42614 22400
rect 42670 22344 42675 22400
rect 42241 22342 42675 22344
rect 42241 22339 42307 22342
rect 42609 22339 42675 22342
rect 58065 22402 58131 22405
rect 59200 22402 60000 22432
rect 58065 22400 60000 22402
rect 58065 22344 58070 22400
rect 58126 22344 60000 22400
rect 58065 22342 60000 22344
rect 58065 22339 58131 22342
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 59200 22312 60000 22342
rect 34930 22271 35246 22272
rect 38745 22266 38811 22269
rect 39389 22266 39455 22269
rect 38745 22264 39455 22266
rect 38745 22208 38750 22264
rect 38806 22208 39394 22264
rect 39450 22208 39455 22264
rect 38745 22206 39455 22208
rect 38745 22203 38811 22206
rect 39389 22203 39455 22206
rect 0 22130 800 22160
rect 933 22130 999 22133
rect 0 22128 999 22130
rect 0 22072 938 22128
rect 994 22072 999 22128
rect 0 22070 999 22072
rect 0 22040 800 22070
rect 933 22067 999 22070
rect 23289 21994 23355 21997
rect 47853 21994 47919 21997
rect 23289 21992 47919 21994
rect 23289 21936 23294 21992
rect 23350 21936 47858 21992
rect 47914 21936 47919 21992
rect 23289 21934 47919 21936
rect 23289 21931 23355 21934
rect 47853 21931 47919 21934
rect 59200 21904 60000 22024
rect 30465 21858 30531 21861
rect 38101 21858 38167 21861
rect 30465 21856 38167 21858
rect 30465 21800 30470 21856
rect 30526 21800 38106 21856
rect 38162 21800 38167 21856
rect 30465 21798 38167 21800
rect 30465 21795 30531 21798
rect 38101 21795 38167 21798
rect 38653 21858 38719 21861
rect 40401 21858 40467 21861
rect 38653 21856 40467 21858
rect 38653 21800 38658 21856
rect 38714 21800 40406 21856
rect 40462 21800 40467 21856
rect 38653 21798 40467 21800
rect 38653 21795 38719 21798
rect 40401 21795 40467 21798
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 50290 21792 50606 21793
rect 50290 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50606 21792
rect 50290 21727 50606 21728
rect 0 21586 800 21616
rect 933 21586 999 21589
rect 0 21584 999 21586
rect 0 21528 938 21584
rect 994 21528 999 21584
rect 0 21526 999 21528
rect 0 21496 800 21526
rect 933 21523 999 21526
rect 29729 21586 29795 21589
rect 31385 21586 31451 21589
rect 29729 21584 31451 21586
rect 29729 21528 29734 21584
rect 29790 21528 31390 21584
rect 31446 21528 31451 21584
rect 29729 21526 31451 21528
rect 29729 21523 29795 21526
rect 31385 21523 31451 21526
rect 58985 21586 59051 21589
rect 59200 21586 60000 21616
rect 58985 21584 60000 21586
rect 58985 21528 58990 21584
rect 59046 21528 60000 21584
rect 58985 21526 60000 21528
rect 58985 21523 59051 21526
rect 59200 21496 60000 21526
rect 30281 21450 30347 21453
rect 36997 21450 37063 21453
rect 46013 21452 46079 21453
rect 46013 21450 46060 21452
rect 30281 21448 37063 21450
rect 30281 21392 30286 21448
rect 30342 21392 37002 21448
rect 37058 21392 37063 21448
rect 30281 21390 37063 21392
rect 45968 21448 46060 21450
rect 45968 21392 46018 21448
rect 45968 21390 46060 21392
rect 30281 21387 30347 21390
rect 36997 21387 37063 21390
rect 46013 21388 46060 21390
rect 46124 21388 46130 21452
rect 48497 21450 48563 21453
rect 48814 21450 48820 21452
rect 48497 21448 48820 21450
rect 48497 21392 48502 21448
rect 48558 21392 48820 21448
rect 48497 21390 48820 21392
rect 46013 21387 46079 21388
rect 48497 21387 48563 21390
rect 48814 21388 48820 21390
rect 48884 21388 48890 21452
rect 42977 21314 43043 21317
rect 48497 21314 48563 21317
rect 42977 21312 48563 21314
rect 42977 21256 42982 21312
rect 43038 21256 48502 21312
rect 48558 21256 48563 21312
rect 42977 21254 48563 21256
rect 42977 21251 43043 21254
rect 48497 21251 48563 21254
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 58065 21178 58131 21181
rect 59200 21178 60000 21208
rect 58065 21176 60000 21178
rect 58065 21120 58070 21176
rect 58126 21120 60000 21176
rect 58065 21118 60000 21120
rect 58065 21115 58131 21118
rect 59200 21088 60000 21118
rect 0 21042 800 21072
rect 933 21042 999 21045
rect 0 21040 999 21042
rect 0 20984 938 21040
rect 994 20984 999 21040
rect 0 20982 999 20984
rect 0 20952 800 20982
rect 933 20979 999 20982
rect 23657 21042 23723 21045
rect 55213 21042 55279 21045
rect 23657 21040 55279 21042
rect 23657 20984 23662 21040
rect 23718 20984 55218 21040
rect 55274 20984 55279 21040
rect 23657 20982 55279 20984
rect 23657 20979 23723 20982
rect 55213 20979 55279 20982
rect 48814 20844 48820 20908
rect 48884 20906 48890 20908
rect 56041 20906 56107 20909
rect 48884 20904 56107 20906
rect 48884 20848 56046 20904
rect 56102 20848 56107 20904
rect 48884 20846 56107 20848
rect 48884 20844 48890 20846
rect 56041 20843 56107 20846
rect 38929 20770 38995 20773
rect 43805 20770 43871 20773
rect 38929 20768 43871 20770
rect 38929 20712 38934 20768
rect 38990 20712 43810 20768
rect 43866 20712 43871 20768
rect 38929 20710 43871 20712
rect 38929 20707 38995 20710
rect 43805 20707 43871 20710
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 50290 20704 50606 20705
rect 50290 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50606 20704
rect 59200 20680 60000 20800
rect 50290 20639 50606 20640
rect 34421 20634 34487 20637
rect 42793 20634 42859 20637
rect 44541 20634 44607 20637
rect 34421 20632 44607 20634
rect 34421 20576 34426 20632
rect 34482 20576 42798 20632
rect 42854 20576 44546 20632
rect 44602 20576 44607 20632
rect 34421 20574 44607 20576
rect 34421 20571 34487 20574
rect 42793 20571 42859 20574
rect 44541 20571 44607 20574
rect 0 20498 800 20528
rect 933 20498 999 20501
rect 0 20496 999 20498
rect 0 20440 938 20496
rect 994 20440 999 20496
rect 0 20438 999 20440
rect 0 20408 800 20438
rect 933 20435 999 20438
rect 35249 20498 35315 20501
rect 40217 20498 40283 20501
rect 35249 20496 40283 20498
rect 35249 20440 35254 20496
rect 35310 20440 40222 20496
rect 40278 20440 40283 20496
rect 35249 20438 40283 20440
rect 35249 20435 35315 20438
rect 40217 20435 40283 20438
rect 46841 20362 46907 20365
rect 48681 20362 48747 20365
rect 56409 20362 56475 20365
rect 46841 20360 56475 20362
rect 46841 20304 46846 20360
rect 46902 20304 48686 20360
rect 48742 20304 56414 20360
rect 56470 20304 56475 20360
rect 46841 20302 56475 20304
rect 46841 20299 46907 20302
rect 48681 20299 48747 20302
rect 56409 20299 56475 20302
rect 58249 20362 58315 20365
rect 59200 20362 60000 20392
rect 58249 20360 60000 20362
rect 58249 20304 58254 20360
rect 58310 20304 60000 20360
rect 58249 20302 60000 20304
rect 58249 20299 58315 20302
rect 59200 20272 60000 20302
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 39573 20090 39639 20093
rect 57605 20090 57671 20093
rect 39573 20088 57671 20090
rect 39573 20032 39578 20088
rect 39634 20032 57610 20088
rect 57666 20032 57671 20088
rect 39573 20030 57671 20032
rect 39573 20027 39639 20030
rect 57605 20027 57671 20030
rect 0 19954 800 19984
rect 933 19954 999 19957
rect 0 19952 999 19954
rect 0 19896 938 19952
rect 994 19896 999 19952
rect 0 19894 999 19896
rect 0 19864 800 19894
rect 933 19891 999 19894
rect 34697 19954 34763 19957
rect 40217 19954 40283 19957
rect 34697 19952 40283 19954
rect 34697 19896 34702 19952
rect 34758 19896 40222 19952
rect 40278 19896 40283 19952
rect 34697 19894 40283 19896
rect 34697 19891 34763 19894
rect 40217 19891 40283 19894
rect 44265 19954 44331 19957
rect 44817 19954 44883 19957
rect 57973 19954 58039 19957
rect 44265 19952 58039 19954
rect 44265 19896 44270 19952
rect 44326 19896 44822 19952
rect 44878 19896 57978 19952
rect 58034 19896 58039 19952
rect 44265 19894 58039 19896
rect 44265 19891 44331 19894
rect 44817 19891 44883 19894
rect 57973 19891 58039 19894
rect 58157 19954 58223 19957
rect 59200 19954 60000 19984
rect 58157 19952 60000 19954
rect 58157 19896 58162 19952
rect 58218 19896 60000 19952
rect 58157 19894 60000 19896
rect 58157 19891 58223 19894
rect 59200 19864 60000 19894
rect 27797 19818 27863 19821
rect 28809 19818 28875 19821
rect 27797 19816 28875 19818
rect 27797 19760 27802 19816
rect 27858 19760 28814 19816
rect 28870 19760 28875 19816
rect 27797 19758 28875 19760
rect 27797 19755 27863 19758
rect 28809 19755 28875 19758
rect 36077 19818 36143 19821
rect 40861 19818 40927 19821
rect 36077 19816 40927 19818
rect 36077 19760 36082 19816
rect 36138 19760 40866 19816
rect 40922 19760 40927 19816
rect 36077 19758 40927 19760
rect 36077 19755 36143 19758
rect 40861 19755 40927 19758
rect 44357 19818 44423 19821
rect 45737 19818 45803 19821
rect 44357 19816 45803 19818
rect 44357 19760 44362 19816
rect 44418 19760 45742 19816
rect 45798 19760 45803 19816
rect 44357 19758 45803 19760
rect 44357 19755 44423 19758
rect 45737 19755 45803 19758
rect 28533 19682 28599 19685
rect 28901 19682 28967 19685
rect 28533 19680 28967 19682
rect 28533 19624 28538 19680
rect 28594 19624 28906 19680
rect 28962 19624 28967 19680
rect 28533 19622 28967 19624
rect 28533 19619 28599 19622
rect 28901 19619 28967 19622
rect 34421 19682 34487 19685
rect 46841 19682 46907 19685
rect 34421 19680 46907 19682
rect 34421 19624 34426 19680
rect 34482 19624 46846 19680
rect 46902 19624 46907 19680
rect 34421 19622 46907 19624
rect 34421 19619 34487 19622
rect 46841 19619 46907 19622
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 50290 19616 50606 19617
rect 50290 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50606 19616
rect 50290 19551 50606 19552
rect 36813 19546 36879 19549
rect 43989 19546 44055 19549
rect 36813 19544 44055 19546
rect 36813 19488 36818 19544
rect 36874 19488 43994 19544
rect 44050 19488 44055 19544
rect 36813 19486 44055 19488
rect 36813 19483 36879 19486
rect 43989 19483 44055 19486
rect 59200 19456 60000 19576
rect 0 19410 800 19440
rect 933 19410 999 19413
rect 0 19408 999 19410
rect 0 19352 938 19408
rect 994 19352 999 19408
rect 0 19350 999 19352
rect 0 19320 800 19350
rect 933 19347 999 19350
rect 58157 19138 58223 19141
rect 59200 19138 60000 19168
rect 58157 19136 60000 19138
rect 58157 19080 58162 19136
rect 58218 19080 60000 19136
rect 58157 19078 60000 19080
rect 58157 19075 58223 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 59200 19048 60000 19078
rect 34930 19007 35246 19008
rect 0 18866 800 18896
rect 1025 18866 1091 18869
rect 0 18864 1091 18866
rect 0 18808 1030 18864
rect 1086 18808 1091 18864
rect 0 18806 1091 18808
rect 0 18776 800 18806
rect 1025 18803 1091 18806
rect 52453 18730 52519 18733
rect 56685 18730 56751 18733
rect 52453 18728 56751 18730
rect 52453 18672 52458 18728
rect 52514 18672 56690 18728
rect 56746 18672 56751 18728
rect 52453 18670 56751 18672
rect 52453 18667 52519 18670
rect 56685 18667 56751 18670
rect 58985 18730 59051 18733
rect 59200 18730 60000 18760
rect 58985 18728 60000 18730
rect 58985 18672 58990 18728
rect 59046 18672 60000 18728
rect 58985 18670 60000 18672
rect 58985 18667 59051 18670
rect 59200 18640 60000 18670
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 50290 18528 50606 18529
rect 50290 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50606 18528
rect 50290 18463 50606 18464
rect 0 18322 800 18352
rect 933 18322 999 18325
rect 0 18320 999 18322
rect 0 18264 938 18320
rect 994 18264 999 18320
rect 0 18262 999 18264
rect 0 18232 800 18262
rect 933 18259 999 18262
rect 59200 18232 60000 18352
rect 26877 18186 26943 18189
rect 31334 18186 31340 18188
rect 26877 18184 31340 18186
rect 26877 18128 26882 18184
rect 26938 18128 31340 18184
rect 26877 18126 31340 18128
rect 26877 18123 26943 18126
rect 31334 18124 31340 18126
rect 31404 18124 31410 18188
rect 43294 17988 43300 18052
rect 43364 18050 43370 18052
rect 43437 18050 43503 18053
rect 43364 18048 43503 18050
rect 43364 17992 43442 18048
rect 43498 17992 43503 18048
rect 43364 17990 43503 17992
rect 43364 17988 43370 17990
rect 43437 17987 43503 17990
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 48405 17916 48471 17917
rect 48405 17912 48452 17916
rect 48516 17914 48522 17916
rect 58985 17914 59051 17917
rect 59200 17914 60000 17944
rect 48405 17856 48410 17912
rect 48405 17852 48452 17856
rect 48516 17854 48562 17914
rect 58985 17912 60000 17914
rect 58985 17856 58990 17912
rect 59046 17856 60000 17912
rect 58985 17854 60000 17856
rect 48516 17852 48522 17854
rect 48405 17851 48471 17852
rect 58985 17851 59051 17854
rect 59200 17824 60000 17854
rect 0 17778 800 17808
rect 933 17778 999 17781
rect 0 17776 999 17778
rect 0 17720 938 17776
rect 994 17720 999 17776
rect 0 17718 999 17720
rect 0 17688 800 17718
rect 933 17715 999 17718
rect 35801 17642 35867 17645
rect 38101 17642 38167 17645
rect 35801 17640 38167 17642
rect 35801 17584 35806 17640
rect 35862 17584 38106 17640
rect 38162 17584 38167 17640
rect 35801 17582 38167 17584
rect 35801 17579 35867 17582
rect 38101 17579 38167 17582
rect 36077 17506 36143 17509
rect 36445 17506 36511 17509
rect 40217 17506 40283 17509
rect 36077 17504 40283 17506
rect 36077 17448 36082 17504
rect 36138 17448 36450 17504
rect 36506 17448 40222 17504
rect 40278 17448 40283 17504
rect 36077 17446 40283 17448
rect 36077 17443 36143 17446
rect 36445 17443 36511 17446
rect 40217 17443 40283 17446
rect 58157 17506 58223 17509
rect 59200 17506 60000 17536
rect 58157 17504 60000 17506
rect 58157 17448 58162 17504
rect 58218 17448 60000 17504
rect 58157 17446 60000 17448
rect 58157 17443 58223 17446
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 50290 17440 50606 17441
rect 50290 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50606 17440
rect 59200 17416 60000 17446
rect 50290 17375 50606 17376
rect 21909 17370 21975 17373
rect 42057 17370 42123 17373
rect 21909 17368 42123 17370
rect 21909 17312 21914 17368
rect 21970 17312 42062 17368
rect 42118 17312 42123 17368
rect 21909 17310 42123 17312
rect 21909 17307 21975 17310
rect 42057 17307 42123 17310
rect 0 17234 800 17264
rect 933 17234 999 17237
rect 0 17232 999 17234
rect 0 17176 938 17232
rect 994 17176 999 17232
rect 0 17174 999 17176
rect 0 17144 800 17174
rect 933 17171 999 17174
rect 24485 17234 24551 17237
rect 44173 17234 44239 17237
rect 24485 17232 44239 17234
rect 24485 17176 24490 17232
rect 24546 17176 44178 17232
rect 44234 17176 44239 17232
rect 24485 17174 44239 17176
rect 24485 17171 24551 17174
rect 44173 17171 44239 17174
rect 31753 17098 31819 17101
rect 32213 17098 32279 17101
rect 35525 17098 35591 17101
rect 31753 17096 35591 17098
rect 31753 17040 31758 17096
rect 31814 17040 32218 17096
rect 32274 17040 35530 17096
rect 35586 17040 35591 17096
rect 31753 17038 35591 17040
rect 31753 17035 31819 17038
rect 32213 17035 32279 17038
rect 35525 17035 35591 17038
rect 35893 17098 35959 17101
rect 48221 17098 48287 17101
rect 35893 17096 48287 17098
rect 35893 17040 35898 17096
rect 35954 17040 48226 17096
rect 48282 17040 48287 17096
rect 35893 17038 48287 17040
rect 35893 17035 35959 17038
rect 48221 17035 48287 17038
rect 48405 17098 48471 17101
rect 52269 17098 52335 17101
rect 48405 17096 52335 17098
rect 48405 17040 48410 17096
rect 48466 17040 52274 17096
rect 52330 17040 52335 17096
rect 48405 17038 52335 17040
rect 48405 17035 48471 17038
rect 52269 17035 52335 17038
rect 59200 17008 60000 17128
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 0 16690 800 16720
rect 933 16690 999 16693
rect 0 16688 999 16690
rect 0 16632 938 16688
rect 994 16632 999 16688
rect 0 16630 999 16632
rect 0 16600 800 16630
rect 933 16627 999 16630
rect 43161 16690 43227 16693
rect 56041 16690 56107 16693
rect 43161 16688 56107 16690
rect 43161 16632 43166 16688
rect 43222 16632 56046 16688
rect 56102 16632 56107 16688
rect 43161 16630 56107 16632
rect 43161 16627 43227 16630
rect 56041 16627 56107 16630
rect 58985 16690 59051 16693
rect 59200 16690 60000 16720
rect 58985 16688 60000 16690
rect 58985 16632 58990 16688
rect 59046 16632 60000 16688
rect 58985 16630 60000 16632
rect 58985 16627 59051 16630
rect 59200 16600 60000 16630
rect 48221 16554 48287 16557
rect 49325 16554 49391 16557
rect 48221 16552 49391 16554
rect 48221 16496 48226 16552
rect 48282 16496 49330 16552
rect 49386 16496 49391 16552
rect 48221 16494 49391 16496
rect 48221 16491 48287 16494
rect 49325 16491 49391 16494
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 50290 16352 50606 16353
rect 50290 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50606 16352
rect 50290 16287 50606 16288
rect 58157 16282 58223 16285
rect 59200 16282 60000 16312
rect 58157 16280 60000 16282
rect 58157 16224 58162 16280
rect 58218 16224 60000 16280
rect 58157 16222 60000 16224
rect 58157 16219 58223 16222
rect 59200 16192 60000 16222
rect 0 16146 800 16176
rect 933 16146 999 16149
rect 0 16144 999 16146
rect 0 16088 938 16144
rect 994 16088 999 16144
rect 0 16086 999 16088
rect 0 16056 800 16086
rect 933 16083 999 16086
rect 46749 16146 46815 16149
rect 59077 16146 59143 16149
rect 46749 16144 59143 16146
rect 46749 16088 46754 16144
rect 46810 16088 59082 16144
rect 59138 16088 59143 16144
rect 46749 16086 59143 16088
rect 46749 16083 46815 16086
rect 59077 16083 59143 16086
rect 36537 16010 36603 16013
rect 38193 16010 38259 16013
rect 36537 16008 38259 16010
rect 36537 15952 36542 16008
rect 36598 15952 38198 16008
rect 38254 15952 38259 16008
rect 36537 15950 38259 15952
rect 36537 15947 36603 15950
rect 38193 15947 38259 15950
rect 20161 15874 20227 15877
rect 34237 15874 34303 15877
rect 20161 15872 34303 15874
rect 20161 15816 20166 15872
rect 20222 15816 34242 15872
rect 34298 15816 34303 15872
rect 20161 15814 34303 15816
rect 20161 15811 20227 15814
rect 34237 15811 34303 15814
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 59200 15784 60000 15904
rect 34930 15743 35246 15744
rect 23197 15738 23263 15741
rect 28717 15738 28783 15741
rect 23197 15736 28783 15738
rect 23197 15680 23202 15736
rect 23258 15680 28722 15736
rect 28778 15680 28783 15736
rect 23197 15678 28783 15680
rect 23197 15675 23263 15678
rect 28717 15675 28783 15678
rect 0 15602 800 15632
rect 933 15602 999 15605
rect 0 15600 999 15602
rect 0 15544 938 15600
rect 994 15544 999 15600
rect 0 15542 999 15544
rect 0 15512 800 15542
rect 933 15539 999 15542
rect 15837 15602 15903 15605
rect 46841 15602 46907 15605
rect 15837 15600 46907 15602
rect 15837 15544 15842 15600
rect 15898 15544 46846 15600
rect 46902 15544 46907 15600
rect 15837 15542 46907 15544
rect 15837 15539 15903 15542
rect 46841 15539 46907 15542
rect 58157 15466 58223 15469
rect 59200 15466 60000 15496
rect 58157 15464 60000 15466
rect 58157 15408 58162 15464
rect 58218 15408 60000 15464
rect 58157 15406 60000 15408
rect 58157 15403 58223 15406
rect 59200 15376 60000 15406
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 50290 15264 50606 15265
rect 50290 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50606 15264
rect 50290 15199 50606 15200
rect 24669 15194 24735 15197
rect 40033 15194 40099 15197
rect 24669 15192 40099 15194
rect 24669 15136 24674 15192
rect 24730 15136 40038 15192
rect 40094 15136 40099 15192
rect 24669 15134 40099 15136
rect 24669 15131 24735 15134
rect 40033 15131 40099 15134
rect 0 15058 800 15088
rect 933 15058 999 15061
rect 0 15056 999 15058
rect 0 15000 938 15056
rect 994 15000 999 15056
rect 0 14998 999 15000
rect 0 14968 800 14998
rect 933 14995 999 14998
rect 30373 15060 30439 15061
rect 30373 15056 30420 15060
rect 30484 15058 30490 15060
rect 58065 15058 58131 15061
rect 59200 15058 60000 15088
rect 30373 15000 30378 15056
rect 30373 14996 30420 15000
rect 30484 14998 30530 15058
rect 58065 15056 60000 15058
rect 58065 15000 58070 15056
rect 58126 15000 60000 15056
rect 58065 14998 60000 15000
rect 30484 14996 30490 14998
rect 30373 14995 30439 14996
rect 58065 14995 58131 14998
rect 59200 14968 60000 14998
rect 23381 14922 23447 14925
rect 39941 14922 40007 14925
rect 23381 14920 40007 14922
rect 23381 14864 23386 14920
rect 23442 14864 39946 14920
rect 40002 14864 40007 14920
rect 23381 14862 40007 14864
rect 23381 14859 23447 14862
rect 39941 14859 40007 14862
rect 29545 14786 29611 14789
rect 32857 14786 32923 14789
rect 29545 14784 32923 14786
rect 29545 14728 29550 14784
rect 29606 14728 32862 14784
rect 32918 14728 32923 14784
rect 29545 14726 32923 14728
rect 29545 14723 29611 14726
rect 32857 14723 32923 14726
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 59200 14560 60000 14680
rect 0 14514 800 14544
rect 933 14514 999 14517
rect 0 14512 999 14514
rect 0 14456 938 14512
rect 994 14456 999 14512
rect 0 14454 999 14456
rect 0 14424 800 14454
rect 933 14451 999 14454
rect 23197 14514 23263 14517
rect 24945 14514 25011 14517
rect 23197 14512 25011 14514
rect 23197 14456 23202 14512
rect 23258 14456 24950 14512
rect 25006 14456 25011 14512
rect 23197 14454 25011 14456
rect 23197 14451 23263 14454
rect 24945 14451 25011 14454
rect 58157 14242 58223 14245
rect 59200 14242 60000 14272
rect 58157 14240 60000 14242
rect 58157 14184 58162 14240
rect 58218 14184 60000 14240
rect 58157 14182 60000 14184
rect 58157 14179 58223 14182
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 50290 14176 50606 14177
rect 50290 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50606 14176
rect 59200 14152 60000 14182
rect 50290 14111 50606 14112
rect 0 13970 800 14000
rect 933 13970 999 13973
rect 0 13968 999 13970
rect 0 13912 938 13968
rect 994 13912 999 13968
rect 0 13910 999 13912
rect 0 13880 800 13910
rect 933 13907 999 13910
rect 28809 13970 28875 13973
rect 58157 13970 58223 13973
rect 28809 13968 58223 13970
rect 28809 13912 28814 13968
rect 28870 13912 58162 13968
rect 58218 13912 58223 13968
rect 28809 13910 58223 13912
rect 28809 13907 28875 13910
rect 58157 13907 58223 13910
rect 29085 13834 29151 13837
rect 34421 13834 34487 13837
rect 29085 13832 34487 13834
rect 29085 13776 29090 13832
rect 29146 13776 34426 13832
rect 34482 13776 34487 13832
rect 29085 13774 34487 13776
rect 29085 13771 29151 13774
rect 34421 13771 34487 13774
rect 39246 13772 39252 13836
rect 39316 13834 39322 13836
rect 42149 13834 42215 13837
rect 39316 13832 42215 13834
rect 39316 13776 42154 13832
rect 42210 13776 42215 13832
rect 39316 13774 42215 13776
rect 39316 13772 39322 13774
rect 42149 13771 42215 13774
rect 58065 13834 58131 13837
rect 59200 13834 60000 13864
rect 58065 13832 60000 13834
rect 58065 13776 58070 13832
rect 58126 13776 60000 13832
rect 58065 13774 60000 13776
rect 58065 13771 58131 13774
rect 59200 13744 60000 13774
rect 31845 13698 31911 13701
rect 33174 13698 33180 13700
rect 31845 13696 33180 13698
rect 31845 13640 31850 13696
rect 31906 13640 33180 13696
rect 31845 13638 33180 13640
rect 31845 13635 31911 13638
rect 33174 13636 33180 13638
rect 33244 13636 33250 13700
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 0 13426 800 13456
rect 933 13426 999 13429
rect 0 13424 999 13426
rect 0 13368 938 13424
rect 994 13368 999 13424
rect 0 13366 999 13368
rect 0 13336 800 13366
rect 933 13363 999 13366
rect 30097 13426 30163 13429
rect 33317 13426 33383 13429
rect 34053 13426 34119 13429
rect 35893 13426 35959 13429
rect 30097 13424 35959 13426
rect 30097 13368 30102 13424
rect 30158 13368 33322 13424
rect 33378 13368 34058 13424
rect 34114 13368 35898 13424
rect 35954 13368 35959 13424
rect 30097 13366 35959 13368
rect 30097 13363 30163 13366
rect 33317 13363 33383 13366
rect 34053 13363 34119 13366
rect 35893 13363 35959 13366
rect 59200 13336 60000 13456
rect 12433 13290 12499 13293
rect 36077 13290 36143 13293
rect 12433 13288 36143 13290
rect 12433 13232 12438 13288
rect 12494 13232 36082 13288
rect 36138 13232 36143 13288
rect 12433 13230 36143 13232
rect 12433 13227 12499 13230
rect 36077 13227 36143 13230
rect 21817 13154 21883 13157
rect 33225 13154 33291 13157
rect 21817 13152 33291 13154
rect 21817 13096 21822 13152
rect 21878 13096 33230 13152
rect 33286 13096 33291 13152
rect 21817 13094 33291 13096
rect 21817 13091 21883 13094
rect 33225 13091 33291 13094
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 50290 13088 50606 13089
rect 50290 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50606 13088
rect 50290 13023 50606 13024
rect 29085 13018 29151 13021
rect 43529 13018 43595 13021
rect 29085 13016 43595 13018
rect 29085 12960 29090 13016
rect 29146 12960 43534 13016
rect 43590 12960 43595 13016
rect 29085 12958 43595 12960
rect 29085 12955 29151 12958
rect 43529 12955 43595 12958
rect 58985 13018 59051 13021
rect 59200 13018 60000 13048
rect 58985 13016 60000 13018
rect 58985 12960 58990 13016
rect 59046 12960 60000 13016
rect 58985 12958 60000 12960
rect 58985 12955 59051 12958
rect 59200 12928 60000 12958
rect 0 12882 800 12912
rect 933 12882 999 12885
rect 0 12880 999 12882
rect 0 12824 938 12880
rect 994 12824 999 12880
rect 0 12822 999 12824
rect 0 12792 800 12822
rect 933 12819 999 12822
rect 40033 12882 40099 12885
rect 55581 12882 55647 12885
rect 40033 12880 55647 12882
rect 40033 12824 40038 12880
rect 40094 12824 55586 12880
rect 55642 12824 55647 12880
rect 40033 12822 55647 12824
rect 40033 12819 40099 12822
rect 55581 12819 55647 12822
rect 58065 12610 58131 12613
rect 59200 12610 60000 12640
rect 58065 12608 60000 12610
rect 58065 12552 58070 12608
rect 58126 12552 60000 12608
rect 58065 12550 60000 12552
rect 58065 12547 58131 12550
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 59200 12520 60000 12550
rect 34930 12479 35246 12480
rect 0 12338 800 12368
rect 933 12338 999 12341
rect 0 12336 999 12338
rect 0 12280 938 12336
rect 994 12280 999 12336
rect 0 12278 999 12280
rect 0 12248 800 12278
rect 933 12275 999 12278
rect 23289 12338 23355 12341
rect 27153 12338 27219 12341
rect 23289 12336 27219 12338
rect 23289 12280 23294 12336
rect 23350 12280 27158 12336
rect 27214 12280 27219 12336
rect 23289 12278 27219 12280
rect 23289 12275 23355 12278
rect 27153 12275 27219 12278
rect 39665 12338 39731 12341
rect 46054 12338 46060 12340
rect 39665 12336 46060 12338
rect 39665 12280 39670 12336
rect 39726 12280 46060 12336
rect 39665 12278 46060 12280
rect 39665 12275 39731 12278
rect 46054 12276 46060 12278
rect 46124 12276 46130 12340
rect 20713 12202 20779 12205
rect 37733 12202 37799 12205
rect 20713 12200 37799 12202
rect 20713 12144 20718 12200
rect 20774 12144 37738 12200
rect 37794 12144 37799 12200
rect 20713 12142 37799 12144
rect 20713 12139 20779 12142
rect 37733 12139 37799 12142
rect 59200 12112 60000 12232
rect 23473 12066 23539 12069
rect 29494 12066 29500 12068
rect 23473 12064 29500 12066
rect 23473 12008 23478 12064
rect 23534 12008 29500 12064
rect 23473 12006 29500 12008
rect 23473 12003 23539 12006
rect 29494 12004 29500 12006
rect 29564 12066 29570 12068
rect 30925 12066 30991 12069
rect 29564 12064 30991 12066
rect 29564 12008 30930 12064
rect 30986 12008 30991 12064
rect 29564 12006 30991 12008
rect 29564 12004 29570 12006
rect 30925 12003 30991 12006
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 50290 12000 50606 12001
rect 50290 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50606 12000
rect 50290 11935 50606 11936
rect 0 11794 800 11824
rect 933 11794 999 11797
rect 0 11792 999 11794
rect 0 11736 938 11792
rect 994 11736 999 11792
rect 0 11734 999 11736
rect 0 11704 800 11734
rect 933 11731 999 11734
rect 40534 11732 40540 11796
rect 40604 11794 40610 11796
rect 43713 11794 43779 11797
rect 40604 11792 43779 11794
rect 40604 11736 43718 11792
rect 43774 11736 43779 11792
rect 40604 11734 43779 11736
rect 40604 11732 40610 11734
rect 43713 11731 43779 11734
rect 58157 11794 58223 11797
rect 59200 11794 60000 11824
rect 58157 11792 60000 11794
rect 58157 11736 58162 11792
rect 58218 11736 60000 11792
rect 58157 11734 60000 11736
rect 58157 11731 58223 11734
rect 59200 11704 60000 11734
rect 22737 11658 22803 11661
rect 26785 11658 26851 11661
rect 34237 11658 34303 11661
rect 22737 11656 34303 11658
rect 22737 11600 22742 11656
rect 22798 11600 26790 11656
rect 26846 11600 34242 11656
rect 34298 11600 34303 11656
rect 22737 11598 34303 11600
rect 22737 11595 22803 11598
rect 26785 11595 26851 11598
rect 34237 11595 34303 11598
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 28993 11386 29059 11389
rect 30741 11386 30807 11389
rect 28993 11384 30807 11386
rect 28993 11328 28998 11384
rect 29054 11328 30746 11384
rect 30802 11328 30807 11384
rect 28993 11326 30807 11328
rect 28993 11323 29059 11326
rect 30741 11323 30807 11326
rect 58065 11386 58131 11389
rect 59200 11386 60000 11416
rect 58065 11384 60000 11386
rect 58065 11328 58070 11384
rect 58126 11328 60000 11384
rect 58065 11326 60000 11328
rect 58065 11323 58131 11326
rect 59200 11296 60000 11326
rect 0 11250 800 11280
rect 933 11250 999 11253
rect 0 11248 999 11250
rect 0 11192 938 11248
rect 994 11192 999 11248
rect 0 11190 999 11192
rect 0 11160 800 11190
rect 933 11187 999 11190
rect 14549 11250 14615 11253
rect 43069 11250 43135 11253
rect 14549 11248 43135 11250
rect 14549 11192 14554 11248
rect 14610 11192 43074 11248
rect 43130 11192 43135 11248
rect 14549 11190 43135 11192
rect 14549 11187 14615 11190
rect 43069 11187 43135 11190
rect 28625 11114 28691 11117
rect 33869 11114 33935 11117
rect 28625 11112 33935 11114
rect 28625 11056 28630 11112
rect 28686 11056 33874 11112
rect 33930 11056 33935 11112
rect 28625 11054 33935 11056
rect 28625 11051 28691 11054
rect 33869 11051 33935 11054
rect 29821 10978 29887 10981
rect 32949 10978 33015 10981
rect 29821 10976 33015 10978
rect 29821 10920 29826 10976
rect 29882 10920 32954 10976
rect 33010 10920 33015 10976
rect 29821 10918 33015 10920
rect 29821 10915 29887 10918
rect 32949 10915 33015 10918
rect 33133 10978 33199 10981
rect 33685 10978 33751 10981
rect 33133 10976 33751 10978
rect 33133 10920 33138 10976
rect 33194 10920 33690 10976
rect 33746 10920 33751 10976
rect 33133 10918 33751 10920
rect 33133 10915 33199 10918
rect 33685 10915 33751 10918
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 50290 10912 50606 10913
rect 50290 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50606 10912
rect 59200 10888 60000 11008
rect 50290 10847 50606 10848
rect 39757 10842 39823 10845
rect 43294 10842 43300 10844
rect 39757 10840 43300 10842
rect 39757 10784 39762 10840
rect 39818 10784 43300 10840
rect 39757 10782 43300 10784
rect 39757 10779 39823 10782
rect 43294 10780 43300 10782
rect 43364 10780 43370 10844
rect 0 10706 800 10736
rect 933 10706 999 10709
rect 0 10704 999 10706
rect 0 10648 938 10704
rect 994 10648 999 10704
rect 0 10646 999 10648
rect 0 10616 800 10646
rect 933 10643 999 10646
rect 22093 10706 22159 10709
rect 38101 10706 38167 10709
rect 22093 10704 38167 10706
rect 22093 10648 22098 10704
rect 22154 10648 38106 10704
rect 38162 10648 38167 10704
rect 22093 10646 38167 10648
rect 22093 10643 22159 10646
rect 38101 10643 38167 10646
rect 22001 10570 22067 10573
rect 43294 10570 43300 10572
rect 22001 10568 43300 10570
rect 22001 10512 22006 10568
rect 22062 10512 43300 10568
rect 22001 10510 43300 10512
rect 22001 10507 22067 10510
rect 43294 10508 43300 10510
rect 43364 10508 43370 10572
rect 58985 10570 59051 10573
rect 59200 10570 60000 10600
rect 58985 10568 60000 10570
rect 58985 10512 58990 10568
rect 59046 10512 60000 10568
rect 58985 10510 60000 10512
rect 58985 10507 59051 10510
rect 59200 10480 60000 10510
rect 27705 10434 27771 10437
rect 28625 10434 28691 10437
rect 27705 10432 28691 10434
rect 27705 10376 27710 10432
rect 27766 10376 28630 10432
rect 28686 10376 28691 10432
rect 27705 10374 28691 10376
rect 27705 10371 27771 10374
rect 28625 10371 28691 10374
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 0 10162 800 10192
rect 933 10162 999 10165
rect 0 10160 999 10162
rect 0 10104 938 10160
rect 994 10104 999 10160
rect 0 10102 999 10104
rect 0 10072 800 10102
rect 933 10099 999 10102
rect 12617 10162 12683 10165
rect 41965 10162 42031 10165
rect 12617 10160 42031 10162
rect 12617 10104 12622 10160
rect 12678 10104 41970 10160
rect 42026 10104 42031 10160
rect 12617 10102 42031 10104
rect 12617 10099 12683 10102
rect 41965 10099 42031 10102
rect 58893 10162 58959 10165
rect 59200 10162 60000 10192
rect 58893 10160 60000 10162
rect 58893 10104 58898 10160
rect 58954 10104 60000 10160
rect 58893 10102 60000 10104
rect 58893 10099 58959 10102
rect 59200 10072 60000 10102
rect 28349 9890 28415 9893
rect 34697 9890 34763 9893
rect 28349 9888 34763 9890
rect 28349 9832 28354 9888
rect 28410 9832 34702 9888
rect 34758 9832 34763 9888
rect 28349 9830 34763 9832
rect 28349 9827 28415 9830
rect 34697 9827 34763 9830
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 50290 9824 50606 9825
rect 50290 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50606 9824
rect 50290 9759 50606 9760
rect 39297 9754 39363 9757
rect 41413 9754 41479 9757
rect 39297 9752 41479 9754
rect 39297 9696 39302 9752
rect 39358 9696 41418 9752
rect 41474 9696 41479 9752
rect 39297 9694 41479 9696
rect 30741 9690 30807 9693
rect 39297 9691 39363 9694
rect 41413 9691 41479 9694
rect 42558 9692 42564 9756
rect 42628 9754 42634 9756
rect 43069 9754 43135 9757
rect 42628 9752 43135 9754
rect 42628 9696 43074 9752
rect 43130 9696 43135 9752
rect 42628 9694 43135 9696
rect 42628 9692 42634 9694
rect 43069 9691 43135 9694
rect 30422 9688 30807 9690
rect 0 9618 800 9648
rect 30422 9632 30746 9688
rect 30802 9632 30807 9688
rect 59200 9664 60000 9784
rect 30422 9630 30807 9632
rect 933 9618 999 9621
rect 30422 9618 30482 9630
rect 30741 9627 30807 9630
rect 0 9616 999 9618
rect 0 9560 938 9616
rect 994 9560 999 9616
rect 0 9558 999 9560
rect 0 9528 800 9558
rect 933 9555 999 9558
rect 30238 9558 30482 9618
rect 22093 9482 22159 9485
rect 26325 9482 26391 9485
rect 27245 9482 27311 9485
rect 22093 9480 27311 9482
rect 22093 9424 22098 9480
rect 22154 9424 26330 9480
rect 26386 9424 27250 9480
rect 27306 9424 27311 9480
rect 22093 9422 27311 9424
rect 22093 9419 22159 9422
rect 26325 9419 26391 9422
rect 27245 9419 27311 9422
rect 27797 9482 27863 9485
rect 28533 9482 28599 9485
rect 27797 9480 28599 9482
rect 27797 9424 27802 9480
rect 27858 9424 28538 9480
rect 28594 9424 28599 9480
rect 27797 9422 28599 9424
rect 27797 9419 27863 9422
rect 28533 9419 28599 9422
rect 30238 9346 30298 9558
rect 31150 9556 31156 9620
rect 31220 9618 31226 9620
rect 31293 9618 31359 9621
rect 31220 9616 31359 9618
rect 31220 9560 31298 9616
rect 31354 9560 31359 9616
rect 31220 9558 31359 9560
rect 31220 9556 31226 9558
rect 31293 9555 31359 9558
rect 33174 9556 33180 9620
rect 33244 9618 33250 9620
rect 33317 9618 33383 9621
rect 33244 9616 33383 9618
rect 33244 9560 33322 9616
rect 33378 9560 33383 9616
rect 33244 9558 33383 9560
rect 33244 9556 33250 9558
rect 33317 9555 33383 9558
rect 37774 9556 37780 9620
rect 37844 9618 37850 9620
rect 41965 9618 42031 9621
rect 37844 9616 42031 9618
rect 37844 9560 41970 9616
rect 42026 9560 42031 9616
rect 37844 9558 42031 9560
rect 37844 9556 37850 9558
rect 41965 9555 42031 9558
rect 30925 9482 30991 9485
rect 36629 9482 36695 9485
rect 30925 9480 36695 9482
rect 30925 9424 30930 9480
rect 30986 9424 36634 9480
rect 36690 9424 36695 9480
rect 30925 9422 36695 9424
rect 30925 9419 30991 9422
rect 36629 9419 36695 9422
rect 30465 9346 30531 9349
rect 30238 9344 30531 9346
rect 30238 9288 30470 9344
rect 30526 9288 30531 9344
rect 30238 9286 30531 9288
rect 30465 9283 30531 9286
rect 30833 9346 30899 9349
rect 31569 9346 31635 9349
rect 30833 9344 31635 9346
rect 30833 9288 30838 9344
rect 30894 9288 31574 9344
rect 31630 9288 31635 9344
rect 30833 9286 31635 9288
rect 30833 9283 30899 9286
rect 31569 9283 31635 9286
rect 58985 9346 59051 9349
rect 59200 9346 60000 9376
rect 58985 9344 60000 9346
rect 58985 9288 58990 9344
rect 59046 9288 60000 9344
rect 58985 9286 60000 9288
rect 58985 9283 59051 9286
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 59200 9256 60000 9286
rect 34930 9215 35246 9216
rect 26969 9210 27035 9213
rect 31477 9210 31543 9213
rect 26969 9208 31543 9210
rect 26969 9152 26974 9208
rect 27030 9152 31482 9208
rect 31538 9152 31543 9208
rect 26969 9150 31543 9152
rect 26969 9147 27035 9150
rect 31477 9147 31543 9150
rect 0 9074 800 9104
rect 933 9074 999 9077
rect 0 9072 999 9074
rect 0 9016 938 9072
rect 994 9016 999 9072
rect 0 9014 999 9016
rect 0 8984 800 9014
rect 933 9011 999 9014
rect 23013 9074 23079 9077
rect 33041 9074 33107 9077
rect 23013 9072 33107 9074
rect 23013 9016 23018 9072
rect 23074 9016 33046 9072
rect 33102 9016 33107 9072
rect 23013 9014 33107 9016
rect 23013 9011 23079 9014
rect 33041 9011 33107 9014
rect 24209 8938 24275 8941
rect 46381 8938 46447 8941
rect 24209 8936 46447 8938
rect 24209 8880 24214 8936
rect 24270 8880 46386 8936
rect 46442 8880 46447 8936
rect 24209 8878 46447 8880
rect 24209 8875 24275 8878
rect 46381 8875 46447 8878
rect 58065 8938 58131 8941
rect 59200 8938 60000 8968
rect 58065 8936 60000 8938
rect 58065 8880 58070 8936
rect 58126 8880 60000 8936
rect 58065 8878 60000 8880
rect 58065 8875 58131 8878
rect 59200 8848 60000 8878
rect 31150 8740 31156 8804
rect 31220 8802 31226 8804
rect 31293 8802 31359 8805
rect 31220 8800 31359 8802
rect 31220 8744 31298 8800
rect 31354 8744 31359 8800
rect 31220 8742 31359 8744
rect 31220 8740 31226 8742
rect 31293 8739 31359 8742
rect 31477 8802 31543 8805
rect 36169 8802 36235 8805
rect 31477 8800 36235 8802
rect 31477 8744 31482 8800
rect 31538 8744 36174 8800
rect 36230 8744 36235 8800
rect 31477 8742 36235 8744
rect 31477 8739 31543 8742
rect 36169 8739 36235 8742
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 50290 8736 50606 8737
rect 50290 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50606 8736
rect 50290 8671 50606 8672
rect 29821 8666 29887 8669
rect 37917 8666 37983 8669
rect 29821 8664 37983 8666
rect 29821 8608 29826 8664
rect 29882 8608 37922 8664
rect 37978 8608 37983 8664
rect 29821 8606 37983 8608
rect 29821 8603 29887 8606
rect 37917 8603 37983 8606
rect 0 8530 800 8560
rect 933 8530 999 8533
rect 0 8528 999 8530
rect 0 8472 938 8528
rect 994 8472 999 8528
rect 0 8470 999 8472
rect 0 8440 800 8470
rect 933 8467 999 8470
rect 28533 8530 28599 8533
rect 28809 8530 28875 8533
rect 28533 8528 28875 8530
rect 28533 8472 28538 8528
rect 28594 8472 28814 8528
rect 28870 8472 28875 8528
rect 28533 8470 28875 8472
rect 28533 8467 28599 8470
rect 28809 8467 28875 8470
rect 29913 8530 29979 8533
rect 32397 8530 32463 8533
rect 29913 8528 32463 8530
rect 29913 8472 29918 8528
rect 29974 8472 32402 8528
rect 32458 8472 32463 8528
rect 29913 8470 32463 8472
rect 29913 8467 29979 8470
rect 32397 8467 32463 8470
rect 33685 8530 33751 8533
rect 58709 8530 58775 8533
rect 33685 8528 58775 8530
rect 33685 8472 33690 8528
rect 33746 8472 58714 8528
rect 58770 8472 58775 8528
rect 33685 8470 58775 8472
rect 33685 8467 33751 8470
rect 58709 8467 58775 8470
rect 59200 8440 60000 8560
rect 27613 8394 27679 8397
rect 36445 8394 36511 8397
rect 27613 8392 36511 8394
rect 27613 8336 27618 8392
rect 27674 8336 36450 8392
rect 36506 8336 36511 8392
rect 27613 8334 36511 8336
rect 27613 8331 27679 8334
rect 36445 8331 36511 8334
rect 43478 8332 43484 8396
rect 43548 8394 43554 8396
rect 44633 8394 44699 8397
rect 43548 8392 44699 8394
rect 43548 8336 44638 8392
rect 44694 8336 44699 8392
rect 43548 8334 44699 8336
rect 43548 8332 43554 8334
rect 44633 8331 44699 8334
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 58157 8122 58223 8125
rect 59200 8122 60000 8152
rect 58157 8120 60000 8122
rect 58157 8064 58162 8120
rect 58218 8064 60000 8120
rect 58157 8062 60000 8064
rect 58157 8059 58223 8062
rect 59200 8032 60000 8062
rect 0 7986 800 8016
rect 933 7986 999 7989
rect 0 7984 999 7986
rect 0 7928 938 7984
rect 994 7928 999 7984
rect 0 7926 999 7928
rect 0 7896 800 7926
rect 933 7923 999 7926
rect 31937 7986 32003 7989
rect 35985 7986 36051 7989
rect 31937 7984 36051 7986
rect 31937 7928 31942 7984
rect 31998 7928 35990 7984
rect 36046 7928 36051 7984
rect 31937 7926 36051 7928
rect 31937 7923 32003 7926
rect 35985 7923 36051 7926
rect 42977 7986 43043 7989
rect 48129 7986 48195 7989
rect 42977 7984 48195 7986
rect 42977 7928 42982 7984
rect 43038 7928 48134 7984
rect 48190 7928 48195 7984
rect 42977 7926 48195 7928
rect 42977 7923 43043 7926
rect 48129 7923 48195 7926
rect 58065 7714 58131 7717
rect 59200 7714 60000 7744
rect 58065 7712 60000 7714
rect 58065 7656 58070 7712
rect 58126 7656 60000 7712
rect 58065 7654 60000 7656
rect 58065 7651 58131 7654
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 50290 7648 50606 7649
rect 50290 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50606 7648
rect 59200 7624 60000 7654
rect 50290 7583 50606 7584
rect 30925 7578 30991 7581
rect 36261 7578 36327 7581
rect 30925 7576 36327 7578
rect 30925 7520 30930 7576
rect 30986 7520 36266 7576
rect 36322 7520 36327 7576
rect 30925 7518 36327 7520
rect 30925 7515 30991 7518
rect 36261 7515 36327 7518
rect 0 7442 800 7472
rect 933 7442 999 7445
rect 0 7440 999 7442
rect 0 7384 938 7440
rect 994 7384 999 7440
rect 0 7382 999 7384
rect 0 7352 800 7382
rect 933 7379 999 7382
rect 11697 7442 11763 7445
rect 38377 7442 38443 7445
rect 11697 7440 38443 7442
rect 11697 7384 11702 7440
rect 11758 7384 38382 7440
rect 38438 7384 38443 7440
rect 11697 7382 38443 7384
rect 11697 7379 11763 7382
rect 38377 7379 38443 7382
rect 28349 7306 28415 7309
rect 58249 7306 58315 7309
rect 28349 7304 58315 7306
rect 28349 7248 28354 7304
rect 28410 7248 58254 7304
rect 58310 7248 58315 7304
rect 28349 7246 58315 7248
rect 28349 7243 28415 7246
rect 58249 7243 58315 7246
rect 59200 7216 60000 7336
rect 30925 7170 30991 7173
rect 34789 7170 34855 7173
rect 30925 7168 34855 7170
rect 30925 7112 30930 7168
rect 30986 7112 34794 7168
rect 34850 7112 34855 7168
rect 30925 7110 34855 7112
rect 30925 7107 30991 7110
rect 34789 7107 34855 7110
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 0 6898 800 6928
rect 933 6898 999 6901
rect 0 6896 999 6898
rect 0 6840 938 6896
rect 994 6840 999 6896
rect 0 6838 999 6840
rect 0 6808 800 6838
rect 933 6835 999 6838
rect 44909 6898 44975 6901
rect 45829 6898 45895 6901
rect 44909 6896 45895 6898
rect 44909 6840 44914 6896
rect 44970 6840 45834 6896
rect 45890 6840 45895 6896
rect 44909 6838 45895 6840
rect 44909 6835 44975 6838
rect 45829 6835 45895 6838
rect 58985 6898 59051 6901
rect 59200 6898 60000 6928
rect 58985 6896 60000 6898
rect 58985 6840 58990 6896
rect 59046 6840 60000 6896
rect 58985 6838 60000 6840
rect 58985 6835 59051 6838
rect 59200 6808 60000 6838
rect 29085 6762 29151 6765
rect 37733 6762 37799 6765
rect 29085 6760 37799 6762
rect 29085 6704 29090 6760
rect 29146 6704 37738 6760
rect 37794 6704 37799 6760
rect 29085 6702 37799 6704
rect 29085 6699 29151 6702
rect 37733 6699 37799 6702
rect 43345 6762 43411 6765
rect 48221 6762 48287 6765
rect 43345 6760 48287 6762
rect 43345 6704 43350 6760
rect 43406 6704 48226 6760
rect 48282 6704 48287 6760
rect 43345 6702 48287 6704
rect 43345 6699 43411 6702
rect 48221 6699 48287 6702
rect 30281 6626 30347 6629
rect 35709 6626 35775 6629
rect 30281 6624 35775 6626
rect 30281 6568 30286 6624
rect 30342 6568 35714 6624
rect 35770 6568 35775 6624
rect 30281 6566 35775 6568
rect 30281 6563 30347 6566
rect 35709 6563 35775 6566
rect 42609 6626 42675 6629
rect 46657 6626 46723 6629
rect 42609 6624 46723 6626
rect 42609 6568 42614 6624
rect 42670 6568 46662 6624
rect 46718 6568 46723 6624
rect 42609 6566 46723 6568
rect 42609 6563 42675 6566
rect 46657 6563 46723 6566
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 50290 6560 50606 6561
rect 50290 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50606 6560
rect 50290 6495 50606 6496
rect 20989 6490 21055 6493
rect 36169 6490 36235 6493
rect 20989 6488 36235 6490
rect 20989 6432 20994 6488
rect 21050 6432 36174 6488
rect 36230 6432 36235 6488
rect 20989 6430 36235 6432
rect 20989 6427 21055 6430
rect 36169 6427 36235 6430
rect 45369 6490 45435 6493
rect 46749 6490 46815 6493
rect 45369 6488 46815 6490
rect 45369 6432 45374 6488
rect 45430 6432 46754 6488
rect 46810 6432 46815 6488
rect 45369 6430 46815 6432
rect 45369 6427 45435 6430
rect 46749 6427 46815 6430
rect 58985 6490 59051 6493
rect 59200 6490 60000 6520
rect 58985 6488 60000 6490
rect 58985 6432 58990 6488
rect 59046 6432 60000 6488
rect 58985 6430 60000 6432
rect 58985 6427 59051 6430
rect 59200 6400 60000 6430
rect 0 6354 800 6384
rect 933 6354 999 6357
rect 0 6352 999 6354
rect 0 6296 938 6352
rect 994 6296 999 6352
rect 0 6294 999 6296
rect 0 6264 800 6294
rect 933 6291 999 6294
rect 25221 6354 25287 6357
rect 33225 6354 33291 6357
rect 43989 6354 44055 6357
rect 25221 6352 44055 6354
rect 25221 6296 25226 6352
rect 25282 6296 33230 6352
rect 33286 6296 43994 6352
rect 44050 6296 44055 6352
rect 25221 6294 44055 6296
rect 25221 6291 25287 6294
rect 33225 6291 33291 6294
rect 43989 6291 44055 6294
rect 25681 6218 25747 6221
rect 27797 6218 27863 6221
rect 25681 6216 27863 6218
rect 25681 6160 25686 6216
rect 25742 6160 27802 6216
rect 27858 6160 27863 6216
rect 25681 6158 27863 6160
rect 25681 6155 25747 6158
rect 27797 6155 27863 6158
rect 28993 6218 29059 6221
rect 35893 6218 35959 6221
rect 28993 6216 35959 6218
rect 28993 6160 28998 6216
rect 29054 6160 35898 6216
rect 35954 6160 35959 6216
rect 28993 6158 35959 6160
rect 28993 6155 29059 6158
rect 35893 6155 35959 6158
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 59200 5992 60000 6112
rect 34930 5951 35246 5952
rect 0 5810 800 5840
rect 933 5810 999 5813
rect 0 5808 999 5810
rect 0 5752 938 5808
rect 994 5752 999 5808
rect 0 5750 999 5752
rect 0 5720 800 5750
rect 933 5747 999 5750
rect 9489 5810 9555 5813
rect 40493 5810 40559 5813
rect 9489 5808 40559 5810
rect 9489 5752 9494 5808
rect 9550 5752 40498 5808
rect 40554 5752 40559 5808
rect 9489 5750 40559 5752
rect 9489 5747 9555 5750
rect 40493 5747 40559 5750
rect 27613 5674 27679 5677
rect 36261 5674 36327 5677
rect 43345 5676 43411 5677
rect 27613 5672 36327 5674
rect 27613 5616 27618 5672
rect 27674 5616 36266 5672
rect 36322 5616 36327 5672
rect 27613 5614 36327 5616
rect 27613 5611 27679 5614
rect 36261 5611 36327 5614
rect 43294 5612 43300 5676
rect 43364 5674 43411 5676
rect 58985 5674 59051 5677
rect 59200 5674 60000 5704
rect 43364 5672 43456 5674
rect 43406 5616 43456 5672
rect 43364 5614 43456 5616
rect 58985 5672 60000 5674
rect 58985 5616 58990 5672
rect 59046 5616 60000 5672
rect 58985 5614 60000 5616
rect 43364 5612 43411 5614
rect 43345 5611 43411 5612
rect 58985 5611 59051 5614
rect 59200 5584 60000 5614
rect 47710 5476 47716 5540
rect 47780 5538 47786 5540
rect 48037 5538 48103 5541
rect 47780 5536 48103 5538
rect 47780 5480 48042 5536
rect 48098 5480 48103 5536
rect 47780 5478 48103 5480
rect 47780 5476 47786 5478
rect 48037 5475 48103 5478
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 50290 5472 50606 5473
rect 50290 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50606 5472
rect 50290 5407 50606 5408
rect 41229 5404 41295 5405
rect 41229 5402 41276 5404
rect 41184 5400 41276 5402
rect 41184 5344 41234 5400
rect 41184 5342 41276 5344
rect 41229 5340 41276 5342
rect 41340 5340 41346 5404
rect 41229 5339 41295 5340
rect 0 5266 800 5296
rect 933 5266 999 5269
rect 0 5264 999 5266
rect 0 5208 938 5264
rect 994 5208 999 5264
rect 0 5206 999 5208
rect 0 5176 800 5206
rect 933 5203 999 5206
rect 19793 5266 19859 5269
rect 27889 5266 27955 5269
rect 19793 5264 27955 5266
rect 19793 5208 19798 5264
rect 19854 5208 27894 5264
rect 27950 5208 27955 5264
rect 19793 5206 27955 5208
rect 19793 5203 19859 5206
rect 27889 5203 27955 5206
rect 58065 5266 58131 5269
rect 59200 5266 60000 5296
rect 58065 5264 60000 5266
rect 58065 5208 58070 5264
rect 58126 5208 60000 5264
rect 58065 5206 60000 5208
rect 58065 5203 58131 5206
rect 59200 5176 60000 5206
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 59200 4768 60000 4888
rect 0 4722 800 4752
rect 933 4722 999 4725
rect 0 4720 999 4722
rect 0 4664 938 4720
rect 994 4664 999 4720
rect 0 4662 999 4664
rect 0 4632 800 4662
rect 933 4659 999 4662
rect 22001 4722 22067 4725
rect 25589 4722 25655 4725
rect 22001 4720 25655 4722
rect 22001 4664 22006 4720
rect 22062 4664 25594 4720
rect 25650 4664 25655 4720
rect 22001 4662 25655 4664
rect 22001 4659 22067 4662
rect 25589 4659 25655 4662
rect 35157 4722 35223 4725
rect 37733 4722 37799 4725
rect 35157 4720 37799 4722
rect 35157 4664 35162 4720
rect 35218 4664 37738 4720
rect 37794 4664 37799 4720
rect 35157 4662 37799 4664
rect 35157 4659 35223 4662
rect 37733 4659 37799 4662
rect 28257 4586 28323 4589
rect 47393 4586 47459 4589
rect 28257 4584 47459 4586
rect 28257 4528 28262 4584
rect 28318 4528 47398 4584
rect 47454 4528 47459 4584
rect 28257 4526 47459 4528
rect 28257 4523 28323 4526
rect 47393 4523 47459 4526
rect 20897 4450 20963 4453
rect 22553 4450 22619 4453
rect 20897 4448 22619 4450
rect 20897 4392 20902 4448
rect 20958 4392 22558 4448
rect 22614 4392 22619 4448
rect 20897 4390 22619 4392
rect 20897 4387 20963 4390
rect 22553 4387 22619 4390
rect 35985 4450 36051 4453
rect 36629 4450 36695 4453
rect 35985 4448 36695 4450
rect 35985 4392 35990 4448
rect 36046 4392 36634 4448
rect 36690 4392 36695 4448
rect 35985 4390 36695 4392
rect 35985 4387 36051 4390
rect 36629 4387 36695 4390
rect 39113 4450 39179 4453
rect 40677 4450 40743 4453
rect 39113 4448 40743 4450
rect 39113 4392 39118 4448
rect 39174 4392 40682 4448
rect 40738 4392 40743 4448
rect 39113 4390 40743 4392
rect 39113 4387 39179 4390
rect 40677 4387 40743 4390
rect 58985 4450 59051 4453
rect 59200 4450 60000 4480
rect 58985 4448 60000 4450
rect 58985 4392 58990 4448
rect 59046 4392 60000 4448
rect 58985 4390 60000 4392
rect 58985 4387 59051 4390
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 50290 4384 50606 4385
rect 50290 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50606 4384
rect 59200 4360 60000 4390
rect 50290 4319 50606 4320
rect 35893 4314 35959 4317
rect 38561 4314 38627 4317
rect 35893 4312 38627 4314
rect 35893 4256 35898 4312
rect 35954 4256 38566 4312
rect 38622 4256 38627 4312
rect 35893 4254 38627 4256
rect 35893 4251 35959 4254
rect 38561 4251 38627 4254
rect 46238 4252 46244 4316
rect 46308 4314 46314 4316
rect 47761 4314 47827 4317
rect 46308 4312 47827 4314
rect 46308 4256 47766 4312
rect 47822 4256 47827 4312
rect 46308 4254 47827 4256
rect 46308 4252 46314 4254
rect 47761 4251 47827 4254
rect 0 4178 800 4208
rect 933 4178 999 4181
rect 0 4176 999 4178
rect 0 4120 938 4176
rect 994 4120 999 4176
rect 0 4118 999 4120
rect 0 4088 800 4118
rect 933 4115 999 4118
rect 19885 4178 19951 4181
rect 22553 4178 22619 4181
rect 19885 4176 22619 4178
rect 19885 4120 19890 4176
rect 19946 4120 22558 4176
rect 22614 4120 22619 4176
rect 19885 4118 22619 4120
rect 19885 4115 19951 4118
rect 22553 4115 22619 4118
rect 37181 4178 37247 4181
rect 53741 4178 53807 4181
rect 37181 4176 53807 4178
rect 37181 4120 37186 4176
rect 37242 4120 53746 4176
rect 53802 4120 53807 4176
rect 37181 4118 53807 4120
rect 37181 4115 37247 4118
rect 53741 4115 53807 4118
rect 10041 4042 10107 4045
rect 20713 4042 20779 4045
rect 10041 4040 20779 4042
rect 10041 3984 10046 4040
rect 10102 3984 20718 4040
rect 20774 3984 20779 4040
rect 10041 3982 20779 3984
rect 10041 3979 10107 3982
rect 20713 3979 20779 3982
rect 31293 4044 31359 4045
rect 31293 4040 31340 4044
rect 31404 4042 31410 4044
rect 43529 4042 43595 4045
rect 31293 3984 31298 4040
rect 31293 3980 31340 3984
rect 31404 3982 31450 4042
rect 31710 4040 43595 4042
rect 31710 3984 43534 4040
rect 43590 3984 43595 4040
rect 31710 3982 43595 3984
rect 31404 3980 31410 3982
rect 31293 3979 31359 3980
rect 27521 3906 27587 3909
rect 31710 3906 31770 3982
rect 43529 3979 43595 3982
rect 44265 4042 44331 4045
rect 47853 4044 47919 4045
rect 48589 4044 48655 4045
rect 44398 4042 44404 4044
rect 44265 4040 44404 4042
rect 44265 3984 44270 4040
rect 44326 3984 44404 4040
rect 44265 3982 44404 3984
rect 44265 3979 44331 3982
rect 44398 3980 44404 3982
rect 44468 3980 44474 4044
rect 47853 4040 47900 4044
rect 47964 4042 47970 4044
rect 48589 4042 48636 4044
rect 47853 3984 47858 4040
rect 47853 3980 47900 3984
rect 47964 3982 48010 4042
rect 48544 4040 48636 4042
rect 48544 3984 48594 4040
rect 48544 3982 48636 3984
rect 47964 3980 47970 3982
rect 48589 3980 48636 3982
rect 48700 3980 48706 4044
rect 58065 4042 58131 4045
rect 59200 4042 60000 4072
rect 58065 4040 60000 4042
rect 58065 3984 58070 4040
rect 58126 3984 60000 4040
rect 58065 3982 60000 3984
rect 47853 3979 47919 3980
rect 48589 3979 48655 3980
rect 58065 3979 58131 3982
rect 59200 3952 60000 3982
rect 27521 3904 31770 3906
rect 27521 3848 27526 3904
rect 27582 3848 31770 3904
rect 27521 3846 31770 3848
rect 39021 3906 39087 3909
rect 40217 3906 40283 3909
rect 39021 3904 40283 3906
rect 39021 3848 39026 3904
rect 39082 3848 40222 3904
rect 40278 3848 40283 3904
rect 39021 3846 40283 3848
rect 27521 3843 27587 3846
rect 39021 3843 39087 3846
rect 40217 3843 40283 3846
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 38469 3770 38535 3773
rect 47393 3770 47459 3773
rect 38469 3768 47459 3770
rect 38469 3712 38474 3768
rect 38530 3712 47398 3768
rect 47454 3712 47459 3768
rect 38469 3710 47459 3712
rect 38469 3707 38535 3710
rect 47393 3707 47459 3710
rect 24945 3634 25011 3637
rect 47669 3634 47735 3637
rect 24945 3632 47735 3634
rect 24945 3576 24950 3632
rect 25006 3576 47674 3632
rect 47730 3576 47735 3632
rect 24945 3574 47735 3576
rect 24945 3571 25011 3574
rect 47669 3571 47735 3574
rect 59200 3544 60000 3664
rect 16757 3498 16823 3501
rect 28901 3498 28967 3501
rect 16757 3496 28967 3498
rect 16757 3440 16762 3496
rect 16818 3440 28906 3496
rect 28962 3440 28967 3496
rect 16757 3438 28967 3440
rect 16757 3435 16823 3438
rect 28901 3435 28967 3438
rect 32857 3498 32923 3501
rect 42701 3498 42767 3501
rect 50429 3498 50495 3501
rect 32857 3496 42626 3498
rect 32857 3440 32862 3496
rect 32918 3440 42626 3496
rect 32857 3438 42626 3440
rect 32857 3435 32923 3438
rect 23105 3362 23171 3365
rect 25681 3362 25747 3365
rect 23105 3360 25747 3362
rect 23105 3304 23110 3360
rect 23166 3304 25686 3360
rect 25742 3304 25747 3360
rect 23105 3302 25747 3304
rect 23105 3299 23171 3302
rect 25681 3299 25747 3302
rect 33726 3300 33732 3364
rect 33796 3362 33802 3364
rect 41873 3362 41939 3365
rect 33796 3360 41939 3362
rect 33796 3304 41878 3360
rect 41934 3304 41939 3360
rect 33796 3302 41939 3304
rect 42566 3362 42626 3438
rect 42701 3496 50495 3498
rect 42701 3440 42706 3496
rect 42762 3440 50434 3496
rect 50490 3440 50495 3496
rect 42701 3438 50495 3440
rect 42701 3435 42767 3438
rect 50429 3435 50495 3438
rect 49877 3362 49943 3365
rect 42566 3360 49943 3362
rect 42566 3304 49882 3360
rect 49938 3304 49943 3360
rect 42566 3302 49943 3304
rect 33796 3300 33802 3302
rect 41873 3299 41939 3302
rect 49877 3299 49943 3302
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 50290 3296 50606 3297
rect 50290 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50606 3296
rect 50290 3231 50606 3232
rect 22829 3226 22895 3229
rect 36261 3226 36327 3229
rect 22829 3224 36327 3226
rect 22829 3168 22834 3224
rect 22890 3168 36266 3224
rect 36322 3168 36327 3224
rect 22829 3166 36327 3168
rect 22829 3163 22895 3166
rect 36261 3163 36327 3166
rect 43621 3226 43687 3229
rect 44449 3226 44515 3229
rect 43621 3224 44515 3226
rect 43621 3168 43626 3224
rect 43682 3168 44454 3224
rect 44510 3168 44515 3224
rect 43621 3166 44515 3168
rect 43621 3163 43687 3166
rect 44449 3163 44515 3166
rect 44633 3226 44699 3229
rect 44766 3226 44772 3228
rect 44633 3224 44772 3226
rect 44633 3168 44638 3224
rect 44694 3168 44772 3224
rect 44633 3166 44772 3168
rect 44633 3163 44699 3166
rect 44766 3164 44772 3166
rect 44836 3164 44842 3228
rect 55213 3226 55279 3229
rect 59200 3226 60000 3256
rect 55213 3224 60000 3226
rect 55213 3168 55218 3224
rect 55274 3168 60000 3224
rect 55213 3166 60000 3168
rect 55213 3163 55279 3166
rect 59200 3136 60000 3166
rect 17953 3090 18019 3093
rect 22553 3090 22619 3093
rect 17953 3088 22619 3090
rect 17953 3032 17958 3088
rect 18014 3032 22558 3088
rect 22614 3032 22619 3088
rect 17953 3030 22619 3032
rect 17953 3027 18019 3030
rect 22553 3027 22619 3030
rect 31017 3090 31083 3093
rect 43897 3090 43963 3093
rect 31017 3088 43963 3090
rect 31017 3032 31022 3088
rect 31078 3032 43902 3088
rect 43958 3032 43963 3088
rect 31017 3030 43963 3032
rect 31017 3027 31083 3030
rect 43897 3027 43963 3030
rect 48405 3090 48471 3093
rect 48589 3090 48655 3093
rect 48405 3088 48655 3090
rect 48405 3032 48410 3088
rect 48466 3032 48594 3088
rect 48650 3032 48655 3088
rect 48405 3030 48655 3032
rect 48405 3027 48471 3030
rect 48589 3027 48655 3030
rect 22645 2954 22711 2957
rect 23565 2954 23631 2957
rect 22645 2952 23631 2954
rect 22645 2896 22650 2952
rect 22706 2896 23570 2952
rect 23626 2896 23631 2952
rect 22645 2894 23631 2896
rect 22645 2891 22711 2894
rect 23565 2891 23631 2894
rect 30782 2892 30788 2956
rect 30852 2954 30858 2956
rect 49233 2954 49299 2957
rect 30852 2952 49299 2954
rect 30852 2896 49238 2952
rect 49294 2896 49299 2952
rect 30852 2894 49299 2896
rect 30852 2892 30858 2894
rect 49233 2891 49299 2894
rect 58893 2818 58959 2821
rect 59200 2818 60000 2848
rect 58893 2816 60000 2818
rect 58893 2760 58898 2816
rect 58954 2760 60000 2816
rect 58893 2758 60000 2760
rect 58893 2755 58959 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 59200 2728 60000 2758
rect 34930 2687 35246 2688
rect 41413 2684 41479 2685
rect 41413 2682 41460 2684
rect 41368 2680 41460 2682
rect 41368 2624 41418 2680
rect 41368 2622 41460 2624
rect 41413 2620 41460 2622
rect 41524 2620 41530 2684
rect 47945 2682 48011 2685
rect 48078 2682 48084 2684
rect 47945 2680 48084 2682
rect 47945 2624 47950 2680
rect 48006 2624 48084 2680
rect 47945 2622 48084 2624
rect 41413 2619 41479 2620
rect 47945 2619 48011 2622
rect 48078 2620 48084 2622
rect 48148 2620 48154 2684
rect 38377 2546 38443 2549
rect 52453 2546 52519 2549
rect 38377 2544 52519 2546
rect 38377 2488 38382 2544
rect 38438 2488 52458 2544
rect 52514 2488 52519 2544
rect 38377 2486 52519 2488
rect 38377 2483 38443 2486
rect 52453 2483 52519 2486
rect 25221 2410 25287 2413
rect 48814 2410 48820 2412
rect 25221 2408 48820 2410
rect 25221 2352 25226 2408
rect 25282 2352 48820 2408
rect 25221 2350 48820 2352
rect 25221 2347 25287 2350
rect 48814 2348 48820 2350
rect 48884 2348 48890 2412
rect 58985 2410 59051 2413
rect 59200 2410 60000 2440
rect 58985 2408 60000 2410
rect 58985 2352 58990 2408
rect 59046 2352 60000 2408
rect 58985 2350 60000 2352
rect 58985 2347 59051 2350
rect 59200 2320 60000 2350
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 50290 2208 50606 2209
rect 50290 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50606 2208
rect 50290 2143 50606 2144
rect 58893 2002 58959 2005
rect 59200 2002 60000 2032
rect 58893 2000 60000 2002
rect 58893 1944 58898 2000
rect 58954 1944 60000 2000
rect 58893 1942 60000 1944
rect 58893 1939 58959 1942
rect 59200 1912 60000 1942
rect 58801 1594 58867 1597
rect 59200 1594 60000 1624
rect 58801 1592 60000 1594
rect 58801 1536 58806 1592
rect 58862 1536 60000 1592
rect 58801 1534 60000 1536
rect 58801 1531 58867 1534
rect 59200 1504 60000 1534
rect 55857 1186 55923 1189
rect 59200 1186 60000 1216
rect 55857 1184 60000 1186
rect 55857 1128 55862 1184
rect 55918 1128 60000 1184
rect 55857 1126 60000 1128
rect 55857 1123 55923 1126
rect 59200 1096 60000 1126
<< via3 >>
rect 19576 57692 19640 57696
rect 19576 57636 19580 57692
rect 19580 57636 19636 57692
rect 19636 57636 19640 57692
rect 19576 57632 19640 57636
rect 19656 57692 19720 57696
rect 19656 57636 19660 57692
rect 19660 57636 19716 57692
rect 19716 57636 19720 57692
rect 19656 57632 19720 57636
rect 19736 57692 19800 57696
rect 19736 57636 19740 57692
rect 19740 57636 19796 57692
rect 19796 57636 19800 57692
rect 19736 57632 19800 57636
rect 19816 57692 19880 57696
rect 19816 57636 19820 57692
rect 19820 57636 19876 57692
rect 19876 57636 19880 57692
rect 19816 57632 19880 57636
rect 50296 57692 50360 57696
rect 50296 57636 50300 57692
rect 50300 57636 50356 57692
rect 50356 57636 50360 57692
rect 50296 57632 50360 57636
rect 50376 57692 50440 57696
rect 50376 57636 50380 57692
rect 50380 57636 50436 57692
rect 50436 57636 50440 57692
rect 50376 57632 50440 57636
rect 50456 57692 50520 57696
rect 50456 57636 50460 57692
rect 50460 57636 50516 57692
rect 50516 57636 50520 57692
rect 50456 57632 50520 57636
rect 50536 57692 50600 57696
rect 50536 57636 50540 57692
rect 50540 57636 50596 57692
rect 50596 57636 50600 57692
rect 50536 57632 50600 57636
rect 4216 57148 4280 57152
rect 4216 57092 4220 57148
rect 4220 57092 4276 57148
rect 4276 57092 4280 57148
rect 4216 57088 4280 57092
rect 4296 57148 4360 57152
rect 4296 57092 4300 57148
rect 4300 57092 4356 57148
rect 4356 57092 4360 57148
rect 4296 57088 4360 57092
rect 4376 57148 4440 57152
rect 4376 57092 4380 57148
rect 4380 57092 4436 57148
rect 4436 57092 4440 57148
rect 4376 57088 4440 57092
rect 4456 57148 4520 57152
rect 4456 57092 4460 57148
rect 4460 57092 4516 57148
rect 4516 57092 4520 57148
rect 4456 57088 4520 57092
rect 34936 57148 35000 57152
rect 34936 57092 34940 57148
rect 34940 57092 34996 57148
rect 34996 57092 35000 57148
rect 34936 57088 35000 57092
rect 35016 57148 35080 57152
rect 35016 57092 35020 57148
rect 35020 57092 35076 57148
rect 35076 57092 35080 57148
rect 35016 57088 35080 57092
rect 35096 57148 35160 57152
rect 35096 57092 35100 57148
rect 35100 57092 35156 57148
rect 35156 57092 35160 57148
rect 35096 57088 35160 57092
rect 35176 57148 35240 57152
rect 35176 57092 35180 57148
rect 35180 57092 35236 57148
rect 35236 57092 35240 57148
rect 35176 57088 35240 57092
rect 48452 56612 48516 56676
rect 19576 56604 19640 56608
rect 19576 56548 19580 56604
rect 19580 56548 19636 56604
rect 19636 56548 19640 56604
rect 19576 56544 19640 56548
rect 19656 56604 19720 56608
rect 19656 56548 19660 56604
rect 19660 56548 19716 56604
rect 19716 56548 19720 56604
rect 19656 56544 19720 56548
rect 19736 56604 19800 56608
rect 19736 56548 19740 56604
rect 19740 56548 19796 56604
rect 19796 56548 19800 56604
rect 19736 56544 19800 56548
rect 19816 56604 19880 56608
rect 19816 56548 19820 56604
rect 19820 56548 19876 56604
rect 19876 56548 19880 56604
rect 19816 56544 19880 56548
rect 50296 56604 50360 56608
rect 50296 56548 50300 56604
rect 50300 56548 50356 56604
rect 50356 56548 50360 56604
rect 50296 56544 50360 56548
rect 50376 56604 50440 56608
rect 50376 56548 50380 56604
rect 50380 56548 50436 56604
rect 50436 56548 50440 56604
rect 50376 56544 50440 56548
rect 50456 56604 50520 56608
rect 50456 56548 50460 56604
rect 50460 56548 50516 56604
rect 50516 56548 50520 56604
rect 50456 56544 50520 56548
rect 50536 56604 50600 56608
rect 50536 56548 50540 56604
rect 50540 56548 50596 56604
rect 50596 56548 50600 56604
rect 50536 56544 50600 56548
rect 4216 56060 4280 56064
rect 4216 56004 4220 56060
rect 4220 56004 4276 56060
rect 4276 56004 4280 56060
rect 4216 56000 4280 56004
rect 4296 56060 4360 56064
rect 4296 56004 4300 56060
rect 4300 56004 4356 56060
rect 4356 56004 4360 56060
rect 4296 56000 4360 56004
rect 4376 56060 4440 56064
rect 4376 56004 4380 56060
rect 4380 56004 4436 56060
rect 4436 56004 4440 56060
rect 4376 56000 4440 56004
rect 4456 56060 4520 56064
rect 4456 56004 4460 56060
rect 4460 56004 4516 56060
rect 4516 56004 4520 56060
rect 4456 56000 4520 56004
rect 34936 56060 35000 56064
rect 34936 56004 34940 56060
rect 34940 56004 34996 56060
rect 34996 56004 35000 56060
rect 34936 56000 35000 56004
rect 35016 56060 35080 56064
rect 35016 56004 35020 56060
rect 35020 56004 35076 56060
rect 35076 56004 35080 56060
rect 35016 56000 35080 56004
rect 35096 56060 35160 56064
rect 35096 56004 35100 56060
rect 35100 56004 35156 56060
rect 35156 56004 35160 56060
rect 35096 56000 35160 56004
rect 35176 56060 35240 56064
rect 35176 56004 35180 56060
rect 35180 56004 35236 56060
rect 35236 56004 35240 56060
rect 35176 56000 35240 56004
rect 19576 55516 19640 55520
rect 19576 55460 19580 55516
rect 19580 55460 19636 55516
rect 19636 55460 19640 55516
rect 19576 55456 19640 55460
rect 19656 55516 19720 55520
rect 19656 55460 19660 55516
rect 19660 55460 19716 55516
rect 19716 55460 19720 55516
rect 19656 55456 19720 55460
rect 19736 55516 19800 55520
rect 19736 55460 19740 55516
rect 19740 55460 19796 55516
rect 19796 55460 19800 55516
rect 19736 55456 19800 55460
rect 19816 55516 19880 55520
rect 19816 55460 19820 55516
rect 19820 55460 19876 55516
rect 19876 55460 19880 55516
rect 19816 55456 19880 55460
rect 50296 55516 50360 55520
rect 50296 55460 50300 55516
rect 50300 55460 50356 55516
rect 50356 55460 50360 55516
rect 50296 55456 50360 55460
rect 50376 55516 50440 55520
rect 50376 55460 50380 55516
rect 50380 55460 50436 55516
rect 50436 55460 50440 55516
rect 50376 55456 50440 55460
rect 50456 55516 50520 55520
rect 50456 55460 50460 55516
rect 50460 55460 50516 55516
rect 50516 55460 50520 55516
rect 50456 55456 50520 55460
rect 50536 55516 50600 55520
rect 50536 55460 50540 55516
rect 50540 55460 50596 55516
rect 50596 55460 50600 55516
rect 50536 55456 50600 55460
rect 4216 54972 4280 54976
rect 4216 54916 4220 54972
rect 4220 54916 4276 54972
rect 4276 54916 4280 54972
rect 4216 54912 4280 54916
rect 4296 54972 4360 54976
rect 4296 54916 4300 54972
rect 4300 54916 4356 54972
rect 4356 54916 4360 54972
rect 4296 54912 4360 54916
rect 4376 54972 4440 54976
rect 4376 54916 4380 54972
rect 4380 54916 4436 54972
rect 4436 54916 4440 54972
rect 4376 54912 4440 54916
rect 4456 54972 4520 54976
rect 4456 54916 4460 54972
rect 4460 54916 4516 54972
rect 4516 54916 4520 54972
rect 4456 54912 4520 54916
rect 34936 54972 35000 54976
rect 34936 54916 34940 54972
rect 34940 54916 34996 54972
rect 34996 54916 35000 54972
rect 34936 54912 35000 54916
rect 35016 54972 35080 54976
rect 35016 54916 35020 54972
rect 35020 54916 35076 54972
rect 35076 54916 35080 54972
rect 35016 54912 35080 54916
rect 35096 54972 35160 54976
rect 35096 54916 35100 54972
rect 35100 54916 35156 54972
rect 35156 54916 35160 54972
rect 35096 54912 35160 54916
rect 35176 54972 35240 54976
rect 35176 54916 35180 54972
rect 35180 54916 35236 54972
rect 35236 54916 35240 54972
rect 35176 54912 35240 54916
rect 19576 54428 19640 54432
rect 19576 54372 19580 54428
rect 19580 54372 19636 54428
rect 19636 54372 19640 54428
rect 19576 54368 19640 54372
rect 19656 54428 19720 54432
rect 19656 54372 19660 54428
rect 19660 54372 19716 54428
rect 19716 54372 19720 54428
rect 19656 54368 19720 54372
rect 19736 54428 19800 54432
rect 19736 54372 19740 54428
rect 19740 54372 19796 54428
rect 19796 54372 19800 54428
rect 19736 54368 19800 54372
rect 19816 54428 19880 54432
rect 19816 54372 19820 54428
rect 19820 54372 19876 54428
rect 19876 54372 19880 54428
rect 19816 54368 19880 54372
rect 50296 54428 50360 54432
rect 50296 54372 50300 54428
rect 50300 54372 50356 54428
rect 50356 54372 50360 54428
rect 50296 54368 50360 54372
rect 50376 54428 50440 54432
rect 50376 54372 50380 54428
rect 50380 54372 50436 54428
rect 50436 54372 50440 54428
rect 50376 54368 50440 54372
rect 50456 54428 50520 54432
rect 50456 54372 50460 54428
rect 50460 54372 50516 54428
rect 50516 54372 50520 54428
rect 50456 54368 50520 54372
rect 50536 54428 50600 54432
rect 50536 54372 50540 54428
rect 50540 54372 50596 54428
rect 50596 54372 50600 54428
rect 50536 54368 50600 54372
rect 4216 53884 4280 53888
rect 4216 53828 4220 53884
rect 4220 53828 4276 53884
rect 4276 53828 4280 53884
rect 4216 53824 4280 53828
rect 4296 53884 4360 53888
rect 4296 53828 4300 53884
rect 4300 53828 4356 53884
rect 4356 53828 4360 53884
rect 4296 53824 4360 53828
rect 4376 53884 4440 53888
rect 4376 53828 4380 53884
rect 4380 53828 4436 53884
rect 4436 53828 4440 53884
rect 4376 53824 4440 53828
rect 4456 53884 4520 53888
rect 4456 53828 4460 53884
rect 4460 53828 4516 53884
rect 4516 53828 4520 53884
rect 4456 53824 4520 53828
rect 34936 53884 35000 53888
rect 34936 53828 34940 53884
rect 34940 53828 34996 53884
rect 34996 53828 35000 53884
rect 34936 53824 35000 53828
rect 35016 53884 35080 53888
rect 35016 53828 35020 53884
rect 35020 53828 35076 53884
rect 35076 53828 35080 53884
rect 35016 53824 35080 53828
rect 35096 53884 35160 53888
rect 35096 53828 35100 53884
rect 35100 53828 35156 53884
rect 35156 53828 35160 53884
rect 35096 53824 35160 53828
rect 35176 53884 35240 53888
rect 35176 53828 35180 53884
rect 35180 53828 35236 53884
rect 35236 53828 35240 53884
rect 35176 53824 35240 53828
rect 19576 53340 19640 53344
rect 19576 53284 19580 53340
rect 19580 53284 19636 53340
rect 19636 53284 19640 53340
rect 19576 53280 19640 53284
rect 19656 53340 19720 53344
rect 19656 53284 19660 53340
rect 19660 53284 19716 53340
rect 19716 53284 19720 53340
rect 19656 53280 19720 53284
rect 19736 53340 19800 53344
rect 19736 53284 19740 53340
rect 19740 53284 19796 53340
rect 19796 53284 19800 53340
rect 19736 53280 19800 53284
rect 19816 53340 19880 53344
rect 19816 53284 19820 53340
rect 19820 53284 19876 53340
rect 19876 53284 19880 53340
rect 19816 53280 19880 53284
rect 50296 53340 50360 53344
rect 50296 53284 50300 53340
rect 50300 53284 50356 53340
rect 50356 53284 50360 53340
rect 50296 53280 50360 53284
rect 50376 53340 50440 53344
rect 50376 53284 50380 53340
rect 50380 53284 50436 53340
rect 50436 53284 50440 53340
rect 50376 53280 50440 53284
rect 50456 53340 50520 53344
rect 50456 53284 50460 53340
rect 50460 53284 50516 53340
rect 50516 53284 50520 53340
rect 50456 53280 50520 53284
rect 50536 53340 50600 53344
rect 50536 53284 50540 53340
rect 50540 53284 50596 53340
rect 50596 53284 50600 53340
rect 50536 53280 50600 53284
rect 4216 52796 4280 52800
rect 4216 52740 4220 52796
rect 4220 52740 4276 52796
rect 4276 52740 4280 52796
rect 4216 52736 4280 52740
rect 4296 52796 4360 52800
rect 4296 52740 4300 52796
rect 4300 52740 4356 52796
rect 4356 52740 4360 52796
rect 4296 52736 4360 52740
rect 4376 52796 4440 52800
rect 4376 52740 4380 52796
rect 4380 52740 4436 52796
rect 4436 52740 4440 52796
rect 4376 52736 4440 52740
rect 4456 52796 4520 52800
rect 4456 52740 4460 52796
rect 4460 52740 4516 52796
rect 4516 52740 4520 52796
rect 4456 52736 4520 52740
rect 34936 52796 35000 52800
rect 34936 52740 34940 52796
rect 34940 52740 34996 52796
rect 34996 52740 35000 52796
rect 34936 52736 35000 52740
rect 35016 52796 35080 52800
rect 35016 52740 35020 52796
rect 35020 52740 35076 52796
rect 35076 52740 35080 52796
rect 35016 52736 35080 52740
rect 35096 52796 35160 52800
rect 35096 52740 35100 52796
rect 35100 52740 35156 52796
rect 35156 52740 35160 52796
rect 35096 52736 35160 52740
rect 35176 52796 35240 52800
rect 35176 52740 35180 52796
rect 35180 52740 35236 52796
rect 35236 52740 35240 52796
rect 35176 52736 35240 52740
rect 48084 52668 48148 52732
rect 47900 52532 47964 52596
rect 19576 52252 19640 52256
rect 19576 52196 19580 52252
rect 19580 52196 19636 52252
rect 19636 52196 19640 52252
rect 19576 52192 19640 52196
rect 19656 52252 19720 52256
rect 19656 52196 19660 52252
rect 19660 52196 19716 52252
rect 19716 52196 19720 52252
rect 19656 52192 19720 52196
rect 19736 52252 19800 52256
rect 19736 52196 19740 52252
rect 19740 52196 19796 52252
rect 19796 52196 19800 52252
rect 19736 52192 19800 52196
rect 19816 52252 19880 52256
rect 19816 52196 19820 52252
rect 19820 52196 19876 52252
rect 19876 52196 19880 52252
rect 19816 52192 19880 52196
rect 50296 52252 50360 52256
rect 50296 52196 50300 52252
rect 50300 52196 50356 52252
rect 50356 52196 50360 52252
rect 50296 52192 50360 52196
rect 50376 52252 50440 52256
rect 50376 52196 50380 52252
rect 50380 52196 50436 52252
rect 50436 52196 50440 52252
rect 50376 52192 50440 52196
rect 50456 52252 50520 52256
rect 50456 52196 50460 52252
rect 50460 52196 50516 52252
rect 50516 52196 50520 52252
rect 50456 52192 50520 52196
rect 50536 52252 50600 52256
rect 50536 52196 50540 52252
rect 50540 52196 50596 52252
rect 50596 52196 50600 52252
rect 50536 52192 50600 52196
rect 4216 51708 4280 51712
rect 4216 51652 4220 51708
rect 4220 51652 4276 51708
rect 4276 51652 4280 51708
rect 4216 51648 4280 51652
rect 4296 51708 4360 51712
rect 4296 51652 4300 51708
rect 4300 51652 4356 51708
rect 4356 51652 4360 51708
rect 4296 51648 4360 51652
rect 4376 51708 4440 51712
rect 4376 51652 4380 51708
rect 4380 51652 4436 51708
rect 4436 51652 4440 51708
rect 4376 51648 4440 51652
rect 4456 51708 4520 51712
rect 4456 51652 4460 51708
rect 4460 51652 4516 51708
rect 4516 51652 4520 51708
rect 4456 51648 4520 51652
rect 34936 51708 35000 51712
rect 34936 51652 34940 51708
rect 34940 51652 34996 51708
rect 34996 51652 35000 51708
rect 34936 51648 35000 51652
rect 35016 51708 35080 51712
rect 35016 51652 35020 51708
rect 35020 51652 35076 51708
rect 35076 51652 35080 51708
rect 35016 51648 35080 51652
rect 35096 51708 35160 51712
rect 35096 51652 35100 51708
rect 35100 51652 35156 51708
rect 35156 51652 35160 51708
rect 35096 51648 35160 51652
rect 35176 51708 35240 51712
rect 35176 51652 35180 51708
rect 35180 51652 35236 51708
rect 35236 51652 35240 51708
rect 35176 51648 35240 51652
rect 19576 51164 19640 51168
rect 19576 51108 19580 51164
rect 19580 51108 19636 51164
rect 19636 51108 19640 51164
rect 19576 51104 19640 51108
rect 19656 51164 19720 51168
rect 19656 51108 19660 51164
rect 19660 51108 19716 51164
rect 19716 51108 19720 51164
rect 19656 51104 19720 51108
rect 19736 51164 19800 51168
rect 19736 51108 19740 51164
rect 19740 51108 19796 51164
rect 19796 51108 19800 51164
rect 19736 51104 19800 51108
rect 19816 51164 19880 51168
rect 19816 51108 19820 51164
rect 19820 51108 19876 51164
rect 19876 51108 19880 51164
rect 19816 51104 19880 51108
rect 50296 51164 50360 51168
rect 50296 51108 50300 51164
rect 50300 51108 50356 51164
rect 50356 51108 50360 51164
rect 50296 51104 50360 51108
rect 50376 51164 50440 51168
rect 50376 51108 50380 51164
rect 50380 51108 50436 51164
rect 50436 51108 50440 51164
rect 50376 51104 50440 51108
rect 50456 51164 50520 51168
rect 50456 51108 50460 51164
rect 50460 51108 50516 51164
rect 50516 51108 50520 51164
rect 50456 51104 50520 51108
rect 50536 51164 50600 51168
rect 50536 51108 50540 51164
rect 50540 51108 50596 51164
rect 50596 51108 50600 51164
rect 50536 51104 50600 51108
rect 47716 51096 47780 51100
rect 47716 51040 47766 51096
rect 47766 51040 47780 51096
rect 47716 51036 47780 51040
rect 4216 50620 4280 50624
rect 4216 50564 4220 50620
rect 4220 50564 4276 50620
rect 4276 50564 4280 50620
rect 4216 50560 4280 50564
rect 4296 50620 4360 50624
rect 4296 50564 4300 50620
rect 4300 50564 4356 50620
rect 4356 50564 4360 50620
rect 4296 50560 4360 50564
rect 4376 50620 4440 50624
rect 4376 50564 4380 50620
rect 4380 50564 4436 50620
rect 4436 50564 4440 50620
rect 4376 50560 4440 50564
rect 4456 50620 4520 50624
rect 4456 50564 4460 50620
rect 4460 50564 4516 50620
rect 4516 50564 4520 50620
rect 4456 50560 4520 50564
rect 34936 50620 35000 50624
rect 34936 50564 34940 50620
rect 34940 50564 34996 50620
rect 34996 50564 35000 50620
rect 34936 50560 35000 50564
rect 35016 50620 35080 50624
rect 35016 50564 35020 50620
rect 35020 50564 35076 50620
rect 35076 50564 35080 50620
rect 35016 50560 35080 50564
rect 35096 50620 35160 50624
rect 35096 50564 35100 50620
rect 35100 50564 35156 50620
rect 35156 50564 35160 50620
rect 35096 50560 35160 50564
rect 35176 50620 35240 50624
rect 35176 50564 35180 50620
rect 35180 50564 35236 50620
rect 35236 50564 35240 50620
rect 35176 50560 35240 50564
rect 19576 50076 19640 50080
rect 19576 50020 19580 50076
rect 19580 50020 19636 50076
rect 19636 50020 19640 50076
rect 19576 50016 19640 50020
rect 19656 50076 19720 50080
rect 19656 50020 19660 50076
rect 19660 50020 19716 50076
rect 19716 50020 19720 50076
rect 19656 50016 19720 50020
rect 19736 50076 19800 50080
rect 19736 50020 19740 50076
rect 19740 50020 19796 50076
rect 19796 50020 19800 50076
rect 19736 50016 19800 50020
rect 19816 50076 19880 50080
rect 19816 50020 19820 50076
rect 19820 50020 19876 50076
rect 19876 50020 19880 50076
rect 19816 50016 19880 50020
rect 50296 50076 50360 50080
rect 50296 50020 50300 50076
rect 50300 50020 50356 50076
rect 50356 50020 50360 50076
rect 50296 50016 50360 50020
rect 50376 50076 50440 50080
rect 50376 50020 50380 50076
rect 50380 50020 50436 50076
rect 50436 50020 50440 50076
rect 50376 50016 50440 50020
rect 50456 50076 50520 50080
rect 50456 50020 50460 50076
rect 50460 50020 50516 50076
rect 50516 50020 50520 50076
rect 50456 50016 50520 50020
rect 50536 50076 50600 50080
rect 50536 50020 50540 50076
rect 50540 50020 50596 50076
rect 50596 50020 50600 50076
rect 50536 50016 50600 50020
rect 42564 49736 42628 49740
rect 42564 49680 42614 49736
rect 42614 49680 42628 49736
rect 42564 49676 42628 49680
rect 4216 49532 4280 49536
rect 4216 49476 4220 49532
rect 4220 49476 4276 49532
rect 4276 49476 4280 49532
rect 4216 49472 4280 49476
rect 4296 49532 4360 49536
rect 4296 49476 4300 49532
rect 4300 49476 4356 49532
rect 4356 49476 4360 49532
rect 4296 49472 4360 49476
rect 4376 49532 4440 49536
rect 4376 49476 4380 49532
rect 4380 49476 4436 49532
rect 4436 49476 4440 49532
rect 4376 49472 4440 49476
rect 4456 49532 4520 49536
rect 4456 49476 4460 49532
rect 4460 49476 4516 49532
rect 4516 49476 4520 49532
rect 4456 49472 4520 49476
rect 34936 49532 35000 49536
rect 34936 49476 34940 49532
rect 34940 49476 34996 49532
rect 34996 49476 35000 49532
rect 34936 49472 35000 49476
rect 35016 49532 35080 49536
rect 35016 49476 35020 49532
rect 35020 49476 35076 49532
rect 35076 49476 35080 49532
rect 35016 49472 35080 49476
rect 35096 49532 35160 49536
rect 35096 49476 35100 49532
rect 35100 49476 35156 49532
rect 35156 49476 35160 49532
rect 35096 49472 35160 49476
rect 35176 49532 35240 49536
rect 35176 49476 35180 49532
rect 35180 49476 35236 49532
rect 35236 49476 35240 49532
rect 35176 49472 35240 49476
rect 19576 48988 19640 48992
rect 19576 48932 19580 48988
rect 19580 48932 19636 48988
rect 19636 48932 19640 48988
rect 19576 48928 19640 48932
rect 19656 48988 19720 48992
rect 19656 48932 19660 48988
rect 19660 48932 19716 48988
rect 19716 48932 19720 48988
rect 19656 48928 19720 48932
rect 19736 48988 19800 48992
rect 19736 48932 19740 48988
rect 19740 48932 19796 48988
rect 19796 48932 19800 48988
rect 19736 48928 19800 48932
rect 19816 48988 19880 48992
rect 19816 48932 19820 48988
rect 19820 48932 19876 48988
rect 19876 48932 19880 48988
rect 19816 48928 19880 48932
rect 50296 48988 50360 48992
rect 50296 48932 50300 48988
rect 50300 48932 50356 48988
rect 50356 48932 50360 48988
rect 50296 48928 50360 48932
rect 50376 48988 50440 48992
rect 50376 48932 50380 48988
rect 50380 48932 50436 48988
rect 50436 48932 50440 48988
rect 50376 48928 50440 48932
rect 50456 48988 50520 48992
rect 50456 48932 50460 48988
rect 50460 48932 50516 48988
rect 50516 48932 50520 48988
rect 50456 48928 50520 48932
rect 50536 48988 50600 48992
rect 50536 48932 50540 48988
rect 50540 48932 50596 48988
rect 50596 48932 50600 48988
rect 50536 48928 50600 48932
rect 4216 48444 4280 48448
rect 4216 48388 4220 48444
rect 4220 48388 4276 48444
rect 4276 48388 4280 48444
rect 4216 48384 4280 48388
rect 4296 48444 4360 48448
rect 4296 48388 4300 48444
rect 4300 48388 4356 48444
rect 4356 48388 4360 48444
rect 4296 48384 4360 48388
rect 4376 48444 4440 48448
rect 4376 48388 4380 48444
rect 4380 48388 4436 48444
rect 4436 48388 4440 48444
rect 4376 48384 4440 48388
rect 4456 48444 4520 48448
rect 4456 48388 4460 48444
rect 4460 48388 4516 48444
rect 4516 48388 4520 48444
rect 4456 48384 4520 48388
rect 34936 48444 35000 48448
rect 34936 48388 34940 48444
rect 34940 48388 34996 48444
rect 34996 48388 35000 48444
rect 34936 48384 35000 48388
rect 35016 48444 35080 48448
rect 35016 48388 35020 48444
rect 35020 48388 35076 48444
rect 35076 48388 35080 48444
rect 35016 48384 35080 48388
rect 35096 48444 35160 48448
rect 35096 48388 35100 48444
rect 35100 48388 35156 48444
rect 35156 48388 35160 48444
rect 35096 48384 35160 48388
rect 35176 48444 35240 48448
rect 35176 48388 35180 48444
rect 35180 48388 35236 48444
rect 35236 48388 35240 48444
rect 35176 48384 35240 48388
rect 19576 47900 19640 47904
rect 19576 47844 19580 47900
rect 19580 47844 19636 47900
rect 19636 47844 19640 47900
rect 19576 47840 19640 47844
rect 19656 47900 19720 47904
rect 19656 47844 19660 47900
rect 19660 47844 19716 47900
rect 19716 47844 19720 47900
rect 19656 47840 19720 47844
rect 19736 47900 19800 47904
rect 19736 47844 19740 47900
rect 19740 47844 19796 47900
rect 19796 47844 19800 47900
rect 19736 47840 19800 47844
rect 19816 47900 19880 47904
rect 19816 47844 19820 47900
rect 19820 47844 19876 47900
rect 19876 47844 19880 47900
rect 19816 47840 19880 47844
rect 50296 47900 50360 47904
rect 50296 47844 50300 47900
rect 50300 47844 50356 47900
rect 50356 47844 50360 47900
rect 50296 47840 50360 47844
rect 50376 47900 50440 47904
rect 50376 47844 50380 47900
rect 50380 47844 50436 47900
rect 50436 47844 50440 47900
rect 50376 47840 50440 47844
rect 50456 47900 50520 47904
rect 50456 47844 50460 47900
rect 50460 47844 50516 47900
rect 50516 47844 50520 47900
rect 50456 47840 50520 47844
rect 50536 47900 50600 47904
rect 50536 47844 50540 47900
rect 50540 47844 50596 47900
rect 50596 47844 50600 47900
rect 50536 47840 50600 47844
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 50296 46812 50360 46816
rect 50296 46756 50300 46812
rect 50300 46756 50356 46812
rect 50356 46756 50360 46812
rect 50296 46752 50360 46756
rect 50376 46812 50440 46816
rect 50376 46756 50380 46812
rect 50380 46756 50436 46812
rect 50436 46756 50440 46812
rect 50376 46752 50440 46756
rect 50456 46812 50520 46816
rect 50456 46756 50460 46812
rect 50460 46756 50516 46812
rect 50516 46756 50520 46812
rect 50456 46752 50520 46756
rect 50536 46812 50600 46816
rect 50536 46756 50540 46812
rect 50540 46756 50596 46812
rect 50596 46756 50600 46812
rect 50536 46752 50600 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 50296 45724 50360 45728
rect 50296 45668 50300 45724
rect 50300 45668 50356 45724
rect 50356 45668 50360 45724
rect 50296 45664 50360 45668
rect 50376 45724 50440 45728
rect 50376 45668 50380 45724
rect 50380 45668 50436 45724
rect 50436 45668 50440 45724
rect 50376 45664 50440 45668
rect 50456 45724 50520 45728
rect 50456 45668 50460 45724
rect 50460 45668 50516 45724
rect 50516 45668 50520 45724
rect 50456 45664 50520 45668
rect 50536 45724 50600 45728
rect 50536 45668 50540 45724
rect 50540 45668 50596 45724
rect 50596 45668 50600 45724
rect 50536 45664 50600 45668
rect 40540 45460 40604 45524
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 50296 44636 50360 44640
rect 50296 44580 50300 44636
rect 50300 44580 50356 44636
rect 50356 44580 50360 44636
rect 50296 44576 50360 44580
rect 50376 44636 50440 44640
rect 50376 44580 50380 44636
rect 50380 44580 50436 44636
rect 50436 44580 50440 44636
rect 50376 44576 50440 44580
rect 50456 44636 50520 44640
rect 50456 44580 50460 44636
rect 50460 44580 50516 44636
rect 50516 44580 50520 44636
rect 50456 44576 50520 44580
rect 50536 44636 50600 44640
rect 50536 44580 50540 44636
rect 50540 44580 50596 44636
rect 50596 44580 50600 44636
rect 50536 44576 50600 44580
rect 48636 44296 48700 44300
rect 48636 44240 48686 44296
rect 48686 44240 48700 44296
rect 48636 44236 48700 44240
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 50296 43548 50360 43552
rect 50296 43492 50300 43548
rect 50300 43492 50356 43548
rect 50356 43492 50360 43548
rect 50296 43488 50360 43492
rect 50376 43548 50440 43552
rect 50376 43492 50380 43548
rect 50380 43492 50436 43548
rect 50436 43492 50440 43548
rect 50376 43488 50440 43492
rect 50456 43548 50520 43552
rect 50456 43492 50460 43548
rect 50460 43492 50516 43548
rect 50516 43492 50520 43548
rect 50456 43488 50520 43492
rect 50536 43548 50600 43552
rect 50536 43492 50540 43548
rect 50540 43492 50596 43548
rect 50596 43492 50600 43548
rect 50536 43488 50600 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 41276 42936 41340 42940
rect 41276 42880 41326 42936
rect 41326 42880 41340 42936
rect 41276 42876 41340 42880
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 50296 42460 50360 42464
rect 50296 42404 50300 42460
rect 50300 42404 50356 42460
rect 50356 42404 50360 42460
rect 50296 42400 50360 42404
rect 50376 42460 50440 42464
rect 50376 42404 50380 42460
rect 50380 42404 50436 42460
rect 50436 42404 50440 42460
rect 50376 42400 50440 42404
rect 50456 42460 50520 42464
rect 50456 42404 50460 42460
rect 50460 42404 50516 42460
rect 50516 42404 50520 42460
rect 50456 42400 50520 42404
rect 50536 42460 50600 42464
rect 50536 42404 50540 42460
rect 50540 42404 50596 42460
rect 50596 42404 50600 42460
rect 50536 42400 50600 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 44404 41380 44468 41444
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 50296 41372 50360 41376
rect 50296 41316 50300 41372
rect 50300 41316 50356 41372
rect 50356 41316 50360 41372
rect 50296 41312 50360 41316
rect 50376 41372 50440 41376
rect 50376 41316 50380 41372
rect 50380 41316 50436 41372
rect 50436 41316 50440 41372
rect 50376 41312 50440 41316
rect 50456 41372 50520 41376
rect 50456 41316 50460 41372
rect 50460 41316 50516 41372
rect 50516 41316 50520 41372
rect 50456 41312 50520 41316
rect 50536 41372 50600 41376
rect 50536 41316 50540 41372
rect 50540 41316 50596 41372
rect 50596 41316 50600 41372
rect 50536 41312 50600 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 50296 40284 50360 40288
rect 50296 40228 50300 40284
rect 50300 40228 50356 40284
rect 50356 40228 50360 40284
rect 50296 40224 50360 40228
rect 50376 40284 50440 40288
rect 50376 40228 50380 40284
rect 50380 40228 50436 40284
rect 50436 40228 50440 40284
rect 50376 40224 50440 40228
rect 50456 40284 50520 40288
rect 50456 40228 50460 40284
rect 50460 40228 50516 40284
rect 50516 40228 50520 40284
rect 50456 40224 50520 40228
rect 50536 40284 50600 40288
rect 50536 40228 50540 40284
rect 50540 40228 50596 40284
rect 50596 40228 50600 40284
rect 50536 40224 50600 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 50296 39196 50360 39200
rect 50296 39140 50300 39196
rect 50300 39140 50356 39196
rect 50356 39140 50360 39196
rect 50296 39136 50360 39140
rect 50376 39196 50440 39200
rect 50376 39140 50380 39196
rect 50380 39140 50436 39196
rect 50436 39140 50440 39196
rect 50376 39136 50440 39140
rect 50456 39196 50520 39200
rect 50456 39140 50460 39196
rect 50460 39140 50516 39196
rect 50516 39140 50520 39196
rect 50456 39136 50520 39140
rect 50536 39196 50600 39200
rect 50536 39140 50540 39196
rect 50540 39140 50596 39196
rect 50596 39140 50600 39196
rect 50536 39136 50600 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 50296 38108 50360 38112
rect 50296 38052 50300 38108
rect 50300 38052 50356 38108
rect 50356 38052 50360 38108
rect 50296 38048 50360 38052
rect 50376 38108 50440 38112
rect 50376 38052 50380 38108
rect 50380 38052 50436 38108
rect 50436 38052 50440 38108
rect 50376 38048 50440 38052
rect 50456 38108 50520 38112
rect 50456 38052 50460 38108
rect 50460 38052 50516 38108
rect 50516 38052 50520 38108
rect 50456 38048 50520 38052
rect 50536 38108 50600 38112
rect 50536 38052 50540 38108
rect 50540 38052 50596 38108
rect 50596 38052 50600 38108
rect 50536 38048 50600 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 50296 37020 50360 37024
rect 50296 36964 50300 37020
rect 50300 36964 50356 37020
rect 50356 36964 50360 37020
rect 50296 36960 50360 36964
rect 50376 37020 50440 37024
rect 50376 36964 50380 37020
rect 50380 36964 50436 37020
rect 50436 36964 50440 37020
rect 50376 36960 50440 36964
rect 50456 37020 50520 37024
rect 50456 36964 50460 37020
rect 50460 36964 50516 37020
rect 50516 36964 50520 37020
rect 50456 36960 50520 36964
rect 50536 37020 50600 37024
rect 50536 36964 50540 37020
rect 50540 36964 50596 37020
rect 50596 36964 50600 37020
rect 50536 36960 50600 36964
rect 41460 36484 41524 36548
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 30420 36000 30484 36004
rect 30420 35944 30470 36000
rect 30470 35944 30484 36000
rect 30420 35940 30484 35944
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 50296 35932 50360 35936
rect 50296 35876 50300 35932
rect 50300 35876 50356 35932
rect 50356 35876 50360 35932
rect 50296 35872 50360 35876
rect 50376 35932 50440 35936
rect 50376 35876 50380 35932
rect 50380 35876 50436 35932
rect 50436 35876 50440 35932
rect 50376 35872 50440 35876
rect 50456 35932 50520 35936
rect 50456 35876 50460 35932
rect 50460 35876 50516 35932
rect 50516 35876 50520 35932
rect 50456 35872 50520 35876
rect 50536 35932 50600 35936
rect 50536 35876 50540 35932
rect 50540 35876 50596 35932
rect 50596 35876 50600 35932
rect 50536 35872 50600 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 50296 34844 50360 34848
rect 50296 34788 50300 34844
rect 50300 34788 50356 34844
rect 50356 34788 50360 34844
rect 50296 34784 50360 34788
rect 50376 34844 50440 34848
rect 50376 34788 50380 34844
rect 50380 34788 50436 34844
rect 50436 34788 50440 34844
rect 50376 34784 50440 34788
rect 50456 34844 50520 34848
rect 50456 34788 50460 34844
rect 50460 34788 50516 34844
rect 50516 34788 50520 34844
rect 50456 34784 50520 34788
rect 50536 34844 50600 34848
rect 50536 34788 50540 34844
rect 50540 34788 50596 34844
rect 50596 34788 50600 34844
rect 50536 34784 50600 34788
rect 30788 34640 30852 34644
rect 30788 34584 30802 34640
rect 30802 34584 30852 34640
rect 30788 34580 30852 34584
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 50296 33756 50360 33760
rect 50296 33700 50300 33756
rect 50300 33700 50356 33756
rect 50356 33700 50360 33756
rect 50296 33696 50360 33700
rect 50376 33756 50440 33760
rect 50376 33700 50380 33756
rect 50380 33700 50436 33756
rect 50436 33700 50440 33756
rect 50376 33696 50440 33700
rect 50456 33756 50520 33760
rect 50456 33700 50460 33756
rect 50460 33700 50516 33756
rect 50516 33700 50520 33756
rect 50456 33696 50520 33700
rect 50536 33756 50600 33760
rect 50536 33700 50540 33756
rect 50540 33700 50596 33756
rect 50596 33700 50600 33756
rect 50536 33696 50600 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 50296 32668 50360 32672
rect 50296 32612 50300 32668
rect 50300 32612 50356 32668
rect 50356 32612 50360 32668
rect 50296 32608 50360 32612
rect 50376 32668 50440 32672
rect 50376 32612 50380 32668
rect 50380 32612 50436 32668
rect 50436 32612 50440 32668
rect 50376 32608 50440 32612
rect 50456 32668 50520 32672
rect 50456 32612 50460 32668
rect 50460 32612 50516 32668
rect 50516 32612 50520 32668
rect 50456 32608 50520 32612
rect 50536 32668 50600 32672
rect 50536 32612 50540 32668
rect 50540 32612 50596 32668
rect 50596 32612 50600 32668
rect 50536 32608 50600 32612
rect 39252 32404 39316 32468
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 29500 32056 29564 32060
rect 29500 32000 29550 32056
rect 29550 32000 29564 32056
rect 29500 31996 29564 32000
rect 37780 31724 37844 31788
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 50296 31580 50360 31584
rect 50296 31524 50300 31580
rect 50300 31524 50356 31580
rect 50356 31524 50360 31580
rect 50296 31520 50360 31524
rect 50376 31580 50440 31584
rect 50376 31524 50380 31580
rect 50380 31524 50436 31580
rect 50436 31524 50440 31580
rect 50376 31520 50440 31524
rect 50456 31580 50520 31584
rect 50456 31524 50460 31580
rect 50460 31524 50516 31580
rect 50516 31524 50520 31580
rect 50456 31520 50520 31524
rect 50536 31580 50600 31584
rect 50536 31524 50540 31580
rect 50540 31524 50596 31580
rect 50596 31524 50600 31580
rect 50536 31520 50600 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 50296 30492 50360 30496
rect 50296 30436 50300 30492
rect 50300 30436 50356 30492
rect 50356 30436 50360 30492
rect 50296 30432 50360 30436
rect 50376 30492 50440 30496
rect 50376 30436 50380 30492
rect 50380 30436 50436 30492
rect 50436 30436 50440 30492
rect 50376 30432 50440 30436
rect 50456 30492 50520 30496
rect 50456 30436 50460 30492
rect 50460 30436 50516 30492
rect 50516 30436 50520 30492
rect 50456 30432 50520 30436
rect 50536 30492 50600 30496
rect 50536 30436 50540 30492
rect 50540 30436 50596 30492
rect 50596 30436 50600 30492
rect 50536 30432 50600 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 46244 29684 46308 29748
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 50296 29404 50360 29408
rect 50296 29348 50300 29404
rect 50300 29348 50356 29404
rect 50356 29348 50360 29404
rect 50296 29344 50360 29348
rect 50376 29404 50440 29408
rect 50376 29348 50380 29404
rect 50380 29348 50436 29404
rect 50436 29348 50440 29404
rect 50376 29344 50440 29348
rect 50456 29404 50520 29408
rect 50456 29348 50460 29404
rect 50460 29348 50516 29404
rect 50516 29348 50520 29404
rect 50456 29344 50520 29348
rect 50536 29404 50600 29408
rect 50536 29348 50540 29404
rect 50540 29348 50596 29404
rect 50596 29348 50600 29404
rect 50536 29344 50600 29348
rect 44772 29004 44836 29068
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 50296 28316 50360 28320
rect 50296 28260 50300 28316
rect 50300 28260 50356 28316
rect 50356 28260 50360 28316
rect 50296 28256 50360 28260
rect 50376 28316 50440 28320
rect 50376 28260 50380 28316
rect 50380 28260 50436 28316
rect 50436 28260 50440 28316
rect 50376 28256 50440 28260
rect 50456 28316 50520 28320
rect 50456 28260 50460 28316
rect 50460 28260 50516 28316
rect 50516 28260 50520 28316
rect 50456 28256 50520 28260
rect 50536 28316 50600 28320
rect 50536 28260 50540 28316
rect 50540 28260 50596 28316
rect 50596 28260 50600 28316
rect 50536 28256 50600 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 50296 27228 50360 27232
rect 50296 27172 50300 27228
rect 50300 27172 50356 27228
rect 50356 27172 50360 27228
rect 50296 27168 50360 27172
rect 50376 27228 50440 27232
rect 50376 27172 50380 27228
rect 50380 27172 50436 27228
rect 50436 27172 50440 27228
rect 50376 27168 50440 27172
rect 50456 27228 50520 27232
rect 50456 27172 50460 27228
rect 50460 27172 50516 27228
rect 50516 27172 50520 27228
rect 50456 27168 50520 27172
rect 50536 27228 50600 27232
rect 50536 27172 50540 27228
rect 50540 27172 50596 27228
rect 50596 27172 50600 27228
rect 50536 27168 50600 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 33732 26344 33796 26348
rect 33732 26288 33782 26344
rect 33782 26288 33796 26344
rect 33732 26284 33796 26288
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 50296 26140 50360 26144
rect 50296 26084 50300 26140
rect 50300 26084 50356 26140
rect 50356 26084 50360 26140
rect 50296 26080 50360 26084
rect 50376 26140 50440 26144
rect 50376 26084 50380 26140
rect 50380 26084 50436 26140
rect 50436 26084 50440 26140
rect 50376 26080 50440 26084
rect 50456 26140 50520 26144
rect 50456 26084 50460 26140
rect 50460 26084 50516 26140
rect 50516 26084 50520 26140
rect 50456 26080 50520 26084
rect 50536 26140 50600 26144
rect 50536 26084 50540 26140
rect 50540 26084 50596 26140
rect 50596 26084 50600 26140
rect 50536 26080 50600 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 50296 25052 50360 25056
rect 50296 24996 50300 25052
rect 50300 24996 50356 25052
rect 50356 24996 50360 25052
rect 50296 24992 50360 24996
rect 50376 25052 50440 25056
rect 50376 24996 50380 25052
rect 50380 24996 50436 25052
rect 50436 24996 50440 25052
rect 50376 24992 50440 24996
rect 50456 25052 50520 25056
rect 50456 24996 50460 25052
rect 50460 24996 50516 25052
rect 50516 24996 50520 25052
rect 50456 24992 50520 24996
rect 50536 25052 50600 25056
rect 50536 24996 50540 25052
rect 50540 24996 50596 25052
rect 50596 24996 50600 25052
rect 50536 24992 50600 24996
rect 43484 24984 43548 24988
rect 43484 24928 43498 24984
rect 43498 24928 43548 24984
rect 43484 24924 43548 24928
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 50296 23964 50360 23968
rect 50296 23908 50300 23964
rect 50300 23908 50356 23964
rect 50356 23908 50360 23964
rect 50296 23904 50360 23908
rect 50376 23964 50440 23968
rect 50376 23908 50380 23964
rect 50380 23908 50436 23964
rect 50436 23908 50440 23964
rect 50376 23904 50440 23908
rect 50456 23964 50520 23968
rect 50456 23908 50460 23964
rect 50460 23908 50516 23964
rect 50516 23908 50520 23964
rect 50456 23904 50520 23908
rect 50536 23964 50600 23968
rect 50536 23908 50540 23964
rect 50540 23908 50596 23964
rect 50596 23908 50600 23964
rect 50536 23904 50600 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 50296 22876 50360 22880
rect 50296 22820 50300 22876
rect 50300 22820 50356 22876
rect 50356 22820 50360 22876
rect 50296 22816 50360 22820
rect 50376 22876 50440 22880
rect 50376 22820 50380 22876
rect 50380 22820 50436 22876
rect 50436 22820 50440 22876
rect 50376 22816 50440 22820
rect 50456 22876 50520 22880
rect 50456 22820 50460 22876
rect 50460 22820 50516 22876
rect 50516 22820 50520 22876
rect 50456 22816 50520 22820
rect 50536 22876 50600 22880
rect 50536 22820 50540 22876
rect 50540 22820 50596 22876
rect 50596 22820 50600 22876
rect 50536 22816 50600 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 50296 21788 50360 21792
rect 50296 21732 50300 21788
rect 50300 21732 50356 21788
rect 50356 21732 50360 21788
rect 50296 21728 50360 21732
rect 50376 21788 50440 21792
rect 50376 21732 50380 21788
rect 50380 21732 50436 21788
rect 50436 21732 50440 21788
rect 50376 21728 50440 21732
rect 50456 21788 50520 21792
rect 50456 21732 50460 21788
rect 50460 21732 50516 21788
rect 50516 21732 50520 21788
rect 50456 21728 50520 21732
rect 50536 21788 50600 21792
rect 50536 21732 50540 21788
rect 50540 21732 50596 21788
rect 50596 21732 50600 21788
rect 50536 21728 50600 21732
rect 46060 21448 46124 21452
rect 46060 21392 46074 21448
rect 46074 21392 46124 21448
rect 46060 21388 46124 21392
rect 48820 21388 48884 21452
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 48820 20844 48884 20908
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 50296 20700 50360 20704
rect 50296 20644 50300 20700
rect 50300 20644 50356 20700
rect 50356 20644 50360 20700
rect 50296 20640 50360 20644
rect 50376 20700 50440 20704
rect 50376 20644 50380 20700
rect 50380 20644 50436 20700
rect 50436 20644 50440 20700
rect 50376 20640 50440 20644
rect 50456 20700 50520 20704
rect 50456 20644 50460 20700
rect 50460 20644 50516 20700
rect 50516 20644 50520 20700
rect 50456 20640 50520 20644
rect 50536 20700 50600 20704
rect 50536 20644 50540 20700
rect 50540 20644 50596 20700
rect 50596 20644 50600 20700
rect 50536 20640 50600 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 50296 19612 50360 19616
rect 50296 19556 50300 19612
rect 50300 19556 50356 19612
rect 50356 19556 50360 19612
rect 50296 19552 50360 19556
rect 50376 19612 50440 19616
rect 50376 19556 50380 19612
rect 50380 19556 50436 19612
rect 50436 19556 50440 19612
rect 50376 19552 50440 19556
rect 50456 19612 50520 19616
rect 50456 19556 50460 19612
rect 50460 19556 50516 19612
rect 50516 19556 50520 19612
rect 50456 19552 50520 19556
rect 50536 19612 50600 19616
rect 50536 19556 50540 19612
rect 50540 19556 50596 19612
rect 50596 19556 50600 19612
rect 50536 19552 50600 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 50296 18524 50360 18528
rect 50296 18468 50300 18524
rect 50300 18468 50356 18524
rect 50356 18468 50360 18524
rect 50296 18464 50360 18468
rect 50376 18524 50440 18528
rect 50376 18468 50380 18524
rect 50380 18468 50436 18524
rect 50436 18468 50440 18524
rect 50376 18464 50440 18468
rect 50456 18524 50520 18528
rect 50456 18468 50460 18524
rect 50460 18468 50516 18524
rect 50516 18468 50520 18524
rect 50456 18464 50520 18468
rect 50536 18524 50600 18528
rect 50536 18468 50540 18524
rect 50540 18468 50596 18524
rect 50596 18468 50600 18524
rect 50536 18464 50600 18468
rect 31340 18124 31404 18188
rect 43300 17988 43364 18052
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 48452 17912 48516 17916
rect 48452 17856 48466 17912
rect 48466 17856 48516 17912
rect 48452 17852 48516 17856
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 50296 17436 50360 17440
rect 50296 17380 50300 17436
rect 50300 17380 50356 17436
rect 50356 17380 50360 17436
rect 50296 17376 50360 17380
rect 50376 17436 50440 17440
rect 50376 17380 50380 17436
rect 50380 17380 50436 17436
rect 50436 17380 50440 17436
rect 50376 17376 50440 17380
rect 50456 17436 50520 17440
rect 50456 17380 50460 17436
rect 50460 17380 50516 17436
rect 50516 17380 50520 17436
rect 50456 17376 50520 17380
rect 50536 17436 50600 17440
rect 50536 17380 50540 17436
rect 50540 17380 50596 17436
rect 50596 17380 50600 17436
rect 50536 17376 50600 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 50296 16348 50360 16352
rect 50296 16292 50300 16348
rect 50300 16292 50356 16348
rect 50356 16292 50360 16348
rect 50296 16288 50360 16292
rect 50376 16348 50440 16352
rect 50376 16292 50380 16348
rect 50380 16292 50436 16348
rect 50436 16292 50440 16348
rect 50376 16288 50440 16292
rect 50456 16348 50520 16352
rect 50456 16292 50460 16348
rect 50460 16292 50516 16348
rect 50516 16292 50520 16348
rect 50456 16288 50520 16292
rect 50536 16348 50600 16352
rect 50536 16292 50540 16348
rect 50540 16292 50596 16348
rect 50596 16292 50600 16348
rect 50536 16288 50600 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 50296 15260 50360 15264
rect 50296 15204 50300 15260
rect 50300 15204 50356 15260
rect 50356 15204 50360 15260
rect 50296 15200 50360 15204
rect 50376 15260 50440 15264
rect 50376 15204 50380 15260
rect 50380 15204 50436 15260
rect 50436 15204 50440 15260
rect 50376 15200 50440 15204
rect 50456 15260 50520 15264
rect 50456 15204 50460 15260
rect 50460 15204 50516 15260
rect 50516 15204 50520 15260
rect 50456 15200 50520 15204
rect 50536 15260 50600 15264
rect 50536 15204 50540 15260
rect 50540 15204 50596 15260
rect 50596 15204 50600 15260
rect 50536 15200 50600 15204
rect 30420 15056 30484 15060
rect 30420 15000 30434 15056
rect 30434 15000 30484 15056
rect 30420 14996 30484 15000
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 50296 14172 50360 14176
rect 50296 14116 50300 14172
rect 50300 14116 50356 14172
rect 50356 14116 50360 14172
rect 50296 14112 50360 14116
rect 50376 14172 50440 14176
rect 50376 14116 50380 14172
rect 50380 14116 50436 14172
rect 50436 14116 50440 14172
rect 50376 14112 50440 14116
rect 50456 14172 50520 14176
rect 50456 14116 50460 14172
rect 50460 14116 50516 14172
rect 50516 14116 50520 14172
rect 50456 14112 50520 14116
rect 50536 14172 50600 14176
rect 50536 14116 50540 14172
rect 50540 14116 50596 14172
rect 50596 14116 50600 14172
rect 50536 14112 50600 14116
rect 39252 13772 39316 13836
rect 33180 13636 33244 13700
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 50296 13084 50360 13088
rect 50296 13028 50300 13084
rect 50300 13028 50356 13084
rect 50356 13028 50360 13084
rect 50296 13024 50360 13028
rect 50376 13084 50440 13088
rect 50376 13028 50380 13084
rect 50380 13028 50436 13084
rect 50436 13028 50440 13084
rect 50376 13024 50440 13028
rect 50456 13084 50520 13088
rect 50456 13028 50460 13084
rect 50460 13028 50516 13084
rect 50516 13028 50520 13084
rect 50456 13024 50520 13028
rect 50536 13084 50600 13088
rect 50536 13028 50540 13084
rect 50540 13028 50596 13084
rect 50596 13028 50600 13084
rect 50536 13024 50600 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 46060 12276 46124 12340
rect 29500 12004 29564 12068
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 50296 11996 50360 12000
rect 50296 11940 50300 11996
rect 50300 11940 50356 11996
rect 50356 11940 50360 11996
rect 50296 11936 50360 11940
rect 50376 11996 50440 12000
rect 50376 11940 50380 11996
rect 50380 11940 50436 11996
rect 50436 11940 50440 11996
rect 50376 11936 50440 11940
rect 50456 11996 50520 12000
rect 50456 11940 50460 11996
rect 50460 11940 50516 11996
rect 50516 11940 50520 11996
rect 50456 11936 50520 11940
rect 50536 11996 50600 12000
rect 50536 11940 50540 11996
rect 50540 11940 50596 11996
rect 50596 11940 50600 11996
rect 50536 11936 50600 11940
rect 40540 11732 40604 11796
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 50296 10908 50360 10912
rect 50296 10852 50300 10908
rect 50300 10852 50356 10908
rect 50356 10852 50360 10908
rect 50296 10848 50360 10852
rect 50376 10908 50440 10912
rect 50376 10852 50380 10908
rect 50380 10852 50436 10908
rect 50436 10852 50440 10908
rect 50376 10848 50440 10852
rect 50456 10908 50520 10912
rect 50456 10852 50460 10908
rect 50460 10852 50516 10908
rect 50516 10852 50520 10908
rect 50456 10848 50520 10852
rect 50536 10908 50600 10912
rect 50536 10852 50540 10908
rect 50540 10852 50596 10908
rect 50596 10852 50600 10908
rect 50536 10848 50600 10852
rect 43300 10780 43364 10844
rect 43300 10508 43364 10572
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 50296 9820 50360 9824
rect 50296 9764 50300 9820
rect 50300 9764 50356 9820
rect 50356 9764 50360 9820
rect 50296 9760 50360 9764
rect 50376 9820 50440 9824
rect 50376 9764 50380 9820
rect 50380 9764 50436 9820
rect 50436 9764 50440 9820
rect 50376 9760 50440 9764
rect 50456 9820 50520 9824
rect 50456 9764 50460 9820
rect 50460 9764 50516 9820
rect 50516 9764 50520 9820
rect 50456 9760 50520 9764
rect 50536 9820 50600 9824
rect 50536 9764 50540 9820
rect 50540 9764 50596 9820
rect 50596 9764 50600 9820
rect 50536 9760 50600 9764
rect 42564 9692 42628 9756
rect 31156 9556 31220 9620
rect 33180 9556 33244 9620
rect 37780 9556 37844 9620
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 31156 8740 31220 8804
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 50296 8732 50360 8736
rect 50296 8676 50300 8732
rect 50300 8676 50356 8732
rect 50356 8676 50360 8732
rect 50296 8672 50360 8676
rect 50376 8732 50440 8736
rect 50376 8676 50380 8732
rect 50380 8676 50436 8732
rect 50436 8676 50440 8732
rect 50376 8672 50440 8676
rect 50456 8732 50520 8736
rect 50456 8676 50460 8732
rect 50460 8676 50516 8732
rect 50516 8676 50520 8732
rect 50456 8672 50520 8676
rect 50536 8732 50600 8736
rect 50536 8676 50540 8732
rect 50540 8676 50596 8732
rect 50596 8676 50600 8732
rect 50536 8672 50600 8676
rect 43484 8332 43548 8396
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 50296 7644 50360 7648
rect 50296 7588 50300 7644
rect 50300 7588 50356 7644
rect 50356 7588 50360 7644
rect 50296 7584 50360 7588
rect 50376 7644 50440 7648
rect 50376 7588 50380 7644
rect 50380 7588 50436 7644
rect 50436 7588 50440 7644
rect 50376 7584 50440 7588
rect 50456 7644 50520 7648
rect 50456 7588 50460 7644
rect 50460 7588 50516 7644
rect 50516 7588 50520 7644
rect 50456 7584 50520 7588
rect 50536 7644 50600 7648
rect 50536 7588 50540 7644
rect 50540 7588 50596 7644
rect 50596 7588 50600 7644
rect 50536 7584 50600 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 50296 6556 50360 6560
rect 50296 6500 50300 6556
rect 50300 6500 50356 6556
rect 50356 6500 50360 6556
rect 50296 6496 50360 6500
rect 50376 6556 50440 6560
rect 50376 6500 50380 6556
rect 50380 6500 50436 6556
rect 50436 6500 50440 6556
rect 50376 6496 50440 6500
rect 50456 6556 50520 6560
rect 50456 6500 50460 6556
rect 50460 6500 50516 6556
rect 50516 6500 50520 6556
rect 50456 6496 50520 6500
rect 50536 6556 50600 6560
rect 50536 6500 50540 6556
rect 50540 6500 50596 6556
rect 50596 6500 50600 6556
rect 50536 6496 50600 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 43300 5672 43364 5676
rect 43300 5616 43350 5672
rect 43350 5616 43364 5672
rect 43300 5612 43364 5616
rect 47716 5476 47780 5540
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 50296 5468 50360 5472
rect 50296 5412 50300 5468
rect 50300 5412 50356 5468
rect 50356 5412 50360 5468
rect 50296 5408 50360 5412
rect 50376 5468 50440 5472
rect 50376 5412 50380 5468
rect 50380 5412 50436 5468
rect 50436 5412 50440 5468
rect 50376 5408 50440 5412
rect 50456 5468 50520 5472
rect 50456 5412 50460 5468
rect 50460 5412 50516 5468
rect 50516 5412 50520 5468
rect 50456 5408 50520 5412
rect 50536 5468 50600 5472
rect 50536 5412 50540 5468
rect 50540 5412 50596 5468
rect 50596 5412 50600 5468
rect 50536 5408 50600 5412
rect 41276 5400 41340 5404
rect 41276 5344 41290 5400
rect 41290 5344 41340 5400
rect 41276 5340 41340 5344
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 50296 4380 50360 4384
rect 50296 4324 50300 4380
rect 50300 4324 50356 4380
rect 50356 4324 50360 4380
rect 50296 4320 50360 4324
rect 50376 4380 50440 4384
rect 50376 4324 50380 4380
rect 50380 4324 50436 4380
rect 50436 4324 50440 4380
rect 50376 4320 50440 4324
rect 50456 4380 50520 4384
rect 50456 4324 50460 4380
rect 50460 4324 50516 4380
rect 50516 4324 50520 4380
rect 50456 4320 50520 4324
rect 50536 4380 50600 4384
rect 50536 4324 50540 4380
rect 50540 4324 50596 4380
rect 50596 4324 50600 4380
rect 50536 4320 50600 4324
rect 46244 4252 46308 4316
rect 31340 4040 31404 4044
rect 31340 3984 31354 4040
rect 31354 3984 31404 4040
rect 31340 3980 31404 3984
rect 44404 3980 44468 4044
rect 47900 4040 47964 4044
rect 47900 3984 47914 4040
rect 47914 3984 47964 4040
rect 47900 3980 47964 3984
rect 48636 4040 48700 4044
rect 48636 3984 48650 4040
rect 48650 3984 48700 4040
rect 48636 3980 48700 3984
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 33732 3300 33796 3364
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 50296 3292 50360 3296
rect 50296 3236 50300 3292
rect 50300 3236 50356 3292
rect 50356 3236 50360 3292
rect 50296 3232 50360 3236
rect 50376 3292 50440 3296
rect 50376 3236 50380 3292
rect 50380 3236 50436 3292
rect 50436 3236 50440 3292
rect 50376 3232 50440 3236
rect 50456 3292 50520 3296
rect 50456 3236 50460 3292
rect 50460 3236 50516 3292
rect 50516 3236 50520 3292
rect 50456 3232 50520 3236
rect 50536 3292 50600 3296
rect 50536 3236 50540 3292
rect 50540 3236 50596 3292
rect 50596 3236 50600 3292
rect 50536 3232 50600 3236
rect 44772 3164 44836 3228
rect 30788 2892 30852 2956
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 41460 2680 41524 2684
rect 41460 2624 41474 2680
rect 41474 2624 41524 2680
rect 41460 2620 41524 2624
rect 48084 2620 48148 2684
rect 48820 2348 48884 2412
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
rect 50296 2204 50360 2208
rect 50296 2148 50300 2204
rect 50300 2148 50356 2204
rect 50356 2148 50360 2204
rect 50296 2144 50360 2148
rect 50376 2204 50440 2208
rect 50376 2148 50380 2204
rect 50380 2148 50436 2204
rect 50436 2148 50440 2204
rect 50376 2144 50440 2148
rect 50456 2204 50520 2208
rect 50456 2148 50460 2204
rect 50460 2148 50516 2204
rect 50516 2148 50520 2204
rect 50456 2144 50520 2148
rect 50536 2204 50600 2208
rect 50536 2148 50540 2204
rect 50540 2148 50596 2204
rect 50596 2148 50600 2204
rect 50536 2144 50600 2148
<< metal4 >>
rect 4208 57152 4528 57712
rect 4208 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4528 57152
rect 4208 56064 4528 57088
rect 4208 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4528 56064
rect 4208 54976 4528 56000
rect 4208 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4528 54976
rect 4208 53888 4528 54912
rect 4208 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4528 53888
rect 4208 52800 4528 53824
rect 4208 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4528 52800
rect 4208 51712 4528 52736
rect 4208 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4528 51712
rect 4208 50624 4528 51648
rect 4208 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4528 50624
rect 4208 49536 4528 50560
rect 4208 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4528 49536
rect 4208 48448 4528 49472
rect 4208 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4528 48448
rect 4208 47360 4528 48384
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 57696 19888 57712
rect 19568 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19888 57696
rect 19568 56608 19888 57632
rect 19568 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19888 56608
rect 19568 55520 19888 56544
rect 19568 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19888 55520
rect 19568 54432 19888 55456
rect 19568 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19888 54432
rect 19568 53344 19888 54368
rect 19568 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19888 53344
rect 19568 52256 19888 53280
rect 19568 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19888 52256
rect 19568 51168 19888 52192
rect 19568 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19888 51168
rect 19568 50080 19888 51104
rect 19568 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19888 50080
rect 19568 48992 19888 50016
rect 19568 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19888 48992
rect 19568 47904 19888 48928
rect 19568 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19888 47904
rect 19568 46816 19888 47840
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 34928 57152 35248 57712
rect 34928 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35248 57152
rect 34928 56064 35248 57088
rect 50288 57696 50608 57712
rect 50288 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50608 57696
rect 48451 56676 48517 56677
rect 48451 56612 48452 56676
rect 48516 56612 48517 56676
rect 48451 56611 48517 56612
rect 34928 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35248 56064
rect 34928 54976 35248 56000
rect 34928 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35248 54976
rect 34928 53888 35248 54912
rect 34928 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35248 53888
rect 34928 52800 35248 53824
rect 34928 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35248 52800
rect 34928 51712 35248 52736
rect 48083 52732 48149 52733
rect 48083 52668 48084 52732
rect 48148 52668 48149 52732
rect 48083 52667 48149 52668
rect 47899 52596 47965 52597
rect 47899 52532 47900 52596
rect 47964 52532 47965 52596
rect 47899 52531 47965 52532
rect 34928 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35248 51712
rect 34928 50624 35248 51648
rect 47715 51100 47781 51101
rect 47715 51036 47716 51100
rect 47780 51036 47781 51100
rect 47715 51035 47781 51036
rect 34928 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35248 50624
rect 34928 49536 35248 50560
rect 42563 49740 42629 49741
rect 42563 49676 42564 49740
rect 42628 49676 42629 49740
rect 42563 49675 42629 49676
rect 34928 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35248 49536
rect 34928 48448 35248 49472
rect 34928 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35248 48448
rect 34928 47360 35248 48384
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 40539 45524 40605 45525
rect 40539 45460 40540 45524
rect 40604 45460 40605 45524
rect 40539 45459 40605 45460
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 30419 36004 30485 36005
rect 30419 35940 30420 36004
rect 30484 35940 30485 36004
rect 30419 35939 30485 35940
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 29499 32060 29565 32061
rect 29499 31996 29500 32060
rect 29564 31996 29565 32060
rect 29499 31995 29565 31996
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 29502 12069 29562 31995
rect 30422 15061 30482 35939
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 30787 34644 30853 34645
rect 30787 34580 30788 34644
rect 30852 34580 30853 34644
rect 30787 34579 30853 34580
rect 30419 15060 30485 15061
rect 30419 14996 30420 15060
rect 30484 14996 30485 15060
rect 30419 14995 30485 14996
rect 29499 12068 29565 12069
rect 29499 12004 29500 12068
rect 29564 12004 29565 12068
rect 29499 12003 29565 12004
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 30790 2957 30850 34579
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 39251 32468 39317 32469
rect 39251 32404 39252 32468
rect 39316 32404 39317 32468
rect 39251 32403 39317 32404
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 37779 31788 37845 31789
rect 37779 31724 37780 31788
rect 37844 31724 37845 31788
rect 37779 31723 37845 31724
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 33731 26348 33797 26349
rect 33731 26284 33732 26348
rect 33796 26284 33797 26348
rect 33731 26283 33797 26284
rect 31339 18188 31405 18189
rect 31339 18124 31340 18188
rect 31404 18124 31405 18188
rect 31339 18123 31405 18124
rect 31155 9620 31221 9621
rect 31155 9556 31156 9620
rect 31220 9556 31221 9620
rect 31155 9555 31221 9556
rect 31158 8805 31218 9555
rect 31155 8804 31221 8805
rect 31155 8740 31156 8804
rect 31220 8740 31221 8804
rect 31155 8739 31221 8740
rect 31342 4045 31402 18123
rect 33179 13700 33245 13701
rect 33179 13636 33180 13700
rect 33244 13636 33245 13700
rect 33179 13635 33245 13636
rect 33182 9621 33242 13635
rect 33179 9620 33245 9621
rect 33179 9556 33180 9620
rect 33244 9556 33245 9620
rect 33179 9555 33245 9556
rect 31339 4044 31405 4045
rect 31339 3980 31340 4044
rect 31404 3980 31405 4044
rect 31339 3979 31405 3980
rect 33734 3365 33794 26283
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 37782 9621 37842 31723
rect 39254 13837 39314 32403
rect 39251 13836 39317 13837
rect 39251 13772 39252 13836
rect 39316 13772 39317 13836
rect 39251 13771 39317 13772
rect 40542 11797 40602 45459
rect 41275 42940 41341 42941
rect 41275 42876 41276 42940
rect 41340 42876 41341 42940
rect 41275 42875 41341 42876
rect 40539 11796 40605 11797
rect 40539 11732 40540 11796
rect 40604 11732 40605 11796
rect 40539 11731 40605 11732
rect 37779 9620 37845 9621
rect 37779 9556 37780 9620
rect 37844 9556 37845 9620
rect 37779 9555 37845 9556
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 41278 5405 41338 42875
rect 41459 36548 41525 36549
rect 41459 36484 41460 36548
rect 41524 36484 41525 36548
rect 41459 36483 41525 36484
rect 41275 5404 41341 5405
rect 41275 5340 41276 5404
rect 41340 5340 41341 5404
rect 41275 5339 41341 5340
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 33731 3364 33797 3365
rect 33731 3300 33732 3364
rect 33796 3300 33797 3364
rect 33731 3299 33797 3300
rect 30787 2956 30853 2957
rect 30787 2892 30788 2956
rect 30852 2892 30853 2956
rect 30787 2891 30853 2892
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 41462 2685 41522 36483
rect 42566 9757 42626 49675
rect 44403 41444 44469 41445
rect 44403 41380 44404 41444
rect 44468 41380 44469 41444
rect 44403 41379 44469 41380
rect 43483 24988 43549 24989
rect 43483 24924 43484 24988
rect 43548 24924 43549 24988
rect 43483 24923 43549 24924
rect 43299 18052 43365 18053
rect 43299 17988 43300 18052
rect 43364 17988 43365 18052
rect 43299 17987 43365 17988
rect 43302 10845 43362 17987
rect 43299 10844 43365 10845
rect 43299 10780 43300 10844
rect 43364 10780 43365 10844
rect 43299 10779 43365 10780
rect 43299 10572 43365 10573
rect 43299 10508 43300 10572
rect 43364 10508 43365 10572
rect 43299 10507 43365 10508
rect 42563 9756 42629 9757
rect 42563 9692 42564 9756
rect 42628 9692 42629 9756
rect 42563 9691 42629 9692
rect 43302 5677 43362 10507
rect 43486 8397 43546 24923
rect 43483 8396 43549 8397
rect 43483 8332 43484 8396
rect 43548 8332 43549 8396
rect 43483 8331 43549 8332
rect 43299 5676 43365 5677
rect 43299 5612 43300 5676
rect 43364 5612 43365 5676
rect 43299 5611 43365 5612
rect 44406 4045 44466 41379
rect 46243 29748 46309 29749
rect 46243 29684 46244 29748
rect 46308 29684 46309 29748
rect 46243 29683 46309 29684
rect 44771 29068 44837 29069
rect 44771 29004 44772 29068
rect 44836 29004 44837 29068
rect 44771 29003 44837 29004
rect 44403 4044 44469 4045
rect 44403 3980 44404 4044
rect 44468 3980 44469 4044
rect 44403 3979 44469 3980
rect 44774 3229 44834 29003
rect 46059 21452 46125 21453
rect 46059 21388 46060 21452
rect 46124 21388 46125 21452
rect 46059 21387 46125 21388
rect 46062 12341 46122 21387
rect 46059 12340 46125 12341
rect 46059 12276 46060 12340
rect 46124 12276 46125 12340
rect 46059 12275 46125 12276
rect 46246 4317 46306 29683
rect 47718 5541 47778 51035
rect 47715 5540 47781 5541
rect 47715 5476 47716 5540
rect 47780 5476 47781 5540
rect 47715 5475 47781 5476
rect 46243 4316 46309 4317
rect 46243 4252 46244 4316
rect 46308 4252 46309 4316
rect 46243 4251 46309 4252
rect 47902 4045 47962 52531
rect 47899 4044 47965 4045
rect 47899 3980 47900 4044
rect 47964 3980 47965 4044
rect 47899 3979 47965 3980
rect 44771 3228 44837 3229
rect 44771 3164 44772 3228
rect 44836 3164 44837 3228
rect 44771 3163 44837 3164
rect 48086 2685 48146 52667
rect 48454 17917 48514 56611
rect 50288 56608 50608 57632
rect 50288 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50608 56608
rect 50288 55520 50608 56544
rect 50288 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50608 55520
rect 50288 54432 50608 55456
rect 50288 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50608 54432
rect 50288 53344 50608 54368
rect 50288 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50608 53344
rect 50288 52256 50608 53280
rect 50288 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50608 52256
rect 50288 51168 50608 52192
rect 50288 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50608 51168
rect 50288 50080 50608 51104
rect 50288 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50608 50080
rect 50288 48992 50608 50016
rect 50288 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50608 48992
rect 50288 47904 50608 48928
rect 50288 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50608 47904
rect 50288 46816 50608 47840
rect 50288 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50608 46816
rect 50288 45728 50608 46752
rect 50288 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50608 45728
rect 50288 44640 50608 45664
rect 50288 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50608 44640
rect 48635 44300 48701 44301
rect 48635 44236 48636 44300
rect 48700 44236 48701 44300
rect 48635 44235 48701 44236
rect 48451 17916 48517 17917
rect 48451 17852 48452 17916
rect 48516 17852 48517 17916
rect 48451 17851 48517 17852
rect 48638 4045 48698 44235
rect 50288 43552 50608 44576
rect 50288 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50608 43552
rect 50288 42464 50608 43488
rect 50288 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50608 42464
rect 50288 41376 50608 42400
rect 50288 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50608 41376
rect 50288 40288 50608 41312
rect 50288 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50608 40288
rect 50288 39200 50608 40224
rect 50288 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50608 39200
rect 50288 38112 50608 39136
rect 50288 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50608 38112
rect 50288 37024 50608 38048
rect 50288 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50608 37024
rect 50288 35936 50608 36960
rect 50288 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50608 35936
rect 50288 34848 50608 35872
rect 50288 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50608 34848
rect 50288 33760 50608 34784
rect 50288 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50608 33760
rect 50288 32672 50608 33696
rect 50288 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50608 32672
rect 50288 31584 50608 32608
rect 50288 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50608 31584
rect 50288 30496 50608 31520
rect 50288 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50608 30496
rect 50288 29408 50608 30432
rect 50288 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50608 29408
rect 50288 28320 50608 29344
rect 50288 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50608 28320
rect 50288 27232 50608 28256
rect 50288 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50608 27232
rect 50288 26144 50608 27168
rect 50288 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50608 26144
rect 50288 25056 50608 26080
rect 50288 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50608 25056
rect 50288 23968 50608 24992
rect 50288 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50608 23968
rect 50288 22880 50608 23904
rect 50288 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50608 22880
rect 50288 21792 50608 22816
rect 50288 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50608 21792
rect 48819 21452 48885 21453
rect 48819 21388 48820 21452
rect 48884 21388 48885 21452
rect 48819 21387 48885 21388
rect 48822 20909 48882 21387
rect 48819 20908 48885 20909
rect 48819 20844 48820 20908
rect 48884 20844 48885 20908
rect 48819 20843 48885 20844
rect 48635 4044 48701 4045
rect 48635 3980 48636 4044
rect 48700 3980 48701 4044
rect 48635 3979 48701 3980
rect 41459 2684 41525 2685
rect 41459 2620 41460 2684
rect 41524 2620 41525 2684
rect 41459 2619 41525 2620
rect 48083 2684 48149 2685
rect 48083 2620 48084 2684
rect 48148 2620 48149 2684
rect 48083 2619 48149 2620
rect 48822 2413 48882 20843
rect 50288 20704 50608 21728
rect 50288 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50608 20704
rect 50288 19616 50608 20640
rect 50288 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50608 19616
rect 50288 18528 50608 19552
rect 50288 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50608 18528
rect 50288 17440 50608 18464
rect 50288 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50608 17440
rect 50288 16352 50608 17376
rect 50288 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50608 16352
rect 50288 15264 50608 16288
rect 50288 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50608 15264
rect 50288 14176 50608 15200
rect 50288 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50608 14176
rect 50288 13088 50608 14112
rect 50288 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50608 13088
rect 50288 12000 50608 13024
rect 50288 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50608 12000
rect 50288 10912 50608 11936
rect 50288 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50608 10912
rect 50288 9824 50608 10848
rect 50288 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50608 9824
rect 50288 8736 50608 9760
rect 50288 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50608 8736
rect 50288 7648 50608 8672
rect 50288 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50608 7648
rect 50288 6560 50608 7584
rect 50288 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50608 6560
rect 50288 5472 50608 6496
rect 50288 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50608 5472
rect 50288 4384 50608 5408
rect 50288 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50608 4384
rect 50288 3296 50608 4320
rect 50288 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50608 3296
rect 48819 2412 48885 2413
rect 48819 2348 48820 2412
rect 48884 2348 48885 2412
rect 48819 2347 48885 2348
rect 50288 2208 50608 3232
rect 50288 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50608 2208
rect 50288 2128 50608 2144
use sky130_fd_sc_hd__diode_2  ANTENNA_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 28060 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1676037725
transform 1 0 33396 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1676037725
transform 1 0 40940 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1676037725
transform 1 0 51244 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1676037725
transform 1 0 49864 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1676037725
transform 1 0 21804 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1676037725
transform 1 0 27232 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1676037725
transform 1 0 33120 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1676037725
transform 1 0 22724 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1676037725
transform 1 0 41124 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1676037725
transform 1 0 49036 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1676037725
transform 1 0 34960 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1676037725
transform 1 0 30544 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1676037725
transform 1 0 27324 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1676037725
transform 1 0 28060 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1676037725
transform 1 0 2944 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1676037725
transform 1 0 2300 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1676037725
transform 1 0 41768 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1676037725
transform 1 0 23092 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1676037725
transform 1 0 24932 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1676037725
transform 1 0 40112 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp 1676037725
transform 1 0 35052 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp 1676037725
transform 1 0 2300 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp 1676037725
transform 1 0 2300 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp 1676037725
transform 1 0 24840 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp 1676037725
transform 1 0 47288 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp 1676037725
transform 1 0 22172 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1676037725
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4876 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49
timestamp 1676037725
transform 1 0 5612 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61
timestamp 1676037725
transform 1 0 6716 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66
timestamp 1676037725
transform 1 0 7176 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_74
timestamp 1676037725
transform 1 0 7912 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1676037725
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_85
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89
timestamp 1676037725
transform 1 0 9292 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_94
timestamp 1676037725
transform 1 0 9752 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_102
timestamp 1676037725
transform 1 0 10488 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1676037725
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_113
timestamp 1676037725
transform 1 0 11500 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117
timestamp 1676037725
transform 1 0 11868 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_122
timestamp 1676037725
transform 1 0 12328 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_130
timestamp 1676037725
transform 1 0 13064 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1676037725
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_146
timestamp 1676037725
transform 1 0 14536 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_156
timestamp 1676037725
transform 1 0 15456 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1676037725
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1676037725
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_174
timestamp 1676037725
transform 1 0 17112 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_184
timestamp 1676037725
transform 1 0 18032 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1676037725
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1676037725
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_202
timestamp 1676037725
transform 1 0 19688 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_212
timestamp 1676037725
transform 1 0 20608 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1676037725
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1676037725
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_230
timestamp 1676037725
transform 1 0 22264 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_240
timestamp 1676037725
transform 1 0 23184 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_250
timestamp 1676037725
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_256
timestamp 1676037725
transform 1 0 24656 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_260
timestamp 1676037725
transform 1 0 25024 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_268
timestamp 1676037725
transform 1 0 25760 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_278
timestamp 1676037725
transform 1 0 26680 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1676037725
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_289
timestamp 1676037725
transform 1 0 27692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_296
timestamp 1676037725
transform 1 0 28336 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_306
timestamp 1676037725
transform 1 0 29256 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_309 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 29532 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_315
timestamp 1676037725
transform 1 0 30084 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_322
timestamp 1676037725
transform 1 0 30728 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_332
timestamp 1676037725
transform 1 0 31648 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1676037725
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_345
timestamp 1676037725
transform 1 0 32844 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_355
timestamp 1676037725
transform 1 0 33764 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_363
timestamp 1676037725
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_365
timestamp 1676037725
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_373
timestamp 1676037725
transform 1 0 35420 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_383
timestamp 1676037725
transform 1 0 36340 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_391
timestamp 1676037725
transform 1 0 37076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_393
timestamp 1676037725
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_401
timestamp 1676037725
transform 1 0 37996 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_411
timestamp 1676037725
transform 1 0 38916 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_419
timestamp 1676037725
transform 1 0 39652 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_421
timestamp 1676037725
transform 1 0 39836 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_429
timestamp 1676037725
transform 1 0 40572 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_433
timestamp 1676037725
transform 1 0 40940 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_440
timestamp 1676037725
transform 1 0 41584 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_449
timestamp 1676037725
transform 1 0 42412 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_457
timestamp 1676037725
transform 1 0 43148 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_465
timestamp 1676037725
transform 1 0 43884 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_473 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 44620 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_477
timestamp 1676037725
transform 1 0 44988 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_483
timestamp 1676037725
transform 1 0 45540 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_491
timestamp 1676037725
transform 1 0 46276 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_499
timestamp 1676037725
transform 1 0 47012 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_503
timestamp 1676037725
transform 1 0 47380 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_505
timestamp 1676037725
transform 1 0 47564 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_518
timestamp 1676037725
transform 1 0 48760 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_528
timestamp 1676037725
transform 1 0 49680 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_533
timestamp 1676037725
transform 1 0 50140 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_541
timestamp 1676037725
transform 1 0 50876 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_551
timestamp 1676037725
transform 1 0 51796 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_559
timestamp 1676037725
transform 1 0 52532 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_561
timestamp 1676037725
transform 1 0 52716 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_567
timestamp 1676037725
transform 1 0 53268 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_581
timestamp 1676037725
transform 1 0 54556 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_587
timestamp 1676037725
transform 1 0 55108 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_589
timestamp 1676037725
transform 1 0 55292 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_595
timestamp 1676037725
transform 1 0 55844 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_603
timestamp 1676037725
transform 1 0 56580 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_607
timestamp 1676037725
transform 1 0 56948 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_614
timestamp 1676037725
transform 1 0 57592 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_617
timestamp 1676037725
transform 1 0 57868 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_623
timestamp 1676037725
transform 1 0 58420 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1676037725
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1676037725
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_39
timestamp 1676037725
transform 1 0 4692 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_47
timestamp 1676037725
transform 1 0 5428 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1676037725
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_65
timestamp 1676037725
transform 1 0 7084 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_73
timestamp 1676037725
transform 1 0 7820 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_81
timestamp 1676037725
transform 1 0 8556 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_89
timestamp 1676037725
transform 1 0 9292 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_99
timestamp 1676037725
transform 1 0 10212 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_105
timestamp 1676037725
transform 1 0 10764 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1676037725
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_121
timestamp 1676037725
transform 1 0 12236 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_127
timestamp 1676037725
transform 1 0 12788 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_132
timestamp 1676037725
transform 1 0 13248 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_140
timestamp 1676037725
transform 1 0 13984 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_148
timestamp 1676037725
transform 1 0 14720 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_156
timestamp 1676037725
transform 1 0 15456 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1676037725
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_174
timestamp 1676037725
transform 1 0 17112 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_184
timestamp 1676037725
transform 1 0 18032 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_194
timestamp 1676037725
transform 1 0 18952 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_204
timestamp 1676037725
transform 1 0 19872 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_215
timestamp 1676037725
transform 1 0 20884 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1676037725
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_225
timestamp 1676037725
transform 1 0 21804 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_231
timestamp 1676037725
transform 1 0 22356 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_239
timestamp 1676037725
transform 1 0 23092 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_249
timestamp 1676037725
transform 1 0 24012 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_269
timestamp 1676037725
transform 1 0 25852 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_278
timestamp 1676037725
transform 1 0 26680 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_281
timestamp 1676037725
transform 1 0 26956 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_289
timestamp 1676037725
transform 1 0 27692 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_297
timestamp 1676037725
transform 1 0 28428 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_302
timestamp 1676037725
transform 1 0 28888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_309
timestamp 1676037725
transform 1 0 29532 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_319
timestamp 1676037725
transform 1 0 30452 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1676037725
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1676037725
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_337
timestamp 1676037725
transform 1 0 32108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_345
timestamp 1676037725
transform 1 0 32844 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_355
timestamp 1676037725
transform 1 0 33764 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_365
timestamp 1676037725
transform 1 0 34684 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_375
timestamp 1676037725
transform 1 0 35604 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 1676037725
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1676037725
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_393
timestamp 1676037725
transform 1 0 37260 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_401
timestamp 1676037725
transform 1 0 37996 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_413
timestamp 1676037725
transform 1 0 39100 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_423
timestamp 1676037725
transform 1 0 40020 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_431
timestamp 1676037725
transform 1 0 40756 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_439
timestamp 1676037725
transform 1 0 41492 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_446
timestamp 1676037725
transform 1 0 42136 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_449
timestamp 1676037725
transform 1 0 42412 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_459
timestamp 1676037725
transform 1 0 43332 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_467
timestamp 1676037725
transform 1 0 44068 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_475
timestamp 1676037725
transform 1 0 44804 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_483
timestamp 1676037725
transform 1 0 45540 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_491
timestamp 1676037725
transform 1 0 46276 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_499
timestamp 1676037725
transform 1 0 47012 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 1676037725
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_505
timestamp 1676037725
transform 1 0 47564 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_517
timestamp 1676037725
transform 1 0 48668 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_527
timestamp 1676037725
transform 1 0 49588 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_535
timestamp 1676037725
transform 1 0 50324 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_543
timestamp 1676037725
transform 1 0 51060 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_551
timestamp 1676037725
transform 1 0 51796 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_559
timestamp 1676037725
transform 1 0 52532 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_561
timestamp 1676037725
transform 1 0 52716 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_567
timestamp 1676037725
transform 1 0 53268 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_575
timestamp 1676037725
transform 1 0 54004 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_583
timestamp 1676037725
transform 1 0 54740 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_591
timestamp 1676037725
transform 1 0 55476 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_599
timestamp 1676037725
transform 1 0 56212 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_608
timestamp 1676037725
transform 1 0 57040 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_617
timestamp 1676037725
transform 1 0 57868 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_623
timestamp 1676037725
transform 1 0 58420 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1676037725
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1676037725
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1676037725
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_53
timestamp 1676037725
transform 1 0 5980 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_61
timestamp 1676037725
transform 1 0 6716 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_66
timestamp 1676037725
transform 1 0 7176 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_74
timestamp 1676037725
transform 1 0 7912 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp 1676037725
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_100
timestamp 1676037725
transform 1 0 10304 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_110
timestamp 1676037725
transform 1 0 11224 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_120
timestamp 1676037725
transform 1 0 12144 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_130
timestamp 1676037725
transform 1 0 13064 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1676037725
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_147
timestamp 1676037725
transform 1 0 14628 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_151
timestamp 1676037725
transform 1 0 14996 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_156
timestamp 1676037725
transform 1 0 15456 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_164
timestamp 1676037725
transform 1 0 16192 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_174
timestamp 1676037725
transform 1 0 17112 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_184
timestamp 1676037725
transform 1 0 18032 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp 1676037725
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1676037725
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_205
timestamp 1676037725
transform 1 0 19964 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_216
timestamp 1676037725
transform 1 0 20976 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_224
timestamp 1676037725
transform 1 0 21712 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_232
timestamp 1676037725
transform 1 0 22448 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_243
timestamp 1676037725
transform 1 0 23460 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_250
timestamp 1676037725
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_253
timestamp 1676037725
transform 1 0 24380 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_265
timestamp 1676037725
transform 1 0 25484 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_285
timestamp 1676037725
transform 1 0 27324 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_293
timestamp 1676037725
transform 1 0 28060 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_298
timestamp 1676037725
transform 1 0 28520 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_306
timestamp 1676037725
transform 1 0 29256 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_309
timestamp 1676037725
transform 1 0 29532 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_321
timestamp 1676037725
transform 1 0 30636 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_332
timestamp 1676037725
transform 1 0 31648 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_342
timestamp 1676037725
transform 1 0 32568 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_352
timestamp 1676037725
transform 1 0 33488 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_362
timestamp 1676037725
transform 1 0 34408 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_365
timestamp 1676037725
transform 1 0 34684 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_373
timestamp 1676037725
transform 1 0 35420 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_381
timestamp 1676037725
transform 1 0 36156 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_398
timestamp 1676037725
transform 1 0 37720 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_406
timestamp 1676037725
transform 1 0 38456 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_418
timestamp 1676037725
transform 1 0 39560 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_421
timestamp 1676037725
transform 1 0 39836 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_427
timestamp 1676037725
transform 1 0 40388 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_435
timestamp 1676037725
transform 1 0 41124 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_457
timestamp 1676037725
transform 1 0 43148 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_470
timestamp 1676037725
transform 1 0 44344 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_477
timestamp 1676037725
transform 1 0 44988 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_483
timestamp 1676037725
transform 1 0 45540 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_489
timestamp 1676037725
transform 1 0 46092 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_494
timestamp 1676037725
transform 1 0 46552 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_507
timestamp 1676037725
transform 1 0 47748 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_525
timestamp 1676037725
transform 1 0 49404 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_531
timestamp 1676037725
transform 1 0 49956 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_533
timestamp 1676037725
transform 1 0 50140 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_539
timestamp 1676037725
transform 1 0 50692 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_547
timestamp 1676037725
transform 1 0 51428 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_555
timestamp 1676037725
transform 1 0 52164 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_563
timestamp 1676037725
transform 1 0 52900 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_571
timestamp 1676037725
transform 1 0 53636 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_579
timestamp 1676037725
transform 1 0 54372 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_586
timestamp 1676037725
transform 1 0 55016 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_589
timestamp 1676037725
transform 1 0 55292 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_608
timestamp 1676037725
transform 1 0 57040 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_618
timestamp 1676037725
transform 1 0 57960 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_624
timestamp 1676037725
transform 1 0 58512 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1676037725
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1676037725
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1676037725
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1676037725
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1676037725
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_69
timestamp 1676037725
transform 1 0 7452 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_81
timestamp 1676037725
transform 1 0 8556 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_85
timestamp 1676037725
transform 1 0 8924 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_90
timestamp 1676037725
transform 1 0 9384 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_101
timestamp 1676037725
transform 1 0 10396 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_105
timestamp 1676037725
transform 1 0 10764 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 1676037725
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_113
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_121
timestamp 1676037725
transform 1 0 12236 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_129
timestamp 1676037725
transform 1 0 12972 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_141
timestamp 1676037725
transform 1 0 14076 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_153
timestamp 1676037725
transform 1 0 15180 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_157
timestamp 1676037725
transform 1 0 15548 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_162
timestamp 1676037725
transform 1 0 16008 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_175
timestamp 1676037725
transform 1 0 17204 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_182
timestamp 1676037725
transform 1 0 17848 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_191
timestamp 1676037725
transform 1 0 18676 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_195
timestamp 1676037725
transform 1 0 19044 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_202
timestamp 1676037725
transform 1 0 19688 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_213
timestamp 1676037725
transform 1 0 20700 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_221
timestamp 1676037725
transform 1 0 21436 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_225
timestamp 1676037725
transform 1 0 21804 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_231
timestamp 1676037725
transform 1 0 22356 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_238
timestamp 1676037725
transform 1 0 23000 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_248
timestamp 1676037725
transform 1 0 23920 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_258
timestamp 1676037725
transform 1 0 24840 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_271
timestamp 1676037725
transform 1 0 26036 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_278
timestamp 1676037725
transform 1 0 26680 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_281
timestamp 1676037725
transform 1 0 26956 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_292
timestamp 1676037725
transform 1 0 27968 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_301
timestamp 1676037725
transform 1 0 28796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_321
timestamp 1676037725
transform 1 0 30636 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_334
timestamp 1676037725
transform 1 0 31832 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_337
timestamp 1676037725
transform 1 0 32108 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_358
timestamp 1676037725
transform 1 0 34040 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_364
timestamp 1676037725
transform 1 0 34592 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_371
timestamp 1676037725
transform 1 0 35236 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_381
timestamp 1676037725
transform 1 0 36156 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_389
timestamp 1676037725
transform 1 0 36892 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_393
timestamp 1676037725
transform 1 0 37260 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_401
timestamp 1676037725
transform 1 0 37996 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_411
timestamp 1676037725
transform 1 0 38916 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_421
timestamp 1676037725
transform 1 0 39836 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_429
timestamp 1676037725
transform 1 0 40572 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_437
timestamp 1676037725
transform 1 0 41308 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_445
timestamp 1676037725
transform 1 0 42044 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_449
timestamp 1676037725
transform 1 0 42412 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_455
timestamp 1676037725
transform 1 0 42964 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_463
timestamp 1676037725
transform 1 0 43700 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_471
timestamp 1676037725
transform 1 0 44436 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_479
timestamp 1676037725
transform 1 0 45172 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_487
timestamp 1676037725
transform 1 0 45908 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_495
timestamp 1676037725
transform 1 0 46644 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1676037725
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_505
timestamp 1676037725
transform 1 0 47564 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_524
timestamp 1676037725
transform 1 0 49312 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_532
timestamp 1676037725
transform 1 0 50048 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_540
timestamp 1676037725
transform 1 0 50784 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_548
timestamp 1676037725
transform 1 0 51520 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_556
timestamp 1676037725
transform 1 0 52256 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_561
timestamp 1676037725
transform 1 0 52716 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_567
timestamp 1676037725
transform 1 0 53268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_579
timestamp 1676037725
transform 1 0 54372 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_584
timestamp 1676037725
transform 1 0 54832 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_592
timestamp 1676037725
transform 1 0 55568 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_605
timestamp 1676037725
transform 1 0 56764 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_614
timestamp 1676037725
transform 1 0 57592 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_617
timestamp 1676037725
transform 1 0 57868 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_623
timestamp 1676037725
transform 1 0 58420 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_11
timestamp 1676037725
transform 1 0 2116 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_23
timestamp 1676037725
transform 1 0 3220 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1676037725
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1676037725
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1676037725
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1676037725
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1676037725
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1676037725
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_97
timestamp 1676037725
transform 1 0 10028 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_105
timestamp 1676037725
transform 1 0 10764 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_117
timestamp 1676037725
transform 1 0 11868 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_129
timestamp 1676037725
transform 1 0 12972 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_137
timestamp 1676037725
transform 1 0 13708 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1676037725
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1676037725
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_183
timestamp 1676037725
transform 1 0 17940 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_190
timestamp 1676037725
transform 1 0 18584 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_197
timestamp 1676037725
transform 1 0 19228 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_205
timestamp 1676037725
transform 1 0 19964 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_215
timestamp 1676037725
transform 1 0 20884 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_223
timestamp 1676037725
transform 1 0 21620 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_227
timestamp 1676037725
transform 1 0 21988 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_238
timestamp 1676037725
transform 1 0 23000 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_248
timestamp 1676037725
transform 1 0 23920 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_253
timestamp 1676037725
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_271
timestamp 1676037725
transform 1 0 26036 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_278
timestamp 1676037725
transform 1 0 26680 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_285
timestamp 1676037725
transform 1 0 27324 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_297
timestamp 1676037725
transform 1 0 28428 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_304
timestamp 1676037725
transform 1 0 29072 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1676037725
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_321
timestamp 1676037725
transform 1 0 30636 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_328
timestamp 1676037725
transform 1 0 31280 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_340
timestamp 1676037725
transform 1 0 32384 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_348
timestamp 1676037725
transform 1 0 33120 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_356
timestamp 1676037725
transform 1 0 33856 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_365
timestamp 1676037725
transform 1 0 34684 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_373
timestamp 1676037725
transform 1 0 35420 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_382
timestamp 1676037725
transform 1 0 36248 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_395
timestamp 1676037725
transform 1 0 37444 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_405
timestamp 1676037725
transform 1 0 38364 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_418
timestamp 1676037725
transform 1 0 39560 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_421
timestamp 1676037725
transform 1 0 39836 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_432
timestamp 1676037725
transform 1 0 40848 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_440
timestamp 1676037725
transform 1 0 41584 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_448
timestamp 1676037725
transform 1 0 42320 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_456
timestamp 1676037725
transform 1 0 43056 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_463
timestamp 1676037725
transform 1 0 43700 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1676037725
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_477
timestamp 1676037725
transform 1 0 44988 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_489
timestamp 1676037725
transform 1 0 46092 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_497
timestamp 1676037725
transform 1 0 46828 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_505
timestamp 1676037725
transform 1 0 47564 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_509
timestamp 1676037725
transform 1 0 47932 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_519
timestamp 1676037725
transform 1 0 48852 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_531
timestamp 1676037725
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_533
timestamp 1676037725
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_545
timestamp 1676037725
transform 1 0 51244 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_557
timestamp 1676037725
transform 1 0 52348 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_569
timestamp 1676037725
transform 1 0 53452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_581
timestamp 1676037725
transform 1 0 54556 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_587
timestamp 1676037725
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_589
timestamp 1676037725
transform 1 0 55292 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_595
timestamp 1676037725
transform 1 0 55844 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_602
timestamp 1676037725
transform 1 0 56488 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_622
timestamp 1676037725
transform 1 0 58328 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_11
timestamp 1676037725
transform 1 0 2116 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_23
timestamp 1676037725
transform 1 0 3220 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_35
timestamp 1676037725
transform 1 0 4324 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_47
timestamp 1676037725
transform 1 0 5428 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1676037725
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1676037725
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1676037725
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1676037725
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1676037725
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1676037725
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1676037725
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1676037725
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1676037725
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1676037725
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1676037725
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1676037725
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_193
timestamp 1676037725
transform 1 0 18860 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_201
timestamp 1676037725
transform 1 0 19596 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_209
timestamp 1676037725
transform 1 0 20332 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_215
timestamp 1676037725
transform 1 0 20884 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_222
timestamp 1676037725
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_225
timestamp 1676037725
transform 1 0 21804 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_229
timestamp 1676037725
transform 1 0 22172 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_239
timestamp 1676037725
transform 1 0 23092 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_247
timestamp 1676037725
transform 1 0 23828 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_266
timestamp 1676037725
transform 1 0 25576 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_270
timestamp 1676037725
transform 1 0 25944 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_278
timestamp 1676037725
transform 1 0 26680 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_281
timestamp 1676037725
transform 1 0 26956 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_289
timestamp 1676037725
transform 1 0 27692 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_309
timestamp 1676037725
transform 1 0 29532 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_5_320
timestamp 1676037725
transform 1 0 30544 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_331
timestamp 1676037725
transform 1 0 31556 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1676037725
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_337
timestamp 1676037725
transform 1 0 32108 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_358
timestamp 1676037725
transform 1 0 34040 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_362
timestamp 1676037725
transform 1 0 34408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_367
timestamp 1676037725
transform 1 0 34868 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_373
timestamp 1676037725
transform 1 0 35420 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_388
timestamp 1676037725
transform 1 0 36800 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_393
timestamp 1676037725
transform 1 0 37260 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_404
timestamp 1676037725
transform 1 0 38272 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_412
timestamp 1676037725
transform 1 0 39008 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_430
timestamp 1676037725
transform 1 0 40664 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_438
timestamp 1676037725
transform 1 0 41400 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_446
timestamp 1676037725
transform 1 0 42136 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_449
timestamp 1676037725
transform 1 0 42412 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_455
timestamp 1676037725
transform 1 0 42964 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1676037725
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_473
timestamp 1676037725
transform 1 0 44620 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_477
timestamp 1676037725
transform 1 0 44988 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_481
timestamp 1676037725
transform 1 0 45356 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_489
timestamp 1676037725
transform 1 0 46092 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_495
timestamp 1676037725
transform 1 0 46644 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1676037725
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_505
timestamp 1676037725
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_517
timestamp 1676037725
transform 1 0 48668 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_529
timestamp 1676037725
transform 1 0 49772 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_541
timestamp 1676037725
transform 1 0 50876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_553
timestamp 1676037725
transform 1 0 51980 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_559
timestamp 1676037725
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_561
timestamp 1676037725
transform 1 0 52716 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_573
timestamp 1676037725
transform 1 0 53820 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_585
timestamp 1676037725
transform 1 0 54924 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_589
timestamp 1676037725
transform 1 0 55292 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_594
timestamp 1676037725
transform 1 0 55752 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_604
timestamp 1676037725
transform 1 0 56672 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_614
timestamp 1676037725
transform 1 0 57592 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_617
timestamp 1676037725
transform 1 0 57868 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_623
timestamp 1676037725
transform 1 0 58420 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_11
timestamp 1676037725
transform 1 0 2116 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_23
timestamp 1676037725
transform 1 0 3220 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1676037725
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1676037725
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1676037725
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1676037725
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1676037725
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1676037725
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_99
timestamp 1676037725
transform 1 0 10212 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1676037725
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1676037725
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1676037725
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1676037725
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1676037725
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1676037725
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_177
timestamp 1676037725
transform 1 0 17388 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_188
timestamp 1676037725
transform 1 0 18400 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_197
timestamp 1676037725
transform 1 0 19228 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_6_212
timestamp 1676037725
transform 1 0 20608 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_224
timestamp 1676037725
transform 1 0 21712 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_232
timestamp 1676037725
transform 1 0 22448 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_241
timestamp 1676037725
transform 1 0 23276 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_249
timestamp 1676037725
transform 1 0 24012 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_253
timestamp 1676037725
transform 1 0 24380 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_261
timestamp 1676037725
transform 1 0 25116 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_280
timestamp 1676037725
transform 1 0 26864 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_288
timestamp 1676037725
transform 1 0 27600 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_294
timestamp 1676037725
transform 1 0 28152 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_306
timestamp 1676037725
transform 1 0 29256 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_309
timestamp 1676037725
transform 1 0 29532 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_313
timestamp 1676037725
transform 1 0 29900 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_320
timestamp 1676037725
transform 1 0 30544 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_330
timestamp 1676037725
transform 1 0 31464 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_338
timestamp 1676037725
transform 1 0 32200 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_349
timestamp 1676037725
transform 1 0 33212 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_357
timestamp 1676037725
transform 1 0 33948 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_362
timestamp 1676037725
transform 1 0 34408 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_365
timestamp 1676037725
transform 1 0 34684 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_373
timestamp 1676037725
transform 1 0 35420 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_388
timestamp 1676037725
transform 1 0 36800 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_398
timestamp 1676037725
transform 1 0 37720 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_406
timestamp 1676037725
transform 1 0 38456 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_414
timestamp 1676037725
transform 1 0 39192 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_421
timestamp 1676037725
transform 1 0 39836 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_427
timestamp 1676037725
transform 1 0 40388 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_439
timestamp 1676037725
transform 1 0 41492 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_451
timestamp 1676037725
transform 1 0 42596 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_455
timestamp 1676037725
transform 1 0 42964 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_467
timestamp 1676037725
transform 1 0 44068 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1676037725
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_477
timestamp 1676037725
transform 1 0 44988 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_484
timestamp 1676037725
transform 1 0 45632 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_491
timestamp 1676037725
transform 1 0 46276 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_498
timestamp 1676037725
transform 1 0 46920 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_510
timestamp 1676037725
transform 1 0 48024 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_522
timestamp 1676037725
transform 1 0 49128 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_530
timestamp 1676037725
transform 1 0 49864 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_533
timestamp 1676037725
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_545
timestamp 1676037725
transform 1 0 51244 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_557
timestamp 1676037725
transform 1 0 52348 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_569
timestamp 1676037725
transform 1 0 53452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_581
timestamp 1676037725
transform 1 0 54556 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_587
timestamp 1676037725
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_589
timestamp 1676037725
transform 1 0 55292 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_597
timestamp 1676037725
transform 1 0 56028 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_601
timestamp 1676037725
transform 1 0 56396 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_621
timestamp 1676037725
transform 1 0 58236 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_11
timestamp 1676037725
transform 1 0 2116 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_23
timestamp 1676037725
transform 1 0 3220 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_35
timestamp 1676037725
transform 1 0 4324 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_47
timestamp 1676037725
transform 1 0 5428 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1676037725
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1676037725
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1676037725
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_93
timestamp 1676037725
transform 1 0 9660 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_108
timestamp 1676037725
transform 1 0 11040 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1676037725
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1676037725
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1676037725
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1676037725
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1676037725
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1676037725
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1676037725
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_205
timestamp 1676037725
transform 1 0 19964 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_219
timestamp 1676037725
transform 1 0 21252 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1676037725
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1676037725
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1676037725
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_249
timestamp 1676037725
transform 1 0 24012 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_257
timestamp 1676037725
transform 1 0 24748 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_267
timestamp 1676037725
transform 1 0 25668 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1676037725
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_281
timestamp 1676037725
transform 1 0 26956 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_292
timestamp 1676037725
transform 1 0 27968 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_304
timestamp 1676037725
transform 1 0 29072 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_308
timestamp 1676037725
transform 1 0 29440 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_314
timestamp 1676037725
transform 1 0 29992 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_325
timestamp 1676037725
transform 1 0 31004 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_333
timestamp 1676037725
transform 1 0 31740 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_337
timestamp 1676037725
transform 1 0 32108 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_341
timestamp 1676037725
transform 1 0 32476 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_347
timestamp 1676037725
transform 1 0 33028 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_359
timestamp 1676037725
transform 1 0 34132 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_366
timestamp 1676037725
transform 1 0 34776 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_384
timestamp 1676037725
transform 1 0 36432 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_393
timestamp 1676037725
transform 1 0 37260 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_401
timestamp 1676037725
transform 1 0 37996 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_409
timestamp 1676037725
transform 1 0 38732 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_416
timestamp 1676037725
transform 1 0 39376 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_423
timestamp 1676037725
transform 1 0 40020 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_430
timestamp 1676037725
transform 1 0 40664 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_442
timestamp 1676037725
transform 1 0 41768 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_449
timestamp 1676037725
transform 1 0 42412 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_453
timestamp 1676037725
transform 1 0 42780 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_471
timestamp 1676037725
transform 1 0 44436 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_484
timestamp 1676037725
transform 1 0 45632 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_496
timestamp 1676037725
transform 1 0 46736 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_505
timestamp 1676037725
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_517
timestamp 1676037725
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_529
timestamp 1676037725
transform 1 0 49772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_541
timestamp 1676037725
transform 1 0 50876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_553
timestamp 1676037725
transform 1 0 51980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_559
timestamp 1676037725
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_561
timestamp 1676037725
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_573
timestamp 1676037725
transform 1 0 53820 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_585
timestamp 1676037725
transform 1 0 54924 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_590
timestamp 1676037725
transform 1 0 55384 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_610
timestamp 1676037725
transform 1 0 57224 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_617
timestamp 1676037725
transform 1 0 57868 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_623
timestamp 1676037725
transform 1 0 58420 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_11
timestamp 1676037725
transform 1 0 2116 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_23
timestamp 1676037725
transform 1 0 3220 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1676037725
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1676037725
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1676037725
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1676037725
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1676037725
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1676037725
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1676037725
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1676037725
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1676037725
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1676037725
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1676037725
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1676037725
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1676037725
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1676037725
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1676037725
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1676037725
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_197
timestamp 1676037725
transform 1 0 19228 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_206
timestamp 1676037725
transform 1 0 20056 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_216
timestamp 1676037725
transform 1 0 20976 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_228
timestamp 1676037725
transform 1 0 22080 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_240
timestamp 1676037725
transform 1 0 23184 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_253
timestamp 1676037725
transform 1 0 24380 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_268
timestamp 1676037725
transform 1 0 25760 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_280
timestamp 1676037725
transform 1 0 26864 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_286
timestamp 1676037725
transform 1 0 27416 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_306
timestamp 1676037725
transform 1 0 29256 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_309
timestamp 1676037725
transform 1 0 29532 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_317
timestamp 1676037725
transform 1 0 30268 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_325
timestamp 1676037725
transform 1 0 31004 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_335
timestamp 1676037725
transform 1 0 31924 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_345
timestamp 1676037725
transform 1 0 32844 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_353
timestamp 1676037725
transform 1 0 33580 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_362
timestamp 1676037725
transform 1 0 34408 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_365
timestamp 1676037725
transform 1 0 34684 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_373
timestamp 1676037725
transform 1 0 35420 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_391
timestamp 1676037725
transform 1 0 37076 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_404
timestamp 1676037725
transform 1 0 38272 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_415
timestamp 1676037725
transform 1 0 39284 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1676037725
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_421
timestamp 1676037725
transform 1 0 39836 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_434
timestamp 1676037725
transform 1 0 41032 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_446
timestamp 1676037725
transform 1 0 42136 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_467
timestamp 1676037725
transform 1 0 44068 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_474
timestamp 1676037725
transform 1 0 44712 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_477
timestamp 1676037725
transform 1 0 44988 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_486
timestamp 1676037725
transform 1 0 45816 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_500
timestamp 1676037725
transform 1 0 47104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_504
timestamp 1676037725
transform 1 0 47472 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_512
timestamp 1676037725
transform 1 0 48208 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_524
timestamp 1676037725
transform 1 0 49312 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_533
timestamp 1676037725
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_545
timestamp 1676037725
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_557
timestamp 1676037725
transform 1 0 52348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_569
timestamp 1676037725
transform 1 0 53452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_581
timestamp 1676037725
transform 1 0 54556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_587
timestamp 1676037725
transform 1 0 55108 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_589
timestamp 1676037725
transform 1 0 55292 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_593
timestamp 1676037725
transform 1 0 55660 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_600
timestamp 1676037725
transform 1 0 56304 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_620
timestamp 1676037725
transform 1 0 58144 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_624
timestamp 1676037725
transform 1 0 58512 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_11
timestamp 1676037725
transform 1 0 2116 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_23
timestamp 1676037725
transform 1 0 3220 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_35
timestamp 1676037725
transform 1 0 4324 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_47
timestamp 1676037725
transform 1 0 5428 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1676037725
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1676037725
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1676037725
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_93
timestamp 1676037725
transform 1 0 9660 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_101
timestamp 1676037725
transform 1 0 10396 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_110
timestamp 1676037725
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_122
timestamp 1676037725
transform 1 0 12328 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_134
timestamp 1676037725
transform 1 0 13432 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_146
timestamp 1676037725
transform 1 0 14536 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_158
timestamp 1676037725
transform 1 0 15640 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_166
timestamp 1676037725
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1676037725
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1676037725
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_205
timestamp 1676037725
transform 1 0 19964 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_212
timestamp 1676037725
transform 1 0 20608 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1676037725
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1676037725
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_249
timestamp 1676037725
transform 1 0 24012 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_266
timestamp 1676037725
transform 1 0 25576 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_278
timestamp 1676037725
transform 1 0 26680 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1676037725
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_293
timestamp 1676037725
transform 1 0 28060 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_319
timestamp 1676037725
transform 1 0 30452 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_323
timestamp 1676037725
transform 1 0 30820 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_331
timestamp 1676037725
transform 1 0 31556 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1676037725
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_337
timestamp 1676037725
transform 1 0 32108 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_348
timestamp 1676037725
transform 1 0 33120 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_354
timestamp 1676037725
transform 1 0 33672 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_375
timestamp 1676037725
transform 1 0 35604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_387
timestamp 1676037725
transform 1 0 36708 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1676037725
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_393
timestamp 1676037725
transform 1 0 37260 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_409
timestamp 1676037725
transform 1 0 38732 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_420
timestamp 1676037725
transform 1 0 39744 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_432
timestamp 1676037725
transform 1 0 40848 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_444
timestamp 1676037725
transform 1 0 41952 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1676037725
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1676037725
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_473
timestamp 1676037725
transform 1 0 44620 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_483
timestamp 1676037725
transform 1 0 45540 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_491
timestamp 1676037725
transform 1 0 46276 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_499
timestamp 1676037725
transform 1 0 47012 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1676037725
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_505
timestamp 1676037725
transform 1 0 47564 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_512
timestamp 1676037725
transform 1 0 48208 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_524
timestamp 1676037725
transform 1 0 49312 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_536
timestamp 1676037725
transform 1 0 50416 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_548
timestamp 1676037725
transform 1 0 51520 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_561
timestamp 1676037725
transform 1 0 52716 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_573
timestamp 1676037725
transform 1 0 53820 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_585
timestamp 1676037725
transform 1 0 54924 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_591
timestamp 1676037725
transform 1 0 55476 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_596
timestamp 1676037725
transform 1 0 55936 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_604
timestamp 1676037725
transform 1 0 56672 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_614
timestamp 1676037725
transform 1 0 57592 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_617
timestamp 1676037725
transform 1 0 57868 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_623
timestamp 1676037725
transform 1 0 58420 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_11
timestamp 1676037725
transform 1 0 2116 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_23
timestamp 1676037725
transform 1 0 3220 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1676037725
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1676037725
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1676037725
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1676037725
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1676037725
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1676037725
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_103
timestamp 1676037725
transform 1 0 10580 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_114
timestamp 1676037725
transform 1 0 11592 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_118
timestamp 1676037725
transform 1 0 11960 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_125
timestamp 1676037725
transform 1 0 12604 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_135
timestamp 1676037725
transform 1 0 13524 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1676037725
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1676037725
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1676037725
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1676037725
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1676037725
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1676037725
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1676037725
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1676037725
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1676037725
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1676037725
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_233
timestamp 1676037725
transform 1 0 22540 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1676037725
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1676037725
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1676037725
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1676037725
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_277
timestamp 1676037725
transform 1 0 26588 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_281
timestamp 1676037725
transform 1 0 26956 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_287
timestamp 1676037725
transform 1 0 27508 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_300
timestamp 1676037725
transform 1 0 28704 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_10_309
timestamp 1676037725
transform 1 0 29532 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_315
timestamp 1676037725
transform 1 0 30084 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_325
timestamp 1676037725
transform 1 0 31004 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_337
timestamp 1676037725
transform 1 0 32108 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_349
timestamp 1676037725
transform 1 0 33212 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_355
timestamp 1676037725
transform 1 0 33764 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_362
timestamp 1676037725
transform 1 0 34408 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_365
timestamp 1676037725
transform 1 0 34684 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_373
timestamp 1676037725
transform 1 0 35420 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_388
timestamp 1676037725
transform 1 0 36800 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_406
timestamp 1676037725
transform 1 0 38456 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_418
timestamp 1676037725
transform 1 0 39560 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1676037725
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1676037725
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_445
timestamp 1676037725
transform 1 0 42044 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_453
timestamp 1676037725
transform 1 0 42780 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_464
timestamp 1676037725
transform 1 0 43792 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_477
timestamp 1676037725
transform 1 0 44988 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_485
timestamp 1676037725
transform 1 0 45724 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_495
timestamp 1676037725
transform 1 0 46644 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_503
timestamp 1676037725
transform 1 0 47380 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_520
timestamp 1676037725
transform 1 0 48944 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_533
timestamp 1676037725
transform 1 0 50140 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_545
timestamp 1676037725
transform 1 0 51244 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_557
timestamp 1676037725
transform 1 0 52348 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_569
timestamp 1676037725
transform 1 0 53452 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_581
timestamp 1676037725
transform 1 0 54556 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_587
timestamp 1676037725
transform 1 0 55108 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_589
timestamp 1676037725
transform 1 0 55292 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_601
timestamp 1676037725
transform 1 0 56396 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_10_610
timestamp 1676037725
transform 1 0 57224 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_616
timestamp 1676037725
transform 1 0 57776 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_623
timestamp 1676037725
transform 1 0 58420 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_11
timestamp 1676037725
transform 1 0 2116 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_23
timestamp 1676037725
transform 1 0 3220 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_35
timestamp 1676037725
transform 1 0 4324 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_47
timestamp 1676037725
transform 1 0 5428 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1676037725
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1676037725
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1676037725
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_93
timestamp 1676037725
transform 1 0 9660 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_101
timestamp 1676037725
transform 1 0 10396 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1676037725
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_113
timestamp 1676037725
transform 1 0 11500 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_119
timestamp 1676037725
transform 1 0 12052 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_127
timestamp 1676037725
transform 1 0 12788 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1676037725
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1676037725
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1676037725
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1676037725
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1676037725
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1676037725
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1676037725
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1676037725
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1676037725
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1676037725
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1676037725
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1676037725
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_249
timestamp 1676037725
transform 1 0 24012 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_267
timestamp 1676037725
transform 1 0 25668 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1676037725
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_281
timestamp 1676037725
transform 1 0 26956 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_289
timestamp 1676037725
transform 1 0 27692 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_300
timestamp 1676037725
transform 1 0 28704 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_310
timestamp 1676037725
transform 1 0 29624 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_333
timestamp 1676037725
transform 1 0 31740 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1676037725
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_349
timestamp 1676037725
transform 1 0 33212 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_358
timestamp 1676037725
transform 1 0 34040 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_362
timestamp 1676037725
transform 1 0 34408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_370
timestamp 1676037725
transform 1 0 35144 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_388
timestamp 1676037725
transform 1 0 36800 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_393
timestamp 1676037725
transform 1 0 37260 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_401
timestamp 1676037725
transform 1 0 37996 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_413
timestamp 1676037725
transform 1 0 39100 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_421
timestamp 1676037725
transform 1 0 39836 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_439
timestamp 1676037725
transform 1 0 41492 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1676037725
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_449
timestamp 1676037725
transform 1 0 42412 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_467
timestamp 1676037725
transform 1 0 44068 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_479
timestamp 1676037725
transform 1 0 45172 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_491
timestamp 1676037725
transform 1 0 46276 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1676037725
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_505
timestamp 1676037725
transform 1 0 47564 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_514
timestamp 1676037725
transform 1 0 48392 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_522
timestamp 1676037725
transform 1 0 49128 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_534
timestamp 1676037725
transform 1 0 50232 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_546
timestamp 1676037725
transform 1 0 51336 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_558
timestamp 1676037725
transform 1 0 52440 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_561
timestamp 1676037725
transform 1 0 52716 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_573
timestamp 1676037725
transform 1 0 53820 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_585
timestamp 1676037725
transform 1 0 54924 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_597
timestamp 1676037725
transform 1 0 56028 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_609
timestamp 1676037725
transform 1 0 57132 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_615
timestamp 1676037725
transform 1 0 57684 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_617
timestamp 1676037725
transform 1 0 57868 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_623
timestamp 1676037725
transform 1 0 58420 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_11
timestamp 1676037725
transform 1 0 2116 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_23
timestamp 1676037725
transform 1 0 3220 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1676037725
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1676037725
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1676037725
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1676037725
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1676037725
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1676037725
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1676037725
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1676037725
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_128
timestamp 1676037725
transform 1 0 12880 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1676037725
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1676037725
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1676037725
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1676037725
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1676037725
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1676037725
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1676037725
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1676037725
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1676037725
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_233
timestamp 1676037725
transform 1 0 22540 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_243
timestamp 1676037725
transform 1 0 23460 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1676037725
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_253
timestamp 1676037725
transform 1 0 24380 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_259
timestamp 1676037725
transform 1 0 24932 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_269
timestamp 1676037725
transform 1 0 25852 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_279
timestamp 1676037725
transform 1 0 26772 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_299
timestamp 1676037725
transform 1 0 28612 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_306
timestamp 1676037725
transform 1 0 29256 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_309
timestamp 1676037725
transform 1 0 29532 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_319
timestamp 1676037725
transform 1 0 30452 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_327
timestamp 1676037725
transform 1 0 31188 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_334
timestamp 1676037725
transform 1 0 31832 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_346
timestamp 1676037725
transform 1 0 32936 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_358
timestamp 1676037725
transform 1 0 34040 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_12_365
timestamp 1676037725
transform 1 0 34684 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_373
timestamp 1676037725
transform 1 0 35420 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_388
timestamp 1676037725
transform 1 0 36800 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_400
timestamp 1676037725
transform 1 0 37904 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_412
timestamp 1676037725
transform 1 0 39008 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_12_421
timestamp 1676037725
transform 1 0 39836 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_429
timestamp 1676037725
transform 1 0 40572 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_439
timestamp 1676037725
transform 1 0 41492 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_451
timestamp 1676037725
transform 1 0 42596 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_463
timestamp 1676037725
transform 1 0 43700 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1676037725
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1676037725
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_477
timestamp 1676037725
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_489
timestamp 1676037725
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_501
timestamp 1676037725
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_513
timestamp 1676037725
transform 1 0 48300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_525
timestamp 1676037725
transform 1 0 49404 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_531
timestamp 1676037725
transform 1 0 49956 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_533
timestamp 1676037725
transform 1 0 50140 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_545
timestamp 1676037725
transform 1 0 51244 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_557
timestamp 1676037725
transform 1 0 52348 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_569
timestamp 1676037725
transform 1 0 53452 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_581
timestamp 1676037725
transform 1 0 54556 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_587
timestamp 1676037725
transform 1 0 55108 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_589
timestamp 1676037725
transform 1 0 55292 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_601
timestamp 1676037725
transform 1 0 56396 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_621
timestamp 1676037725
transform 1 0 58236 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_11
timestamp 1676037725
transform 1 0 2116 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_23
timestamp 1676037725
transform 1 0 3220 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_35
timestamp 1676037725
transform 1 0 4324 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_47
timestamp 1676037725
transform 1 0 5428 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1676037725
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1676037725
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1676037725
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1676037725
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1676037725
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1676037725
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_113
timestamp 1676037725
transform 1 0 11500 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_121
timestamp 1676037725
transform 1 0 12236 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_129
timestamp 1676037725
transform 1 0 12972 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_139
timestamp 1676037725
transform 1 0 13892 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_151
timestamp 1676037725
transform 1 0 14996 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_163
timestamp 1676037725
transform 1 0 16100 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1676037725
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1676037725
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1676037725
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1676037725
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1676037725
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1676037725
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1676037725
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_225
timestamp 1676037725
transform 1 0 21804 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_233
timestamp 1676037725
transform 1 0 22540 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_244
timestamp 1676037725
transform 1 0 23552 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_264
timestamp 1676037725
transform 1 0 25392 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_272
timestamp 1676037725
transform 1 0 26128 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_278
timestamp 1676037725
transform 1 0 26680 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_281
timestamp 1676037725
transform 1 0 26956 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_299
timestamp 1676037725
transform 1 0 28612 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_311
timestamp 1676037725
transform 1 0 29716 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_320
timestamp 1676037725
transform 1 0 30544 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_324
timestamp 1676037725
transform 1 0 30912 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_334
timestamp 1676037725
transform 1 0 31832 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_337
timestamp 1676037725
transform 1 0 32108 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_345
timestamp 1676037725
transform 1 0 32844 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_354
timestamp 1676037725
transform 1 0 33672 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_374
timestamp 1676037725
transform 1 0 35512 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_387
timestamp 1676037725
transform 1 0 36708 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1676037725
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1676037725
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_405
timestamp 1676037725
transform 1 0 38364 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_409
timestamp 1676037725
transform 1 0 38732 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_417
timestamp 1676037725
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_429
timestamp 1676037725
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1676037725
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1676037725
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1676037725
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_461
timestamp 1676037725
transform 1 0 43516 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_476
timestamp 1676037725
transform 1 0 44896 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_480
timestamp 1676037725
transform 1 0 45264 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_490
timestamp 1676037725
transform 1 0 46184 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_502
timestamp 1676037725
transform 1 0 47288 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_505
timestamp 1676037725
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_517
timestamp 1676037725
transform 1 0 48668 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_529
timestamp 1676037725
transform 1 0 49772 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_541
timestamp 1676037725
transform 1 0 50876 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_553
timestamp 1676037725
transform 1 0 51980 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_559
timestamp 1676037725
transform 1 0 52532 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_561
timestamp 1676037725
transform 1 0 52716 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_573
timestamp 1676037725
transform 1 0 53820 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_585
timestamp 1676037725
transform 1 0 54924 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_597
timestamp 1676037725
transform 1 0 56028 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_604
timestamp 1676037725
transform 1 0 56672 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_614
timestamp 1676037725
transform 1 0 57592 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_617
timestamp 1676037725
transform 1 0 57868 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1676037725
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_11
timestamp 1676037725
transform 1 0 2116 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_23
timestamp 1676037725
transform 1 0 3220 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1676037725
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1676037725
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1676037725
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1676037725
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1676037725
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1676037725
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1676037725
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1676037725
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1676037725
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1676037725
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_121
timestamp 1676037725
transform 1 0 12236 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_129
timestamp 1676037725
transform 1 0 12972 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_137
timestamp 1676037725
transform 1 0 13708 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1676037725
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1676037725
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1676037725
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1676037725
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1676037725
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1676037725
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1676037725
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1676037725
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1676037725
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_233
timestamp 1676037725
transform 1 0 22540 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_247
timestamp 1676037725
transform 1 0 23828 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1676037725
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1676037725
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_271
timestamp 1676037725
transform 1 0 26036 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_279
timestamp 1676037725
transform 1 0 26772 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_14_286
timestamp 1676037725
transform 1 0 27416 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_292
timestamp 1676037725
transform 1 0 27968 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_297
timestamp 1676037725
transform 1 0 28428 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_305
timestamp 1676037725
transform 1 0 29164 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1676037725
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_321
timestamp 1676037725
transform 1 0 30636 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_347
timestamp 1676037725
transform 1 0 33028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_359
timestamp 1676037725
transform 1 0 34132 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1676037725
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_365
timestamp 1676037725
transform 1 0 34684 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_378
timestamp 1676037725
transform 1 0 35880 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_391
timestamp 1676037725
transform 1 0 37076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_403
timestamp 1676037725
transform 1 0 38180 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_416
timestamp 1676037725
transform 1 0 39376 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_421
timestamp 1676037725
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_433
timestamp 1676037725
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_445
timestamp 1676037725
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_457
timestamp 1676037725
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1676037725
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1676037725
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_477
timestamp 1676037725
transform 1 0 44988 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_495
timestamp 1676037725
transform 1 0 46644 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_507
timestamp 1676037725
transform 1 0 47748 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_519
timestamp 1676037725
transform 1 0 48852 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_531
timestamp 1676037725
transform 1 0 49956 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_533
timestamp 1676037725
transform 1 0 50140 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_545
timestamp 1676037725
transform 1 0 51244 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_557
timestamp 1676037725
transform 1 0 52348 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_569
timestamp 1676037725
transform 1 0 53452 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_581
timestamp 1676037725
transform 1 0 54556 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_587
timestamp 1676037725
transform 1 0 55108 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_589
timestamp 1676037725
transform 1 0 55292 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_601
timestamp 1676037725
transform 1 0 56396 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_621
timestamp 1676037725
transform 1 0 58236 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1676037725
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_11
timestamp 1676037725
transform 1 0 2116 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_23
timestamp 1676037725
transform 1 0 3220 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_35
timestamp 1676037725
transform 1 0 4324 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_47
timestamp 1676037725
transform 1 0 5428 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1676037725
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1676037725
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1676037725
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1676037725
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1676037725
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1676037725
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_113
timestamp 1676037725
transform 1 0 11500 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_121
timestamp 1676037725
transform 1 0 12236 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_129
timestamp 1676037725
transform 1 0 12972 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_139
timestamp 1676037725
transform 1 0 13892 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_151
timestamp 1676037725
transform 1 0 14996 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_163
timestamp 1676037725
transform 1 0 16100 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1676037725
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1676037725
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1676037725
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1676037725
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_205
timestamp 1676037725
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1676037725
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1676037725
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1676037725
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_237
timestamp 1676037725
transform 1 0 22908 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_241
timestamp 1676037725
transform 1 0 23276 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_252
timestamp 1676037725
transform 1 0 24288 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_260
timestamp 1676037725
transform 1 0 25024 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_272
timestamp 1676037725
transform 1 0 26128 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_281
timestamp 1676037725
transform 1 0 26956 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_289
timestamp 1676037725
transform 1 0 27692 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_299
timestamp 1676037725
transform 1 0 28612 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_320
timestamp 1676037725
transform 1 0 30544 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_332
timestamp 1676037725
transform 1 0 31648 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_337
timestamp 1676037725
transform 1 0 32108 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_15_360
timestamp 1676037725
transform 1 0 34224 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_368
timestamp 1676037725
transform 1 0 34960 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_371
timestamp 1676037725
transform 1 0 35236 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_382
timestamp 1676037725
transform 1 0 36248 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_390
timestamp 1676037725
transform 1 0 36984 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_393
timestamp 1676037725
transform 1 0 37260 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_401
timestamp 1676037725
transform 1 0 37996 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_420
timestamp 1676037725
transform 1 0 39744 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_427
timestamp 1676037725
transform 1 0 40388 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_439
timestamp 1676037725
transform 1 0 41492 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1676037725
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_449
timestamp 1676037725
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_461
timestamp 1676037725
transform 1 0 43516 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_469
timestamp 1676037725
transform 1 0 44252 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_488
timestamp 1676037725
transform 1 0 46000 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_501
timestamp 1676037725
transform 1 0 47196 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_505
timestamp 1676037725
transform 1 0 47564 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_517
timestamp 1676037725
transform 1 0 48668 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_529
timestamp 1676037725
transform 1 0 49772 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_541
timestamp 1676037725
transform 1 0 50876 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_553
timestamp 1676037725
transform 1 0 51980 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_559
timestamp 1676037725
transform 1 0 52532 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_561
timestamp 1676037725
transform 1 0 52716 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_573
timestamp 1676037725
transform 1 0 53820 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_585
timestamp 1676037725
transform 1 0 54924 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_597
timestamp 1676037725
transform 1 0 56028 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_604
timestamp 1676037725
transform 1 0 56672 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_614
timestamp 1676037725
transform 1 0 57592 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_617
timestamp 1676037725
transform 1 0 57868 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_622
timestamp 1676037725
transform 1 0 58328 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1676037725
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_11
timestamp 1676037725
transform 1 0 2116 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_23
timestamp 1676037725
transform 1 0 3220 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1676037725
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1676037725
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1676037725
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1676037725
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1676037725
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1676037725
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1676037725
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1676037725
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1676037725
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1676037725
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_121
timestamp 1676037725
transform 1 0 12236 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_129
timestamp 1676037725
transform 1 0 12972 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_136
timestamp 1676037725
transform 1 0 13616 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1676037725
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_150
timestamp 1676037725
transform 1 0 14904 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_160
timestamp 1676037725
transform 1 0 15824 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_168
timestamp 1676037725
transform 1 0 16560 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_176
timestamp 1676037725
transform 1 0 17296 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_188
timestamp 1676037725
transform 1 0 18400 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_197
timestamp 1676037725
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_205
timestamp 1676037725
transform 1 0 19964 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_217
timestamp 1676037725
transform 1 0 21068 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_229
timestamp 1676037725
transform 1 0 22172 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_250
timestamp 1676037725
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_253
timestamp 1676037725
transform 1 0 24380 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_259
timestamp 1676037725
transform 1 0 24932 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_271
timestamp 1676037725
transform 1 0 26036 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_283
timestamp 1676037725
transform 1 0 27140 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_295
timestamp 1676037725
transform 1 0 28244 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_306
timestamp 1676037725
transform 1 0 29256 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_309
timestamp 1676037725
transform 1 0 29532 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_319
timestamp 1676037725
transform 1 0 30452 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_325
timestamp 1676037725
transform 1 0 31004 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_347
timestamp 1676037725
transform 1 0 33028 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_359
timestamp 1676037725
transform 1 0 34132 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1676037725
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_365
timestamp 1676037725
transform 1 0 34684 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_369
timestamp 1676037725
transform 1 0 35052 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_386
timestamp 1676037725
transform 1 0 36616 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_397
timestamp 1676037725
transform 1 0 37628 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_409
timestamp 1676037725
transform 1 0 38732 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_418
timestamp 1676037725
transform 1 0 39560 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_421
timestamp 1676037725
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_433
timestamp 1676037725
transform 1 0 40940 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_458
timestamp 1676037725
transform 1 0 43240 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_470
timestamp 1676037725
transform 1 0 44344 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_477
timestamp 1676037725
transform 1 0 44988 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_488
timestamp 1676037725
transform 1 0 46000 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_501
timestamp 1676037725
transform 1 0 47196 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_509
timestamp 1676037725
transform 1 0 47932 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_519
timestamp 1676037725
transform 1 0 48852 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_531
timestamp 1676037725
transform 1 0 49956 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_533
timestamp 1676037725
transform 1 0 50140 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_545
timestamp 1676037725
transform 1 0 51244 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_557
timestamp 1676037725
transform 1 0 52348 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_569
timestamp 1676037725
transform 1 0 53452 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_581
timestamp 1676037725
transform 1 0 54556 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_587
timestamp 1676037725
transform 1 0 55108 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_589
timestamp 1676037725
transform 1 0 55292 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_601
timestamp 1676037725
transform 1 0 56396 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_613
timestamp 1676037725
transform 1 0 57500 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_623
timestamp 1676037725
transform 1 0 58420 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1676037725
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_11
timestamp 1676037725
transform 1 0 2116 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_23
timestamp 1676037725
transform 1 0 3220 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_35
timestamp 1676037725
transform 1 0 4324 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_47
timestamp 1676037725
transform 1 0 5428 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1676037725
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1676037725
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1676037725
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1676037725
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1676037725
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1676037725
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1676037725
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1676037725
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_125
timestamp 1676037725
transform 1 0 12604 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_129
timestamp 1676037725
transform 1 0 12972 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1676037725
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1676037725
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1676037725
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1676037725
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_169
timestamp 1676037725
transform 1 0 16652 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_177
timestamp 1676037725
transform 1 0 17388 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_187
timestamp 1676037725
transform 1 0 18308 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_199
timestamp 1676037725
transform 1 0 19412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_211
timestamp 1676037725
transform 1 0 20516 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1676037725
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1676037725
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_237
timestamp 1676037725
transform 1 0 22908 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_245
timestamp 1676037725
transform 1 0 23644 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_253
timestamp 1676037725
transform 1 0 24380 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_17_265
timestamp 1676037725
transform 1 0 25484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_277
timestamp 1676037725
transform 1 0 26588 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_281
timestamp 1676037725
transform 1 0 26956 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_287
timestamp 1676037725
transform 1 0 27508 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_299
timestamp 1676037725
transform 1 0 28612 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_307
timestamp 1676037725
transform 1 0 29348 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_325
timestamp 1676037725
transform 1 0 31004 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_334
timestamp 1676037725
transform 1 0 31832 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_337
timestamp 1676037725
transform 1 0 32108 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_348
timestamp 1676037725
transform 1 0 33120 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_360
timestamp 1676037725
transform 1 0 34224 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_364
timestamp 1676037725
transform 1 0 34592 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_370
timestamp 1676037725
transform 1 0 35144 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_390
timestamp 1676037725
transform 1 0 36984 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_393
timestamp 1676037725
transform 1 0 37260 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_404
timestamp 1676037725
transform 1 0 38272 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_416
timestamp 1676037725
transform 1 0 39376 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_428
timestamp 1676037725
transform 1 0 40480 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_446
timestamp 1676037725
transform 1 0 42136 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_449
timestamp 1676037725
transform 1 0 42412 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_457
timestamp 1676037725
transform 1 0 43148 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_465
timestamp 1676037725
transform 1 0 43884 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_483
timestamp 1676037725
transform 1 0 45540 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_493
timestamp 1676037725
transform 1 0 46460 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_501
timestamp 1676037725
transform 1 0 47196 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_505
timestamp 1676037725
transform 1 0 47564 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_513
timestamp 1676037725
transform 1 0 48300 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_529
timestamp 1676037725
transform 1 0 49772 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_541
timestamp 1676037725
transform 1 0 50876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_553
timestamp 1676037725
transform 1 0 51980 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_559
timestamp 1676037725
transform 1 0 52532 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_561
timestamp 1676037725
transform 1 0 52716 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_573
timestamp 1676037725
transform 1 0 53820 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_585
timestamp 1676037725
transform 1 0 54924 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_597
timestamp 1676037725
transform 1 0 56028 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_605
timestamp 1676037725
transform 1 0 56764 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_613
timestamp 1676037725
transform 1 0 57500 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_617
timestamp 1676037725
transform 1 0 57868 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_623
timestamp 1676037725
transform 1 0 58420 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1676037725
transform 1 0 1380 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_11
timestamp 1676037725
transform 1 0 2116 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_23
timestamp 1676037725
transform 1 0 3220 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1676037725
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1676037725
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1676037725
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1676037725
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1676037725
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1676037725
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1676037725
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1676037725
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1676037725
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1676037725
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_121
timestamp 1676037725
transform 1 0 12236 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_129
timestamp 1676037725
transform 1 0 12972 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1676037725
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1676037725
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1676037725
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1676037725
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1676037725
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1676037725
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1676037725
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1676037725
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1676037725
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_221
timestamp 1676037725
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_237
timestamp 1676037725
transform 1 0 22908 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1676037725
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1676037725
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_271
timestamp 1676037725
transform 1 0 26036 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_283
timestamp 1676037725
transform 1 0 27140 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_295
timestamp 1676037725
transform 1 0 28244 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_301
timestamp 1676037725
transform 1 0 28796 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_306
timestamp 1676037725
transform 1 0 29256 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_309
timestamp 1676037725
transform 1 0 29532 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_317
timestamp 1676037725
transform 1 0 30268 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_335
timestamp 1676037725
transform 1 0 31924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_347
timestamp 1676037725
transform 1 0 33028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_359
timestamp 1676037725
transform 1 0 34132 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1676037725
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1676037725
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_377
timestamp 1676037725
transform 1 0 35788 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_400
timestamp 1676037725
transform 1 0 37904 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_412
timestamp 1676037725
transform 1 0 39008 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_18_421
timestamp 1676037725
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_433
timestamp 1676037725
transform 1 0 40940 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_448
timestamp 1676037725
transform 1 0 42320 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_461
timestamp 1676037725
transform 1 0 43516 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_473
timestamp 1676037725
transform 1 0 44620 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_477
timestamp 1676037725
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_489
timestamp 1676037725
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_501
timestamp 1676037725
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_513
timestamp 1676037725
transform 1 0 48300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_530
timestamp 1676037725
transform 1 0 49864 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_533
timestamp 1676037725
transform 1 0 50140 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_551
timestamp 1676037725
transform 1 0 51796 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_563
timestamp 1676037725
transform 1 0 52900 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_575
timestamp 1676037725
transform 1 0 54004 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_587
timestamp 1676037725
transform 1 0 55108 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_589
timestamp 1676037725
transform 1 0 55292 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_601
timestamp 1676037725
transform 1 0 56396 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_621
timestamp 1676037725
transform 1 0 58236 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1676037725
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_11
timestamp 1676037725
transform 1 0 2116 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_23
timestamp 1676037725
transform 1 0 3220 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_35
timestamp 1676037725
transform 1 0 4324 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_47
timestamp 1676037725
transform 1 0 5428 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1676037725
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1676037725
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1676037725
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1676037725
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1676037725
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1676037725
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1676037725
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1676037725
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1676037725
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1676037725
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1676037725
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1676037725
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1676037725
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1676037725
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1676037725
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1676037725
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_205
timestamp 1676037725
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1676037725
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1676037725
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1676037725
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_246
timestamp 1676037725
transform 1 0 23736 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_266
timestamp 1676037725
transform 1 0 25576 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_274
timestamp 1676037725
transform 1 0 26312 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1676037725
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_293
timestamp 1676037725
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_305
timestamp 1676037725
transform 1 0 29164 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_309
timestamp 1676037725
transform 1 0 29532 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_314
timestamp 1676037725
transform 1 0 29992 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_326
timestamp 1676037725
transform 1 0 31096 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_334
timestamp 1676037725
transform 1 0 31832 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1676037725
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_349
timestamp 1676037725
transform 1 0 33212 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_375
timestamp 1676037725
transform 1 0 35604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_387
timestamp 1676037725
transform 1 0 36708 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1676037725
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_393
timestamp 1676037725
transform 1 0 37260 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_404
timestamp 1676037725
transform 1 0 38272 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_416
timestamp 1676037725
transform 1 0 39376 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_428
timestamp 1676037725
transform 1 0 40480 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_440
timestamp 1676037725
transform 1 0 41584 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_449
timestamp 1676037725
transform 1 0 42412 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_460
timestamp 1676037725
transform 1 0 43424 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_472
timestamp 1676037725
transform 1 0 44528 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_484
timestamp 1676037725
transform 1 0 45632 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_496
timestamp 1676037725
transform 1 0 46736 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_19_505
timestamp 1676037725
transform 1 0 47564 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_517
timestamp 1676037725
transform 1 0 48668 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_545
timestamp 1676037725
transform 1 0 51244 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_555
timestamp 1676037725
transform 1 0 52164 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_559
timestamp 1676037725
transform 1 0 52532 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_561
timestamp 1676037725
transform 1 0 52716 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_573
timestamp 1676037725
transform 1 0 53820 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_585
timestamp 1676037725
transform 1 0 54924 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_591
timestamp 1676037725
transform 1 0 55476 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_599
timestamp 1676037725
transform 1 0 56212 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_612
timestamp 1676037725
transform 1 0 57408 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_617
timestamp 1676037725
transform 1 0 57868 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_623
timestamp 1676037725
transform 1 0 58420 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1676037725
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_11
timestamp 1676037725
transform 1 0 2116 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_23
timestamp 1676037725
transform 1 0 3220 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1676037725
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1676037725
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1676037725
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1676037725
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1676037725
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1676037725
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1676037725
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1676037725
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1676037725
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1676037725
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1676037725
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1676037725
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1676037725
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1676037725
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_153
timestamp 1676037725
transform 1 0 15180 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1676037725
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1676037725
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1676037725
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1676037725
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1676037725
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_209
timestamp 1676037725
transform 1 0 20332 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_221
timestamp 1676037725
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_233
timestamp 1676037725
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_249
timestamp 1676037725
transform 1 0 24012 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_253
timestamp 1676037725
transform 1 0 24380 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_261
timestamp 1676037725
transform 1 0 25116 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_278
timestamp 1676037725
transform 1 0 26680 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_291
timestamp 1676037725
transform 1 0 27876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_303
timestamp 1676037725
transform 1 0 28980 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1676037725
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_309
timestamp 1676037725
transform 1 0 29532 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_319
timestamp 1676037725
transform 1 0 30452 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_327
timestamp 1676037725
transform 1 0 31188 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_339
timestamp 1676037725
transform 1 0 32292 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_346
timestamp 1676037725
transform 1 0 32936 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_362
timestamp 1676037725
transform 1 0 34408 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1676037725
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_377
timestamp 1676037725
transform 1 0 35788 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_398
timestamp 1676037725
transform 1 0 37720 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_410
timestamp 1676037725
transform 1 0 38824 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_418
timestamp 1676037725
transform 1 0 39560 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_421
timestamp 1676037725
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_433
timestamp 1676037725
transform 1 0 40940 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_441
timestamp 1676037725
transform 1 0 41676 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_462
timestamp 1676037725
transform 1 0 43608 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_474
timestamp 1676037725
transform 1 0 44712 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_477
timestamp 1676037725
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_489
timestamp 1676037725
transform 1 0 46092 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_517
timestamp 1676037725
transform 1 0 48668 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_529
timestamp 1676037725
transform 1 0 49772 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_533
timestamp 1676037725
transform 1 0 50140 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_543
timestamp 1676037725
transform 1 0 51060 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_547
timestamp 1676037725
transform 1 0 51428 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_559
timestamp 1676037725
transform 1 0 52532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_571
timestamp 1676037725
transform 1 0 53636 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_583
timestamp 1676037725
transform 1 0 54740 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_587
timestamp 1676037725
transform 1 0 55108 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_589
timestamp 1676037725
transform 1 0 55292 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_601
timestamp 1676037725
transform 1 0 56396 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_622
timestamp 1676037725
transform 1 0 58328 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1676037725
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_11
timestamp 1676037725
transform 1 0 2116 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_23
timestamp 1676037725
transform 1 0 3220 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_35
timestamp 1676037725
transform 1 0 4324 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_47
timestamp 1676037725
transform 1 0 5428 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1676037725
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1676037725
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1676037725
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1676037725
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1676037725
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1676037725
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1676037725
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1676037725
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1676037725
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1676037725
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_149
timestamp 1676037725
transform 1 0 14812 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_158
timestamp 1676037725
transform 1 0 15640 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1676037725
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1676037725
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1676037725
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_193
timestamp 1676037725
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_205
timestamp 1676037725
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_217
timestamp 1676037725
transform 1 0 21068 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1676037725
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1676037725
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_237
timestamp 1676037725
transform 1 0 22908 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_245
timestamp 1676037725
transform 1 0 23644 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_256
timestamp 1676037725
transform 1 0 24656 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_278
timestamp 1676037725
transform 1 0 26680 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_281
timestamp 1676037725
transform 1 0 26956 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_291
timestamp 1676037725
transform 1 0 27876 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_303
timestamp 1676037725
transform 1 0 28980 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_312
timestamp 1676037725
transform 1 0 29808 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_318
timestamp 1676037725
transform 1 0 30360 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_323
timestamp 1676037725
transform 1 0 30820 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_21_333
timestamp 1676037725
transform 1 0 31740 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_337
timestamp 1676037725
transform 1 0 32108 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_346
timestamp 1676037725
transform 1 0 32936 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_353
timestamp 1676037725
transform 1 0 33580 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1676037725
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1676037725
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1676037725
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_393
timestamp 1676037725
transform 1 0 37260 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_404
timestamp 1676037725
transform 1 0 38272 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_416
timestamp 1676037725
transform 1 0 39376 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_428
timestamp 1676037725
transform 1 0 40480 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_440
timestamp 1676037725
transform 1 0 41584 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_449
timestamp 1676037725
transform 1 0 42412 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_467
timestamp 1676037725
transform 1 0 44068 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_479
timestamp 1676037725
transform 1 0 45172 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_491
timestamp 1676037725
transform 1 0 46276 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1676037725
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_505
timestamp 1676037725
transform 1 0 47564 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_517
timestamp 1676037725
transform 1 0 48668 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_529
timestamp 1676037725
transform 1 0 49772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_532
timestamp 1676037725
transform 1 0 50048 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_542
timestamp 1676037725
transform 1 0 50968 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_554
timestamp 1676037725
transform 1 0 52072 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_561
timestamp 1676037725
transform 1 0 52716 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_573
timestamp 1676037725
transform 1 0 53820 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_585
timestamp 1676037725
transform 1 0 54924 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_597
timestamp 1676037725
transform 1 0 56028 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_604
timestamp 1676037725
transform 1 0 56672 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_614
timestamp 1676037725
transform 1 0 57592 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_617
timestamp 1676037725
transform 1 0 57868 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_623
timestamp 1676037725
transform 1 0 58420 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1676037725
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_11
timestamp 1676037725
transform 1 0 2116 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_23
timestamp 1676037725
transform 1 0 3220 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1676037725
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1676037725
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1676037725
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1676037725
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1676037725
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1676037725
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1676037725
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1676037725
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1676037725
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1676037725
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1676037725
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1676037725
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1676037725
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_141
timestamp 1676037725
transform 1 0 14076 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_156
timestamp 1676037725
transform 1 0 15456 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_166
timestamp 1676037725
transform 1 0 16376 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_182
timestamp 1676037725
transform 1 0 17848 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1676037725
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_197
timestamp 1676037725
transform 1 0 19228 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_205
timestamp 1676037725
transform 1 0 19964 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_213
timestamp 1676037725
transform 1 0 20700 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_221
timestamp 1676037725
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_233
timestamp 1676037725
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_249
timestamp 1676037725
transform 1 0 24012 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_253
timestamp 1676037725
transform 1 0 24380 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_259
timestamp 1676037725
transform 1 0 24932 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_264
timestamp 1676037725
transform 1 0 25392 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_272
timestamp 1676037725
transform 1 0 26128 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_282
timestamp 1676037725
transform 1 0 27048 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_294
timestamp 1676037725
transform 1 0 28152 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_298
timestamp 1676037725
transform 1 0 28520 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_306
timestamp 1676037725
transform 1 0 29256 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_309
timestamp 1676037725
transform 1 0 29532 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_327
timestamp 1676037725
transform 1 0 31188 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_335
timestamp 1676037725
transform 1 0 31924 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_342
timestamp 1676037725
transform 1 0 32568 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_346
timestamp 1676037725
transform 1 0 32936 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_354
timestamp 1676037725
transform 1 0 33672 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_362
timestamp 1676037725
transform 1 0 34408 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_365
timestamp 1676037725
transform 1 0 34684 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_371
timestamp 1676037725
transform 1 0 35236 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_378
timestamp 1676037725
transform 1 0 35880 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_390
timestamp 1676037725
transform 1 0 36984 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_402
timestamp 1676037725
transform 1 0 38088 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_414
timestamp 1676037725
transform 1 0 39192 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_22_421
timestamp 1676037725
transform 1 0 39836 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_426
timestamp 1676037725
transform 1 0 40296 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_437
timestamp 1676037725
transform 1 0 41308 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_449
timestamp 1676037725
transform 1 0 42412 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_461
timestamp 1676037725
transform 1 0 43516 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_473
timestamp 1676037725
transform 1 0 44620 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_477
timestamp 1676037725
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_489
timestamp 1676037725
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_501
timestamp 1676037725
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_513
timestamp 1676037725
transform 1 0 48300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_525
timestamp 1676037725
transform 1 0 49404 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_530
timestamp 1676037725
transform 1 0 49864 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_533
timestamp 1676037725
transform 1 0 50140 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_551
timestamp 1676037725
transform 1 0 51796 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_563
timestamp 1676037725
transform 1 0 52900 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_575
timestamp 1676037725
transform 1 0 54004 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_587
timestamp 1676037725
transform 1 0 55108 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_589
timestamp 1676037725
transform 1 0 55292 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_601
timestamp 1676037725
transform 1 0 56396 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_613
timestamp 1676037725
transform 1 0 57500 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_623
timestamp 1676037725
transform 1 0 58420 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1676037725
transform 1 0 1380 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_11
timestamp 1676037725
transform 1 0 2116 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_23
timestamp 1676037725
transform 1 0 3220 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_35
timestamp 1676037725
transform 1 0 4324 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_47
timestamp 1676037725
transform 1 0 5428 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1676037725
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1676037725
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1676037725
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1676037725
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1676037725
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1676037725
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1676037725
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1676037725
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1676037725
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1676037725
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_149
timestamp 1676037725
transform 1 0 14812 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_159
timestamp 1676037725
transform 1 0 15732 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1676037725
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_169
timestamp 1676037725
transform 1 0 16652 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_177
timestamp 1676037725
transform 1 0 17388 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_184
timestamp 1676037725
transform 1 0 18032 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_192
timestamp 1676037725
transform 1 0 18768 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_204
timestamp 1676037725
transform 1 0 19872 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_212
timestamp 1676037725
transform 1 0 20608 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_220
timestamp 1676037725
transform 1 0 21344 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_225
timestamp 1676037725
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_236
timestamp 1676037725
transform 1 0 22816 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_244
timestamp 1676037725
transform 1 0 23552 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_256
timestamp 1676037725
transform 1 0 24656 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_265
timestamp 1676037725
transform 1 0 25484 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_278
timestamp 1676037725
transform 1 0 26680 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1676037725
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_293
timestamp 1676037725
transform 1 0 28060 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_301
timestamp 1676037725
transform 1 0 28796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_309
timestamp 1676037725
transform 1 0 29532 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_317
timestamp 1676037725
transform 1 0 30268 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_325
timestamp 1676037725
transform 1 0 31004 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_330
timestamp 1676037725
transform 1 0 31464 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_337
timestamp 1676037725
transform 1 0 32108 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_343
timestamp 1676037725
transform 1 0 32660 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_358
timestamp 1676037725
transform 1 0 34040 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_366
timestamp 1676037725
transform 1 0 34776 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_378
timestamp 1676037725
transform 1 0 35880 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_390
timestamp 1676037725
transform 1 0 36984 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_393
timestamp 1676037725
transform 1 0 37260 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_414
timestamp 1676037725
transform 1 0 39192 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_23_438
timestamp 1676037725
transform 1 0 41400 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_446
timestamp 1676037725
transform 1 0 42136 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_449
timestamp 1676037725
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_470
timestamp 1676037725
transform 1 0 44344 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_482
timestamp 1676037725
transform 1 0 45448 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_494
timestamp 1676037725
transform 1 0 46552 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_502
timestamp 1676037725
transform 1 0 47288 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_505
timestamp 1676037725
transform 1 0 47564 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_512
timestamp 1676037725
transform 1 0 48208 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_524
timestamp 1676037725
transform 1 0 49312 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_532
timestamp 1676037725
transform 1 0 50048 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_536
timestamp 1676037725
transform 1 0 50416 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_546
timestamp 1676037725
transform 1 0 51336 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_558
timestamp 1676037725
transform 1 0 52440 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_561
timestamp 1676037725
transform 1 0 52716 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_573
timestamp 1676037725
transform 1 0 53820 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_586
timestamp 1676037725
transform 1 0 55016 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_598
timestamp 1676037725
transform 1 0 56120 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_610
timestamp 1676037725
transform 1 0 57224 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_617
timestamp 1676037725
transform 1 0 57868 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_623
timestamp 1676037725
transform 1 0 58420 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1676037725
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_11
timestamp 1676037725
transform 1 0 2116 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_23
timestamp 1676037725
transform 1 0 3220 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1676037725
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1676037725
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1676037725
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1676037725
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1676037725
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1676037725
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1676037725
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1676037725
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_97
timestamp 1676037725
transform 1 0 10028 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_103
timestamp 1676037725
transform 1 0 10580 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_118
timestamp 1676037725
transform 1 0 11960 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_130
timestamp 1676037725
transform 1 0 13064 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1676037725
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_141
timestamp 1676037725
transform 1 0 14076 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_145
timestamp 1676037725
transform 1 0 14444 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_153
timestamp 1676037725
transform 1 0 15180 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_164
timestamp 1676037725
transform 1 0 16192 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_172
timestamp 1676037725
transform 1 0 16928 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_182
timestamp 1676037725
transform 1 0 17848 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_191
timestamp 1676037725
transform 1 0 18676 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1676037725
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_197
timestamp 1676037725
transform 1 0 19228 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_24_211
timestamp 1676037725
transform 1 0 20516 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_217
timestamp 1676037725
transform 1 0 21068 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_225
timestamp 1676037725
transform 1 0 21804 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_229
timestamp 1676037725
transform 1 0 22172 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_239
timestamp 1676037725
transform 1 0 23092 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_247
timestamp 1676037725
transform 1 0 23828 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1676037725
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_253
timestamp 1676037725
transform 1 0 24380 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_268
timestamp 1676037725
transform 1 0 25760 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_280
timestamp 1676037725
transform 1 0 26864 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_292
timestamp 1676037725
transform 1 0 27968 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_298
timestamp 1676037725
transform 1 0 28520 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_306
timestamp 1676037725
transform 1 0 29256 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_309
timestamp 1676037725
transform 1 0 29532 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_318
timestamp 1676037725
transform 1 0 30360 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_327
timestamp 1676037725
transform 1 0 31188 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_331
timestamp 1676037725
transform 1 0 31556 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_340
timestamp 1676037725
transform 1 0 32384 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_348
timestamp 1676037725
transform 1 0 33120 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_352
timestamp 1676037725
transform 1 0 33488 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_358
timestamp 1676037725
transform 1 0 34040 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1676037725
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1676037725
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1676037725
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_401
timestamp 1676037725
transform 1 0 37996 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_412
timestamp 1676037725
transform 1 0 39008 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_24_421
timestamp 1676037725
transform 1 0 39836 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_429
timestamp 1676037725
transform 1 0 40572 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_447
timestamp 1676037725
transform 1 0 42228 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_472
timestamp 1676037725
transform 1 0 44528 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_477
timestamp 1676037725
transform 1 0 44988 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_500
timestamp 1676037725
transform 1 0 47104 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_512
timestamp 1676037725
transform 1 0 48208 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_524
timestamp 1676037725
transform 1 0 49312 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_533
timestamp 1676037725
transform 1 0 50140 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_544
timestamp 1676037725
transform 1 0 51152 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_555
timestamp 1676037725
transform 1 0 52164 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_567
timestamp 1676037725
transform 1 0 53268 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_579
timestamp 1676037725
transform 1 0 54372 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_587
timestamp 1676037725
transform 1 0 55108 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_589
timestamp 1676037725
transform 1 0 55292 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_601
timestamp 1676037725
transform 1 0 56396 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_613
timestamp 1676037725
transform 1 0 57500 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_623
timestamp 1676037725
transform 1 0 58420 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1676037725
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_11
timestamp 1676037725
transform 1 0 2116 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_23
timestamp 1676037725
transform 1 0 3220 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_35
timestamp 1676037725
transform 1 0 4324 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_47
timestamp 1676037725
transform 1 0 5428 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1676037725
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1676037725
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1676037725
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1676037725
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1676037725
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1676037725
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1676037725
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1676037725
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1676037725
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1676037725
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1676037725
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_161
timestamp 1676037725
transform 1 0 15916 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1676037725
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_169
timestamp 1676037725
transform 1 0 16652 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_192
timestamp 1676037725
transform 1 0 18768 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_200
timestamp 1676037725
transform 1 0 19504 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_220
timestamp 1676037725
transform 1 0 21344 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_225
timestamp 1676037725
transform 1 0 21804 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_235
timestamp 1676037725
transform 1 0 22724 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_245
timestamp 1676037725
transform 1 0 23644 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_256
timestamp 1676037725
transform 1 0 24656 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1676037725
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1676037725
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_281
timestamp 1676037725
transform 1 0 26956 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_289
timestamp 1676037725
transform 1 0 27692 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_296
timestamp 1676037725
transform 1 0 28336 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_316
timestamp 1676037725
transform 1 0 30176 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_325
timestamp 1676037725
transform 1 0 31004 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_334
timestamp 1676037725
transform 1 0 31832 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_337
timestamp 1676037725
transform 1 0 32108 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_359
timestamp 1676037725
transform 1 0 34132 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_366
timestamp 1676037725
transform 1 0 34776 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_372
timestamp 1676037725
transform 1 0 35328 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_377
timestamp 1676037725
transform 1 0 35788 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_385
timestamp 1676037725
transform 1 0 36524 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_390
timestamp 1676037725
transform 1 0 36984 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_393
timestamp 1676037725
transform 1 0 37260 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_404
timestamp 1676037725
transform 1 0 38272 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_425
timestamp 1676037725
transform 1 0 40204 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_433
timestamp 1676037725
transform 1 0 40940 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_445
timestamp 1676037725
transform 1 0 42044 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_449
timestamp 1676037725
transform 1 0 42412 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_457
timestamp 1676037725
transform 1 0 43148 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_464
timestamp 1676037725
transform 1 0 43792 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_488
timestamp 1676037725
transform 1 0 46000 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_501
timestamp 1676037725
transform 1 0 47196 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_505
timestamp 1676037725
transform 1 0 47564 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_523
timestamp 1676037725
transform 1 0 49220 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_531
timestamp 1676037725
transform 1 0 49956 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_548
timestamp 1676037725
transform 1 0 51520 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_561
timestamp 1676037725
transform 1 0 52716 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_573
timestamp 1676037725
transform 1 0 53820 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_594
timestamp 1676037725
transform 1 0 55752 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_606
timestamp 1676037725
transform 1 0 56856 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_614
timestamp 1676037725
transform 1 0 57592 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_617
timestamp 1676037725
transform 1 0 57868 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_623
timestamp 1676037725
transform 1 0 58420 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1676037725
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_11
timestamp 1676037725
transform 1 0 2116 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_23
timestamp 1676037725
transform 1 0 3220 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1676037725
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1676037725
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1676037725
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1676037725
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1676037725
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1676037725
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1676037725
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1676037725
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1676037725
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1676037725
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1676037725
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1676037725
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1676037725
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1676037725
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1676037725
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_165
timestamp 1676037725
transform 1 0 16284 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_171
timestamp 1676037725
transform 1 0 16836 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1676037725
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_197
timestamp 1676037725
transform 1 0 19228 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_205
timestamp 1676037725
transform 1 0 19964 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_225
timestamp 1676037725
transform 1 0 21804 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_246
timestamp 1676037725
transform 1 0 23736 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_26_253
timestamp 1676037725
transform 1 0 24380 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_259
timestamp 1676037725
transform 1 0 24932 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_268
timestamp 1676037725
transform 1 0 25760 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_283
timestamp 1676037725
transform 1 0 27140 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_296
timestamp 1676037725
transform 1 0 28336 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_306
timestamp 1676037725
transform 1 0 29256 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_309
timestamp 1676037725
transform 1 0 29532 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_327
timestamp 1676037725
transform 1 0 31188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_333
timestamp 1676037725
transform 1 0 31740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_350
timestamp 1676037725
transform 1 0 33304 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_358
timestamp 1676037725
transform 1 0 34040 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_365
timestamp 1676037725
transform 1 0 34684 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_375
timestamp 1676037725
transform 1 0 35604 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_383
timestamp 1676037725
transform 1 0 36340 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_391
timestamp 1676037725
transform 1 0 37076 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_398
timestamp 1676037725
transform 1 0 37720 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_418
timestamp 1676037725
transform 1 0 39560 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_421
timestamp 1676037725
transform 1 0 39836 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_432
timestamp 1676037725
transform 1 0 40848 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_444
timestamp 1676037725
transform 1 0 41952 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_456
timestamp 1676037725
transform 1 0 43056 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_462
timestamp 1676037725
transform 1 0 43608 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_474
timestamp 1676037725
transform 1 0 44712 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_477
timestamp 1676037725
transform 1 0 44988 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_496
timestamp 1676037725
transform 1 0 46736 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_505
timestamp 1676037725
transform 1 0 47564 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_513
timestamp 1676037725
transform 1 0 48300 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_522
timestamp 1676037725
transform 1 0 49128 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_530
timestamp 1676037725
transform 1 0 49864 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_533
timestamp 1676037725
transform 1 0 50140 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_26_545
timestamp 1676037725
transform 1 0 51244 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_567
timestamp 1676037725
transform 1 0 53268 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_579
timestamp 1676037725
transform 1 0 54372 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_585
timestamp 1676037725
transform 1 0 54924 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_589
timestamp 1676037725
transform 1 0 55292 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_602
timestamp 1676037725
transform 1 0 56488 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_622
timestamp 1676037725
transform 1 0 58328 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1676037725
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_11
timestamp 1676037725
transform 1 0 2116 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_23
timestamp 1676037725
transform 1 0 3220 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_35
timestamp 1676037725
transform 1 0 4324 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_47
timestamp 1676037725
transform 1 0 5428 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1676037725
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1676037725
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1676037725
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1676037725
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1676037725
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1676037725
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1676037725
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1676037725
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1676037725
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1676037725
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1676037725
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1676037725
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1676037725
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_169
timestamp 1676037725
transform 1 0 16652 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_177
timestamp 1676037725
transform 1 0 17388 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_183
timestamp 1676037725
transform 1 0 17940 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_191
timestamp 1676037725
transform 1 0 18676 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_210
timestamp 1676037725
transform 1 0 20424 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_218
timestamp 1676037725
transform 1 0 21160 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_225
timestamp 1676037725
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_231
timestamp 1676037725
transform 1 0 22356 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_241
timestamp 1676037725
transform 1 0 23276 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_252
timestamp 1676037725
transform 1 0 24288 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_268
timestamp 1676037725
transform 1 0 25760 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_278
timestamp 1676037725
transform 1 0 26680 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_281
timestamp 1676037725
transform 1 0 26956 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_290
timestamp 1676037725
transform 1 0 27784 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_298
timestamp 1676037725
transform 1 0 28520 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_317
timestamp 1676037725
transform 1 0 30268 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_325
timestamp 1676037725
transform 1 0 31004 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_329
timestamp 1676037725
transform 1 0 31372 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_334
timestamp 1676037725
transform 1 0 31832 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_337
timestamp 1676037725
transform 1 0 32108 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_343
timestamp 1676037725
transform 1 0 32660 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_351
timestamp 1676037725
transform 1 0 33396 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_369
timestamp 1676037725
transform 1 0 35052 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_390
timestamp 1676037725
transform 1 0 36984 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_393
timestamp 1676037725
transform 1 0 37260 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_399
timestamp 1676037725
transform 1 0 37812 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_412
timestamp 1676037725
transform 1 0 39008 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_420
timestamp 1676037725
transform 1 0 39744 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_428
timestamp 1676037725
transform 1 0 40480 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_436
timestamp 1676037725
transform 1 0 41216 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_442
timestamp 1676037725
transform 1 0 41768 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_449
timestamp 1676037725
transform 1 0 42412 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_459
timestamp 1676037725
transform 1 0 43332 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_463
timestamp 1676037725
transform 1 0 43700 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_470
timestamp 1676037725
transform 1 0 44344 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_485
timestamp 1676037725
transform 1 0 45724 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_495
timestamp 1676037725
transform 1 0 46644 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1676037725
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_505
timestamp 1676037725
transform 1 0 47564 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_525
timestamp 1676037725
transform 1 0 49404 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_537
timestamp 1676037725
transform 1 0 50508 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_549
timestamp 1676037725
transform 1 0 51612 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_558
timestamp 1676037725
transform 1 0 52440 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_561
timestamp 1676037725
transform 1 0 52716 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_573
timestamp 1676037725
transform 1 0 53820 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_585
timestamp 1676037725
transform 1 0 54924 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_593
timestamp 1676037725
transform 1 0 55660 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_603
timestamp 1676037725
transform 1 0 56580 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_607
timestamp 1676037725
transform 1 0 56948 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_614
timestamp 1676037725
transform 1 0 57592 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_617
timestamp 1676037725
transform 1 0 57868 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_623
timestamp 1676037725
transform 1 0 58420 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1676037725
transform 1 0 1380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_11
timestamp 1676037725
transform 1 0 2116 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1676037725
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1676037725
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1676037725
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1676037725
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1676037725
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1676037725
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1676037725
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1676037725
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1676037725
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1676037725
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1676037725
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1676037725
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1676037725
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1676037725
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1676037725
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1676037725
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1676037725
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_177
timestamp 1676037725
transform 1 0 17388 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_181
timestamp 1676037725
transform 1 0 17756 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_185
timestamp 1676037725
transform 1 0 18124 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_193
timestamp 1676037725
transform 1 0 18860 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1676037725
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_209
timestamp 1676037725
transform 1 0 20332 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_215
timestamp 1676037725
transform 1 0 20884 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_222
timestamp 1676037725
transform 1 0 21528 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_234
timestamp 1676037725
transform 1 0 22632 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_246
timestamp 1676037725
transform 1 0 23736 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1676037725
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_264
timestamp 1676037725
transform 1 0 25392 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_275
timestamp 1676037725
transform 1 0 26404 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_282
timestamp 1676037725
transform 1 0 27048 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_294
timestamp 1676037725
transform 1 0 28152 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_303
timestamp 1676037725
transform 1 0 28980 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1676037725
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_309
timestamp 1676037725
transform 1 0 29532 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_315
timestamp 1676037725
transform 1 0 30084 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_323
timestamp 1676037725
transform 1 0 30820 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_329
timestamp 1676037725
transform 1 0 31372 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_333
timestamp 1676037725
transform 1 0 31740 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_341
timestamp 1676037725
transform 1 0 32476 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_362
timestamp 1676037725
transform 1 0 34408 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_365
timestamp 1676037725
transform 1 0 34684 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_371
timestamp 1676037725
transform 1 0 35236 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_375
timestamp 1676037725
transform 1 0 35604 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_383
timestamp 1676037725
transform 1 0 36340 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_391
timestamp 1676037725
transform 1 0 37076 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_399
timestamp 1676037725
transform 1 0 37812 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_405
timestamp 1676037725
transform 1 0 38364 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_410
timestamp 1676037725
transform 1 0 38824 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_418
timestamp 1676037725
transform 1 0 39560 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_421
timestamp 1676037725
transform 1 0 39836 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_428
timestamp 1676037725
transform 1 0 40480 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_28_438
timestamp 1676037725
transform 1 0 41400 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_446
timestamp 1676037725
transform 1 0 42136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_464
timestamp 1676037725
transform 1 0 43792 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_474
timestamp 1676037725
transform 1 0 44712 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_477
timestamp 1676037725
transform 1 0 44988 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_485
timestamp 1676037725
transform 1 0 45724 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_493
timestamp 1676037725
transform 1 0 46460 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_501
timestamp 1676037725
transform 1 0 47196 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_517
timestamp 1676037725
transform 1 0 48668 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_524
timestamp 1676037725
transform 1 0 49312 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_28_533
timestamp 1676037725
transform 1 0 50140 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_545
timestamp 1676037725
transform 1 0 51244 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_551
timestamp 1676037725
transform 1 0 51796 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_555
timestamp 1676037725
transform 1 0 52164 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_567
timestamp 1676037725
transform 1 0 53268 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_579
timestamp 1676037725
transform 1 0 54372 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_587
timestamp 1676037725
transform 1 0 55108 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_589
timestamp 1676037725
transform 1 0 55292 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_597
timestamp 1676037725
transform 1 0 56028 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_602
timestamp 1676037725
transform 1 0 56488 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_28_622
timestamp 1676037725
transform 1 0 58328 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1676037725
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_11
timestamp 1676037725
transform 1 0 2116 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1676037725
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1676037725
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1676037725
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1676037725
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1676037725
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1676037725
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1676037725
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1676037725
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1676037725
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1676037725
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1676037725
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1676037725
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1676037725
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1676037725
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1676037725
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1676037725
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1676037725
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1676037725
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1676037725
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1676037725
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_205
timestamp 1676037725
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1676037725
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1676037725
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1676037725
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_237
timestamp 1676037725
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_249
timestamp 1676037725
transform 1 0 24012 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_257
timestamp 1676037725
transform 1 0 24748 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_261
timestamp 1676037725
transform 1 0 25116 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_268
timestamp 1676037725
transform 1 0 25760 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_276
timestamp 1676037725
transform 1 0 26496 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1676037725
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_293
timestamp 1676037725
transform 1 0 28060 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_299
timestamp 1676037725
transform 1 0 28612 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_304
timestamp 1676037725
transform 1 0 29072 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_312
timestamp 1676037725
transform 1 0 29808 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_319
timestamp 1676037725
transform 1 0 30452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_331
timestamp 1676037725
transform 1 0 31556 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1676037725
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_337
timestamp 1676037725
transform 1 0 32108 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_344
timestamp 1676037725
transform 1 0 32752 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_352
timestamp 1676037725
transform 1 0 33488 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_360
timestamp 1676037725
transform 1 0 34224 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_364
timestamp 1676037725
transform 1 0 34592 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_369
timestamp 1676037725
transform 1 0 35052 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_375
timestamp 1676037725
transform 1 0 35604 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_382
timestamp 1676037725
transform 1 0 36248 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_390
timestamp 1676037725
transform 1 0 36984 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_393
timestamp 1676037725
transform 1 0 37260 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_399
timestamp 1676037725
transform 1 0 37812 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_407
timestamp 1676037725
transform 1 0 38548 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_415
timestamp 1676037725
transform 1 0 39284 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_423
timestamp 1676037725
transform 1 0 40020 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_428
timestamp 1676037725
transform 1 0 40480 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_436
timestamp 1676037725
transform 1 0 41216 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_440
timestamp 1676037725
transform 1 0 41584 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_446
timestamp 1676037725
transform 1 0 42136 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_449
timestamp 1676037725
transform 1 0 42412 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_457
timestamp 1676037725
transform 1 0 43148 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_473
timestamp 1676037725
transform 1 0 44620 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_486
timestamp 1676037725
transform 1 0 45816 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_498
timestamp 1676037725
transform 1 0 46920 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_505
timestamp 1676037725
transform 1 0 47564 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_521
timestamp 1676037725
transform 1 0 49036 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_545
timestamp 1676037725
transform 1 0 51244 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_557
timestamp 1676037725
transform 1 0 52348 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_561
timestamp 1676037725
transform 1 0 52716 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_573
timestamp 1676037725
transform 1 0 53820 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_585
timestamp 1676037725
transform 1 0 54924 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_593
timestamp 1676037725
transform 1 0 55660 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_597
timestamp 1676037725
transform 1 0 56028 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_603
timestamp 1676037725
transform 1 0 56580 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_610
timestamp 1676037725
transform 1 0 57224 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_617
timestamp 1676037725
transform 1 0 57868 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_623
timestamp 1676037725
transform 1 0 58420 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1676037725
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_11
timestamp 1676037725
transform 1 0 2116 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_23
timestamp 1676037725
transform 1 0 3220 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1676037725
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1676037725
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1676037725
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1676037725
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1676037725
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1676037725
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1676037725
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1676037725
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1676037725
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1676037725
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1676037725
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1676037725
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1676037725
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1676037725
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1676037725
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1676037725
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1676037725
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1676037725
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1676037725
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1676037725
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_209
timestamp 1676037725
transform 1 0 20332 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_219
timestamp 1676037725
transform 1 0 21252 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_242
timestamp 1676037725
transform 1 0 23368 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1676037725
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1676037725
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_263
timestamp 1676037725
transform 1 0 25300 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_273
timestamp 1676037725
transform 1 0 26220 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_279
timestamp 1676037725
transform 1 0 26772 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_284
timestamp 1676037725
transform 1 0 27232 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_292
timestamp 1676037725
transform 1 0 27968 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_304
timestamp 1676037725
transform 1 0 29072 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_309
timestamp 1676037725
transform 1 0 29532 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_317
timestamp 1676037725
transform 1 0 30268 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_329
timestamp 1676037725
transform 1 0 31372 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_337
timestamp 1676037725
transform 1 0 32108 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_342
timestamp 1676037725
transform 1 0 32568 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_354
timestamp 1676037725
transform 1 0 33672 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_362
timestamp 1676037725
transform 1 0 34408 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_365
timestamp 1676037725
transform 1 0 34684 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_372
timestamp 1676037725
transform 1 0 35328 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_379
timestamp 1676037725
transform 1 0 35972 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_388
timestamp 1676037725
transform 1 0 36800 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_396
timestamp 1676037725
transform 1 0 37536 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_404
timestamp 1676037725
transform 1 0 38272 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_413
timestamp 1676037725
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1676037725
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_421
timestamp 1676037725
transform 1 0 39836 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_427
timestamp 1676037725
transform 1 0 40388 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_435
timestamp 1676037725
transform 1 0 41124 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_453
timestamp 1676037725
transform 1 0 42780 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_466
timestamp 1676037725
transform 1 0 43976 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_474
timestamp 1676037725
transform 1 0 44712 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_477
timestamp 1676037725
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_489
timestamp 1676037725
transform 1 0 46092 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_497
timestamp 1676037725
transform 1 0 46828 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_503
timestamp 1676037725
transform 1 0 47380 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_30_523
timestamp 1676037725
transform 1 0 49220 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_531
timestamp 1676037725
transform 1 0 49956 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_533
timestamp 1676037725
transform 1 0 50140 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_545
timestamp 1676037725
transform 1 0 51244 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_557
timestamp 1676037725
transform 1 0 52348 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_569
timestamp 1676037725
transform 1 0 53452 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_581
timestamp 1676037725
transform 1 0 54556 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_587
timestamp 1676037725
transform 1 0 55108 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_589
timestamp 1676037725
transform 1 0 55292 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_599
timestamp 1676037725
transform 1 0 56212 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_613
timestamp 1676037725
transform 1 0 57500 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_623
timestamp 1676037725
transform 1 0 58420 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1676037725
transform 1 0 1380 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_11
timestamp 1676037725
transform 1 0 2116 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_23
timestamp 1676037725
transform 1 0 3220 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_35
timestamp 1676037725
transform 1 0 4324 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_47
timestamp 1676037725
transform 1 0 5428 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1676037725
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1676037725
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1676037725
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1676037725
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1676037725
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1676037725
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1676037725
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1676037725
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1676037725
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1676037725
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1676037725
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1676037725
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1676037725
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1676037725
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1676037725
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_193
timestamp 1676037725
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_205
timestamp 1676037725
transform 1 0 19964 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_209
timestamp 1676037725
transform 1 0 20332 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_214
timestamp 1676037725
transform 1 0 20792 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1676037725
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1676037725
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_231
timestamp 1676037725
transform 1 0 22356 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_235
timestamp 1676037725
transform 1 0 22724 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_245
timestamp 1676037725
transform 1 0 23644 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_254
timestamp 1676037725
transform 1 0 24472 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_266
timestamp 1676037725
transform 1 0 25576 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_278
timestamp 1676037725
transform 1 0 26680 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_281
timestamp 1676037725
transform 1 0 26956 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_290
timestamp 1676037725
transform 1 0 27784 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_294
timestamp 1676037725
transform 1 0 28152 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_299
timestamp 1676037725
transform 1 0 28612 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_311
timestamp 1676037725
transform 1 0 29716 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_323
timestamp 1676037725
transform 1 0 30820 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1676037725
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1676037725
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_365
timestamp 1676037725
transform 1 0 34684 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_373
timestamp 1676037725
transform 1 0 35420 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_384
timestamp 1676037725
transform 1 0 36432 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_393
timestamp 1676037725
transform 1 0 37260 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_399
timestamp 1676037725
transform 1 0 37812 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_419
timestamp 1676037725
transform 1 0 39652 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_427
timestamp 1676037725
transform 1 0 40388 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_31_441
timestamp 1676037725
transform 1 0 41676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1676037725
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_449
timestamp 1676037725
transform 1 0 42412 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_455
timestamp 1676037725
transform 1 0 42964 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_463
timestamp 1676037725
transform 1 0 43700 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_469
timestamp 1676037725
transform 1 0 44252 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_489
timestamp 1676037725
transform 1 0 46092 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_493
timestamp 1676037725
transform 1 0 46460 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_502
timestamp 1676037725
transform 1 0 47288 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_505
timestamp 1676037725
transform 1 0 47564 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_529
timestamp 1676037725
transform 1 0 49772 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_536
timestamp 1676037725
transform 1 0 50416 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_548
timestamp 1676037725
transform 1 0 51520 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_552
timestamp 1676037725
transform 1 0 51888 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_556
timestamp 1676037725
transform 1 0 52256 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_561
timestamp 1676037725
transform 1 0 52716 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_579
timestamp 1676037725
transform 1 0 54372 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_591
timestamp 1676037725
transform 1 0 55476 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_610
timestamp 1676037725
transform 1 0 57224 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_617
timestamp 1676037725
transform 1 0 57868 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_623
timestamp 1676037725
transform 1 0 58420 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1676037725
transform 1 0 1380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_11
timestamp 1676037725
transform 1 0 2116 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_19
timestamp 1676037725
transform 1 0 2852 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1676037725
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1676037725
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1676037725
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1676037725
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1676037725
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1676037725
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1676037725
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1676037725
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1676037725
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1676037725
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1676037725
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1676037725
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1676037725
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1676037725
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1676037725
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1676037725
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_177
timestamp 1676037725
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1676037725
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1676037725
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1676037725
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1676037725
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_221
timestamp 1676037725
transform 1 0 21436 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_231
timestamp 1676037725
transform 1 0 22356 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_243
timestamp 1676037725
transform 1 0 23460 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1676037725
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_253
timestamp 1676037725
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_265
timestamp 1676037725
transform 1 0 25484 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_273
timestamp 1676037725
transform 1 0 26220 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_291
timestamp 1676037725
transform 1 0 27876 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_304
timestamp 1676037725
transform 1 0 29072 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_309
timestamp 1676037725
transform 1 0 29532 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_321
timestamp 1676037725
transform 1 0 30636 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_329
timestamp 1676037725
transform 1 0 31372 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_337
timestamp 1676037725
transform 1 0 32108 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_345
timestamp 1676037725
transform 1 0 32844 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_362
timestamp 1676037725
transform 1 0 34408 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_365
timestamp 1676037725
transform 1 0 34684 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_379
timestamp 1676037725
transform 1 0 35972 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_391
timestamp 1676037725
transform 1 0 37076 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_402
timestamp 1676037725
transform 1 0 38088 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_410
timestamp 1676037725
transform 1 0 38824 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_418
timestamp 1676037725
transform 1 0 39560 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_421
timestamp 1676037725
transform 1 0 39836 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_428
timestamp 1676037725
transform 1 0 40480 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_436
timestamp 1676037725
transform 1 0 41216 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_444
timestamp 1676037725
transform 1 0 41952 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_452
timestamp 1676037725
transform 1 0 42688 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_462
timestamp 1676037725
transform 1 0 43608 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_474
timestamp 1676037725
transform 1 0 44712 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_477
timestamp 1676037725
transform 1 0 44988 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_485
timestamp 1676037725
transform 1 0 45724 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_497
timestamp 1676037725
transform 1 0 46828 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_505
timestamp 1676037725
transform 1 0 47564 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_516
timestamp 1676037725
transform 1 0 48576 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_525
timestamp 1676037725
transform 1 0 49404 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_531
timestamp 1676037725
transform 1 0 49956 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_533
timestamp 1676037725
transform 1 0 50140 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_543
timestamp 1676037725
transform 1 0 51060 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_551
timestamp 1676037725
transform 1 0 51796 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_569
timestamp 1676037725
transform 1 0 53452 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_581
timestamp 1676037725
transform 1 0 54556 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_587
timestamp 1676037725
transform 1 0 55108 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_589
timestamp 1676037725
transform 1 0 55292 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_32_600
timestamp 1676037725
transform 1 0 56304 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_612
timestamp 1676037725
transform 1 0 57408 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_616
timestamp 1676037725
transform 1 0 57776 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_623
timestamp 1676037725
transform 1 0 58420 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1676037725
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_11
timestamp 1676037725
transform 1 0 2116 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_23
timestamp 1676037725
transform 1 0 3220 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_35
timestamp 1676037725
transform 1 0 4324 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_47
timestamp 1676037725
transform 1 0 5428 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1676037725
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1676037725
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1676037725
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1676037725
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1676037725
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1676037725
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1676037725
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1676037725
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1676037725
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1676037725
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1676037725
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1676037725
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1676037725
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1676037725
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1676037725
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_193
timestamp 1676037725
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_205
timestamp 1676037725
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1676037725
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1676037725
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1676037725
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_237
timestamp 1676037725
transform 1 0 22908 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_33_259
timestamp 1676037725
transform 1 0 24932 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_278
timestamp 1676037725
transform 1 0 26680 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_281
timestamp 1676037725
transform 1 0 26956 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_287
timestamp 1676037725
transform 1 0 27508 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_308
timestamp 1676037725
transform 1 0 29440 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_33_333
timestamp 1676037725
transform 1 0 31740 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_337
timestamp 1676037725
transform 1 0 32108 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_341
timestamp 1676037725
transform 1 0 32476 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_346
timestamp 1676037725
transform 1 0 32936 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_367
timestamp 1676037725
transform 1 0 34868 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_375
timestamp 1676037725
transform 1 0 35604 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_383
timestamp 1676037725
transform 1 0 36340 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_390
timestamp 1676037725
transform 1 0 36984 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_393
timestamp 1676037725
transform 1 0 37260 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_399
timestamp 1676037725
transform 1 0 37812 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_407
timestamp 1676037725
transform 1 0 38548 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_416
timestamp 1676037725
transform 1 0 39376 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_437
timestamp 1676037725
transform 1 0 41308 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_445
timestamp 1676037725
transform 1 0 42044 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_449
timestamp 1676037725
transform 1 0 42412 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_454
timestamp 1676037725
transform 1 0 42872 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_475
timestamp 1676037725
transform 1 0 44804 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_483
timestamp 1676037725
transform 1 0 45540 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_491
timestamp 1676037725
transform 1 0 46276 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1676037725
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_505
timestamp 1676037725
transform 1 0 47564 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_515
timestamp 1676037725
transform 1 0 48484 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_519
timestamp 1676037725
transform 1 0 48852 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_528
timestamp 1676037725
transform 1 0 49680 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_548
timestamp 1676037725
transform 1 0 51520 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_554
timestamp 1676037725
transform 1 0 52072 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_558
timestamp 1676037725
transform 1 0 52440 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_561
timestamp 1676037725
transform 1 0 52716 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_571
timestamp 1676037725
transform 1 0 53636 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_583
timestamp 1676037725
transform 1 0 54740 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_603
timestamp 1676037725
transform 1 0 56580 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_615
timestamp 1676037725
transform 1 0 57684 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_617
timestamp 1676037725
transform 1 0 57868 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_623
timestamp 1676037725
transform 1 0 58420 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1676037725
transform 1 0 1380 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_11
timestamp 1676037725
transform 1 0 2116 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_23
timestamp 1676037725
transform 1 0 3220 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1676037725
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1676037725
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1676037725
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1676037725
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1676037725
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1676037725
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1676037725
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1676037725
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1676037725
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1676037725
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1676037725
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1676037725
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1676037725
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1676037725
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1676037725
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1676037725
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1676037725
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1676037725
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1676037725
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1676037725
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_209
timestamp 1676037725
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_221
timestamp 1676037725
transform 1 0 21436 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_225
timestamp 1676037725
transform 1 0 21804 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_233
timestamp 1676037725
transform 1 0 22540 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_237
timestamp 1676037725
transform 1 0 22908 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_242
timestamp 1676037725
transform 1 0 23368 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_250
timestamp 1676037725
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_253
timestamp 1676037725
transform 1 0 24380 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_261
timestamp 1676037725
transform 1 0 25116 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_266
timestamp 1676037725
transform 1 0 25576 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_287
timestamp 1676037725
transform 1 0 27508 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_294
timestamp 1676037725
transform 1 0 28152 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_306
timestamp 1676037725
transform 1 0 29256 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_309
timestamp 1676037725
transform 1 0 29532 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_328
timestamp 1676037725
transform 1 0 31280 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_348
timestamp 1676037725
transform 1 0 33120 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_356
timestamp 1676037725
transform 1 0 33856 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_365
timestamp 1676037725
transform 1 0 34684 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_383
timestamp 1676037725
transform 1 0 36340 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_391
timestamp 1676037725
transform 1 0 37076 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_399
timestamp 1676037725
transform 1 0 37812 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_407
timestamp 1676037725
transform 1 0 38548 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_415
timestamp 1676037725
transform 1 0 39284 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 1676037725
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_421
timestamp 1676037725
transform 1 0 39836 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_427
timestamp 1676037725
transform 1 0 40388 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_435
timestamp 1676037725
transform 1 0 41124 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_443
timestamp 1676037725
transform 1 0 41860 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_34_456
timestamp 1676037725
transform 1 0 43056 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_34_470
timestamp 1676037725
transform 1 0 44344 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_34_477
timestamp 1676037725
transform 1 0 44988 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_487
timestamp 1676037725
transform 1 0 45908 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_499
timestamp 1676037725
transform 1 0 47012 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_511
timestamp 1676037725
transform 1 0 48116 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_530
timestamp 1676037725
transform 1 0 49864 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_533
timestamp 1676037725
transform 1 0 50140 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_545
timestamp 1676037725
transform 1 0 51244 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_557
timestamp 1676037725
transform 1 0 52348 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_569
timestamp 1676037725
transform 1 0 53452 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_581
timestamp 1676037725
transform 1 0 54556 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_587
timestamp 1676037725
transform 1 0 55108 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_589
timestamp 1676037725
transform 1 0 55292 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_593
timestamp 1676037725
transform 1 0 55660 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_602
timestamp 1676037725
transform 1 0 56488 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_622
timestamp 1676037725
transform 1 0 58328 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1676037725
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_11
timestamp 1676037725
transform 1 0 2116 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_23
timestamp 1676037725
transform 1 0 3220 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_35
timestamp 1676037725
transform 1 0 4324 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_47
timestamp 1676037725
transform 1 0 5428 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1676037725
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1676037725
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1676037725
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1676037725
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1676037725
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1676037725
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1676037725
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1676037725
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1676037725
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1676037725
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 1676037725
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1676037725
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1676037725
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1676037725
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1676037725
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_193
timestamp 1676037725
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_205
timestamp 1676037725
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1676037725
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1676037725
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1676037725
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_236
timestamp 1676037725
transform 1 0 22816 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_251
timestamp 1676037725
transform 1 0 24196 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_261
timestamp 1676037725
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_273
timestamp 1676037725
transform 1 0 26220 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_278
timestamp 1676037725
transform 1 0 26680 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_281
timestamp 1676037725
transform 1 0 26956 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_289
timestamp 1676037725
transform 1 0 27692 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_296
timestamp 1676037725
transform 1 0 28336 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_307
timestamp 1676037725
transform 1 0 29348 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_318
timestamp 1676037725
transform 1 0 30360 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_331
timestamp 1676037725
transform 1 0 31556 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1676037725
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_337
timestamp 1676037725
transform 1 0 32108 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_343
timestamp 1676037725
transform 1 0 32660 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_363
timestamp 1676037725
transform 1 0 34500 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_373
timestamp 1676037725
transform 1 0 35420 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_381
timestamp 1676037725
transform 1 0 36156 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_35_389
timestamp 1676037725
transform 1 0 36892 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_393
timestamp 1676037725
transform 1 0 37260 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_399
timestamp 1676037725
transform 1 0 37812 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_407
timestamp 1676037725
transform 1 0 38548 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_35_430
timestamp 1676037725
transform 1 0 40664 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_436
timestamp 1676037725
transform 1 0 41216 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_442
timestamp 1676037725
transform 1 0 41768 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_35_449
timestamp 1676037725
transform 1 0 42412 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_468
timestamp 1676037725
transform 1 0 44160 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_477
timestamp 1676037725
transform 1 0 44988 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_492
timestamp 1676037725
transform 1 0 46368 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_505
timestamp 1676037725
transform 1 0 47564 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_517
timestamp 1676037725
transform 1 0 48668 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_521
timestamp 1676037725
transform 1 0 49036 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_533
timestamp 1676037725
transform 1 0 50140 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_545
timestamp 1676037725
transform 1 0 51244 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_557
timestamp 1676037725
transform 1 0 52348 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_561
timestamp 1676037725
transform 1 0 52716 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_579
timestamp 1676037725
transform 1 0 54372 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_587
timestamp 1676037725
transform 1 0 55108 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_594
timestamp 1676037725
transform 1 0 55752 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_614
timestamp 1676037725
transform 1 0 57592 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_617
timestamp 1676037725
transform 1 0 57868 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_623
timestamp 1676037725
transform 1 0 58420 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_3
timestamp 1676037725
transform 1 0 1380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_11
timestamp 1676037725
transform 1 0 2116 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_20
timestamp 1676037725
transform 1 0 2944 0 1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1676037725
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1676037725
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1676037725
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1676037725
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1676037725
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1676037725
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1676037725
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1676037725
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1676037725
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1676037725
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1676037725
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1676037725
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1676037725
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1676037725
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_165
timestamp 1676037725
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_177
timestamp 1676037725
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1676037725
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1676037725
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1676037725
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_209
timestamp 1676037725
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_221
timestamp 1676037725
transform 1 0 21436 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_225
timestamp 1676037725
transform 1 0 21804 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_233
timestamp 1676037725
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1676037725
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1676037725
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1676037725
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_265
timestamp 1676037725
transform 1 0 25484 0 1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_36_277
timestamp 1676037725
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_289
timestamp 1676037725
transform 1 0 27692 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_36_296
timestamp 1676037725
transform 1 0 28336 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_36_306
timestamp 1676037725
transform 1 0 29256 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_309
timestamp 1676037725
transform 1 0 29532 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_321
timestamp 1676037725
transform 1 0 30636 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_332
timestamp 1676037725
transform 1 0 31648 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_340
timestamp 1676037725
transform 1 0 32384 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_348
timestamp 1676037725
transform 1 0 33120 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_356
timestamp 1676037725
transform 1 0 33856 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_36_365
timestamp 1676037725
transform 1 0 34684 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_381
timestamp 1676037725
transform 1 0 36156 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_389
timestamp 1676037725
transform 1 0 36892 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_396
timestamp 1676037725
transform 1 0 37536 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_405
timestamp 1676037725
transform 1 0 38364 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_417
timestamp 1676037725
transform 1 0 39468 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_421
timestamp 1676037725
transform 1 0 39836 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_427
timestamp 1676037725
transform 1 0 40388 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_36_438
timestamp 1676037725
transform 1 0 41400 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_444
timestamp 1676037725
transform 1 0 41952 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_464
timestamp 1676037725
transform 1 0 43792 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_473
timestamp 1676037725
transform 1 0 44620 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_477
timestamp 1676037725
transform 1 0 44988 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_496
timestamp 1676037725
transform 1 0 46736 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_509
timestamp 1676037725
transform 1 0 47932 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_36_520
timestamp 1676037725
transform 1 0 48944 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_533
timestamp 1676037725
transform 1 0 50140 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_545
timestamp 1676037725
transform 1 0 51244 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_549
timestamp 1676037725
transform 1 0 51612 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_566
timestamp 1676037725
transform 1 0 53176 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_577
timestamp 1676037725
transform 1 0 54188 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_585
timestamp 1676037725
transform 1 0 54924 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_36_589
timestamp 1676037725
transform 1 0 55292 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_611
timestamp 1676037725
transform 1 0 57316 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_622
timestamp 1676037725
transform 1 0 58328 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_37_3
timestamp 1676037725
transform 1 0 1380 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_37_17
timestamp 1676037725
transform 1 0 2668 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_29
timestamp 1676037725
transform 1 0 3772 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_41
timestamp 1676037725
transform 1 0 4876 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_53
timestamp 1676037725
transform 1 0 5980 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1676037725
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1676037725
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1676037725
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1676037725
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1676037725
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1676037725
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1676037725
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1676037725
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1676037725
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1676037725
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1676037725
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1676037725
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1676037725
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_181
timestamp 1676037725
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_193
timestamp 1676037725
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_205
timestamp 1676037725
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1676037725
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1676037725
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_225
timestamp 1676037725
transform 1 0 21804 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_37_251
timestamp 1676037725
transform 1 0 24196 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_263
timestamp 1676037725
transform 1 0 25300 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_275
timestamp 1676037725
transform 1 0 26404 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1676037725
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1676037725
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_293
timestamp 1676037725
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_305
timestamp 1676037725
transform 1 0 29164 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_313
timestamp 1676037725
transform 1 0 29900 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_321
timestamp 1676037725
transform 1 0 30636 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_331
timestamp 1676037725
transform 1 0 31556 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1676037725
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_337
timestamp 1676037725
transform 1 0 32108 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_341
timestamp 1676037725
transform 1 0 32476 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_349
timestamp 1676037725
transform 1 0 33212 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_357
timestamp 1676037725
transform 1 0 33948 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_370
timestamp 1676037725
transform 1 0 35144 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_390
timestamp 1676037725
transform 1 0 36984 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_393
timestamp 1676037725
transform 1 0 37260 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_399
timestamp 1676037725
transform 1 0 37812 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_405
timestamp 1676037725
transform 1 0 38364 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_422
timestamp 1676037725
transform 1 0 39928 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_430
timestamp 1676037725
transform 1 0 40664 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_436
timestamp 1676037725
transform 1 0 41216 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_37_445
timestamp 1676037725
transform 1 0 42044 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_449
timestamp 1676037725
transform 1 0 42412 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_455
timestamp 1676037725
transform 1 0 42964 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_463
timestamp 1676037725
transform 1 0 43700 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_483
timestamp 1676037725
transform 1 0 45540 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_489
timestamp 1676037725
transform 1 0 46092 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_499
timestamp 1676037725
transform 1 0 47012 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 1676037725
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_505
timestamp 1676037725
transform 1 0 47564 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_513
timestamp 1676037725
transform 1 0 48300 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_531
timestamp 1676037725
transform 1 0 49956 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_550
timestamp 1676037725
transform 1 0 51704 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_558
timestamp 1676037725
transform 1 0 52440 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_561
timestamp 1676037725
transform 1 0 52716 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_568
timestamp 1676037725
transform 1 0 53360 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_580
timestamp 1676037725
transform 1 0 54464 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_592
timestamp 1676037725
transform 1 0 55568 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_37_607
timestamp 1676037725
transform 1 0 56948 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_615
timestamp 1676037725
transform 1 0 57684 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_617
timestamp 1676037725
transform 1 0 57868 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_623
timestamp 1676037725
transform 1 0 58420 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_3
timestamp 1676037725
transform 1 0 1380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_11
timestamp 1676037725
transform 1 0 2116 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_20
timestamp 1676037725
transform 1 0 2944 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1676037725
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1676037725
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1676037725
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1676037725
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1676037725
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1676037725
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1676037725
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1676037725
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1676037725
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 1676037725
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1676037725
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1676037725
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1676037725
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1676037725
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_165
timestamp 1676037725
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_177
timestamp 1676037725
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1676037725
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1676037725
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1676037725
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_209
timestamp 1676037725
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_221
timestamp 1676037725
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_233
timestamp 1676037725
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1676037725
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1676037725
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1676037725
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 1676037725
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_277
timestamp 1676037725
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_289
timestamp 1676037725
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1676037725
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1676037725
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_309
timestamp 1676037725
transform 1 0 29532 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_315
timestamp 1676037725
transform 1 0 30084 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_322
timestamp 1676037725
transform 1 0 30728 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_334
timestamp 1676037725
transform 1 0 31832 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_346
timestamp 1676037725
transform 1 0 32936 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_353
timestamp 1676037725
transform 1 0 33580 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_38_361
timestamp 1676037725
transform 1 0 34316 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_365
timestamp 1676037725
transform 1 0 34684 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_371
timestamp 1676037725
transform 1 0 35236 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_377
timestamp 1676037725
transform 1 0 35788 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_382
timestamp 1676037725
transform 1 0 36248 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_395
timestamp 1676037725
transform 1 0 37444 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_403
timestamp 1676037725
transform 1 0 38180 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_409
timestamp 1676037725
transform 1 0 38732 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_418
timestamp 1676037725
transform 1 0 39560 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_421
timestamp 1676037725
transform 1 0 39836 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_427
timestamp 1676037725
transform 1 0 40388 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_435
timestamp 1676037725
transform 1 0 41124 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_439
timestamp 1676037725
transform 1 0 41492 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_448
timestamp 1676037725
transform 1 0 42320 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_456
timestamp 1676037725
transform 1 0 43056 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_468
timestamp 1676037725
transform 1 0 44160 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_38_477
timestamp 1676037725
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_489
timestamp 1676037725
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_501
timestamp 1676037725
transform 1 0 47196 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_509
timestamp 1676037725
transform 1 0 47932 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_519
timestamp 1676037725
transform 1 0 48852 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_531
timestamp 1676037725
transform 1 0 49956 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_533
timestamp 1676037725
transform 1 0 50140 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_545
timestamp 1676037725
transform 1 0 51244 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_553
timestamp 1676037725
transform 1 0 51980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_565
timestamp 1676037725
transform 1 0 53084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_577
timestamp 1676037725
transform 1 0 54188 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_585
timestamp 1676037725
transform 1 0 54924 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_589
timestamp 1676037725
transform 1 0 55292 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_597
timestamp 1676037725
transform 1 0 56028 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_603
timestamp 1676037725
transform 1 0 56580 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_613
timestamp 1676037725
transform 1 0 57500 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_623
timestamp 1676037725
transform 1 0 58420 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_3
timestamp 1676037725
transform 1 0 1380 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_11
timestamp 1676037725
transform 1 0 2116 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_23
timestamp 1676037725
transform 1 0 3220 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_35
timestamp 1676037725
transform 1 0 4324 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_47
timestamp 1676037725
transform 1 0 5428 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1676037725
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1676037725
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1676037725
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1676037725
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1676037725
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1676037725
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1676037725
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1676037725
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1676037725
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1676037725
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_149
timestamp 1676037725
transform 1 0 14812 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_157
timestamp 1676037725
transform 1 0 15548 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_164
timestamp 1676037725
transform 1 0 16192 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1676037725
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1676037725
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_193
timestamp 1676037725
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_205
timestamp 1676037725
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1676037725
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1676037725
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1676037725
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_237
timestamp 1676037725
transform 1 0 22908 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_257
timestamp 1676037725
transform 1 0 24748 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_269
timestamp 1676037725
transform 1 0 25852 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_277
timestamp 1676037725
transform 1 0 26588 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1676037725
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_293
timestamp 1676037725
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_305
timestamp 1676037725
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_317
timestamp 1676037725
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1676037725
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1676037725
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1676037725
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_349
timestamp 1676037725
transform 1 0 33212 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_357
timestamp 1676037725
transform 1 0 33948 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_362
timestamp 1676037725
transform 1 0 34408 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_374
timestamp 1676037725
transform 1 0 35512 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_390
timestamp 1676037725
transform 1 0 36984 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1676037725
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_409
timestamp 1676037725
transform 1 0 38732 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_417
timestamp 1676037725
transform 1 0 39468 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_429
timestamp 1676037725
transform 1 0 40572 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_437
timestamp 1676037725
transform 1 0 41308 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_444
timestamp 1676037725
transform 1 0 41952 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_449
timestamp 1676037725
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_461
timestamp 1676037725
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_473
timestamp 1676037725
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_485
timestamp 1676037725
transform 1 0 45724 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_497
timestamp 1676037725
transform 1 0 46828 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 1676037725
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_505
timestamp 1676037725
transform 1 0 47564 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_517
timestamp 1676037725
transform 1 0 48668 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_529
timestamp 1676037725
transform 1 0 49772 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_541
timestamp 1676037725
transform 1 0 50876 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_553
timestamp 1676037725
transform 1 0 51980 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_559
timestamp 1676037725
transform 1 0 52532 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_561
timestamp 1676037725
transform 1 0 52716 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_573
timestamp 1676037725
transform 1 0 53820 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_585
timestamp 1676037725
transform 1 0 54924 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_597
timestamp 1676037725
transform 1 0 56028 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_609
timestamp 1676037725
transform 1 0 57132 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_615
timestamp 1676037725
transform 1 0 57684 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_617
timestamp 1676037725
transform 1 0 57868 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_623
timestamp 1676037725
transform 1 0 58420 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_3
timestamp 1676037725
transform 1 0 1380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_11
timestamp 1676037725
transform 1 0 2116 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_20
timestamp 1676037725
transform 1 0 2944 0 1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1676037725
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1676037725
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1676037725
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1676037725
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1676037725
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1676037725
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1676037725
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1676037725
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1676037725
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1676037725
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1676037725
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1676037725
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1676037725
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1676037725
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_165
timestamp 1676037725
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_177
timestamp 1676037725
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1676037725
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1676037725
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1676037725
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_209
timestamp 1676037725
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_221
timestamp 1676037725
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_233
timestamp 1676037725
transform 1 0 22540 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_250
timestamp 1676037725
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1676037725
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1676037725
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_277
timestamp 1676037725
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_289
timestamp 1676037725
transform 1 0 27692 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_293
timestamp 1676037725
transform 1 0 28060 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_302
timestamp 1676037725
transform 1 0 28888 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_40_309
timestamp 1676037725
transform 1 0 29532 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_319
timestamp 1676037725
transform 1 0 30452 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_331
timestamp 1676037725
transform 1 0 31556 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_343
timestamp 1676037725
transform 1 0 32660 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_355
timestamp 1676037725
transform 1 0 33764 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1676037725
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1676037725
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1676037725
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_389
timestamp 1676037725
transform 1 0 36892 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_400
timestamp 1676037725
transform 1 0 37904 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_412
timestamp 1676037725
transform 1 0 39008 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_40_421
timestamp 1676037725
transform 1 0 39836 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_429
timestamp 1676037725
transform 1 0 40572 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_435
timestamp 1676037725
transform 1 0 41124 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_447
timestamp 1676037725
transform 1 0 42228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_459
timestamp 1676037725
transform 1 0 43332 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_471
timestamp 1676037725
transform 1 0 44436 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1676037725
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_477
timestamp 1676037725
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_489
timestamp 1676037725
transform 1 0 46092 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_497
timestamp 1676037725
transform 1 0 46828 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_508
timestamp 1676037725
transform 1 0 47840 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_520
timestamp 1676037725
transform 1 0 48944 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_533
timestamp 1676037725
transform 1 0 50140 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_545
timestamp 1676037725
transform 1 0 51244 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_557
timestamp 1676037725
transform 1 0 52348 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_569
timestamp 1676037725
transform 1 0 53452 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_581
timestamp 1676037725
transform 1 0 54556 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_587
timestamp 1676037725
transform 1 0 55108 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_589
timestamp 1676037725
transform 1 0 55292 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_601
timestamp 1676037725
transform 1 0 56396 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_613
timestamp 1676037725
transform 1 0 57500 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_623
timestamp 1676037725
transform 1 0 58420 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_3
timestamp 1676037725
transform 1 0 1380 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_11
timestamp 1676037725
transform 1 0 2116 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_20
timestamp 1676037725
transform 1 0 2944 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_32
timestamp 1676037725
transform 1 0 4048 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_44
timestamp 1676037725
transform 1 0 5152 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1676037725
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1676037725
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1676037725
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1676037725
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1676037725
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1676037725
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1676037725
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1676037725
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1676037725
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1676037725
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1676037725
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1676037725
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1676037725
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1676037725
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_193
timestamp 1676037725
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_205
timestamp 1676037725
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1676037725
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1676037725
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_225
timestamp 1676037725
transform 1 0 21804 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_234
timestamp 1676037725
transform 1 0 22632 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_257
timestamp 1676037725
transform 1 0 24748 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_270
timestamp 1676037725
transform 1 0 25944 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_278
timestamp 1676037725
transform 1 0 26680 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_281
timestamp 1676037725
transform 1 0 26956 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_41_294
timestamp 1676037725
transform 1 0 28152 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_41_320
timestamp 1676037725
transform 1 0 30544 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_332
timestamp 1676037725
transform 1 0 31648 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1676037725
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1676037725
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_361
timestamp 1676037725
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_373
timestamp 1676037725
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1676037725
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1676037725
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_393
timestamp 1676037725
transform 1 0 37260 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_402
timestamp 1676037725
transform 1 0 38088 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_414
timestamp 1676037725
transform 1 0 39192 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_426
timestamp 1676037725
transform 1 0 40296 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_438
timestamp 1676037725
transform 1 0 41400 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_446
timestamp 1676037725
transform 1 0 42136 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_449
timestamp 1676037725
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_461
timestamp 1676037725
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_473
timestamp 1676037725
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_485
timestamp 1676037725
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_497
timestamp 1676037725
transform 1 0 46828 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_503
timestamp 1676037725
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_505
timestamp 1676037725
transform 1 0 47564 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_514
timestamp 1676037725
transform 1 0 48392 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_526
timestamp 1676037725
transform 1 0 49496 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_538
timestamp 1676037725
transform 1 0 50600 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_550
timestamp 1676037725
transform 1 0 51704 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_558
timestamp 1676037725
transform 1 0 52440 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_561
timestamp 1676037725
transform 1 0 52716 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_573
timestamp 1676037725
transform 1 0 53820 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_585
timestamp 1676037725
transform 1 0 54924 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_597
timestamp 1676037725
transform 1 0 56028 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_609
timestamp 1676037725
transform 1 0 57132 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_615
timestamp 1676037725
transform 1 0 57684 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_617
timestamp 1676037725
transform 1 0 57868 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_623
timestamp 1676037725
transform 1 0 58420 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_3
timestamp 1676037725
transform 1 0 1380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_11
timestamp 1676037725
transform 1 0 2116 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_20
timestamp 1676037725
transform 1 0 2944 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1676037725
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1676037725
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1676037725
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1676037725
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1676037725
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1676037725
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1676037725
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1676037725
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1676037725
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1676037725
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1676037725
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1676037725
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1676037725
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1676037725
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_165
timestamp 1676037725
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_177
timestamp 1676037725
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1676037725
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1676037725
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1676037725
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_209
timestamp 1676037725
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_221
timestamp 1676037725
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_233
timestamp 1676037725
transform 1 0 22540 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_244
timestamp 1676037725
transform 1 0 23552 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_253
timestamp 1676037725
transform 1 0 24380 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_264
timestamp 1676037725
transform 1 0 25392 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_276
timestamp 1676037725
transform 1 0 26496 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_282
timestamp 1676037725
transform 1 0 27048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_290
timestamp 1676037725
transform 1 0 27784 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_303
timestamp 1676037725
transform 1 0 28980 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1676037725
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_309
timestamp 1676037725
transform 1 0 29532 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_331
timestamp 1676037725
transform 1 0 31556 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_343
timestamp 1676037725
transform 1 0 32660 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_355
timestamp 1676037725
transform 1 0 33764 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1676037725
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1676037725
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_377
timestamp 1676037725
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_389
timestamp 1676037725
transform 1 0 36892 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_401
timestamp 1676037725
transform 1 0 37996 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_413
timestamp 1676037725
transform 1 0 39100 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_419
timestamp 1676037725
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_421
timestamp 1676037725
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_433
timestamp 1676037725
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_445
timestamp 1676037725
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_457
timestamp 1676037725
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 1676037725
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1676037725
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_477
timestamp 1676037725
transform 1 0 44988 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_485
timestamp 1676037725
transform 1 0 45724 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_496
timestamp 1676037725
transform 1 0 46736 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_508
timestamp 1676037725
transform 1 0 47840 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_519
timestamp 1676037725
transform 1 0 48852 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_531
timestamp 1676037725
transform 1 0 49956 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_533
timestamp 1676037725
transform 1 0 50140 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_545
timestamp 1676037725
transform 1 0 51244 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_557
timestamp 1676037725
transform 1 0 52348 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_569
timestamp 1676037725
transform 1 0 53452 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_581
timestamp 1676037725
transform 1 0 54556 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_587
timestamp 1676037725
transform 1 0 55108 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_589
timestamp 1676037725
transform 1 0 55292 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_601
timestamp 1676037725
transform 1 0 56396 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_613
timestamp 1676037725
transform 1 0 57500 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_623
timestamp 1676037725
transform 1 0 58420 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_3
timestamp 1676037725
transform 1 0 1380 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_11
timestamp 1676037725
transform 1 0 2116 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_23
timestamp 1676037725
transform 1 0 3220 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_35
timestamp 1676037725
transform 1 0 4324 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_47
timestamp 1676037725
transform 1 0 5428 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1676037725
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1676037725
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1676037725
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1676037725
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1676037725
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1676037725
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1676037725
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1676037725
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1676037725
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1676037725
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1676037725
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1676037725
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1676037725
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1676037725
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1676037725
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_193
timestamp 1676037725
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_205
timestamp 1676037725
transform 1 0 19964 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_213
timestamp 1676037725
transform 1 0 20700 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_222
timestamp 1676037725
transform 1 0 21528 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_225
timestamp 1676037725
transform 1 0 21804 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_233
timestamp 1676037725
transform 1 0 22540 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_249
timestamp 1676037725
transform 1 0 24012 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_257
timestamp 1676037725
transform 1 0 24748 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_269
timestamp 1676037725
transform 1 0 25852 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_277
timestamp 1676037725
transform 1 0 26588 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_281
timestamp 1676037725
transform 1 0 26956 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_289
timestamp 1676037725
transform 1 0 27692 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_302
timestamp 1676037725
transform 1 0 28888 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_314
timestamp 1676037725
transform 1 0 29992 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_324
timestamp 1676037725
transform 1 0 30912 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1676037725
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1676037725
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_361
timestamp 1676037725
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_373
timestamp 1676037725
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1676037725
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1676037725
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_393
timestamp 1676037725
transform 1 0 37260 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_403
timestamp 1676037725
transform 1 0 38180 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_413
timestamp 1676037725
transform 1 0 39100 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_425
timestamp 1676037725
transform 1 0 40204 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_437
timestamp 1676037725
transform 1 0 41308 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_445
timestamp 1676037725
transform 1 0 42044 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_43_449
timestamp 1676037725
transform 1 0 42412 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_457
timestamp 1676037725
transform 1 0 43148 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_467
timestamp 1676037725
transform 1 0 44068 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_479
timestamp 1676037725
transform 1 0 45172 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_491
timestamp 1676037725
transform 1 0 46276 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1676037725
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_505
timestamp 1676037725
transform 1 0 47564 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_517
timestamp 1676037725
transform 1 0 48668 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_529
timestamp 1676037725
transform 1 0 49772 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_541
timestamp 1676037725
transform 1 0 50876 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_553
timestamp 1676037725
transform 1 0 51980 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_559
timestamp 1676037725
transform 1 0 52532 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_561
timestamp 1676037725
transform 1 0 52716 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_573
timestamp 1676037725
transform 1 0 53820 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_585
timestamp 1676037725
transform 1 0 54924 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_597
timestamp 1676037725
transform 1 0 56028 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_609
timestamp 1676037725
transform 1 0 57132 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_615
timestamp 1676037725
transform 1 0 57684 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_617
timestamp 1676037725
transform 1 0 57868 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_623
timestamp 1676037725
transform 1 0 58420 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_3
timestamp 1676037725
transform 1 0 1380 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_11
timestamp 1676037725
transform 1 0 2116 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_23
timestamp 1676037725
transform 1 0 3220 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1676037725
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1676037725
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1676037725
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1676037725
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1676037725
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1676037725
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1676037725
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1676037725
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1676037725
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1676037725
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1676037725
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1676037725
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1676037725
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1676037725
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1676037725
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1676037725
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_177
timestamp 1676037725
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1676037725
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1676037725
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1676037725
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_209
timestamp 1676037725
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_221
timestamp 1676037725
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_233
timestamp 1676037725
transform 1 0 22540 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1676037725
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1676037725
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_253
timestamp 1676037725
transform 1 0 24380 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_259
timestamp 1676037725
transform 1 0 24932 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_267
timestamp 1676037725
transform 1 0 25668 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_273
timestamp 1676037725
transform 1 0 26220 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_281
timestamp 1676037725
transform 1 0 26956 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1676037725
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1676037725
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_309
timestamp 1676037725
transform 1 0 29532 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_318
timestamp 1676037725
transform 1 0 30360 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_322
timestamp 1676037725
transform 1 0 30728 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_44_337
timestamp 1676037725
transform 1 0 32108 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_349
timestamp 1676037725
transform 1 0 33212 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_361
timestamp 1676037725
transform 1 0 34316 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1676037725
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_377
timestamp 1676037725
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_389
timestamp 1676037725
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_401
timestamp 1676037725
transform 1 0 37996 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_413
timestamp 1676037725
transform 1 0 39100 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_419
timestamp 1676037725
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_421
timestamp 1676037725
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_433
timestamp 1676037725
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_445
timestamp 1676037725
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_457
timestamp 1676037725
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_469
timestamp 1676037725
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 1676037725
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_477
timestamp 1676037725
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_489
timestamp 1676037725
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_501
timestamp 1676037725
transform 1 0 47196 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_507
timestamp 1676037725
transform 1 0 47748 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_516
timestamp 1676037725
transform 1 0 48576 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_528
timestamp 1676037725
transform 1 0 49680 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_533
timestamp 1676037725
transform 1 0 50140 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_545
timestamp 1676037725
transform 1 0 51244 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_557
timestamp 1676037725
transform 1 0 52348 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_569
timestamp 1676037725
transform 1 0 53452 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_581
timestamp 1676037725
transform 1 0 54556 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_587
timestamp 1676037725
transform 1 0 55108 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_589
timestamp 1676037725
transform 1 0 55292 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_601
timestamp 1676037725
transform 1 0 56396 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_613
timestamp 1676037725
transform 1 0 57500 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_623
timestamp 1676037725
transform 1 0 58420 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_3
timestamp 1676037725
transform 1 0 1380 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_9
timestamp 1676037725
transform 1 0 1932 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_17
timestamp 1676037725
transform 1 0 2668 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_29
timestamp 1676037725
transform 1 0 3772 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_41
timestamp 1676037725
transform 1 0 4876 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_53
timestamp 1676037725
transform 1 0 5980 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1676037725
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1676037725
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1676037725
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_93
timestamp 1676037725
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1676037725
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1676037725
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1676037725
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1676037725
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1676037725
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1676037725
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1676037725
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1676037725
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1676037725
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1676037725
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_193
timestamp 1676037725
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_205
timestamp 1676037725
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1676037725
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1676037725
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_225
timestamp 1676037725
transform 1 0 21804 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_233
timestamp 1676037725
transform 1 0 22540 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_45_249
timestamp 1676037725
transform 1 0 24012 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_257
timestamp 1676037725
transform 1 0 24748 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_266
timestamp 1676037725
transform 1 0 25576 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_45_277
timestamp 1676037725
transform 1 0 26588 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_45_281
timestamp 1676037725
transform 1 0 26956 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_289
timestamp 1676037725
transform 1 0 27692 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_300
timestamp 1676037725
transform 1 0 28704 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_312
timestamp 1676037725
transform 1 0 29808 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_318
timestamp 1676037725
transform 1 0 30360 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_326
timestamp 1676037725
transform 1 0 31096 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_334
timestamp 1676037725
transform 1 0 31832 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_337
timestamp 1676037725
transform 1 0 32108 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_351
timestamp 1676037725
transform 1 0 33396 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_363
timestamp 1676037725
transform 1 0 34500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_375
timestamp 1676037725
transform 1 0 35604 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_387
timestamp 1676037725
transform 1 0 36708 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1676037725
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_393
timestamp 1676037725
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_405
timestamp 1676037725
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_417
timestamp 1676037725
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_429
timestamp 1676037725
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_441
timestamp 1676037725
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1676037725
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_449
timestamp 1676037725
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_461
timestamp 1676037725
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_473
timestamp 1676037725
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_485
timestamp 1676037725
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1676037725
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1676037725
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_505
timestamp 1676037725
transform 1 0 47564 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_517
timestamp 1676037725
transform 1 0 48668 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_529
timestamp 1676037725
transform 1 0 49772 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_541
timestamp 1676037725
transform 1 0 50876 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_553
timestamp 1676037725
transform 1 0 51980 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_559
timestamp 1676037725
transform 1 0 52532 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_561
timestamp 1676037725
transform 1 0 52716 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_573
timestamp 1676037725
transform 1 0 53820 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_585
timestamp 1676037725
transform 1 0 54924 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_597
timestamp 1676037725
transform 1 0 56028 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_609
timestamp 1676037725
transform 1 0 57132 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_615
timestamp 1676037725
transform 1 0 57684 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_617
timestamp 1676037725
transform 1 0 57868 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_623
timestamp 1676037725
transform 1 0 58420 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_3
timestamp 1676037725
transform 1 0 1380 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_9
timestamp 1676037725
transform 1 0 1932 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_21
timestamp 1676037725
transform 1 0 3036 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1676037725
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1676037725
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1676037725
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1676037725
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1676037725
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1676037725
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1676037725
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1676037725
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1676037725
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_109
timestamp 1676037725
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_121
timestamp 1676037725
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1676037725
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1676037725
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1676037725
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1676037725
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_165
timestamp 1676037725
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_177
timestamp 1676037725
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1676037725
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1676037725
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1676037725
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1676037725
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_221
timestamp 1676037725
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_233
timestamp 1676037725
transform 1 0 22540 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_250
timestamp 1676037725
transform 1 0 24104 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_253
timestamp 1676037725
transform 1 0 24380 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_261
timestamp 1676037725
transform 1 0 25116 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_272
timestamp 1676037725
transform 1 0 26128 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_283
timestamp 1676037725
transform 1 0 27140 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_287
timestamp 1676037725
transform 1 0 27508 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_296
timestamp 1676037725
transform 1 0 28336 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_309
timestamp 1676037725
transform 1 0 29532 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_313
timestamp 1676037725
transform 1 0 29900 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_326
timestamp 1676037725
transform 1 0 31096 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_334
timestamp 1676037725
transform 1 0 31832 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_342
timestamp 1676037725
transform 1 0 32568 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_362
timestamp 1676037725
transform 1 0 34408 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1676037725
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1676037725
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_389
timestamp 1676037725
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_401
timestamp 1676037725
transform 1 0 37996 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_413
timestamp 1676037725
transform 1 0 39100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_419
timestamp 1676037725
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_421
timestamp 1676037725
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_433
timestamp 1676037725
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_445
timestamp 1676037725
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_457
timestamp 1676037725
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 1676037725
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1676037725
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_477
timestamp 1676037725
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_489
timestamp 1676037725
transform 1 0 46092 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_501
timestamp 1676037725
transform 1 0 47196 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_513
timestamp 1676037725
transform 1 0 48300 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_529
timestamp 1676037725
transform 1 0 49772 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_533
timestamp 1676037725
transform 1 0 50140 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_545
timestamp 1676037725
transform 1 0 51244 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_557
timestamp 1676037725
transform 1 0 52348 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_569
timestamp 1676037725
transform 1 0 53452 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_581
timestamp 1676037725
transform 1 0 54556 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_587
timestamp 1676037725
transform 1 0 55108 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_589
timestamp 1676037725
transform 1 0 55292 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_601
timestamp 1676037725
transform 1 0 56396 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_613
timestamp 1676037725
transform 1 0 57500 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_623
timestamp 1676037725
transform 1 0 58420 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_3
timestamp 1676037725
transform 1 0 1380 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_9
timestamp 1676037725
transform 1 0 1932 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_21
timestamp 1676037725
transform 1 0 3036 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_33
timestamp 1676037725
transform 1 0 4140 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_45
timestamp 1676037725
transform 1 0 5244 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_53
timestamp 1676037725
transform 1 0 5980 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1676037725
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1676037725
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1676037725
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_93
timestamp 1676037725
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1676037725
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1676037725
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1676037725
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1676037725
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_137
timestamp 1676037725
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_149
timestamp 1676037725
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1676037725
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1676037725
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1676037725
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_181
timestamp 1676037725
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_193
timestamp 1676037725
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_205
timestamp 1676037725
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1676037725
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1676037725
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1676037725
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_256
timestamp 1676037725
transform 1 0 24656 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_272
timestamp 1676037725
transform 1 0 26128 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_281
timestamp 1676037725
transform 1 0 26956 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_289
timestamp 1676037725
transform 1 0 27692 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_297
timestamp 1676037725
transform 1 0 28428 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_305
timestamp 1676037725
transform 1 0 29164 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_318
timestamp 1676037725
transform 1 0 30360 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_331
timestamp 1676037725
transform 1 0 31556 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1676037725
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1676037725
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1676037725
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1676037725
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_373
timestamp 1676037725
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1676037725
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1676037725
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_393
timestamp 1676037725
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_405
timestamp 1676037725
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_417
timestamp 1676037725
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_429
timestamp 1676037725
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_441
timestamp 1676037725
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1676037725
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_449
timestamp 1676037725
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_461
timestamp 1676037725
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_473
timestamp 1676037725
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_485
timestamp 1676037725
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_497
timestamp 1676037725
transform 1 0 46828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 1676037725
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_505
timestamp 1676037725
transform 1 0 47564 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_517
timestamp 1676037725
transform 1 0 48668 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_529
timestamp 1676037725
transform 1 0 49772 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_541
timestamp 1676037725
transform 1 0 50876 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_553
timestamp 1676037725
transform 1 0 51980 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_559
timestamp 1676037725
transform 1 0 52532 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_561
timestamp 1676037725
transform 1 0 52716 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_573
timestamp 1676037725
transform 1 0 53820 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_585
timestamp 1676037725
transform 1 0 54924 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_597
timestamp 1676037725
transform 1 0 56028 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_609
timestamp 1676037725
transform 1 0 57132 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_615
timestamp 1676037725
transform 1 0 57684 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_617
timestamp 1676037725
transform 1 0 57868 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_623
timestamp 1676037725
transform 1 0 58420 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_3
timestamp 1676037725
transform 1 0 1380 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_9
timestamp 1676037725
transform 1 0 1932 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_21
timestamp 1676037725
transform 1 0 3036 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1676037725
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1676037725
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1676037725
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1676037725
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1676037725
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1676037725
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1676037725
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1676037725
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1676037725
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1676037725
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_121
timestamp 1676037725
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1676037725
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1676037725
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1676037725
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_153
timestamp 1676037725
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_165
timestamp 1676037725
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_177
timestamp 1676037725
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1676037725
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1676037725
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1676037725
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_209
timestamp 1676037725
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_221
timestamp 1676037725
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_233
timestamp 1676037725
transform 1 0 22540 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_250
timestamp 1676037725
transform 1 0 24104 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_253
timestamp 1676037725
transform 1 0 24380 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_261
timestamp 1676037725
transform 1 0 25116 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_270
timestamp 1676037725
transform 1 0 25944 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_282
timestamp 1676037725
transform 1 0 27048 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_294
timestamp 1676037725
transform 1 0 28152 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_298
timestamp 1676037725
transform 1 0 28520 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_306
timestamp 1676037725
transform 1 0 29256 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_309
timestamp 1676037725
transform 1 0 29532 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_320
timestamp 1676037725
transform 1 0 30544 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_328
timestamp 1676037725
transform 1 0 31280 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_338
timestamp 1676037725
transform 1 0 32200 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_350
timestamp 1676037725
transform 1 0 33304 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_362
timestamp 1676037725
transform 1 0 34408 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1676037725
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1676037725
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_389
timestamp 1676037725
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_401
timestamp 1676037725
transform 1 0 37996 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_413
timestamp 1676037725
transform 1 0 39100 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 1676037725
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_421
timestamp 1676037725
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_433
timestamp 1676037725
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_445
timestamp 1676037725
transform 1 0 42044 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_454
timestamp 1676037725
transform 1 0 42872 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_466
timestamp 1676037725
transform 1 0 43976 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_474
timestamp 1676037725
transform 1 0 44712 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_477
timestamp 1676037725
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_489
timestamp 1676037725
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_501
timestamp 1676037725
transform 1 0 47196 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_513
timestamp 1676037725
transform 1 0 48300 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_522
timestamp 1676037725
transform 1 0 49128 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_530
timestamp 1676037725
transform 1 0 49864 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_533
timestamp 1676037725
transform 1 0 50140 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_545
timestamp 1676037725
transform 1 0 51244 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_557
timestamp 1676037725
transform 1 0 52348 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_569
timestamp 1676037725
transform 1 0 53452 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_581
timestamp 1676037725
transform 1 0 54556 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_587
timestamp 1676037725
transform 1 0 55108 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_589
timestamp 1676037725
transform 1 0 55292 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_601
timestamp 1676037725
transform 1 0 56396 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_613
timestamp 1676037725
transform 1 0 57500 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_623
timestamp 1676037725
transform 1 0 58420 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_3
timestamp 1676037725
transform 1 0 1380 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_9
timestamp 1676037725
transform 1 0 1932 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_18
timestamp 1676037725
transform 1 0 2760 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_30
timestamp 1676037725
transform 1 0 3864 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_42
timestamp 1676037725
transform 1 0 4968 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_54
timestamp 1676037725
transform 1 0 6072 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1676037725
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1676037725
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_81
timestamp 1676037725
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_93
timestamp 1676037725
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1676037725
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1676037725
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1676037725
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1676037725
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_137
timestamp 1676037725
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_149
timestamp 1676037725
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1676037725
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1676037725
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1676037725
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_181
timestamp 1676037725
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_193
timestamp 1676037725
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_205
timestamp 1676037725
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1676037725
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1676037725
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_49_225
timestamp 1676037725
transform 1 0 21804 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_233
timestamp 1676037725
transform 1 0 22540 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_256
timestamp 1676037725
transform 1 0 24656 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_268
timestamp 1676037725
transform 1 0 25760 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1676037725
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_295
timestamp 1676037725
transform 1 0 28244 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_304
timestamp 1676037725
transform 1 0 29072 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_324
timestamp 1676037725
transform 1 0 30912 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_334
timestamp 1676037725
transform 1 0 31832 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1676037725
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1676037725
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1676037725
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1676037725
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1676037725
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1676037725
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_393
timestamp 1676037725
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_405
timestamp 1676037725
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_417
timestamp 1676037725
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_429
timestamp 1676037725
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_441
timestamp 1676037725
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1676037725
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_449
timestamp 1676037725
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_461
timestamp 1676037725
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_473
timestamp 1676037725
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_485
timestamp 1676037725
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 1676037725
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1676037725
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_505
timestamp 1676037725
transform 1 0 47564 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_517
timestamp 1676037725
transform 1 0 48668 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_529
timestamp 1676037725
transform 1 0 49772 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_541
timestamp 1676037725
transform 1 0 50876 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_553
timestamp 1676037725
transform 1 0 51980 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_559
timestamp 1676037725
transform 1 0 52532 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_561
timestamp 1676037725
transform 1 0 52716 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_573
timestamp 1676037725
transform 1 0 53820 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_585
timestamp 1676037725
transform 1 0 54924 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_597
timestamp 1676037725
transform 1 0 56028 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_609
timestamp 1676037725
transform 1 0 57132 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_615
timestamp 1676037725
transform 1 0 57684 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_617
timestamp 1676037725
transform 1 0 57868 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_623
timestamp 1676037725
transform 1 0 58420 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_3
timestamp 1676037725
transform 1 0 1380 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_9
timestamp 1676037725
transform 1 0 1932 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_17
timestamp 1676037725
transform 1 0 2668 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_25
timestamp 1676037725
transform 1 0 3404 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1676037725
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1676037725
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1676037725
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1676037725
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1676037725
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1676037725
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1676037725
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1676037725
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_109
timestamp 1676037725
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_121
timestamp 1676037725
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1676037725
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1676037725
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1676037725
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1676037725
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_165
timestamp 1676037725
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_177
timestamp 1676037725
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1676037725
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1676037725
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1676037725
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_209
timestamp 1676037725
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_221
timestamp 1676037725
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_233
timestamp 1676037725
transform 1 0 22540 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_237
timestamp 1676037725
transform 1 0 22908 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_250
timestamp 1676037725
transform 1 0 24104 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1676037725
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_265
timestamp 1676037725
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_277
timestamp 1676037725
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_289
timestamp 1676037725
transform 1 0 27692 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_295
timestamp 1676037725
transform 1 0 28244 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_306
timestamp 1676037725
transform 1 0 29256 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_309
timestamp 1676037725
transform 1 0 29532 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_320
timestamp 1676037725
transform 1 0 30544 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_332
timestamp 1676037725
transform 1 0 31648 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_50_348
timestamp 1676037725
transform 1 0 33120 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_360
timestamp 1676037725
transform 1 0 34224 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1676037725
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_377
timestamp 1676037725
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_389
timestamp 1676037725
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_401
timestamp 1676037725
transform 1 0 37996 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_413
timestamp 1676037725
transform 1 0 39100 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_419
timestamp 1676037725
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_421
timestamp 1676037725
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_433
timestamp 1676037725
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_445
timestamp 1676037725
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_457
timestamp 1676037725
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1676037725
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1676037725
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_477
timestamp 1676037725
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_489
timestamp 1676037725
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_501
timestamp 1676037725
transform 1 0 47196 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_513
timestamp 1676037725
transform 1 0 48300 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_525
timestamp 1676037725
transform 1 0 49404 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_531
timestamp 1676037725
transform 1 0 49956 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_533
timestamp 1676037725
transform 1 0 50140 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_545
timestamp 1676037725
transform 1 0 51244 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_557
timestamp 1676037725
transform 1 0 52348 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_569
timestamp 1676037725
transform 1 0 53452 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_581
timestamp 1676037725
transform 1 0 54556 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_587
timestamp 1676037725
transform 1 0 55108 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_589
timestamp 1676037725
transform 1 0 55292 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_601
timestamp 1676037725
transform 1 0 56396 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_613
timestamp 1676037725
transform 1 0 57500 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_623
timestamp 1676037725
transform 1 0 58420 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_3
timestamp 1676037725
transform 1 0 1380 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_9
timestamp 1676037725
transform 1 0 1932 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_20
timestamp 1676037725
transform 1 0 2944 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_32
timestamp 1676037725
transform 1 0 4048 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_44
timestamp 1676037725
transform 1 0 5152 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1676037725
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1676037725
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1676037725
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_93
timestamp 1676037725
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1676037725
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1676037725
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1676037725
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1676037725
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_137
timestamp 1676037725
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_149
timestamp 1676037725
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1676037725
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1676037725
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_169
timestamp 1676037725
transform 1 0 16652 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_178
timestamp 1676037725
transform 1 0 17480 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_190
timestamp 1676037725
transform 1 0 18584 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_202
timestamp 1676037725
transform 1 0 19688 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_214
timestamp 1676037725
transform 1 0 20792 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_222
timestamp 1676037725
transform 1 0 21528 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_225
timestamp 1676037725
transform 1 0 21804 0 -1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_51_241
timestamp 1676037725
transform 1 0 23276 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_253
timestamp 1676037725
transform 1 0 24380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_265
timestamp 1676037725
transform 1 0 25484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_277
timestamp 1676037725
transform 1 0 26588 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1676037725
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_293
timestamp 1676037725
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_305
timestamp 1676037725
transform 1 0 29164 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_313
timestamp 1676037725
transform 1 0 29900 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_331
timestamp 1676037725
transform 1 0 31556 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1676037725
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1676037725
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1676037725
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1676037725
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_373
timestamp 1676037725
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1676037725
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1676037725
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_393
timestamp 1676037725
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_405
timestamp 1676037725
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_417
timestamp 1676037725
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_429
timestamp 1676037725
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_441
timestamp 1676037725
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1676037725
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_449
timestamp 1676037725
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_461
timestamp 1676037725
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_473
timestamp 1676037725
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_485
timestamp 1676037725
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1676037725
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1676037725
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_505
timestamp 1676037725
transform 1 0 47564 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_517
timestamp 1676037725
transform 1 0 48668 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_529
timestamp 1676037725
transform 1 0 49772 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_541
timestamp 1676037725
transform 1 0 50876 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_553
timestamp 1676037725
transform 1 0 51980 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_559
timestamp 1676037725
transform 1 0 52532 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_561
timestamp 1676037725
transform 1 0 52716 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_573
timestamp 1676037725
transform 1 0 53820 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_585
timestamp 1676037725
transform 1 0 54924 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_597
timestamp 1676037725
transform 1 0 56028 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_609
timestamp 1676037725
transform 1 0 57132 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_615
timestamp 1676037725
transform 1 0 57684 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_617
timestamp 1676037725
transform 1 0 57868 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_623
timestamp 1676037725
transform 1 0 58420 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_3
timestamp 1676037725
transform 1 0 1380 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_9
timestamp 1676037725
transform 1 0 1932 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_21
timestamp 1676037725
transform 1 0 3036 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1676037725
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1676037725
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1676037725
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1676037725
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1676037725
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1676037725
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1676037725
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1676037725
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1676037725
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_109
timestamp 1676037725
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_121
timestamp 1676037725
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1676037725
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1676037725
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1676037725
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_153
timestamp 1676037725
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_165
timestamp 1676037725
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_177
timestamp 1676037725
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1676037725
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1676037725
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1676037725
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_209
timestamp 1676037725
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_221
timestamp 1676037725
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_233
timestamp 1676037725
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1676037725
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1676037725
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1676037725
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_265
timestamp 1676037725
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_277
timestamp 1676037725
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_289
timestamp 1676037725
transform 1 0 27692 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_304
timestamp 1676037725
transform 1 0 29072 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_309
timestamp 1676037725
transform 1 0 29532 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_320
timestamp 1676037725
transform 1 0 30544 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_328
timestamp 1676037725
transform 1 0 31280 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_339
timestamp 1676037725
transform 1 0 32292 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_351
timestamp 1676037725
transform 1 0 33396 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1676037725
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1676037725
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_377
timestamp 1676037725
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_389
timestamp 1676037725
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_401
timestamp 1676037725
transform 1 0 37996 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_413
timestamp 1676037725
transform 1 0 39100 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_419
timestamp 1676037725
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_421
timestamp 1676037725
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_433
timestamp 1676037725
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_445
timestamp 1676037725
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_457
timestamp 1676037725
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1676037725
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1676037725
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_477
timestamp 1676037725
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_489
timestamp 1676037725
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_501
timestamp 1676037725
transform 1 0 47196 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_512
timestamp 1676037725
transform 1 0 48208 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_524
timestamp 1676037725
transform 1 0 49312 0 1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_52_533
timestamp 1676037725
transform 1 0 50140 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_545
timestamp 1676037725
transform 1 0 51244 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_557
timestamp 1676037725
transform 1 0 52348 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_569
timestamp 1676037725
transform 1 0 53452 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_581
timestamp 1676037725
transform 1 0 54556 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_587
timestamp 1676037725
transform 1 0 55108 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_589
timestamp 1676037725
transform 1 0 55292 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_601
timestamp 1676037725
transform 1 0 56396 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_613
timestamp 1676037725
transform 1 0 57500 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_52_623
timestamp 1676037725
transform 1 0 58420 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_3
timestamp 1676037725
transform 1 0 1380 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_9
timestamp 1676037725
transform 1 0 1932 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_17
timestamp 1676037725
transform 1 0 2668 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_29
timestamp 1676037725
transform 1 0 3772 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_41
timestamp 1676037725
transform 1 0 4876 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_53
timestamp 1676037725
transform 1 0 5980 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1676037725
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1676037725
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1676037725
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1676037725
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1676037725
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1676037725
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1676037725
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1676037725
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1676037725
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_149
timestamp 1676037725
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1676037725
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1676037725
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1676037725
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_181
timestamp 1676037725
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_193
timestamp 1676037725
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_205
timestamp 1676037725
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1676037725
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1676037725
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1676037725
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_237
timestamp 1676037725
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_249
timestamp 1676037725
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_261
timestamp 1676037725
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1676037725
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1676037725
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1676037725
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1676037725
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1676037725
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_317
timestamp 1676037725
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1676037725
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1676037725
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1676037725
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1676037725
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_361
timestamp 1676037725
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_373
timestamp 1676037725
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1676037725
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1676037725
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1676037725
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_405
timestamp 1676037725
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_417
timestamp 1676037725
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_429
timestamp 1676037725
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 1676037725
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1676037725
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_449
timestamp 1676037725
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_461
timestamp 1676037725
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_473
timestamp 1676037725
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_485
timestamp 1676037725
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_497
timestamp 1676037725
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 1676037725
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_505
timestamp 1676037725
transform 1 0 47564 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_514
timestamp 1676037725
transform 1 0 48392 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_526
timestamp 1676037725
transform 1 0 49496 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_538
timestamp 1676037725
transform 1 0 50600 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_550
timestamp 1676037725
transform 1 0 51704 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_558
timestamp 1676037725
transform 1 0 52440 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_561
timestamp 1676037725
transform 1 0 52716 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_573
timestamp 1676037725
transform 1 0 53820 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_585
timestamp 1676037725
transform 1 0 54924 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_597
timestamp 1676037725
transform 1 0 56028 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_609
timestamp 1676037725
transform 1 0 57132 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_615
timestamp 1676037725
transform 1 0 57684 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_617
timestamp 1676037725
transform 1 0 57868 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_623
timestamp 1676037725
transform 1 0 58420 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_3
timestamp 1676037725
transform 1 0 1380 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_9
timestamp 1676037725
transform 1 0 1932 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_17
timestamp 1676037725
transform 1 0 2668 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_25
timestamp 1676037725
transform 1 0 3404 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1676037725
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1676037725
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1676037725
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1676037725
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1676037725
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1676037725
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1676037725
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1676037725
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1676037725
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1676037725
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1676037725
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1676037725
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1676037725
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1676037725
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_165
timestamp 1676037725
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_177
timestamp 1676037725
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1676037725
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1676037725
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1676037725
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_209
timestamp 1676037725
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_221
timestamp 1676037725
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_233
timestamp 1676037725
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1676037725
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1676037725
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1676037725
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_265
timestamp 1676037725
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_277
timestamp 1676037725
transform 1 0 26588 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_283
timestamp 1676037725
transform 1 0 27140 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_286
timestamp 1676037725
transform 1 0 27416 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_295
timestamp 1676037725
transform 1 0 28244 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1676037725
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1676037725
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1676037725
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1676037725
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1676037725
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1676037725
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1676037725
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1676037725
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_377
timestamp 1676037725
transform 1 0 35788 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_383
timestamp 1676037725
transform 1 0 36340 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_393
timestamp 1676037725
transform 1 0 37260 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_405
timestamp 1676037725
transform 1 0 38364 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_417
timestamp 1676037725
transform 1 0 39468 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_54_421
timestamp 1676037725
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_433
timestamp 1676037725
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_445
timestamp 1676037725
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_457
timestamp 1676037725
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 1676037725
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1676037725
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_477
timestamp 1676037725
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_489
timestamp 1676037725
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_501
timestamp 1676037725
transform 1 0 47196 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_513
timestamp 1676037725
transform 1 0 48300 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_525
timestamp 1676037725
transform 1 0 49404 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_531
timestamp 1676037725
transform 1 0 49956 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_533
timestamp 1676037725
transform 1 0 50140 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_545
timestamp 1676037725
transform 1 0 51244 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_557
timestamp 1676037725
transform 1 0 52348 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_569
timestamp 1676037725
transform 1 0 53452 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_581
timestamp 1676037725
transform 1 0 54556 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_587
timestamp 1676037725
transform 1 0 55108 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_589
timestamp 1676037725
transform 1 0 55292 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_601
timestamp 1676037725
transform 1 0 56396 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_613
timestamp 1676037725
transform 1 0 57500 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_623
timestamp 1676037725
transform 1 0 58420 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_55_3
timestamp 1676037725
transform 1 0 1380 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_9
timestamp 1676037725
transform 1 0 1932 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_55_17
timestamp 1676037725
transform 1 0 2668 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_55_22
timestamp 1676037725
transform 1 0 3128 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_33
timestamp 1676037725
transform 1 0 4140 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_45
timestamp 1676037725
transform 1 0 5244 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_53
timestamp 1676037725
transform 1 0 5980 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1676037725
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1676037725
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1676037725
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1676037725
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1676037725
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1676037725
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1676037725
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1676037725
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1676037725
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1676037725
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1676037725
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1676037725
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1676037725
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_181
timestamp 1676037725
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_193
timestamp 1676037725
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_205
timestamp 1676037725
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1676037725
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1676037725
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1676037725
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_237
timestamp 1676037725
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_249
timestamp 1676037725
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_261
timestamp 1676037725
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1676037725
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1676037725
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_281
timestamp 1676037725
transform 1 0 26956 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_289
timestamp 1676037725
transform 1 0 27692 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_299
timestamp 1676037725
transform 1 0 28612 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_312
timestamp 1676037725
transform 1 0 29808 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_324
timestamp 1676037725
transform 1 0 30912 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1676037725
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1676037725
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1676037725
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_373
timestamp 1676037725
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1676037725
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1676037725
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_393
timestamp 1676037725
transform 1 0 37260 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_401
timestamp 1676037725
transform 1 0 37996 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_413
timestamp 1676037725
transform 1 0 39100 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_425
timestamp 1676037725
transform 1 0 40204 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_437
timestamp 1676037725
transform 1 0 41308 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_445
timestamp 1676037725
transform 1 0 42044 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_449
timestamp 1676037725
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_461
timestamp 1676037725
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_473
timestamp 1676037725
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_485
timestamp 1676037725
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_497
timestamp 1676037725
transform 1 0 46828 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_503
timestamp 1676037725
transform 1 0 47380 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_505
timestamp 1676037725
transform 1 0 47564 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_517
timestamp 1676037725
transform 1 0 48668 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_529
timestamp 1676037725
transform 1 0 49772 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_541
timestamp 1676037725
transform 1 0 50876 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_553
timestamp 1676037725
transform 1 0 51980 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_559
timestamp 1676037725
transform 1 0 52532 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_561
timestamp 1676037725
transform 1 0 52716 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_573
timestamp 1676037725
transform 1 0 53820 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_585
timestamp 1676037725
transform 1 0 54924 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_597
timestamp 1676037725
transform 1 0 56028 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_609
timestamp 1676037725
transform 1 0 57132 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_615
timestamp 1676037725
transform 1 0 57684 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_617
timestamp 1676037725
transform 1 0 57868 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_623
timestamp 1676037725
transform 1 0 58420 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_3
timestamp 1676037725
transform 1 0 1380 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_9
timestamp 1676037725
transform 1 0 1932 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_21
timestamp 1676037725
transform 1 0 3036 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1676037725
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1676037725
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1676037725
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1676037725
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1676037725
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1676037725
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1676037725
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1676037725
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1676037725
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1676037725
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1676037725
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1676037725
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1676037725
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1676037725
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1676037725
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1676037725
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1676037725
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1676037725
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1676037725
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1676037725
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1676037725
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_221
timestamp 1676037725
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_233
timestamp 1676037725
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1676037725
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1676037725
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1676037725
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_265
timestamp 1676037725
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_277
timestamp 1676037725
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_289
timestamp 1676037725
transform 1 0 27692 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_299
timestamp 1676037725
transform 1 0 28612 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1676037725
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1676037725
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1676037725
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1676037725
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1676037725
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1676037725
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1676037725
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1676037725
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1676037725
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_389
timestamp 1676037725
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_401
timestamp 1676037725
transform 1 0 37996 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_413
timestamp 1676037725
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1676037725
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_421
timestamp 1676037725
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_433
timestamp 1676037725
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_445
timestamp 1676037725
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_457
timestamp 1676037725
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 1676037725
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1676037725
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_477
timestamp 1676037725
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_489
timestamp 1676037725
transform 1 0 46092 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_501
timestamp 1676037725
transform 1 0 47196 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_513
timestamp 1676037725
transform 1 0 48300 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_525
timestamp 1676037725
transform 1 0 49404 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_531
timestamp 1676037725
transform 1 0 49956 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_533
timestamp 1676037725
transform 1 0 50140 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_545
timestamp 1676037725
transform 1 0 51244 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_557
timestamp 1676037725
transform 1 0 52348 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_569
timestamp 1676037725
transform 1 0 53452 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_581
timestamp 1676037725
transform 1 0 54556 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_587
timestamp 1676037725
transform 1 0 55108 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_589
timestamp 1676037725
transform 1 0 55292 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_601
timestamp 1676037725
transform 1 0 56396 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_613
timestamp 1676037725
transform 1 0 57500 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_623
timestamp 1676037725
transform 1 0 58420 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_3
timestamp 1676037725
transform 1 0 1380 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_9
timestamp 1676037725
transform 1 0 1932 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_21
timestamp 1676037725
transform 1 0 3036 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_33
timestamp 1676037725
transform 1 0 4140 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_45
timestamp 1676037725
transform 1 0 5244 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_53
timestamp 1676037725
transform 1 0 5980 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1676037725
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1676037725
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1676037725
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1676037725
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1676037725
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1676037725
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1676037725
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1676037725
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1676037725
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1676037725
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1676037725
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1676037725
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1676037725
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1676037725
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_193
timestamp 1676037725
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_205
timestamp 1676037725
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1676037725
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1676037725
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1676037725
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_237
timestamp 1676037725
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_249
timestamp 1676037725
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_261
timestamp 1676037725
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1676037725
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1676037725
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1676037725
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1676037725
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_305
timestamp 1676037725
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_317
timestamp 1676037725
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1676037725
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1676037725
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_337
timestamp 1676037725
transform 1 0 32108 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_345
timestamp 1676037725
transform 1 0 32844 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_367
timestamp 1676037725
transform 1 0 34868 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_379
timestamp 1676037725
transform 1 0 35972 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1676037725
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_393
timestamp 1676037725
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_405
timestamp 1676037725
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_417
timestamp 1676037725
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_429
timestamp 1676037725
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 1676037725
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1676037725
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_449
timestamp 1676037725
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_461
timestamp 1676037725
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_473
timestamp 1676037725
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_485
timestamp 1676037725
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_497
timestamp 1676037725
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 1676037725
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_505
timestamp 1676037725
transform 1 0 47564 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_517
timestamp 1676037725
transform 1 0 48668 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_529
timestamp 1676037725
transform 1 0 49772 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_541
timestamp 1676037725
transform 1 0 50876 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_553
timestamp 1676037725
transform 1 0 51980 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_559
timestamp 1676037725
transform 1 0 52532 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_561
timestamp 1676037725
transform 1 0 52716 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_573
timestamp 1676037725
transform 1 0 53820 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_585
timestamp 1676037725
transform 1 0 54924 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_597
timestamp 1676037725
transform 1 0 56028 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_609
timestamp 1676037725
transform 1 0 57132 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_615
timestamp 1676037725
transform 1 0 57684 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_617
timestamp 1676037725
transform 1 0 57868 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_623
timestamp 1676037725
transform 1 0 58420 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_3
timestamp 1676037725
transform 1 0 1380 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_9
timestamp 1676037725
transform 1 0 1932 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_21
timestamp 1676037725
transform 1 0 3036 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1676037725
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_29
timestamp 1676037725
transform 1 0 3772 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_39
timestamp 1676037725
transform 1 0 4692 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_51
timestamp 1676037725
transform 1 0 5796 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_63
timestamp 1676037725
transform 1 0 6900 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_75
timestamp 1676037725
transform 1 0 8004 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1676037725
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1676037725
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1676037725
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1676037725
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1676037725
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1676037725
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1676037725
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1676037725
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1676037725
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1676037725
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1676037725
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1676037725
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1676037725
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1676037725
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1676037725
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_221
timestamp 1676037725
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_233
timestamp 1676037725
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1676037725
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1676037725
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 1676037725
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_265
timestamp 1676037725
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_277
timestamp 1676037725
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_289
timestamp 1676037725
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1676037725
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1676037725
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1676037725
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1676037725
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1676037725
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_345
timestamp 1676037725
transform 1 0 32844 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_353
timestamp 1676037725
transform 1 0 33580 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_360
timestamp 1676037725
transform 1 0 34224 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_365
timestamp 1676037725
transform 1 0 34684 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_372
timestamp 1676037725
transform 1 0 35328 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_384
timestamp 1676037725
transform 1 0 36432 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_396
timestamp 1676037725
transform 1 0 37536 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_408
timestamp 1676037725
transform 1 0 38640 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_421
timestamp 1676037725
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_433
timestamp 1676037725
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_445
timestamp 1676037725
transform 1 0 42044 0 1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_58_460
timestamp 1676037725
transform 1 0 43424 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_472
timestamp 1676037725
transform 1 0 44528 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_477
timestamp 1676037725
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_489
timestamp 1676037725
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_515
timestamp 1676037725
transform 1 0 48484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_527
timestamp 1676037725
transform 1 0 49588 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_531
timestamp 1676037725
transform 1 0 49956 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_533
timestamp 1676037725
transform 1 0 50140 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_545
timestamp 1676037725
transform 1 0 51244 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_557
timestamp 1676037725
transform 1 0 52348 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_569
timestamp 1676037725
transform 1 0 53452 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_581
timestamp 1676037725
transform 1 0 54556 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_587
timestamp 1676037725
transform 1 0 55108 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_589
timestamp 1676037725
transform 1 0 55292 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_601
timestamp 1676037725
transform 1 0 56396 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_613
timestamp 1676037725
transform 1 0 57500 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_623
timestamp 1676037725
transform 1 0 58420 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_3
timestamp 1676037725
transform 1 0 1380 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_9
timestamp 1676037725
transform 1 0 1932 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_21
timestamp 1676037725
transform 1 0 3036 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_33
timestamp 1676037725
transform 1 0 4140 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_45
timestamp 1676037725
transform 1 0 5244 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_53
timestamp 1676037725
transform 1 0 5980 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1676037725
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1676037725
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1676037725
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1676037725
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1676037725
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1676037725
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1676037725
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1676037725
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1676037725
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1676037725
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1676037725
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1676037725
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1676037725
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1676037725
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1676037725
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1676037725
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1676037725
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1676037725
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1676037725
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1676037725
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_249
timestamp 1676037725
transform 1 0 24012 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_260
timestamp 1676037725
transform 1 0 25024 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_272
timestamp 1676037725
transform 1 0 26128 0 -1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1676037725
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_293
timestamp 1676037725
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_305
timestamp 1676037725
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_317
timestamp 1676037725
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1676037725
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1676037725
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_337
timestamp 1676037725
transform 1 0 32108 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_349
timestamp 1676037725
transform 1 0 33212 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_353
timestamp 1676037725
transform 1 0 33580 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_364
timestamp 1676037725
transform 1 0 34592 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_376
timestamp 1676037725
transform 1 0 35696 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_388
timestamp 1676037725
transform 1 0 36800 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_393
timestamp 1676037725
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_405
timestamp 1676037725
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_417
timestamp 1676037725
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_429
timestamp 1676037725
transform 1 0 40572 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_59_437
timestamp 1676037725
transform 1 0 41308 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_446
timestamp 1676037725
transform 1 0 42136 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_449
timestamp 1676037725
transform 1 0 42412 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_465
timestamp 1676037725
transform 1 0 43884 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_477
timestamp 1676037725
transform 1 0 44988 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_489
timestamp 1676037725
transform 1 0 46092 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_59_501
timestamp 1676037725
transform 1 0 47196 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_505
timestamp 1676037725
transform 1 0 47564 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_517
timestamp 1676037725
transform 1 0 48668 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_529
timestamp 1676037725
transform 1 0 49772 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_541
timestamp 1676037725
transform 1 0 50876 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_553
timestamp 1676037725
transform 1 0 51980 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_559
timestamp 1676037725
transform 1 0 52532 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_561
timestamp 1676037725
transform 1 0 52716 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_573
timestamp 1676037725
transform 1 0 53820 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_585
timestamp 1676037725
transform 1 0 54924 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_597
timestamp 1676037725
transform 1 0 56028 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_609
timestamp 1676037725
transform 1 0 57132 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_615
timestamp 1676037725
transform 1 0 57684 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_617
timestamp 1676037725
transform 1 0 57868 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_623
timestamp 1676037725
transform 1 0 58420 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_3
timestamp 1676037725
transform 1 0 1380 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_9
timestamp 1676037725
transform 1 0 1932 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_21
timestamp 1676037725
transform 1 0 3036 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1676037725
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1676037725
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1676037725
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1676037725
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1676037725
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1676037725
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1676037725
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1676037725
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1676037725
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1676037725
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1676037725
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1676037725
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1676037725
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1676037725
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1676037725
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1676037725
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1676037725
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1676037725
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1676037725
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1676037725
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_209
timestamp 1676037725
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_221
timestamp 1676037725
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_233
timestamp 1676037725
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1676037725
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1676037725
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1676037725
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_265
timestamp 1676037725
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_277
timestamp 1676037725
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_289
timestamp 1676037725
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1676037725
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1676037725
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_309
timestamp 1676037725
transform 1 0 29532 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_317
timestamp 1676037725
transform 1 0 30268 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_326
timestamp 1676037725
transform 1 0 31096 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_341
timestamp 1676037725
transform 1 0 32476 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_354
timestamp 1676037725
transform 1 0 33672 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_362
timestamp 1676037725
transform 1 0 34408 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1676037725
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1676037725
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_389
timestamp 1676037725
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_401
timestamp 1676037725
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_413
timestamp 1676037725
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1676037725
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_421
timestamp 1676037725
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_433
timestamp 1676037725
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_445
timestamp 1676037725
transform 1 0 42044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_455
timestamp 1676037725
transform 1 0 42964 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_467
timestamp 1676037725
transform 1 0 44068 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1676037725
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_477
timestamp 1676037725
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_489
timestamp 1676037725
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_501
timestamp 1676037725
transform 1 0 47196 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_513
timestamp 1676037725
transform 1 0 48300 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_525
timestamp 1676037725
transform 1 0 49404 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_531
timestamp 1676037725
transform 1 0 49956 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_533
timestamp 1676037725
transform 1 0 50140 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_545
timestamp 1676037725
transform 1 0 51244 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_557
timestamp 1676037725
transform 1 0 52348 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_569
timestamp 1676037725
transform 1 0 53452 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_581
timestamp 1676037725
transform 1 0 54556 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_587
timestamp 1676037725
transform 1 0 55108 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_589
timestamp 1676037725
transform 1 0 55292 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_601
timestamp 1676037725
transform 1 0 56396 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_613
timestamp 1676037725
transform 1 0 57500 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_623
timestamp 1676037725
transform 1 0 58420 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_3
timestamp 1676037725
transform 1 0 1380 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_9
timestamp 1676037725
transform 1 0 1932 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_15
timestamp 1676037725
transform 1 0 2484 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_24
timestamp 1676037725
transform 1 0 3312 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_36
timestamp 1676037725
transform 1 0 4416 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_48
timestamp 1676037725
transform 1 0 5520 0 -1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1676037725
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1676037725
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1676037725
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1676037725
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1676037725
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1676037725
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1676037725
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1676037725
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1676037725
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1676037725
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1676037725
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1676037725
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1676037725
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1676037725
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1676037725
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_205
timestamp 1676037725
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1676037725
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1676037725
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1676037725
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_237
timestamp 1676037725
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_249
timestamp 1676037725
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_261
timestamp 1676037725
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1676037725
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1676037725
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_281
timestamp 1676037725
transform 1 0 26956 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_289
timestamp 1676037725
transform 1 0 27692 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_299
timestamp 1676037725
transform 1 0 28612 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_312
timestamp 1676037725
transform 1 0 29808 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_324
timestamp 1676037725
transform 1 0 30912 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_337
timestamp 1676037725
transform 1 0 32108 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_345
timestamp 1676037725
transform 1 0 32844 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_354
timestamp 1676037725
transform 1 0 33672 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_366
timestamp 1676037725
transform 1 0 34776 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_378
timestamp 1676037725
transform 1 0 35880 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_390
timestamp 1676037725
transform 1 0 36984 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_393
timestamp 1676037725
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_405
timestamp 1676037725
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_417
timestamp 1676037725
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_429
timestamp 1676037725
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 1676037725
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1676037725
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_449
timestamp 1676037725
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_461
timestamp 1676037725
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_473
timestamp 1676037725
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_485
timestamp 1676037725
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 1676037725
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1676037725
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_505
timestamp 1676037725
transform 1 0 47564 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_517
timestamp 1676037725
transform 1 0 48668 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_529
timestamp 1676037725
transform 1 0 49772 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_541
timestamp 1676037725
transform 1 0 50876 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_553
timestamp 1676037725
transform 1 0 51980 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_559
timestamp 1676037725
transform 1 0 52532 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_561
timestamp 1676037725
transform 1 0 52716 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_573
timestamp 1676037725
transform 1 0 53820 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_585
timestamp 1676037725
transform 1 0 54924 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_597
timestamp 1676037725
transform 1 0 56028 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_609
timestamp 1676037725
transform 1 0 57132 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_615
timestamp 1676037725
transform 1 0 57684 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_617
timestamp 1676037725
transform 1 0 57868 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_623
timestamp 1676037725
transform 1 0 58420 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_3
timestamp 1676037725
transform 1 0 1380 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_9
timestamp 1676037725
transform 1 0 1932 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_21
timestamp 1676037725
transform 1 0 3036 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1676037725
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1676037725
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1676037725
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1676037725
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1676037725
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1676037725
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1676037725
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1676037725
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1676037725
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1676037725
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1676037725
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1676037725
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1676037725
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1676037725
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1676037725
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1676037725
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1676037725
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1676037725
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1676037725
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_197
timestamp 1676037725
transform 1 0 19228 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_203
timestamp 1676037725
transform 1 0 19780 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_211
timestamp 1676037725
transform 1 0 20516 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_223
timestamp 1676037725
transform 1 0 21620 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_235
timestamp 1676037725
transform 1 0 22724 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_247
timestamp 1676037725
transform 1 0 23828 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1676037725
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1676037725
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_265
timestamp 1676037725
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_277
timestamp 1676037725
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_289
timestamp 1676037725
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1676037725
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1676037725
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_309
timestamp 1676037725
transform 1 0 29532 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_315
timestamp 1676037725
transform 1 0 30084 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1676037725
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1676037725
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1676037725
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1676037725
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1676037725
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_377
timestamp 1676037725
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_389
timestamp 1676037725
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_401
timestamp 1676037725
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_413
timestamp 1676037725
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 1676037725
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_421
timestamp 1676037725
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_433
timestamp 1676037725
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_445
timestamp 1676037725
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_457
timestamp 1676037725
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1676037725
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1676037725
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_477
timestamp 1676037725
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_489
timestamp 1676037725
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_501
timestamp 1676037725
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_513
timestamp 1676037725
transform 1 0 48300 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_525
timestamp 1676037725
transform 1 0 49404 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_531
timestamp 1676037725
transform 1 0 49956 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_533
timestamp 1676037725
transform 1 0 50140 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_545
timestamp 1676037725
transform 1 0 51244 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_557
timestamp 1676037725
transform 1 0 52348 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_569
timestamp 1676037725
transform 1 0 53452 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_581
timestamp 1676037725
transform 1 0 54556 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_587
timestamp 1676037725
transform 1 0 55108 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_589
timestamp 1676037725
transform 1 0 55292 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_601
timestamp 1676037725
transform 1 0 56396 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_613
timestamp 1676037725
transform 1 0 57500 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_623
timestamp 1676037725
transform 1 0 58420 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_3
timestamp 1676037725
transform 1 0 1380 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_9
timestamp 1676037725
transform 1 0 1932 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_21
timestamp 1676037725
transform 1 0 3036 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_39
timestamp 1676037725
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1676037725
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1676037725
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1676037725
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1676037725
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1676037725
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 1676037725
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1676037725
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1676037725
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1676037725
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1676037725
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1676037725
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_149
timestamp 1676037725
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1676037725
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1676037725
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1676037725
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_181
timestamp 1676037725
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_193
timestamp 1676037725
transform 1 0 18860 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_201
timestamp 1676037725
transform 1 0 19596 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_222
timestamp 1676037725
transform 1 0 21528 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_225
timestamp 1676037725
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_237
timestamp 1676037725
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_249
timestamp 1676037725
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_261
timestamp 1676037725
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_273
timestamp 1676037725
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1676037725
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_281
timestamp 1676037725
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_293
timestamp 1676037725
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_305
timestamp 1676037725
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_317
timestamp 1676037725
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1676037725
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1676037725
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_337
timestamp 1676037725
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_349
timestamp 1676037725
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_361
timestamp 1676037725
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_373
timestamp 1676037725
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1676037725
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1676037725
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_393
timestamp 1676037725
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_405
timestamp 1676037725
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_417
timestamp 1676037725
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_429
timestamp 1676037725
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1676037725
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1676037725
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_449
timestamp 1676037725
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_461
timestamp 1676037725
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_473
timestamp 1676037725
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_485
timestamp 1676037725
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1676037725
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1676037725
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_505
timestamp 1676037725
transform 1 0 47564 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_517
timestamp 1676037725
transform 1 0 48668 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_529
timestamp 1676037725
transform 1 0 49772 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_541
timestamp 1676037725
transform 1 0 50876 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_553
timestamp 1676037725
transform 1 0 51980 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_559
timestamp 1676037725
transform 1 0 52532 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_561
timestamp 1676037725
transform 1 0 52716 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_573
timestamp 1676037725
transform 1 0 53820 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_585
timestamp 1676037725
transform 1 0 54924 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_597
timestamp 1676037725
transform 1 0 56028 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_609
timestamp 1676037725
transform 1 0 57132 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_615
timestamp 1676037725
transform 1 0 57684 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_617
timestamp 1676037725
transform 1 0 57868 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_623
timestamp 1676037725
transform 1 0 58420 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_3
timestamp 1676037725
transform 1 0 1380 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_9
timestamp 1676037725
transform 1 0 1932 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_21
timestamp 1676037725
transform 1 0 3036 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1676037725
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1676037725
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1676037725
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_53
timestamp 1676037725
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_65
timestamp 1676037725
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1676037725
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1676037725
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1676037725
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_97
timestamp 1676037725
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_109
timestamp 1676037725
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_121
timestamp 1676037725
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1676037725
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1676037725
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_141
timestamp 1676037725
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_153
timestamp 1676037725
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_165
timestamp 1676037725
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_177
timestamp 1676037725
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1676037725
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1676037725
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_197
timestamp 1676037725
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_209
timestamp 1676037725
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_221
timestamp 1676037725
transform 1 0 21436 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_233
timestamp 1676037725
transform 1 0 22540 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_245
timestamp 1676037725
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1676037725
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_253
timestamp 1676037725
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_265
timestamp 1676037725
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_277
timestamp 1676037725
transform 1 0 26588 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_289
timestamp 1676037725
transform 1 0 27692 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_301
timestamp 1676037725
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1676037725
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_309
timestamp 1676037725
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_321
timestamp 1676037725
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_333
timestamp 1676037725
transform 1 0 31740 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_345
timestamp 1676037725
transform 1 0 32844 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1676037725
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1676037725
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_365
timestamp 1676037725
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_377
timestamp 1676037725
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_389
timestamp 1676037725
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_401
timestamp 1676037725
transform 1 0 37996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_413
timestamp 1676037725
transform 1 0 39100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_419
timestamp 1676037725
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_421
timestamp 1676037725
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_433
timestamp 1676037725
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_445
timestamp 1676037725
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_457
timestamp 1676037725
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_469
timestamp 1676037725
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1676037725
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_477
timestamp 1676037725
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_489
timestamp 1676037725
transform 1 0 46092 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_501
timestamp 1676037725
transform 1 0 47196 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_513
timestamp 1676037725
transform 1 0 48300 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_525
timestamp 1676037725
transform 1 0 49404 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_531
timestamp 1676037725
transform 1 0 49956 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_533
timestamp 1676037725
transform 1 0 50140 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_545
timestamp 1676037725
transform 1 0 51244 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_557
timestamp 1676037725
transform 1 0 52348 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_569
timestamp 1676037725
transform 1 0 53452 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_581
timestamp 1676037725
transform 1 0 54556 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_587
timestamp 1676037725
transform 1 0 55108 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_589
timestamp 1676037725
transform 1 0 55292 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_601
timestamp 1676037725
transform 1 0 56396 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_613
timestamp 1676037725
transform 1 0 57500 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_623
timestamp 1676037725
transform 1 0 58420 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_3
timestamp 1676037725
transform 1 0 1380 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_9
timestamp 1676037725
transform 1 0 1932 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_21
timestamp 1676037725
transform 1 0 3036 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_33
timestamp 1676037725
transform 1 0 4140 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_45
timestamp 1676037725
transform 1 0 5244 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_53
timestamp 1676037725
transform 1 0 5980 0 -1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_65_57
timestamp 1676037725
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_69
timestamp 1676037725
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_81
timestamp 1676037725
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_93
timestamp 1676037725
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1676037725
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1676037725
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_113
timestamp 1676037725
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_125
timestamp 1676037725
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_137
timestamp 1676037725
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_149
timestamp 1676037725
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1676037725
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1676037725
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_169
timestamp 1676037725
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_181
timestamp 1676037725
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_193
timestamp 1676037725
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_205
timestamp 1676037725
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_217
timestamp 1676037725
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1676037725
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_225
timestamp 1676037725
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_237
timestamp 1676037725
transform 1 0 22908 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_249
timestamp 1676037725
transform 1 0 24012 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_261
timestamp 1676037725
transform 1 0 25116 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_273
timestamp 1676037725
transform 1 0 26220 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_279
timestamp 1676037725
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_281
timestamp 1676037725
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_293
timestamp 1676037725
transform 1 0 28060 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_305
timestamp 1676037725
transform 1 0 29164 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_317
timestamp 1676037725
transform 1 0 30268 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_329
timestamp 1676037725
transform 1 0 31372 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_335
timestamp 1676037725
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_65_337
timestamp 1676037725
transform 1 0 32108 0 -1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_65_351
timestamp 1676037725
transform 1 0 33396 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_363
timestamp 1676037725
transform 1 0 34500 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_375
timestamp 1676037725
transform 1 0 35604 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_387
timestamp 1676037725
transform 1 0 36708 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1676037725
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_393
timestamp 1676037725
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_405
timestamp 1676037725
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_417
timestamp 1676037725
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_429
timestamp 1676037725
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_441
timestamp 1676037725
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1676037725
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_449
timestamp 1676037725
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_461
timestamp 1676037725
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_473
timestamp 1676037725
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_485
timestamp 1676037725
transform 1 0 45724 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_497
timestamp 1676037725
transform 1 0 46828 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_503
timestamp 1676037725
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_505
timestamp 1676037725
transform 1 0 47564 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_517
timestamp 1676037725
transform 1 0 48668 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_529
timestamp 1676037725
transform 1 0 49772 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_541
timestamp 1676037725
transform 1 0 50876 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_553
timestamp 1676037725
transform 1 0 51980 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_559
timestamp 1676037725
transform 1 0 52532 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_561
timestamp 1676037725
transform 1 0 52716 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_573
timestamp 1676037725
transform 1 0 53820 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_585
timestamp 1676037725
transform 1 0 54924 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_597
timestamp 1676037725
transform 1 0 56028 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_609
timestamp 1676037725
transform 1 0 57132 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_615
timestamp 1676037725
transform 1 0 57684 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_617
timestamp 1676037725
transform 1 0 57868 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_3
timestamp 1676037725
transform 1 0 1380 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_9
timestamp 1676037725
transform 1 0 1932 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_21
timestamp 1676037725
transform 1 0 3036 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1676037725
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_29
timestamp 1676037725
transform 1 0 3772 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_37
timestamp 1676037725
transform 1 0 4508 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_47
timestamp 1676037725
transform 1 0 5428 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_59
timestamp 1676037725
transform 1 0 6532 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_71
timestamp 1676037725
transform 1 0 7636 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1676037725
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_85
timestamp 1676037725
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_97
timestamp 1676037725
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_109
timestamp 1676037725
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_121
timestamp 1676037725
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1676037725
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1676037725
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_141
timestamp 1676037725
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_153
timestamp 1676037725
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_165
timestamp 1676037725
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_177
timestamp 1676037725
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1676037725
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1676037725
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_197
timestamp 1676037725
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_209
timestamp 1676037725
transform 1 0 20332 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_221
timestamp 1676037725
transform 1 0 21436 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_233
timestamp 1676037725
transform 1 0 22540 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_245
timestamp 1676037725
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1676037725
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_253
timestamp 1676037725
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_265
timestamp 1676037725
transform 1 0 25484 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_277
timestamp 1676037725
transform 1 0 26588 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_289
timestamp 1676037725
transform 1 0 27692 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_301
timestamp 1676037725
transform 1 0 28796 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_307
timestamp 1676037725
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_309
timestamp 1676037725
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_321
timestamp 1676037725
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_333
timestamp 1676037725
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_66_345
timestamp 1676037725
transform 1 0 32844 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_66_356
timestamp 1676037725
transform 1 0 33856 0 1 38080
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_66_365
timestamp 1676037725
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_377
timestamp 1676037725
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_389
timestamp 1676037725
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_401
timestamp 1676037725
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_413
timestamp 1676037725
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_419
timestamp 1676037725
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_421
timestamp 1676037725
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_433
timestamp 1676037725
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_445
timestamp 1676037725
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_457
timestamp 1676037725
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_469
timestamp 1676037725
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 1676037725
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_477
timestamp 1676037725
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_489
timestamp 1676037725
transform 1 0 46092 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_501
timestamp 1676037725
transform 1 0 47196 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_513
timestamp 1676037725
transform 1 0 48300 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_525
timestamp 1676037725
transform 1 0 49404 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_531
timestamp 1676037725
transform 1 0 49956 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_533
timestamp 1676037725
transform 1 0 50140 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_545
timestamp 1676037725
transform 1 0 51244 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_557
timestamp 1676037725
transform 1 0 52348 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_569
timestamp 1676037725
transform 1 0 53452 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_581
timestamp 1676037725
transform 1 0 54556 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_587
timestamp 1676037725
transform 1 0 55108 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_589
timestamp 1676037725
transform 1 0 55292 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_601
timestamp 1676037725
transform 1 0 56396 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_613
timestamp 1676037725
transform 1 0 57500 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_67_3
timestamp 1676037725
transform 1 0 1380 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_67_9
timestamp 1676037725
transform 1 0 1932 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_21
timestamp 1676037725
transform 1 0 3036 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_33
timestamp 1676037725
transform 1 0 4140 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_45
timestamp 1676037725
transform 1 0 5244 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_53
timestamp 1676037725
transform 1 0 5980 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1676037725
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_69
timestamp 1676037725
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_81
timestamp 1676037725
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_93
timestamp 1676037725
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1676037725
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1676037725
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_113
timestamp 1676037725
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_125
timestamp 1676037725
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_137
timestamp 1676037725
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_149
timestamp 1676037725
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1676037725
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1676037725
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_169
timestamp 1676037725
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_181
timestamp 1676037725
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_193
timestamp 1676037725
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_205
timestamp 1676037725
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1676037725
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1676037725
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_225
timestamp 1676037725
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_237
timestamp 1676037725
transform 1 0 22908 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_249
timestamp 1676037725
transform 1 0 24012 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_261
timestamp 1676037725
transform 1 0 25116 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_273
timestamp 1676037725
transform 1 0 26220 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_279
timestamp 1676037725
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_281
timestamp 1676037725
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_293
timestamp 1676037725
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_305
timestamp 1676037725
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_317
timestamp 1676037725
transform 1 0 30268 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_329
timestamp 1676037725
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1676037725
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_67_337
timestamp 1676037725
transform 1 0 32108 0 -1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_67_350
timestamp 1676037725
transform 1 0 33304 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_362
timestamp 1676037725
transform 1 0 34408 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_374
timestamp 1676037725
transform 1 0 35512 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_386
timestamp 1676037725
transform 1 0 36616 0 -1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_67_393
timestamp 1676037725
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_405
timestamp 1676037725
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_417
timestamp 1676037725
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_429
timestamp 1676037725
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_441
timestamp 1676037725
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1676037725
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_449
timestamp 1676037725
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_461
timestamp 1676037725
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_473
timestamp 1676037725
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_485
timestamp 1676037725
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_497
timestamp 1676037725
transform 1 0 46828 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_503
timestamp 1676037725
transform 1 0 47380 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_505
timestamp 1676037725
transform 1 0 47564 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_517
timestamp 1676037725
transform 1 0 48668 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_529
timestamp 1676037725
transform 1 0 49772 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_541
timestamp 1676037725
transform 1 0 50876 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_553
timestamp 1676037725
transform 1 0 51980 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_559
timestamp 1676037725
transform 1 0 52532 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_561
timestamp 1676037725
transform 1 0 52716 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_573
timestamp 1676037725
transform 1 0 53820 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_585
timestamp 1676037725
transform 1 0 54924 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_597
timestamp 1676037725
transform 1 0 56028 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_609
timestamp 1676037725
transform 1 0 57132 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_615
timestamp 1676037725
transform 1 0 57684 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_67_617
timestamp 1676037725
transform 1 0 57868 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_67_623
timestamp 1676037725
transform 1 0 58420 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_3
timestamp 1676037725
transform 1 0 1380 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_68_9
timestamp 1676037725
transform 1 0 1932 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_21
timestamp 1676037725
transform 1 0 3036 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1676037725
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1676037725
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1676037725
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_53
timestamp 1676037725
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_65
timestamp 1676037725
transform 1 0 7084 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_68_76
timestamp 1676037725
transform 1 0 8096 0 1 39168
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_68_85
timestamp 1676037725
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_97
timestamp 1676037725
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_109
timestamp 1676037725
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_121
timestamp 1676037725
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1676037725
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1676037725
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_141
timestamp 1676037725
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_153
timestamp 1676037725
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_165
timestamp 1676037725
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_177
timestamp 1676037725
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1676037725
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1676037725
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_197
timestamp 1676037725
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_209
timestamp 1676037725
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_221
timestamp 1676037725
transform 1 0 21436 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_233
timestamp 1676037725
transform 1 0 22540 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_245
timestamp 1676037725
transform 1 0 23644 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_251
timestamp 1676037725
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_253
timestamp 1676037725
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_265
timestamp 1676037725
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_277
timestamp 1676037725
transform 1 0 26588 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_289
timestamp 1676037725
transform 1 0 27692 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_301
timestamp 1676037725
transform 1 0 28796 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 1676037725
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_309
timestamp 1676037725
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_321
timestamp 1676037725
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_333
timestamp 1676037725
transform 1 0 31740 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_345
timestamp 1676037725
transform 1 0 32844 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_357
timestamp 1676037725
transform 1 0 33948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_363
timestamp 1676037725
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_365
timestamp 1676037725
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_377
timestamp 1676037725
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_389
timestamp 1676037725
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_401
timestamp 1676037725
transform 1 0 37996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_413
timestamp 1676037725
transform 1 0 39100 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_419
timestamp 1676037725
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_421
timestamp 1676037725
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_433
timestamp 1676037725
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_445
timestamp 1676037725
transform 1 0 42044 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_457
timestamp 1676037725
transform 1 0 43148 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_469
timestamp 1676037725
transform 1 0 44252 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_475
timestamp 1676037725
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_477
timestamp 1676037725
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_489
timestamp 1676037725
transform 1 0 46092 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_501
timestamp 1676037725
transform 1 0 47196 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_513
timestamp 1676037725
transform 1 0 48300 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_525
timestamp 1676037725
transform 1 0 49404 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_531
timestamp 1676037725
transform 1 0 49956 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_533
timestamp 1676037725
transform 1 0 50140 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_545
timestamp 1676037725
transform 1 0 51244 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_557
timestamp 1676037725
transform 1 0 52348 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_569
timestamp 1676037725
transform 1 0 53452 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_581
timestamp 1676037725
transform 1 0 54556 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_587
timestamp 1676037725
transform 1 0 55108 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_589
timestamp 1676037725
transform 1 0 55292 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_601
timestamp 1676037725
transform 1 0 56396 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_613
timestamp 1676037725
transform 1 0 57500 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_69_3
timestamp 1676037725
transform 1 0 1380 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_69_9
timestamp 1676037725
transform 1 0 1932 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_21
timestamp 1676037725
transform 1 0 3036 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_33
timestamp 1676037725
transform 1 0 4140 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_45
timestamp 1676037725
transform 1 0 5244 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_69_53
timestamp 1676037725
transform 1 0 5980 0 -1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_69_57
timestamp 1676037725
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_69
timestamp 1676037725
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_81
timestamp 1676037725
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_93
timestamp 1676037725
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1676037725
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1676037725
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_113
timestamp 1676037725
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_125
timestamp 1676037725
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_137
timestamp 1676037725
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_149
timestamp 1676037725
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1676037725
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1676037725
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_169
timestamp 1676037725
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_181
timestamp 1676037725
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_193
timestamp 1676037725
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_205
timestamp 1676037725
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_217
timestamp 1676037725
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1676037725
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_225
timestamp 1676037725
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_237
timestamp 1676037725
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_249
timestamp 1676037725
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_261
timestamp 1676037725
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_273
timestamp 1676037725
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1676037725
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_281
timestamp 1676037725
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_293
timestamp 1676037725
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_305
timestamp 1676037725
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_317
timestamp 1676037725
transform 1 0 30268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_329
timestamp 1676037725
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_335
timestamp 1676037725
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_337
timestamp 1676037725
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_349
timestamp 1676037725
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_361
timestamp 1676037725
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_373
timestamp 1676037725
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_385
timestamp 1676037725
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 1676037725
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_393
timestamp 1676037725
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_405
timestamp 1676037725
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_417
timestamp 1676037725
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_429
timestamp 1676037725
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_441
timestamp 1676037725
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 1676037725
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_449
timestamp 1676037725
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_461
timestamp 1676037725
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_473
timestamp 1676037725
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_485
timestamp 1676037725
transform 1 0 45724 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_497
timestamp 1676037725
transform 1 0 46828 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_503
timestamp 1676037725
transform 1 0 47380 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_505
timestamp 1676037725
transform 1 0 47564 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_517
timestamp 1676037725
transform 1 0 48668 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_529
timestamp 1676037725
transform 1 0 49772 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_541
timestamp 1676037725
transform 1 0 50876 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_553
timestamp 1676037725
transform 1 0 51980 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_559
timestamp 1676037725
transform 1 0 52532 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_561
timestamp 1676037725
transform 1 0 52716 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_573
timestamp 1676037725
transform 1 0 53820 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_585
timestamp 1676037725
transform 1 0 54924 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_597
timestamp 1676037725
transform 1 0 56028 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_609
timestamp 1676037725
transform 1 0 57132 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_615
timestamp 1676037725
transform 1 0 57684 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_69_617
timestamp 1676037725
transform 1 0 57868 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_69_623
timestamp 1676037725
transform 1 0 58420 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_3
timestamp 1676037725
transform 1 0 1380 0 1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_70_9
timestamp 1676037725
transform 1 0 1932 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_21
timestamp 1676037725
transform 1 0 3036 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1676037725
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1676037725
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1676037725
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_53
timestamp 1676037725
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_65
timestamp 1676037725
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1676037725
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1676037725
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_70_85
timestamp 1676037725
transform 1 0 8924 0 1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_70_95
timestamp 1676037725
transform 1 0 9844 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_107
timestamp 1676037725
transform 1 0 10948 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_119
timestamp 1676037725
transform 1 0 12052 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_131
timestamp 1676037725
transform 1 0 13156 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1676037725
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_141
timestamp 1676037725
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_153
timestamp 1676037725
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_165
timestamp 1676037725
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_177
timestamp 1676037725
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1676037725
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1676037725
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_197
timestamp 1676037725
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_209
timestamp 1676037725
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_221
timestamp 1676037725
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_233
timestamp 1676037725
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_245
timestamp 1676037725
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1676037725
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_253
timestamp 1676037725
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_265
timestamp 1676037725
transform 1 0 25484 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_277
timestamp 1676037725
transform 1 0 26588 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_289
timestamp 1676037725
transform 1 0 27692 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_301
timestamp 1676037725
transform 1 0 28796 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_307
timestamp 1676037725
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_309
timestamp 1676037725
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_321
timestamp 1676037725
transform 1 0 30636 0 1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_70_334
timestamp 1676037725
transform 1 0 31832 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_346
timestamp 1676037725
transform 1 0 32936 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_358
timestamp 1676037725
transform 1 0 34040 0 1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_70_365
timestamp 1676037725
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_377
timestamp 1676037725
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_389
timestamp 1676037725
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_401
timestamp 1676037725
transform 1 0 37996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_413
timestamp 1676037725
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_419
timestamp 1676037725
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_70_421
timestamp 1676037725
transform 1 0 39836 0 1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_70_430
timestamp 1676037725
transform 1 0 40664 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_442
timestamp 1676037725
transform 1 0 41768 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_454
timestamp 1676037725
transform 1 0 42872 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_466
timestamp 1676037725
transform 1 0 43976 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_70_474
timestamp 1676037725
transform 1 0 44712 0 1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_70_477
timestamp 1676037725
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_489
timestamp 1676037725
transform 1 0 46092 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_501
timestamp 1676037725
transform 1 0 47196 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_513
timestamp 1676037725
transform 1 0 48300 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_525
timestamp 1676037725
transform 1 0 49404 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_531
timestamp 1676037725
transform 1 0 49956 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_533
timestamp 1676037725
transform 1 0 50140 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_545
timestamp 1676037725
transform 1 0 51244 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_557
timestamp 1676037725
transform 1 0 52348 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_569
timestamp 1676037725
transform 1 0 53452 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_581
timestamp 1676037725
transform 1 0 54556 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_587
timestamp 1676037725
transform 1 0 55108 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_589
timestamp 1676037725
transform 1 0 55292 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_601
timestamp 1676037725
transform 1 0 56396 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_613
timestamp 1676037725
transform 1 0 57500 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_3
timestamp 1676037725
transform 1 0 1380 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_9
timestamp 1676037725
transform 1 0 1932 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_21
timestamp 1676037725
transform 1 0 3036 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_33
timestamp 1676037725
transform 1 0 4140 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_45
timestamp 1676037725
transform 1 0 5244 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_71_53
timestamp 1676037725
transform 1 0 5980 0 -1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1676037725
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_69
timestamp 1676037725
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_81
timestamp 1676037725
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_93
timestamp 1676037725
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1676037725
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1676037725
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_113
timestamp 1676037725
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_125
timestamp 1676037725
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_137
timestamp 1676037725
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_149
timestamp 1676037725
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1676037725
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1676037725
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_169
timestamp 1676037725
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_181
timestamp 1676037725
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_193
timestamp 1676037725
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_205
timestamp 1676037725
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_217
timestamp 1676037725
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1676037725
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_225
timestamp 1676037725
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_237
timestamp 1676037725
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_249
timestamp 1676037725
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_261
timestamp 1676037725
transform 1 0 25116 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_273
timestamp 1676037725
transform 1 0 26220 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_279
timestamp 1676037725
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_281
timestamp 1676037725
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_293
timestamp 1676037725
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_305
timestamp 1676037725
transform 1 0 29164 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_317
timestamp 1676037725
transform 1 0 30268 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_329
timestamp 1676037725
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_335
timestamp 1676037725
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_337
timestamp 1676037725
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_349
timestamp 1676037725
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_361
timestamp 1676037725
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_373
timestamp 1676037725
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_385
timestamp 1676037725
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_391
timestamp 1676037725
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_393
timestamp 1676037725
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_405
timestamp 1676037725
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_417
timestamp 1676037725
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_429
timestamp 1676037725
transform 1 0 40572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_441
timestamp 1676037725
transform 1 0 41676 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_447
timestamp 1676037725
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_449
timestamp 1676037725
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_461
timestamp 1676037725
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_473
timestamp 1676037725
transform 1 0 44620 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_485
timestamp 1676037725
transform 1 0 45724 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_497
timestamp 1676037725
transform 1 0 46828 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_503
timestamp 1676037725
transform 1 0 47380 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_505
timestamp 1676037725
transform 1 0 47564 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_517
timestamp 1676037725
transform 1 0 48668 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_529
timestamp 1676037725
transform 1 0 49772 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_541
timestamp 1676037725
transform 1 0 50876 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_553
timestamp 1676037725
transform 1 0 51980 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_559
timestamp 1676037725
transform 1 0 52532 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_561
timestamp 1676037725
transform 1 0 52716 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_573
timestamp 1676037725
transform 1 0 53820 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_585
timestamp 1676037725
transform 1 0 54924 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_597
timestamp 1676037725
transform 1 0 56028 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_609
timestamp 1676037725
transform 1 0 57132 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_615
timestamp 1676037725
transform 1 0 57684 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_617
timestamp 1676037725
transform 1 0 57868 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_72_3
timestamp 1676037725
transform 1 0 1380 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_9
timestamp 1676037725
transform 1 0 1932 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_21
timestamp 1676037725
transform 1 0 3036 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1676037725
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1676037725
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_41
timestamp 1676037725
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_53
timestamp 1676037725
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_65
timestamp 1676037725
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1676037725
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1676037725
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_85
timestamp 1676037725
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_97
timestamp 1676037725
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_109
timestamp 1676037725
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_121
timestamp 1676037725
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1676037725
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1676037725
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_141
timestamp 1676037725
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_153
timestamp 1676037725
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_165
timestamp 1676037725
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_177
timestamp 1676037725
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1676037725
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1676037725
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_197
timestamp 1676037725
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_209
timestamp 1676037725
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_221
timestamp 1676037725
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_233
timestamp 1676037725
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_245
timestamp 1676037725
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1676037725
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_253
timestamp 1676037725
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_265
timestamp 1676037725
transform 1 0 25484 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_72_273
timestamp 1676037725
transform 1 0 26220 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_283
timestamp 1676037725
transform 1 0 27140 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_295
timestamp 1676037725
transform 1 0 28244 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 1676037725
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_309
timestamp 1676037725
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_321
timestamp 1676037725
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_333
timestamp 1676037725
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_345
timestamp 1676037725
transform 1 0 32844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_357
timestamp 1676037725
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 1676037725
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_365
timestamp 1676037725
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_377
timestamp 1676037725
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_389
timestamp 1676037725
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_401
timestamp 1676037725
transform 1 0 37996 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_413
timestamp 1676037725
transform 1 0 39100 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_419
timestamp 1676037725
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_421
timestamp 1676037725
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_433
timestamp 1676037725
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_445
timestamp 1676037725
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_457
timestamp 1676037725
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_469
timestamp 1676037725
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 1676037725
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_477
timestamp 1676037725
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_489
timestamp 1676037725
transform 1 0 46092 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_501
timestamp 1676037725
transform 1 0 47196 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_513
timestamp 1676037725
transform 1 0 48300 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_525
timestamp 1676037725
transform 1 0 49404 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_531
timestamp 1676037725
transform 1 0 49956 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_533
timestamp 1676037725
transform 1 0 50140 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_545
timestamp 1676037725
transform 1 0 51244 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_557
timestamp 1676037725
transform 1 0 52348 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_569
timestamp 1676037725
transform 1 0 53452 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_581
timestamp 1676037725
transform 1 0 54556 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_587
timestamp 1676037725
transform 1 0 55108 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_589
timestamp 1676037725
transform 1 0 55292 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_601
timestamp 1676037725
transform 1 0 56396 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_613
timestamp 1676037725
transform 1 0 57500 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_619
timestamp 1676037725
transform 1 0 58052 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_72_623
timestamp 1676037725
transform 1 0 58420 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_3
timestamp 1676037725
transform 1 0 1380 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_9
timestamp 1676037725
transform 1 0 1932 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_21
timestamp 1676037725
transform 1 0 3036 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_33
timestamp 1676037725
transform 1 0 4140 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_45
timestamp 1676037725
transform 1 0 5244 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_73_53
timestamp 1676037725
transform 1 0 5980 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1676037725
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_69
timestamp 1676037725
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_81
timestamp 1676037725
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_93
timestamp 1676037725
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1676037725
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1676037725
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_113
timestamp 1676037725
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_125
timestamp 1676037725
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_137
timestamp 1676037725
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_149
timestamp 1676037725
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1676037725
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1676037725
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_169
timestamp 1676037725
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_181
timestamp 1676037725
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_193
timestamp 1676037725
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_205
timestamp 1676037725
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1676037725
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1676037725
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_225
timestamp 1676037725
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_237
timestamp 1676037725
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_249
timestamp 1676037725
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_261
timestamp 1676037725
transform 1 0 25116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_273
timestamp 1676037725
transform 1 0 26220 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1676037725
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_281
timestamp 1676037725
transform 1 0 26956 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_289
timestamp 1676037725
transform 1 0 27692 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_298
timestamp 1676037725
transform 1 0 28520 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_310
timestamp 1676037725
transform 1 0 29624 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_322
timestamp 1676037725
transform 1 0 30728 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_73_334
timestamp 1676037725
transform 1 0 31832 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_337
timestamp 1676037725
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_349
timestamp 1676037725
transform 1 0 33212 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_361
timestamp 1676037725
transform 1 0 34316 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_373
timestamp 1676037725
transform 1 0 35420 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_385
timestamp 1676037725
transform 1 0 36524 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_391
timestamp 1676037725
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_393
timestamp 1676037725
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_405
timestamp 1676037725
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_417
timestamp 1676037725
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_429
timestamp 1676037725
transform 1 0 40572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_441
timestamp 1676037725
transform 1 0 41676 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_447
timestamp 1676037725
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_449
timestamp 1676037725
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_461
timestamp 1676037725
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_473
timestamp 1676037725
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_485
timestamp 1676037725
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_497
timestamp 1676037725
transform 1 0 46828 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_503
timestamp 1676037725
transform 1 0 47380 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_505
timestamp 1676037725
transform 1 0 47564 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_517
timestamp 1676037725
transform 1 0 48668 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_529
timestamp 1676037725
transform 1 0 49772 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_541
timestamp 1676037725
transform 1 0 50876 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_553
timestamp 1676037725
transform 1 0 51980 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_559
timestamp 1676037725
transform 1 0 52532 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_561
timestamp 1676037725
transform 1 0 52716 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_573
timestamp 1676037725
transform 1 0 53820 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_585
timestamp 1676037725
transform 1 0 54924 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_597
timestamp 1676037725
transform 1 0 56028 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_609
timestamp 1676037725
transform 1 0 57132 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_615
timestamp 1676037725
transform 1 0 57684 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_73_617
timestamp 1676037725
transform 1 0 57868 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_73_623
timestamp 1676037725
transform 1 0 58420 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_74_3
timestamp 1676037725
transform 1 0 1380 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_74_9
timestamp 1676037725
transform 1 0 1932 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_21
timestamp 1676037725
transform 1 0 3036 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1676037725
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1676037725
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_41
timestamp 1676037725
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_53
timestamp 1676037725
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_65
timestamp 1676037725
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1676037725
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1676037725
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_85
timestamp 1676037725
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_97
timestamp 1676037725
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_109
timestamp 1676037725
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_121
timestamp 1676037725
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1676037725
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1676037725
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_141
timestamp 1676037725
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_153
timestamp 1676037725
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_165
timestamp 1676037725
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_177
timestamp 1676037725
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1676037725
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1676037725
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_197
timestamp 1676037725
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_209
timestamp 1676037725
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_221
timestamp 1676037725
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_233
timestamp 1676037725
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1676037725
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1676037725
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_253
timestamp 1676037725
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_265
timestamp 1676037725
transform 1 0 25484 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_277
timestamp 1676037725
transform 1 0 26588 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_289
timestamp 1676037725
transform 1 0 27692 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_301
timestamp 1676037725
transform 1 0 28796 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_307
timestamp 1676037725
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_309
timestamp 1676037725
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_321
timestamp 1676037725
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_333
timestamp 1676037725
transform 1 0 31740 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_345
timestamp 1676037725
transform 1 0 32844 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_357
timestamp 1676037725
transform 1 0 33948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1676037725
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_365
timestamp 1676037725
transform 1 0 34684 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_377
timestamp 1676037725
transform 1 0 35788 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_389
timestamp 1676037725
transform 1 0 36892 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_401
timestamp 1676037725
transform 1 0 37996 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_413
timestamp 1676037725
transform 1 0 39100 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_419
timestamp 1676037725
transform 1 0 39652 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_421
timestamp 1676037725
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_433
timestamp 1676037725
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_445
timestamp 1676037725
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_457
timestamp 1676037725
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_469
timestamp 1676037725
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_475
timestamp 1676037725
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_477
timestamp 1676037725
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_489
timestamp 1676037725
transform 1 0 46092 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_501
timestamp 1676037725
transform 1 0 47196 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_513
timestamp 1676037725
transform 1 0 48300 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_525
timestamp 1676037725
transform 1 0 49404 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_531
timestamp 1676037725
transform 1 0 49956 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_533
timestamp 1676037725
transform 1 0 50140 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_545
timestamp 1676037725
transform 1 0 51244 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_557
timestamp 1676037725
transform 1 0 52348 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_569
timestamp 1676037725
transform 1 0 53452 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_581
timestamp 1676037725
transform 1 0 54556 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_587
timestamp 1676037725
transform 1 0 55108 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_589
timestamp 1676037725
transform 1 0 55292 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_601
timestamp 1676037725
transform 1 0 56396 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_613
timestamp 1676037725
transform 1 0 57500 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_74_623
timestamp 1676037725
transform 1 0 58420 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_75_3
timestamp 1676037725
transform 1 0 1380 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_9
timestamp 1676037725
transform 1 0 1932 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_21
timestamp 1676037725
transform 1 0 3036 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_33
timestamp 1676037725
transform 1 0 4140 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_45
timestamp 1676037725
transform 1 0 5244 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_75_53
timestamp 1676037725
transform 1 0 5980 0 -1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1676037725
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_69
timestamp 1676037725
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_81
timestamp 1676037725
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_93
timestamp 1676037725
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1676037725
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1676037725
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_113
timestamp 1676037725
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_125
timestamp 1676037725
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_137
timestamp 1676037725
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_149
timestamp 1676037725
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1676037725
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1676037725
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_169
timestamp 1676037725
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_181
timestamp 1676037725
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_193
timestamp 1676037725
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_205
timestamp 1676037725
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1676037725
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1676037725
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_225
timestamp 1676037725
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_237
timestamp 1676037725
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_249
timestamp 1676037725
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_261
timestamp 1676037725
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_273
timestamp 1676037725
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_279
timestamp 1676037725
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_281
timestamp 1676037725
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_293
timestamp 1676037725
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_305
timestamp 1676037725
transform 1 0 29164 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_317
timestamp 1676037725
transform 1 0 30268 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_329
timestamp 1676037725
transform 1 0 31372 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 1676037725
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_337
timestamp 1676037725
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_349
timestamp 1676037725
transform 1 0 33212 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_361
timestamp 1676037725
transform 1 0 34316 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_373
timestamp 1676037725
transform 1 0 35420 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_385
timestamp 1676037725
transform 1 0 36524 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_391
timestamp 1676037725
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_393
timestamp 1676037725
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_405
timestamp 1676037725
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_417
timestamp 1676037725
transform 1 0 39468 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_429
timestamp 1676037725
transform 1 0 40572 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_441
timestamp 1676037725
transform 1 0 41676 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_447
timestamp 1676037725
transform 1 0 42228 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_449
timestamp 1676037725
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_461
timestamp 1676037725
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_473
timestamp 1676037725
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_485
timestamp 1676037725
transform 1 0 45724 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_497
timestamp 1676037725
transform 1 0 46828 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_503
timestamp 1676037725
transform 1 0 47380 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_505
timestamp 1676037725
transform 1 0 47564 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_517
timestamp 1676037725
transform 1 0 48668 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_529
timestamp 1676037725
transform 1 0 49772 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_541
timestamp 1676037725
transform 1 0 50876 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_553
timestamp 1676037725
transform 1 0 51980 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_559
timestamp 1676037725
transform 1 0 52532 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_561
timestamp 1676037725
transform 1 0 52716 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_573
timestamp 1676037725
transform 1 0 53820 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_585
timestamp 1676037725
transform 1 0 54924 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_597
timestamp 1676037725
transform 1 0 56028 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_609
timestamp 1676037725
transform 1 0 57132 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_615
timestamp 1676037725
transform 1 0 57684 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_75_617
timestamp 1676037725
transform 1 0 57868 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_75_623
timestamp 1676037725
transform 1 0 58420 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_3
timestamp 1676037725
transform 1 0 1380 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_9
timestamp 1676037725
transform 1 0 1932 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_21
timestamp 1676037725
transform 1 0 3036 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1676037725
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1676037725
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1676037725
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_53
timestamp 1676037725
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_65
timestamp 1676037725
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1676037725
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1676037725
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_85
timestamp 1676037725
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_97
timestamp 1676037725
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_109
timestamp 1676037725
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_121
timestamp 1676037725
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1676037725
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1676037725
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_141
timestamp 1676037725
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_153
timestamp 1676037725
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_165
timestamp 1676037725
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_177
timestamp 1676037725
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1676037725
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1676037725
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_197
timestamp 1676037725
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_209
timestamp 1676037725
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_221
timestamp 1676037725
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_233
timestamp 1676037725
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1676037725
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1676037725
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_253
timestamp 1676037725
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_265
timestamp 1676037725
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_277
timestamp 1676037725
transform 1 0 26588 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_289
timestamp 1676037725
transform 1 0 27692 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_301
timestamp 1676037725
transform 1 0 28796 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_307
timestamp 1676037725
transform 1 0 29348 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_309
timestamp 1676037725
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_321
timestamp 1676037725
transform 1 0 30636 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_333
timestamp 1676037725
transform 1 0 31740 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_345
timestamp 1676037725
transform 1 0 32844 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_357
timestamp 1676037725
transform 1 0 33948 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_363
timestamp 1676037725
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_365
timestamp 1676037725
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_377
timestamp 1676037725
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_389
timestamp 1676037725
transform 1 0 36892 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_401
timestamp 1676037725
transform 1 0 37996 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_413
timestamp 1676037725
transform 1 0 39100 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_419
timestamp 1676037725
transform 1 0 39652 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_421
timestamp 1676037725
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_433
timestamp 1676037725
transform 1 0 40940 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_444
timestamp 1676037725
transform 1 0 41952 0 1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_76_455
timestamp 1676037725
transform 1 0 42964 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_467
timestamp 1676037725
transform 1 0 44068 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_76_475
timestamp 1676037725
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_477
timestamp 1676037725
transform 1 0 44988 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_489
timestamp 1676037725
transform 1 0 46092 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_501
timestamp 1676037725
transform 1 0 47196 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_513
timestamp 1676037725
transform 1 0 48300 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_525
timestamp 1676037725
transform 1 0 49404 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_531
timestamp 1676037725
transform 1 0 49956 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_533
timestamp 1676037725
transform 1 0 50140 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_545
timestamp 1676037725
transform 1 0 51244 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_557
timestamp 1676037725
transform 1 0 52348 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_569
timestamp 1676037725
transform 1 0 53452 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_581
timestamp 1676037725
transform 1 0 54556 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_587
timestamp 1676037725
transform 1 0 55108 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_589
timestamp 1676037725
transform 1 0 55292 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_601
timestamp 1676037725
transform 1 0 56396 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_613
timestamp 1676037725
transform 1 0 57500 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_76_623
timestamp 1676037725
transform 1 0 58420 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_3
timestamp 1676037725
transform 1 0 1380 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_77_9
timestamp 1676037725
transform 1 0 1932 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_21
timestamp 1676037725
transform 1 0 3036 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_33
timestamp 1676037725
transform 1 0 4140 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_45
timestamp 1676037725
transform 1 0 5244 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_77_53
timestamp 1676037725
transform 1 0 5980 0 -1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_77_57
timestamp 1676037725
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_69
timestamp 1676037725
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_81
timestamp 1676037725
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_93
timestamp 1676037725
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1676037725
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1676037725
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_113
timestamp 1676037725
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_125
timestamp 1676037725
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_137
timestamp 1676037725
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_149
timestamp 1676037725
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1676037725
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1676037725
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_169
timestamp 1676037725
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_181
timestamp 1676037725
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_193
timestamp 1676037725
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_205
timestamp 1676037725
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1676037725
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1676037725
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_225
timestamp 1676037725
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_237
timestamp 1676037725
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_249
timestamp 1676037725
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_261
timestamp 1676037725
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_273
timestamp 1676037725
transform 1 0 26220 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_279
timestamp 1676037725
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_281
timestamp 1676037725
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_293
timestamp 1676037725
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_305
timestamp 1676037725
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_317
timestamp 1676037725
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_329
timestamp 1676037725
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_335
timestamp 1676037725
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_337
timestamp 1676037725
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_349
timestamp 1676037725
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_361
timestamp 1676037725
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_373
timestamp 1676037725
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_385
timestamp 1676037725
transform 1 0 36524 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_391
timestamp 1676037725
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_393
timestamp 1676037725
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_405
timestamp 1676037725
transform 1 0 38364 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_417
timestamp 1676037725
transform 1 0 39468 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_429
timestamp 1676037725
transform 1 0 40572 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_77_446
timestamp 1676037725
transform 1 0 42136 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_77_449
timestamp 1676037725
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_461
timestamp 1676037725
transform 1 0 43516 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_473
timestamp 1676037725
transform 1 0 44620 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_485
timestamp 1676037725
transform 1 0 45724 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_497
timestamp 1676037725
transform 1 0 46828 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_503
timestamp 1676037725
transform 1 0 47380 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_505
timestamp 1676037725
transform 1 0 47564 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_517
timestamp 1676037725
transform 1 0 48668 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_529
timestamp 1676037725
transform 1 0 49772 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_541
timestamp 1676037725
transform 1 0 50876 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_553
timestamp 1676037725
transform 1 0 51980 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_559
timestamp 1676037725
transform 1 0 52532 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_561
timestamp 1676037725
transform 1 0 52716 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_573
timestamp 1676037725
transform 1 0 53820 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_585
timestamp 1676037725
transform 1 0 54924 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_597
timestamp 1676037725
transform 1 0 56028 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_609
timestamp 1676037725
transform 1 0 57132 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_615
timestamp 1676037725
transform 1 0 57684 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_77_617
timestamp 1676037725
transform 1 0 57868 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_623
timestamp 1676037725
transform 1 0 58420 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_3
timestamp 1676037725
transform 1 0 1380 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_9
timestamp 1676037725
transform 1 0 1932 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_21
timestamp 1676037725
transform 1 0 3036 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1676037725
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1676037725
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_41
timestamp 1676037725
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_53
timestamp 1676037725
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_65
timestamp 1676037725
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1676037725
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1676037725
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_85
timestamp 1676037725
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_97
timestamp 1676037725
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_109
timestamp 1676037725
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_121
timestamp 1676037725
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1676037725
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1676037725
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_141
timestamp 1676037725
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_153
timestamp 1676037725
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_165
timestamp 1676037725
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_177
timestamp 1676037725
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1676037725
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1676037725
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_197
timestamp 1676037725
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_209
timestamp 1676037725
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_221
timestamp 1676037725
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_233
timestamp 1676037725
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1676037725
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1676037725
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_253
timestamp 1676037725
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_265
timestamp 1676037725
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_277
timestamp 1676037725
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_289
timestamp 1676037725
transform 1 0 27692 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_301
timestamp 1676037725
transform 1 0 28796 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_307
timestamp 1676037725
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_309
timestamp 1676037725
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_321
timestamp 1676037725
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_333
timestamp 1676037725
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_345
timestamp 1676037725
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_357
timestamp 1676037725
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_363
timestamp 1676037725
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_365
timestamp 1676037725
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_377
timestamp 1676037725
transform 1 0 35788 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_389
timestamp 1676037725
transform 1 0 36892 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_401
timestamp 1676037725
transform 1 0 37996 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_413
timestamp 1676037725
transform 1 0 39100 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_419
timestamp 1676037725
transform 1 0 39652 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_421
timestamp 1676037725
transform 1 0 39836 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_433
timestamp 1676037725
transform 1 0 40940 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_445
timestamp 1676037725
transform 1 0 42044 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_457
timestamp 1676037725
transform 1 0 43148 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_469
timestamp 1676037725
transform 1 0 44252 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_475
timestamp 1676037725
transform 1 0 44804 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_477
timestamp 1676037725
transform 1 0 44988 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_489
timestamp 1676037725
transform 1 0 46092 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_501
timestamp 1676037725
transform 1 0 47196 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_513
timestamp 1676037725
transform 1 0 48300 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_528
timestamp 1676037725
transform 1 0 49680 0 1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_78_533
timestamp 1676037725
transform 1 0 50140 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_545
timestamp 1676037725
transform 1 0 51244 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_557
timestamp 1676037725
transform 1 0 52348 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_569
timestamp 1676037725
transform 1 0 53452 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_581
timestamp 1676037725
transform 1 0 54556 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_587
timestamp 1676037725
transform 1 0 55108 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_589
timestamp 1676037725
transform 1 0 55292 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_601
timestamp 1676037725
transform 1 0 56396 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_78_613
timestamp 1676037725
transform 1 0 57500 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_78_623
timestamp 1676037725
transform 1 0 58420 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_3
timestamp 1676037725
transform 1 0 1380 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_9
timestamp 1676037725
transform 1 0 1932 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_21
timestamp 1676037725
transform 1 0 3036 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_33
timestamp 1676037725
transform 1 0 4140 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_45
timestamp 1676037725
transform 1 0 5244 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_79_53
timestamp 1676037725
transform 1 0 5980 0 -1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 1676037725
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_69
timestamp 1676037725
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_81
timestamp 1676037725
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_93
timestamp 1676037725
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1676037725
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1676037725
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_113
timestamp 1676037725
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_125
timestamp 1676037725
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_137
timestamp 1676037725
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_149
timestamp 1676037725
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_161
timestamp 1676037725
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1676037725
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_169
timestamp 1676037725
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_181
timestamp 1676037725
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_193
timestamp 1676037725
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_205
timestamp 1676037725
transform 1 0 19964 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_217
timestamp 1676037725
transform 1 0 21068 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1676037725
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_225
timestamp 1676037725
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_237
timestamp 1676037725
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_249
timestamp 1676037725
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_261
timestamp 1676037725
transform 1 0 25116 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_273
timestamp 1676037725
transform 1 0 26220 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_279
timestamp 1676037725
transform 1 0 26772 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_281
timestamp 1676037725
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_293
timestamp 1676037725
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_305
timestamp 1676037725
transform 1 0 29164 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_317
timestamp 1676037725
transform 1 0 30268 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_329
timestamp 1676037725
transform 1 0 31372 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_335
timestamp 1676037725
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_79_337
timestamp 1676037725
transform 1 0 32108 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_347
timestamp 1676037725
transform 1 0 33028 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_359
timestamp 1676037725
transform 1 0 34132 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_367
timestamp 1676037725
transform 1 0 34868 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_79_370
timestamp 1676037725
transform 1 0 35144 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_379
timestamp 1676037725
transform 1 0 35972 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_79_391
timestamp 1676037725
transform 1 0 37076 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_393
timestamp 1676037725
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_405
timestamp 1676037725
transform 1 0 38364 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_417
timestamp 1676037725
transform 1 0 39468 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_429
timestamp 1676037725
transform 1 0 40572 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_441
timestamp 1676037725
transform 1 0 41676 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_447
timestamp 1676037725
transform 1 0 42228 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_449
timestamp 1676037725
transform 1 0 42412 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_461
timestamp 1676037725
transform 1 0 43516 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_473
timestamp 1676037725
transform 1 0 44620 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_485
timestamp 1676037725
transform 1 0 45724 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_497
timestamp 1676037725
transform 1 0 46828 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_503
timestamp 1676037725
transform 1 0 47380 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_505
timestamp 1676037725
transform 1 0 47564 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_517
timestamp 1676037725
transform 1 0 48668 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_529
timestamp 1676037725
transform 1 0 49772 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_541
timestamp 1676037725
transform 1 0 50876 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_553
timestamp 1676037725
transform 1 0 51980 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_559
timestamp 1676037725
transform 1 0 52532 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_561
timestamp 1676037725
transform 1 0 52716 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_573
timestamp 1676037725
transform 1 0 53820 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_585
timestamp 1676037725
transform 1 0 54924 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_597
timestamp 1676037725
transform 1 0 56028 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_609
timestamp 1676037725
transform 1 0 57132 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_615
timestamp 1676037725
transform 1 0 57684 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_79_617
timestamp 1676037725
transform 1 0 57868 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_623
timestamp 1676037725
transform 1 0 58420 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_3
timestamp 1676037725
transform 1 0 1380 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_80_9
timestamp 1676037725
transform 1 0 1932 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_21
timestamp 1676037725
transform 1 0 3036 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1676037725
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1676037725
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_41
timestamp 1676037725
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_53
timestamp 1676037725
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_65
timestamp 1676037725
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1676037725
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1676037725
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_85
timestamp 1676037725
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_97
timestamp 1676037725
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_109
timestamp 1676037725
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_121
timestamp 1676037725
transform 1 0 12236 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_133
timestamp 1676037725
transform 1 0 13340 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1676037725
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_141
timestamp 1676037725
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_153
timestamp 1676037725
transform 1 0 15180 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_165
timestamp 1676037725
transform 1 0 16284 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_177
timestamp 1676037725
transform 1 0 17388 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_189
timestamp 1676037725
transform 1 0 18492 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_195
timestamp 1676037725
transform 1 0 19044 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_197
timestamp 1676037725
transform 1 0 19228 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_209
timestamp 1676037725
transform 1 0 20332 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_221
timestamp 1676037725
transform 1 0 21436 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_233
timestamp 1676037725
transform 1 0 22540 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_245
timestamp 1676037725
transform 1 0 23644 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_251
timestamp 1676037725
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_253
timestamp 1676037725
transform 1 0 24380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_265
timestamp 1676037725
transform 1 0 25484 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_277
timestamp 1676037725
transform 1 0 26588 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_289
timestamp 1676037725
transform 1 0 27692 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_301
timestamp 1676037725
transform 1 0 28796 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_307
timestamp 1676037725
transform 1 0 29348 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_309
timestamp 1676037725
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_321
timestamp 1676037725
transform 1 0 30636 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_333
timestamp 1676037725
transform 1 0 31740 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_345
timestamp 1676037725
transform 1 0 32844 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_357
timestamp 1676037725
transform 1 0 33948 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_363
timestamp 1676037725
transform 1 0 34500 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_365
timestamp 1676037725
transform 1 0 34684 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_377
timestamp 1676037725
transform 1 0 35788 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_383
timestamp 1676037725
transform 1 0 36340 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_391
timestamp 1676037725
transform 1 0 37076 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_403
timestamp 1676037725
transform 1 0 38180 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_415
timestamp 1676037725
transform 1 0 39284 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_419
timestamp 1676037725
transform 1 0 39652 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_421
timestamp 1676037725
transform 1 0 39836 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_433
timestamp 1676037725
transform 1 0 40940 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_445
timestamp 1676037725
transform 1 0 42044 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_457
timestamp 1676037725
transform 1 0 43148 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_469
timestamp 1676037725
transform 1 0 44252 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_475
timestamp 1676037725
transform 1 0 44804 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_477
timestamp 1676037725
transform 1 0 44988 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_489
timestamp 1676037725
transform 1 0 46092 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_501
timestamp 1676037725
transform 1 0 47196 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_513
timestamp 1676037725
transform 1 0 48300 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_525
timestamp 1676037725
transform 1 0 49404 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_531
timestamp 1676037725
transform 1 0 49956 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_533
timestamp 1676037725
transform 1 0 50140 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_545
timestamp 1676037725
transform 1 0 51244 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_557
timestamp 1676037725
transform 1 0 52348 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_569
timestamp 1676037725
transform 1 0 53452 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_581
timestamp 1676037725
transform 1 0 54556 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_587
timestamp 1676037725
transform 1 0 55108 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_589
timestamp 1676037725
transform 1 0 55292 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_601
timestamp 1676037725
transform 1 0 56396 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_613
timestamp 1676037725
transform 1 0 57500 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_623
timestamp 1676037725
transform 1 0 58420 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_3
timestamp 1676037725
transform 1 0 1380 0 -1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_81_9
timestamp 1676037725
transform 1 0 1932 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_21
timestamp 1676037725
transform 1 0 3036 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_33
timestamp 1676037725
transform 1 0 4140 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_45
timestamp 1676037725
transform 1 0 5244 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_81_53
timestamp 1676037725
transform 1 0 5980 0 -1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_81_57
timestamp 1676037725
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_69
timestamp 1676037725
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_81
timestamp 1676037725
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_93
timestamp 1676037725
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_105
timestamp 1676037725
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1676037725
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_113
timestamp 1676037725
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_125
timestamp 1676037725
transform 1 0 12604 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_137
timestamp 1676037725
transform 1 0 13708 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_149
timestamp 1676037725
transform 1 0 14812 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_161
timestamp 1676037725
transform 1 0 15916 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1676037725
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_169
timestamp 1676037725
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_181
timestamp 1676037725
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_193
timestamp 1676037725
transform 1 0 18860 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_205
timestamp 1676037725
transform 1 0 19964 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_217
timestamp 1676037725
transform 1 0 21068 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_223
timestamp 1676037725
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_225
timestamp 1676037725
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_237
timestamp 1676037725
transform 1 0 22908 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_249
timestamp 1676037725
transform 1 0 24012 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_261
timestamp 1676037725
transform 1 0 25116 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_273
timestamp 1676037725
transform 1 0 26220 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_279
timestamp 1676037725
transform 1 0 26772 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_281
timestamp 1676037725
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_293
timestamp 1676037725
transform 1 0 28060 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_305
timestamp 1676037725
transform 1 0 29164 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_317
timestamp 1676037725
transform 1 0 30268 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_329
timestamp 1676037725
transform 1 0 31372 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_335
timestamp 1676037725
transform 1 0 31924 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_81_337
timestamp 1676037725
transform 1 0 32108 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_346
timestamp 1676037725
transform 1 0 32936 0 -1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_81_350
timestamp 1676037725
transform 1 0 33304 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_362
timestamp 1676037725
transform 1 0 34408 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_374
timestamp 1676037725
transform 1 0 35512 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_386
timestamp 1676037725
transform 1 0 36616 0 -1 46784
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_81_393
timestamp 1676037725
transform 1 0 37260 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_405
timestamp 1676037725
transform 1 0 38364 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_417
timestamp 1676037725
transform 1 0 39468 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_429
timestamp 1676037725
transform 1 0 40572 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_441
timestamp 1676037725
transform 1 0 41676 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_447
timestamp 1676037725
transform 1 0 42228 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_449
timestamp 1676037725
transform 1 0 42412 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_461
timestamp 1676037725
transform 1 0 43516 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_473
timestamp 1676037725
transform 1 0 44620 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_485
timestamp 1676037725
transform 1 0 45724 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_497
timestamp 1676037725
transform 1 0 46828 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_503
timestamp 1676037725
transform 1 0 47380 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_505
timestamp 1676037725
transform 1 0 47564 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_517
timestamp 1676037725
transform 1 0 48668 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_529
timestamp 1676037725
transform 1 0 49772 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_541
timestamp 1676037725
transform 1 0 50876 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_553
timestamp 1676037725
transform 1 0 51980 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_559
timestamp 1676037725
transform 1 0 52532 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_561
timestamp 1676037725
transform 1 0 52716 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_573
timestamp 1676037725
transform 1 0 53820 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_585
timestamp 1676037725
transform 1 0 54924 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_597
timestamp 1676037725
transform 1 0 56028 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_609
timestamp 1676037725
transform 1 0 57132 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_615
timestamp 1676037725
transform 1 0 57684 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_81_617
timestamp 1676037725
transform 1 0 57868 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_623
timestamp 1676037725
transform 1 0 58420 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_3
timestamp 1676037725
transform 1 0 1380 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_9
timestamp 1676037725
transform 1 0 1932 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_21
timestamp 1676037725
transform 1 0 3036 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1676037725
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_29
timestamp 1676037725
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_41
timestamp 1676037725
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_53
timestamp 1676037725
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_65
timestamp 1676037725
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_77
timestamp 1676037725
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1676037725
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_85
timestamp 1676037725
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_97
timestamp 1676037725
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_109
timestamp 1676037725
transform 1 0 11132 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_121
timestamp 1676037725
transform 1 0 12236 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_133
timestamp 1676037725
transform 1 0 13340 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_139
timestamp 1676037725
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_141
timestamp 1676037725
transform 1 0 14076 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_153
timestamp 1676037725
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_165
timestamp 1676037725
transform 1 0 16284 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_177
timestamp 1676037725
transform 1 0 17388 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_189
timestamp 1676037725
transform 1 0 18492 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_195
timestamp 1676037725
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_197
timestamp 1676037725
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_209
timestamp 1676037725
transform 1 0 20332 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_221
timestamp 1676037725
transform 1 0 21436 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_233
timestamp 1676037725
transform 1 0 22540 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_245
timestamp 1676037725
transform 1 0 23644 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_251
timestamp 1676037725
transform 1 0 24196 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_253
timestamp 1676037725
transform 1 0 24380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_265
timestamp 1676037725
transform 1 0 25484 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_277
timestamp 1676037725
transform 1 0 26588 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_289
timestamp 1676037725
transform 1 0 27692 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_301
timestamp 1676037725
transform 1 0 28796 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_307
timestamp 1676037725
transform 1 0 29348 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_309
timestamp 1676037725
transform 1 0 29532 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_321
timestamp 1676037725
transform 1 0 30636 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_333
timestamp 1676037725
transform 1 0 31740 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_345
timestamp 1676037725
transform 1 0 32844 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_357
timestamp 1676037725
transform 1 0 33948 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_363
timestamp 1676037725
transform 1 0 34500 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_365
timestamp 1676037725
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_377
timestamp 1676037725
transform 1 0 35788 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_389
timestamp 1676037725
transform 1 0 36892 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_401
timestamp 1676037725
transform 1 0 37996 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_413
timestamp 1676037725
transform 1 0 39100 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_419
timestamp 1676037725
transform 1 0 39652 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_421
timestamp 1676037725
transform 1 0 39836 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_433
timestamp 1676037725
transform 1 0 40940 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_445
timestamp 1676037725
transform 1 0 42044 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_457
timestamp 1676037725
transform 1 0 43148 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_469
timestamp 1676037725
transform 1 0 44252 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_475
timestamp 1676037725
transform 1 0 44804 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_477
timestamp 1676037725
transform 1 0 44988 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_489
timestamp 1676037725
transform 1 0 46092 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_501
timestamp 1676037725
transform 1 0 47196 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_513
timestamp 1676037725
transform 1 0 48300 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_525
timestamp 1676037725
transform 1 0 49404 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_531
timestamp 1676037725
transform 1 0 49956 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_533
timestamp 1676037725
transform 1 0 50140 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_545
timestamp 1676037725
transform 1 0 51244 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_557
timestamp 1676037725
transform 1 0 52348 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_569
timestamp 1676037725
transform 1 0 53452 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_581
timestamp 1676037725
transform 1 0 54556 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_587
timestamp 1676037725
transform 1 0 55108 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_589
timestamp 1676037725
transform 1 0 55292 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_601
timestamp 1676037725
transform 1 0 56396 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_613
timestamp 1676037725
transform 1 0 57500 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_82_623
timestamp 1676037725
transform 1 0 58420 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_83_3
timestamp 1676037725
transform 1 0 1380 0 -1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_83_9
timestamp 1676037725
transform 1 0 1932 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_21
timestamp 1676037725
transform 1 0 3036 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_33
timestamp 1676037725
transform 1 0 4140 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_45
timestamp 1676037725
transform 1 0 5244 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_83_53
timestamp 1676037725
transform 1 0 5980 0 -1 47872
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_83_57
timestamp 1676037725
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_69
timestamp 1676037725
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_81
timestamp 1676037725
transform 1 0 8556 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_93
timestamp 1676037725
transform 1 0 9660 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_105
timestamp 1676037725
transform 1 0 10764 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_111
timestamp 1676037725
transform 1 0 11316 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_113
timestamp 1676037725
transform 1 0 11500 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_125
timestamp 1676037725
transform 1 0 12604 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_137
timestamp 1676037725
transform 1 0 13708 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_149
timestamp 1676037725
transform 1 0 14812 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_161
timestamp 1676037725
transform 1 0 15916 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_167
timestamp 1676037725
transform 1 0 16468 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_169
timestamp 1676037725
transform 1 0 16652 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_181
timestamp 1676037725
transform 1 0 17756 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_193
timestamp 1676037725
transform 1 0 18860 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_205
timestamp 1676037725
transform 1 0 19964 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_217
timestamp 1676037725
transform 1 0 21068 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_223
timestamp 1676037725
transform 1 0 21620 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_225
timestamp 1676037725
transform 1 0 21804 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_237
timestamp 1676037725
transform 1 0 22908 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_249
timestamp 1676037725
transform 1 0 24012 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_261
timestamp 1676037725
transform 1 0 25116 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_273
timestamp 1676037725
transform 1 0 26220 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_279
timestamp 1676037725
transform 1 0 26772 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_281
timestamp 1676037725
transform 1 0 26956 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_293
timestamp 1676037725
transform 1 0 28060 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_305
timestamp 1676037725
transform 1 0 29164 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_317
timestamp 1676037725
transform 1 0 30268 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_321
timestamp 1676037725
transform 1 0 30636 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_83_330
timestamp 1676037725
transform 1 0 31464 0 -1 47872
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_83_337
timestamp 1676037725
transform 1 0 32108 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_349
timestamp 1676037725
transform 1 0 33212 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_361
timestamp 1676037725
transform 1 0 34316 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_373
timestamp 1676037725
transform 1 0 35420 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_385
timestamp 1676037725
transform 1 0 36524 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_391
timestamp 1676037725
transform 1 0 37076 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_393
timestamp 1676037725
transform 1 0 37260 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_405
timestamp 1676037725
transform 1 0 38364 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_417
timestamp 1676037725
transform 1 0 39468 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_429
timestamp 1676037725
transform 1 0 40572 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_83_435
timestamp 1676037725
transform 1 0 41124 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_83_446
timestamp 1676037725
transform 1 0 42136 0 -1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_83_449
timestamp 1676037725
transform 1 0 42412 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_461
timestamp 1676037725
transform 1 0 43516 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_473
timestamp 1676037725
transform 1 0 44620 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_485
timestamp 1676037725
transform 1 0 45724 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_497
timestamp 1676037725
transform 1 0 46828 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_503
timestamp 1676037725
transform 1 0 47380 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_505
timestamp 1676037725
transform 1 0 47564 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_517
timestamp 1676037725
transform 1 0 48668 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_529
timestamp 1676037725
transform 1 0 49772 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_541
timestamp 1676037725
transform 1 0 50876 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_553
timestamp 1676037725
transform 1 0 51980 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_559
timestamp 1676037725
transform 1 0 52532 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_561
timestamp 1676037725
transform 1 0 52716 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_573
timestamp 1676037725
transform 1 0 53820 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_585
timestamp 1676037725
transform 1 0 54924 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_597
timestamp 1676037725
transform 1 0 56028 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_83_609
timestamp 1676037725
transform 1 0 57132 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_83_614
timestamp 1676037725
transform 1 0 57592 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_83_617
timestamp 1676037725
transform 1 0 57868 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_83_623
timestamp 1676037725
transform 1 0 58420 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_84_3
timestamp 1676037725
transform 1 0 1380 0 1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_84_9
timestamp 1676037725
transform 1 0 1932 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_21
timestamp 1676037725
transform 1 0 3036 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_27
timestamp 1676037725
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_29
timestamp 1676037725
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_41
timestamp 1676037725
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_53
timestamp 1676037725
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_65
timestamp 1676037725
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_77
timestamp 1676037725
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 1676037725
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_85
timestamp 1676037725
transform 1 0 8924 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_97
timestamp 1676037725
transform 1 0 10028 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_109
timestamp 1676037725
transform 1 0 11132 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_121
timestamp 1676037725
transform 1 0 12236 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_133
timestamp 1676037725
transform 1 0 13340 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_139
timestamp 1676037725
transform 1 0 13892 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_141
timestamp 1676037725
transform 1 0 14076 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_153
timestamp 1676037725
transform 1 0 15180 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_165
timestamp 1676037725
transform 1 0 16284 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_177
timestamp 1676037725
transform 1 0 17388 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_189
timestamp 1676037725
transform 1 0 18492 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_195
timestamp 1676037725
transform 1 0 19044 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_197
timestamp 1676037725
transform 1 0 19228 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_209
timestamp 1676037725
transform 1 0 20332 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_221
timestamp 1676037725
transform 1 0 21436 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_233
timestamp 1676037725
transform 1 0 22540 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_245
timestamp 1676037725
transform 1 0 23644 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_251
timestamp 1676037725
transform 1 0 24196 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_253
timestamp 1676037725
transform 1 0 24380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_265
timestamp 1676037725
transform 1 0 25484 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_277
timestamp 1676037725
transform 1 0 26588 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_289
timestamp 1676037725
transform 1 0 27692 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_301
timestamp 1676037725
transform 1 0 28796 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_307
timestamp 1676037725
transform 1 0 29348 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_309
timestamp 1676037725
transform 1 0 29532 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_84_321
timestamp 1676037725
transform 1 0 30636 0 1 47872
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_84_334
timestamp 1676037725
transform 1 0 31832 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_346
timestamp 1676037725
transform 1 0 32936 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_358
timestamp 1676037725
transform 1 0 34040 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_84_365
timestamp 1676037725
transform 1 0 34684 0 1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_84_374
timestamp 1676037725
transform 1 0 35512 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_386
timestamp 1676037725
transform 1 0 36616 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_398
timestamp 1676037725
transform 1 0 37720 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_410
timestamp 1676037725
transform 1 0 38824 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_84_418
timestamp 1676037725
transform 1 0 39560 0 1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_84_421
timestamp 1676037725
transform 1 0 39836 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_433
timestamp 1676037725
transform 1 0 40940 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_445
timestamp 1676037725
transform 1 0 42044 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_457
timestamp 1676037725
transform 1 0 43148 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_469
timestamp 1676037725
transform 1 0 44252 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_475
timestamp 1676037725
transform 1 0 44804 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_477
timestamp 1676037725
transform 1 0 44988 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_489
timestamp 1676037725
transform 1 0 46092 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_501
timestamp 1676037725
transform 1 0 47196 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_513
timestamp 1676037725
transform 1 0 48300 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_525
timestamp 1676037725
transform 1 0 49404 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_531
timestamp 1676037725
transform 1 0 49956 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_533
timestamp 1676037725
transform 1 0 50140 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_545
timestamp 1676037725
transform 1 0 51244 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_557
timestamp 1676037725
transform 1 0 52348 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_569
timestamp 1676037725
transform 1 0 53452 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_581
timestamp 1676037725
transform 1 0 54556 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_587
timestamp 1676037725
transform 1 0 55108 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_589
timestamp 1676037725
transform 1 0 55292 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_601
timestamp 1676037725
transform 1 0 56396 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_84_613
timestamp 1676037725
transform 1 0 57500 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_84_623
timestamp 1676037725
transform 1 0 58420 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_85_3
timestamp 1676037725
transform 1 0 1380 0 -1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_85_9
timestamp 1676037725
transform 1 0 1932 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_21
timestamp 1676037725
transform 1 0 3036 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_33
timestamp 1676037725
transform 1 0 4140 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_85_45
timestamp 1676037725
transform 1 0 5244 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_85_53
timestamp 1676037725
transform 1 0 5980 0 -1 48960
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_85_57
timestamp 1676037725
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_69
timestamp 1676037725
transform 1 0 7452 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_81
timestamp 1676037725
transform 1 0 8556 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_85_93
timestamp 1676037725
transform 1 0 9660 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_85_104
timestamp 1676037725
transform 1 0 10672 0 -1 48960
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_85_113
timestamp 1676037725
transform 1 0 11500 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_125
timestamp 1676037725
transform 1 0 12604 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_137
timestamp 1676037725
transform 1 0 13708 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_149
timestamp 1676037725
transform 1 0 14812 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_161
timestamp 1676037725
transform 1 0 15916 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_167
timestamp 1676037725
transform 1 0 16468 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_169
timestamp 1676037725
transform 1 0 16652 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_181
timestamp 1676037725
transform 1 0 17756 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_193
timestamp 1676037725
transform 1 0 18860 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_205
timestamp 1676037725
transform 1 0 19964 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_217
timestamp 1676037725
transform 1 0 21068 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_223
timestamp 1676037725
transform 1 0 21620 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_225
timestamp 1676037725
transform 1 0 21804 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_237
timestamp 1676037725
transform 1 0 22908 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_249
timestamp 1676037725
transform 1 0 24012 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_261
timestamp 1676037725
transform 1 0 25116 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_273
timestamp 1676037725
transform 1 0 26220 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_279
timestamp 1676037725
transform 1 0 26772 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_281
timestamp 1676037725
transform 1 0 26956 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_293
timestamp 1676037725
transform 1 0 28060 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_305
timestamp 1676037725
transform 1 0 29164 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_85_334
timestamp 1676037725
transform 1 0 31832 0 -1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_85_337
timestamp 1676037725
transform 1 0 32108 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_349
timestamp 1676037725
transform 1 0 33212 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_361
timestamp 1676037725
transform 1 0 34316 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_373
timestamp 1676037725
transform 1 0 35420 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_385
timestamp 1676037725
transform 1 0 36524 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_391
timestamp 1676037725
transform 1 0 37076 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_393
timestamp 1676037725
transform 1 0 37260 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_405
timestamp 1676037725
transform 1 0 38364 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_417
timestamp 1676037725
transform 1 0 39468 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_429
timestamp 1676037725
transform 1 0 40572 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_441
timestamp 1676037725
transform 1 0 41676 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_447
timestamp 1676037725
transform 1 0 42228 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_449
timestamp 1676037725
transform 1 0 42412 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_461
timestamp 1676037725
transform 1 0 43516 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_473
timestamp 1676037725
transform 1 0 44620 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_485
timestamp 1676037725
transform 1 0 45724 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_497
timestamp 1676037725
transform 1 0 46828 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_503
timestamp 1676037725
transform 1 0 47380 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_505
timestamp 1676037725
transform 1 0 47564 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_517
timestamp 1676037725
transform 1 0 48668 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_529
timestamp 1676037725
transform 1 0 49772 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_541
timestamp 1676037725
transform 1 0 50876 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_553
timestamp 1676037725
transform 1 0 51980 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_559
timestamp 1676037725
transform 1 0 52532 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_561
timestamp 1676037725
transform 1 0 52716 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_573
timestamp 1676037725
transform 1 0 53820 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_585
timestamp 1676037725
transform 1 0 54924 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_597
timestamp 1676037725
transform 1 0 56028 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_609
timestamp 1676037725
transform 1 0 57132 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_615
timestamp 1676037725
transform 1 0 57684 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_85_617
timestamp 1676037725
transform 1 0 57868 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_85_623
timestamp 1676037725
transform 1 0 58420 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_86_3
timestamp 1676037725
transform 1 0 1380 0 1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_86_11
timestamp 1676037725
transform 1 0 2116 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_23
timestamp 1676037725
transform 1 0 3220 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 1676037725
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_29
timestamp 1676037725
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_41
timestamp 1676037725
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_53
timestamp 1676037725
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_65
timestamp 1676037725
transform 1 0 7084 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_77
timestamp 1676037725
transform 1 0 8188 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_83
timestamp 1676037725
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_85
timestamp 1676037725
transform 1 0 8924 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_97
timestamp 1676037725
transform 1 0 10028 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_109
timestamp 1676037725
transform 1 0 11132 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_121
timestamp 1676037725
transform 1 0 12236 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_133
timestamp 1676037725
transform 1 0 13340 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_139
timestamp 1676037725
transform 1 0 13892 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_141
timestamp 1676037725
transform 1 0 14076 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_153
timestamp 1676037725
transform 1 0 15180 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_165
timestamp 1676037725
transform 1 0 16284 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_177
timestamp 1676037725
transform 1 0 17388 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_189
timestamp 1676037725
transform 1 0 18492 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_195
timestamp 1676037725
transform 1 0 19044 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_197
timestamp 1676037725
transform 1 0 19228 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_209
timestamp 1676037725
transform 1 0 20332 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_221
timestamp 1676037725
transform 1 0 21436 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_233
timestamp 1676037725
transform 1 0 22540 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_245
timestamp 1676037725
transform 1 0 23644 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_251
timestamp 1676037725
transform 1 0 24196 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_253
timestamp 1676037725
transform 1 0 24380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_265
timestamp 1676037725
transform 1 0 25484 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_277
timestamp 1676037725
transform 1 0 26588 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_289
timestamp 1676037725
transform 1 0 27692 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_301
timestamp 1676037725
transform 1 0 28796 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_307
timestamp 1676037725
transform 1 0 29348 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_86_309
timestamp 1676037725
transform 1 0 29532 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_315
timestamp 1676037725
transform 1 0 30084 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_323
timestamp 1676037725
transform 1 0 30820 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_335
timestamp 1676037725
transform 1 0 31924 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_347
timestamp 1676037725
transform 1 0 33028 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_359
timestamp 1676037725
transform 1 0 34132 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_363
timestamp 1676037725
transform 1 0 34500 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_365
timestamp 1676037725
transform 1 0 34684 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_377
timestamp 1676037725
transform 1 0 35788 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_389
timestamp 1676037725
transform 1 0 36892 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_401
timestamp 1676037725
transform 1 0 37996 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_413
timestamp 1676037725
transform 1 0 39100 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_419
timestamp 1676037725
transform 1 0 39652 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_421
timestamp 1676037725
transform 1 0 39836 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_433
timestamp 1676037725
transform 1 0 40940 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_445
timestamp 1676037725
transform 1 0 42044 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_457
timestamp 1676037725
transform 1 0 43148 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_469
timestamp 1676037725
transform 1 0 44252 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_475
timestamp 1676037725
transform 1 0 44804 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_477
timestamp 1676037725
transform 1 0 44988 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_489
timestamp 1676037725
transform 1 0 46092 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_501
timestamp 1676037725
transform 1 0 47196 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_513
timestamp 1676037725
transform 1 0 48300 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_525
timestamp 1676037725
transform 1 0 49404 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_531
timestamp 1676037725
transform 1 0 49956 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_533
timestamp 1676037725
transform 1 0 50140 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_545
timestamp 1676037725
transform 1 0 51244 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_557
timestamp 1676037725
transform 1 0 52348 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_569
timestamp 1676037725
transform 1 0 53452 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_581
timestamp 1676037725
transform 1 0 54556 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_587
timestamp 1676037725
transform 1 0 55108 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_589
timestamp 1676037725
transform 1 0 55292 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_601
timestamp 1676037725
transform 1 0 56396 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_613
timestamp 1676037725
transform 1 0 57500 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_86_623
timestamp 1676037725
transform 1 0 58420 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_87_3
timestamp 1676037725
transform 1 0 1380 0 -1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_87_11
timestamp 1676037725
transform 1 0 2116 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_23
timestamp 1676037725
transform 1 0 3220 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_35
timestamp 1676037725
transform 1 0 4324 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_87_47
timestamp 1676037725
transform 1 0 5428 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_87_55
timestamp 1676037725
transform 1 0 6164 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_57
timestamp 1676037725
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_69
timestamp 1676037725
transform 1 0 7452 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_81
timestamp 1676037725
transform 1 0 8556 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_93
timestamp 1676037725
transform 1 0 9660 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_105
timestamp 1676037725
transform 1 0 10764 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_111
timestamp 1676037725
transform 1 0 11316 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_113
timestamp 1676037725
transform 1 0 11500 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_125
timestamp 1676037725
transform 1 0 12604 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_137
timestamp 1676037725
transform 1 0 13708 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_149
timestamp 1676037725
transform 1 0 14812 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_161
timestamp 1676037725
transform 1 0 15916 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_167
timestamp 1676037725
transform 1 0 16468 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_169
timestamp 1676037725
transform 1 0 16652 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_181
timestamp 1676037725
transform 1 0 17756 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_193
timestamp 1676037725
transform 1 0 18860 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_205
timestamp 1676037725
transform 1 0 19964 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_217
timestamp 1676037725
transform 1 0 21068 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_223
timestamp 1676037725
transform 1 0 21620 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_225
timestamp 1676037725
transform 1 0 21804 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_237
timestamp 1676037725
transform 1 0 22908 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_249
timestamp 1676037725
transform 1 0 24012 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_261
timestamp 1676037725
transform 1 0 25116 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_273
timestamp 1676037725
transform 1 0 26220 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_279
timestamp 1676037725
transform 1 0 26772 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_281
timestamp 1676037725
transform 1 0 26956 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_293
timestamp 1676037725
transform 1 0 28060 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_305
timestamp 1676037725
transform 1 0 29164 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_317
timestamp 1676037725
transform 1 0 30268 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_329
timestamp 1676037725
transform 1 0 31372 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_335
timestamp 1676037725
transform 1 0 31924 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_337
timestamp 1676037725
transform 1 0 32108 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_349
timestamp 1676037725
transform 1 0 33212 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_361
timestamp 1676037725
transform 1 0 34316 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_373
timestamp 1676037725
transform 1 0 35420 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_385
timestamp 1676037725
transform 1 0 36524 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_391
timestamp 1676037725
transform 1 0 37076 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_393
timestamp 1676037725
transform 1 0 37260 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_405
timestamp 1676037725
transform 1 0 38364 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_417
timestamp 1676037725
transform 1 0 39468 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_429
timestamp 1676037725
transform 1 0 40572 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_441
timestamp 1676037725
transform 1 0 41676 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_447
timestamp 1676037725
transform 1 0 42228 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_87_449
timestamp 1676037725
transform 1 0 42412 0 -1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_87_465
timestamp 1676037725
transform 1 0 43884 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_477
timestamp 1676037725
transform 1 0 44988 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_489
timestamp 1676037725
transform 1 0 46092 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_87_501
timestamp 1676037725
transform 1 0 47196 0 -1 50048
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_87_505
timestamp 1676037725
transform 1 0 47564 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_517
timestamp 1676037725
transform 1 0 48668 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_529
timestamp 1676037725
transform 1 0 49772 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_541
timestamp 1676037725
transform 1 0 50876 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_553
timestamp 1676037725
transform 1 0 51980 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_559
timestamp 1676037725
transform 1 0 52532 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_561
timestamp 1676037725
transform 1 0 52716 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_573
timestamp 1676037725
transform 1 0 53820 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_585
timestamp 1676037725
transform 1 0 54924 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_597
timestamp 1676037725
transform 1 0 56028 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_609
timestamp 1676037725
transform 1 0 57132 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_615
timestamp 1676037725
transform 1 0 57684 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_87_617
timestamp 1676037725
transform 1 0 57868 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_87_623
timestamp 1676037725
transform 1 0 58420 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_88_3
timestamp 1676037725
transform 1 0 1380 0 1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_88_11
timestamp 1676037725
transform 1 0 2116 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_23
timestamp 1676037725
transform 1 0 3220 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_27
timestamp 1676037725
transform 1 0 3588 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_29
timestamp 1676037725
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_41
timestamp 1676037725
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_53
timestamp 1676037725
transform 1 0 5980 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_65
timestamp 1676037725
transform 1 0 7084 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_77
timestamp 1676037725
transform 1 0 8188 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_83
timestamp 1676037725
transform 1 0 8740 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_85
timestamp 1676037725
transform 1 0 8924 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_97
timestamp 1676037725
transform 1 0 10028 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_109
timestamp 1676037725
transform 1 0 11132 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_121
timestamp 1676037725
transform 1 0 12236 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_133
timestamp 1676037725
transform 1 0 13340 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_139
timestamp 1676037725
transform 1 0 13892 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_141
timestamp 1676037725
transform 1 0 14076 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_153
timestamp 1676037725
transform 1 0 15180 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_165
timestamp 1676037725
transform 1 0 16284 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_177
timestamp 1676037725
transform 1 0 17388 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_189
timestamp 1676037725
transform 1 0 18492 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_195
timestamp 1676037725
transform 1 0 19044 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_197
timestamp 1676037725
transform 1 0 19228 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_209
timestamp 1676037725
transform 1 0 20332 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_221
timestamp 1676037725
transform 1 0 21436 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_233
timestamp 1676037725
transform 1 0 22540 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_245
timestamp 1676037725
transform 1 0 23644 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_251
timestamp 1676037725
transform 1 0 24196 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_253
timestamp 1676037725
transform 1 0 24380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_265
timestamp 1676037725
transform 1 0 25484 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_277
timestamp 1676037725
transform 1 0 26588 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_289
timestamp 1676037725
transform 1 0 27692 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_301
timestamp 1676037725
transform 1 0 28796 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_307
timestamp 1676037725
transform 1 0 29348 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_309
timestamp 1676037725
transform 1 0 29532 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_321
timestamp 1676037725
transform 1 0 30636 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_333
timestamp 1676037725
transform 1 0 31740 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_345
timestamp 1676037725
transform 1 0 32844 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_357
timestamp 1676037725
transform 1 0 33948 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_363
timestamp 1676037725
transform 1 0 34500 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_365
timestamp 1676037725
transform 1 0 34684 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_377
timestamp 1676037725
transform 1 0 35788 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_389
timestamp 1676037725
transform 1 0 36892 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_401
timestamp 1676037725
transform 1 0 37996 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_413
timestamp 1676037725
transform 1 0 39100 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_419
timestamp 1676037725
transform 1 0 39652 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_421
timestamp 1676037725
transform 1 0 39836 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_433
timestamp 1676037725
transform 1 0 40940 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_445
timestamp 1676037725
transform 1 0 42044 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_457
timestamp 1676037725
transform 1 0 43148 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_469
timestamp 1676037725
transform 1 0 44252 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_475
timestamp 1676037725
transform 1 0 44804 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_477
timestamp 1676037725
transform 1 0 44988 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_489
timestamp 1676037725
transform 1 0 46092 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_501
timestamp 1676037725
transform 1 0 47196 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_527
timestamp 1676037725
transform 1 0 49588 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_531
timestamp 1676037725
transform 1 0 49956 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_533
timestamp 1676037725
transform 1 0 50140 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_545
timestamp 1676037725
transform 1 0 51244 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_557
timestamp 1676037725
transform 1 0 52348 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_569
timestamp 1676037725
transform 1 0 53452 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_581
timestamp 1676037725
transform 1 0 54556 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_587
timestamp 1676037725
transform 1 0 55108 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_589
timestamp 1676037725
transform 1 0 55292 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_601
timestamp 1676037725
transform 1 0 56396 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_613
timestamp 1676037725
transform 1 0 57500 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_88_623
timestamp 1676037725
transform 1 0 58420 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_89_3
timestamp 1676037725
transform 1 0 1380 0 -1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_89_11
timestamp 1676037725
transform 1 0 2116 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_23
timestamp 1676037725
transform 1 0 3220 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_35
timestamp 1676037725
transform 1 0 4324 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_89_47
timestamp 1676037725
transform 1 0 5428 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_89_55
timestamp 1676037725
transform 1 0 6164 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_57
timestamp 1676037725
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_69
timestamp 1676037725
transform 1 0 7452 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_81
timestamp 1676037725
transform 1 0 8556 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_93
timestamp 1676037725
transform 1 0 9660 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_105
timestamp 1676037725
transform 1 0 10764 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_111
timestamp 1676037725
transform 1 0 11316 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_113
timestamp 1676037725
transform 1 0 11500 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_125
timestamp 1676037725
transform 1 0 12604 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_137
timestamp 1676037725
transform 1 0 13708 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_149
timestamp 1676037725
transform 1 0 14812 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_161
timestamp 1676037725
transform 1 0 15916 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_167
timestamp 1676037725
transform 1 0 16468 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_169
timestamp 1676037725
transform 1 0 16652 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_181
timestamp 1676037725
transform 1 0 17756 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_193
timestamp 1676037725
transform 1 0 18860 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_205
timestamp 1676037725
transform 1 0 19964 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_217
timestamp 1676037725
transform 1 0 21068 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_223
timestamp 1676037725
transform 1 0 21620 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_225
timestamp 1676037725
transform 1 0 21804 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_237
timestamp 1676037725
transform 1 0 22908 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_249
timestamp 1676037725
transform 1 0 24012 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_261
timestamp 1676037725
transform 1 0 25116 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_273
timestamp 1676037725
transform 1 0 26220 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_279
timestamp 1676037725
transform 1 0 26772 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_281
timestamp 1676037725
transform 1 0 26956 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_293
timestamp 1676037725
transform 1 0 28060 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_305
timestamp 1676037725
transform 1 0 29164 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_317
timestamp 1676037725
transform 1 0 30268 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_329
timestamp 1676037725
transform 1 0 31372 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_335
timestamp 1676037725
transform 1 0 31924 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_337
timestamp 1676037725
transform 1 0 32108 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_349
timestamp 1676037725
transform 1 0 33212 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_361
timestamp 1676037725
transform 1 0 34316 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_373
timestamp 1676037725
transform 1 0 35420 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_385
timestamp 1676037725
transform 1 0 36524 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_391
timestamp 1676037725
transform 1 0 37076 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_393
timestamp 1676037725
transform 1 0 37260 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_405
timestamp 1676037725
transform 1 0 38364 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_417
timestamp 1676037725
transform 1 0 39468 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_429
timestamp 1676037725
transform 1 0 40572 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_441
timestamp 1676037725
transform 1 0 41676 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_447
timestamp 1676037725
transform 1 0 42228 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_449
timestamp 1676037725
transform 1 0 42412 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_461
timestamp 1676037725
transform 1 0 43516 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_473
timestamp 1676037725
transform 1 0 44620 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_485
timestamp 1676037725
transform 1 0 45724 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_497
timestamp 1676037725
transform 1 0 46828 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_503
timestamp 1676037725
transform 1 0 47380 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_89_519
timestamp 1676037725
transform 1 0 48852 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_89_523
timestamp 1676037725
transform 1 0 49220 0 -1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_89_533
timestamp 1676037725
transform 1 0 50140 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_545
timestamp 1676037725
transform 1 0 51244 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_89_557
timestamp 1676037725
transform 1 0 52348 0 -1 51136
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_89_561
timestamp 1676037725
transform 1 0 52716 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_573
timestamp 1676037725
transform 1 0 53820 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_585
timestamp 1676037725
transform 1 0 54924 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_597
timestamp 1676037725
transform 1 0 56028 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_609
timestamp 1676037725
transform 1 0 57132 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_615
timestamp 1676037725
transform 1 0 57684 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_89_617
timestamp 1676037725
transform 1 0 57868 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_89_623
timestamp 1676037725
transform 1 0 58420 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_90_3
timestamp 1676037725
transform 1 0 1380 0 1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_90_11
timestamp 1676037725
transform 1 0 2116 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_90_23
timestamp 1676037725
transform 1 0 3220 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_27
timestamp 1676037725
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_29
timestamp 1676037725
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_41
timestamp 1676037725
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_53
timestamp 1676037725
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_65
timestamp 1676037725
transform 1 0 7084 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_77
timestamp 1676037725
transform 1 0 8188 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_83
timestamp 1676037725
transform 1 0 8740 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_85
timestamp 1676037725
transform 1 0 8924 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_97
timestamp 1676037725
transform 1 0 10028 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_109
timestamp 1676037725
transform 1 0 11132 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_121
timestamp 1676037725
transform 1 0 12236 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_133
timestamp 1676037725
transform 1 0 13340 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_139
timestamp 1676037725
transform 1 0 13892 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_141
timestamp 1676037725
transform 1 0 14076 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_153
timestamp 1676037725
transform 1 0 15180 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_165
timestamp 1676037725
transform 1 0 16284 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_177
timestamp 1676037725
transform 1 0 17388 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_189
timestamp 1676037725
transform 1 0 18492 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_195
timestamp 1676037725
transform 1 0 19044 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_197
timestamp 1676037725
transform 1 0 19228 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_209
timestamp 1676037725
transform 1 0 20332 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_221
timestamp 1676037725
transform 1 0 21436 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_233
timestamp 1676037725
transform 1 0 22540 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_245
timestamp 1676037725
transform 1 0 23644 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_251
timestamp 1676037725
transform 1 0 24196 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_253
timestamp 1676037725
transform 1 0 24380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_265
timestamp 1676037725
transform 1 0 25484 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_277
timestamp 1676037725
transform 1 0 26588 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_289
timestamp 1676037725
transform 1 0 27692 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_301
timestamp 1676037725
transform 1 0 28796 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_307
timestamp 1676037725
transform 1 0 29348 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_309
timestamp 1676037725
transform 1 0 29532 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_321
timestamp 1676037725
transform 1 0 30636 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_333
timestamp 1676037725
transform 1 0 31740 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_345
timestamp 1676037725
transform 1 0 32844 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_357
timestamp 1676037725
transform 1 0 33948 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_363
timestamp 1676037725
transform 1 0 34500 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_365
timestamp 1676037725
transform 1 0 34684 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_377
timestamp 1676037725
transform 1 0 35788 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_398
timestamp 1676037725
transform 1 0 37720 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_90_410
timestamp 1676037725
transform 1 0 38824 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_90_418
timestamp 1676037725
transform 1 0 39560 0 1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_90_421
timestamp 1676037725
transform 1 0 39836 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_433
timestamp 1676037725
transform 1 0 40940 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_445
timestamp 1676037725
transform 1 0 42044 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_457
timestamp 1676037725
transform 1 0 43148 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_469
timestamp 1676037725
transform 1 0 44252 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_475
timestamp 1676037725
transform 1 0 44804 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_477
timestamp 1676037725
transform 1 0 44988 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_90_489
timestamp 1676037725
transform 1 0 46092 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_90_505
timestamp 1676037725
transform 1 0 47564 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_90_526
timestamp 1676037725
transform 1 0 49496 0 1 51136
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_90_533
timestamp 1676037725
transform 1 0 50140 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_545
timestamp 1676037725
transform 1 0 51244 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_557
timestamp 1676037725
transform 1 0 52348 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_569
timestamp 1676037725
transform 1 0 53452 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_581
timestamp 1676037725
transform 1 0 54556 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_587
timestamp 1676037725
transform 1 0 55108 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_589
timestamp 1676037725
transform 1 0 55292 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_90_601
timestamp 1676037725
transform 1 0 56396 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_90_609
timestamp 1676037725
transform 1 0 57132 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_90_615
timestamp 1676037725
transform 1 0 57684 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_90_623
timestamp 1676037725
transform 1 0 58420 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_91_3
timestamp 1676037725
transform 1 0 1380 0 -1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_91_9
timestamp 1676037725
transform 1 0 1932 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_21
timestamp 1676037725
transform 1 0 3036 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_33
timestamp 1676037725
transform 1 0 4140 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_45
timestamp 1676037725
transform 1 0 5244 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_91_53
timestamp 1676037725
transform 1 0 5980 0 -1 52224
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_91_57
timestamp 1676037725
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_69
timestamp 1676037725
transform 1 0 7452 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_81
timestamp 1676037725
transform 1 0 8556 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_93
timestamp 1676037725
transform 1 0 9660 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_105
timestamp 1676037725
transform 1 0 10764 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_111
timestamp 1676037725
transform 1 0 11316 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_113
timestamp 1676037725
transform 1 0 11500 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_125
timestamp 1676037725
transform 1 0 12604 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_137
timestamp 1676037725
transform 1 0 13708 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_149
timestamp 1676037725
transform 1 0 14812 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_161
timestamp 1676037725
transform 1 0 15916 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_167
timestamp 1676037725
transform 1 0 16468 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_169
timestamp 1676037725
transform 1 0 16652 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_181
timestamp 1676037725
transform 1 0 17756 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_193
timestamp 1676037725
transform 1 0 18860 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_205
timestamp 1676037725
transform 1 0 19964 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_217
timestamp 1676037725
transform 1 0 21068 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_223
timestamp 1676037725
transform 1 0 21620 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_225
timestamp 1676037725
transform 1 0 21804 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_237
timestamp 1676037725
transform 1 0 22908 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_249
timestamp 1676037725
transform 1 0 24012 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_261
timestamp 1676037725
transform 1 0 25116 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_273
timestamp 1676037725
transform 1 0 26220 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_279
timestamp 1676037725
transform 1 0 26772 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_281
timestamp 1676037725
transform 1 0 26956 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_293
timestamp 1676037725
transform 1 0 28060 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_305
timestamp 1676037725
transform 1 0 29164 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_317
timestamp 1676037725
transform 1 0 30268 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_329
timestamp 1676037725
transform 1 0 31372 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_335
timestamp 1676037725
transform 1 0 31924 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_337
timestamp 1676037725
transform 1 0 32108 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_349
timestamp 1676037725
transform 1 0 33212 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_361
timestamp 1676037725
transform 1 0 34316 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_373
timestamp 1676037725
transform 1 0 35420 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_385
timestamp 1676037725
transform 1 0 36524 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_391
timestamp 1676037725
transform 1 0 37076 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_393
timestamp 1676037725
transform 1 0 37260 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_405
timestamp 1676037725
transform 1 0 38364 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_417
timestamp 1676037725
transform 1 0 39468 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_429
timestamp 1676037725
transform 1 0 40572 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_441
timestamp 1676037725
transform 1 0 41676 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_447
timestamp 1676037725
transform 1 0 42228 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_449
timestamp 1676037725
transform 1 0 42412 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_461
timestamp 1676037725
transform 1 0 43516 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_473
timestamp 1676037725
transform 1 0 44620 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_485
timestamp 1676037725
transform 1 0 45724 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_497
timestamp 1676037725
transform 1 0 46828 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_503
timestamp 1676037725
transform 1 0 47380 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_91_505
timestamp 1676037725
transform 1 0 47564 0 -1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_91_521
timestamp 1676037725
transform 1 0 49036 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_533
timestamp 1676037725
transform 1 0 50140 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_545
timestamp 1676037725
transform 1 0 51244 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_91_557
timestamp 1676037725
transform 1 0 52348 0 -1 52224
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_91_561
timestamp 1676037725
transform 1 0 52716 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_573
timestamp 1676037725
transform 1 0 53820 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_585
timestamp 1676037725
transform 1 0 54924 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_597
timestamp 1676037725
transform 1 0 56028 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_91_609
timestamp 1676037725
transform 1 0 57132 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_91_614
timestamp 1676037725
transform 1 0 57592 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_91_617
timestamp 1676037725
transform 1 0 57868 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_91_623
timestamp 1676037725
transform 1 0 58420 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_92_3
timestamp 1676037725
transform 1 0 1380 0 1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_92_11
timestamp 1676037725
transform 1 0 2116 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_23
timestamp 1676037725
transform 1 0 3220 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_27
timestamp 1676037725
transform 1 0 3588 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_29
timestamp 1676037725
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_41
timestamp 1676037725
transform 1 0 4876 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_53
timestamp 1676037725
transform 1 0 5980 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_65
timestamp 1676037725
transform 1 0 7084 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_77
timestamp 1676037725
transform 1 0 8188 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_83
timestamp 1676037725
transform 1 0 8740 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_85
timestamp 1676037725
transform 1 0 8924 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_97
timestamp 1676037725
transform 1 0 10028 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_109
timestamp 1676037725
transform 1 0 11132 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_121
timestamp 1676037725
transform 1 0 12236 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_133
timestamp 1676037725
transform 1 0 13340 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_139
timestamp 1676037725
transform 1 0 13892 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_141
timestamp 1676037725
transform 1 0 14076 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_153
timestamp 1676037725
transform 1 0 15180 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_165
timestamp 1676037725
transform 1 0 16284 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_177
timestamp 1676037725
transform 1 0 17388 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_189
timestamp 1676037725
transform 1 0 18492 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_195
timestamp 1676037725
transform 1 0 19044 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_197
timestamp 1676037725
transform 1 0 19228 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_209
timestamp 1676037725
transform 1 0 20332 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_221
timestamp 1676037725
transform 1 0 21436 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_233
timestamp 1676037725
transform 1 0 22540 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_245
timestamp 1676037725
transform 1 0 23644 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_251
timestamp 1676037725
transform 1 0 24196 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_253
timestamp 1676037725
transform 1 0 24380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_265
timestamp 1676037725
transform 1 0 25484 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_277
timestamp 1676037725
transform 1 0 26588 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_289
timestamp 1676037725
transform 1 0 27692 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_301
timestamp 1676037725
transform 1 0 28796 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_307
timestamp 1676037725
transform 1 0 29348 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_309
timestamp 1676037725
transform 1 0 29532 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_321
timestamp 1676037725
transform 1 0 30636 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_333
timestamp 1676037725
transform 1 0 31740 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_345
timestamp 1676037725
transform 1 0 32844 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_357
timestamp 1676037725
transform 1 0 33948 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_363
timestamp 1676037725
transform 1 0 34500 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_365
timestamp 1676037725
transform 1 0 34684 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_377
timestamp 1676037725
transform 1 0 35788 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_389
timestamp 1676037725
transform 1 0 36892 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_401
timestamp 1676037725
transform 1 0 37996 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_413
timestamp 1676037725
transform 1 0 39100 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_419
timestamp 1676037725
transform 1 0 39652 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_421
timestamp 1676037725
transform 1 0 39836 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_433
timestamp 1676037725
transform 1 0 40940 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_92_441
timestamp 1676037725
transform 1 0 41676 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_92_444
timestamp 1676037725
transform 1 0 41952 0 1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_92_453
timestamp 1676037725
transform 1 0 42780 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_465
timestamp 1676037725
transform 1 0 43884 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_92_473
timestamp 1676037725
transform 1 0 44620 0 1 52224
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_92_477
timestamp 1676037725
transform 1 0 44988 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_489
timestamp 1676037725
transform 1 0 46092 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_92_501
timestamp 1676037725
transform 1 0 47196 0 1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_92_517
timestamp 1676037725
transform 1 0 48668 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_92_529
timestamp 1676037725
transform 1 0 49772 0 1 52224
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_92_533
timestamp 1676037725
transform 1 0 50140 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_545
timestamp 1676037725
transform 1 0 51244 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_557
timestamp 1676037725
transform 1 0 52348 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_569
timestamp 1676037725
transform 1 0 53452 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_581
timestamp 1676037725
transform 1 0 54556 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_587
timestamp 1676037725
transform 1 0 55108 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_589
timestamp 1676037725
transform 1 0 55292 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_601
timestamp 1676037725
transform 1 0 56396 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_613
timestamp 1676037725
transform 1 0 57500 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_92_623
timestamp 1676037725
transform 1 0 58420 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_93_3
timestamp 1676037725
transform 1 0 1380 0 -1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_93_11
timestamp 1676037725
transform 1 0 2116 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_23
timestamp 1676037725
transform 1 0 3220 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_35
timestamp 1676037725
transform 1 0 4324 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_47
timestamp 1676037725
transform 1 0 5428 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_93_55
timestamp 1676037725
transform 1 0 6164 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_57
timestamp 1676037725
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_69
timestamp 1676037725
transform 1 0 7452 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_81
timestamp 1676037725
transform 1 0 8556 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_93
timestamp 1676037725
transform 1 0 9660 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_105
timestamp 1676037725
transform 1 0 10764 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_111
timestamp 1676037725
transform 1 0 11316 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_113
timestamp 1676037725
transform 1 0 11500 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_125
timestamp 1676037725
transform 1 0 12604 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_137
timestamp 1676037725
transform 1 0 13708 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_149
timestamp 1676037725
transform 1 0 14812 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_161
timestamp 1676037725
transform 1 0 15916 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_167
timestamp 1676037725
transform 1 0 16468 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_169
timestamp 1676037725
transform 1 0 16652 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_181
timestamp 1676037725
transform 1 0 17756 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_193
timestamp 1676037725
transform 1 0 18860 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_205
timestamp 1676037725
transform 1 0 19964 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_217
timestamp 1676037725
transform 1 0 21068 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_223
timestamp 1676037725
transform 1 0 21620 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_225
timestamp 1676037725
transform 1 0 21804 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_237
timestamp 1676037725
transform 1 0 22908 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_249
timestamp 1676037725
transform 1 0 24012 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_261
timestamp 1676037725
transform 1 0 25116 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_273
timestamp 1676037725
transform 1 0 26220 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_279
timestamp 1676037725
transform 1 0 26772 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_281
timestamp 1676037725
transform 1 0 26956 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_293
timestamp 1676037725
transform 1 0 28060 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_305
timestamp 1676037725
transform 1 0 29164 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_317
timestamp 1676037725
transform 1 0 30268 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_329
timestamp 1676037725
transform 1 0 31372 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_335
timestamp 1676037725
transform 1 0 31924 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_337
timestamp 1676037725
transform 1 0 32108 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_349
timestamp 1676037725
transform 1 0 33212 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_361
timestamp 1676037725
transform 1 0 34316 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_373
timestamp 1676037725
transform 1 0 35420 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_385
timestamp 1676037725
transform 1 0 36524 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_391
timestamp 1676037725
transform 1 0 37076 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_393
timestamp 1676037725
transform 1 0 37260 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_405
timestamp 1676037725
transform 1 0 38364 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_417
timestamp 1676037725
transform 1 0 39468 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_429
timestamp 1676037725
transform 1 0 40572 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_441
timestamp 1676037725
transform 1 0 41676 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_447
timestamp 1676037725
transform 1 0 42228 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_449
timestamp 1676037725
transform 1 0 42412 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_461
timestamp 1676037725
transform 1 0 43516 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_473
timestamp 1676037725
transform 1 0 44620 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_485
timestamp 1676037725
transform 1 0 45724 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_497
timestamp 1676037725
transform 1 0 46828 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_503
timestamp 1676037725
transform 1 0 47380 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_93_505
timestamp 1676037725
transform 1 0 47564 0 -1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_93_521
timestamp 1676037725
transform 1 0 49036 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_533
timestamp 1676037725
transform 1 0 50140 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_545
timestamp 1676037725
transform 1 0 51244 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_93_557
timestamp 1676037725
transform 1 0 52348 0 -1 53312
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_93_561
timestamp 1676037725
transform 1 0 52716 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_573
timestamp 1676037725
transform 1 0 53820 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_585
timestamp 1676037725
transform 1 0 54924 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_597
timestamp 1676037725
transform 1 0 56028 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_609
timestamp 1676037725
transform 1 0 57132 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_615
timestamp 1676037725
transform 1 0 57684 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_93_617
timestamp 1676037725
transform 1 0 57868 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_93_623
timestamp 1676037725
transform 1 0 58420 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_3
timestamp 1676037725
transform 1 0 1380 0 1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_94_11
timestamp 1676037725
transform 1 0 2116 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_23
timestamp 1676037725
transform 1 0 3220 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_27
timestamp 1676037725
transform 1 0 3588 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_29
timestamp 1676037725
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_41
timestamp 1676037725
transform 1 0 4876 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_53
timestamp 1676037725
transform 1 0 5980 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_65
timestamp 1676037725
transform 1 0 7084 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_77
timestamp 1676037725
transform 1 0 8188 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_83
timestamp 1676037725
transform 1 0 8740 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_85
timestamp 1676037725
transform 1 0 8924 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_97
timestamp 1676037725
transform 1 0 10028 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_109
timestamp 1676037725
transform 1 0 11132 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_121
timestamp 1676037725
transform 1 0 12236 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_133
timestamp 1676037725
transform 1 0 13340 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_139
timestamp 1676037725
transform 1 0 13892 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_141
timestamp 1676037725
transform 1 0 14076 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_153
timestamp 1676037725
transform 1 0 15180 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_165
timestamp 1676037725
transform 1 0 16284 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_177
timestamp 1676037725
transform 1 0 17388 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_189
timestamp 1676037725
transform 1 0 18492 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_195
timestamp 1676037725
transform 1 0 19044 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_197
timestamp 1676037725
transform 1 0 19228 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_209
timestamp 1676037725
transform 1 0 20332 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_221
timestamp 1676037725
transform 1 0 21436 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_233
timestamp 1676037725
transform 1 0 22540 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_245
timestamp 1676037725
transform 1 0 23644 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_251
timestamp 1676037725
transform 1 0 24196 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_253
timestamp 1676037725
transform 1 0 24380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_265
timestamp 1676037725
transform 1 0 25484 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_277
timestamp 1676037725
transform 1 0 26588 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_289
timestamp 1676037725
transform 1 0 27692 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_301
timestamp 1676037725
transform 1 0 28796 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_307
timestamp 1676037725
transform 1 0 29348 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_309
timestamp 1676037725
transform 1 0 29532 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_321
timestamp 1676037725
transform 1 0 30636 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_333
timestamp 1676037725
transform 1 0 31740 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_345
timestamp 1676037725
transform 1 0 32844 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_357
timestamp 1676037725
transform 1 0 33948 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_363
timestamp 1676037725
transform 1 0 34500 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_365
timestamp 1676037725
transform 1 0 34684 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_377
timestamp 1676037725
transform 1 0 35788 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_389
timestamp 1676037725
transform 1 0 36892 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_401
timestamp 1676037725
transform 1 0 37996 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_413
timestamp 1676037725
transform 1 0 39100 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_419
timestamp 1676037725
transform 1 0 39652 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_421
timestamp 1676037725
transform 1 0 39836 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_433
timestamp 1676037725
transform 1 0 40940 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_445
timestamp 1676037725
transform 1 0 42044 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_457
timestamp 1676037725
transform 1 0 43148 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_469
timestamp 1676037725
transform 1 0 44252 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_475
timestamp 1676037725
transform 1 0 44804 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_477
timestamp 1676037725
transform 1 0 44988 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_489
timestamp 1676037725
transform 1 0 46092 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_501
timestamp 1676037725
transform 1 0 47196 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_513
timestamp 1676037725
transform 1 0 48300 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_525
timestamp 1676037725
transform 1 0 49404 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_531
timestamp 1676037725
transform 1 0 49956 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_533
timestamp 1676037725
transform 1 0 50140 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_545
timestamp 1676037725
transform 1 0 51244 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_557
timestamp 1676037725
transform 1 0 52348 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_569
timestamp 1676037725
transform 1 0 53452 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_581
timestamp 1676037725
transform 1 0 54556 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_587
timestamp 1676037725
transform 1 0 55108 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_589
timestamp 1676037725
transform 1 0 55292 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_601
timestamp 1676037725
transform 1 0 56396 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_613
timestamp 1676037725
transform 1 0 57500 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_94_623
timestamp 1676037725
transform 1 0 58420 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_3
timestamp 1676037725
transform 1 0 1380 0 -1 54400
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_95_11
timestamp 1676037725
transform 1 0 2116 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_23
timestamp 1676037725
transform 1 0 3220 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_35
timestamp 1676037725
transform 1 0 4324 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_95_47
timestamp 1676037725
transform 1 0 5428 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_55
timestamp 1676037725
transform 1 0 6164 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_57
timestamp 1676037725
transform 1 0 6348 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_69
timestamp 1676037725
transform 1 0 7452 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_81
timestamp 1676037725
transform 1 0 8556 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_93
timestamp 1676037725
transform 1 0 9660 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_105
timestamp 1676037725
transform 1 0 10764 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_111
timestamp 1676037725
transform 1 0 11316 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_113
timestamp 1676037725
transform 1 0 11500 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_125
timestamp 1676037725
transform 1 0 12604 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_137
timestamp 1676037725
transform 1 0 13708 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_149
timestamp 1676037725
transform 1 0 14812 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_161
timestamp 1676037725
transform 1 0 15916 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_167
timestamp 1676037725
transform 1 0 16468 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_169
timestamp 1676037725
transform 1 0 16652 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_181
timestamp 1676037725
transform 1 0 17756 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_193
timestamp 1676037725
transform 1 0 18860 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_205
timestamp 1676037725
transform 1 0 19964 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_217
timestamp 1676037725
transform 1 0 21068 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_223
timestamp 1676037725
transform 1 0 21620 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_225
timestamp 1676037725
transform 1 0 21804 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_237
timestamp 1676037725
transform 1 0 22908 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_249
timestamp 1676037725
transform 1 0 24012 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_261
timestamp 1676037725
transform 1 0 25116 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_273
timestamp 1676037725
transform 1 0 26220 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_279
timestamp 1676037725
transform 1 0 26772 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_281
timestamp 1676037725
transform 1 0 26956 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_293
timestamp 1676037725
transform 1 0 28060 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_305
timestamp 1676037725
transform 1 0 29164 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_317
timestamp 1676037725
transform 1 0 30268 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_329
timestamp 1676037725
transform 1 0 31372 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_335
timestamp 1676037725
transform 1 0 31924 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_337
timestamp 1676037725
transform 1 0 32108 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_349
timestamp 1676037725
transform 1 0 33212 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_361
timestamp 1676037725
transform 1 0 34316 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_373
timestamp 1676037725
transform 1 0 35420 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_385
timestamp 1676037725
transform 1 0 36524 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_391
timestamp 1676037725
transform 1 0 37076 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_393
timestamp 1676037725
transform 1 0 37260 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_405
timestamp 1676037725
transform 1 0 38364 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_417
timestamp 1676037725
transform 1 0 39468 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_429
timestamp 1676037725
transform 1 0 40572 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_441
timestamp 1676037725
transform 1 0 41676 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_447
timestamp 1676037725
transform 1 0 42228 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_449
timestamp 1676037725
transform 1 0 42412 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_461
timestamp 1676037725
transform 1 0 43516 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_473
timestamp 1676037725
transform 1 0 44620 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_485
timestamp 1676037725
transform 1 0 45724 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_497
timestamp 1676037725
transform 1 0 46828 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_503
timestamp 1676037725
transform 1 0 47380 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_505
timestamp 1676037725
transform 1 0 47564 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_517
timestamp 1676037725
transform 1 0 48668 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_529
timestamp 1676037725
transform 1 0 49772 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_541
timestamp 1676037725
transform 1 0 50876 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_553
timestamp 1676037725
transform 1 0 51980 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_559
timestamp 1676037725
transform 1 0 52532 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_561
timestamp 1676037725
transform 1 0 52716 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_573
timestamp 1676037725
transform 1 0 53820 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_585
timestamp 1676037725
transform 1 0 54924 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_597
timestamp 1676037725
transform 1 0 56028 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_609
timestamp 1676037725
transform 1 0 57132 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_615
timestamp 1676037725
transform 1 0 57684 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_617
timestamp 1676037725
transform 1 0 57868 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_623
timestamp 1676037725
transform 1 0 58420 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_96_3
timestamp 1676037725
transform 1 0 1380 0 1 54400
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_96_11
timestamp 1676037725
transform 1 0 2116 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_96_23
timestamp 1676037725
transform 1 0 3220 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_96_27
timestamp 1676037725
transform 1 0 3588 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_29
timestamp 1676037725
transform 1 0 3772 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_41
timestamp 1676037725
transform 1 0 4876 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_53
timestamp 1676037725
transform 1 0 5980 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_65
timestamp 1676037725
transform 1 0 7084 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_77
timestamp 1676037725
transform 1 0 8188 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_83
timestamp 1676037725
transform 1 0 8740 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_85
timestamp 1676037725
transform 1 0 8924 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_97
timestamp 1676037725
transform 1 0 10028 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_109
timestamp 1676037725
transform 1 0 11132 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_121
timestamp 1676037725
transform 1 0 12236 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_133
timestamp 1676037725
transform 1 0 13340 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_139
timestamp 1676037725
transform 1 0 13892 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_141
timestamp 1676037725
transform 1 0 14076 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_153
timestamp 1676037725
transform 1 0 15180 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_165
timestamp 1676037725
transform 1 0 16284 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_177
timestamp 1676037725
transform 1 0 17388 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_189
timestamp 1676037725
transform 1 0 18492 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_195
timestamp 1676037725
transform 1 0 19044 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_197
timestamp 1676037725
transform 1 0 19228 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_209
timestamp 1676037725
transform 1 0 20332 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_221
timestamp 1676037725
transform 1 0 21436 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_233
timestamp 1676037725
transform 1 0 22540 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_245
timestamp 1676037725
transform 1 0 23644 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_251
timestamp 1676037725
transform 1 0 24196 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_253
timestamp 1676037725
transform 1 0 24380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_265
timestamp 1676037725
transform 1 0 25484 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_277
timestamp 1676037725
transform 1 0 26588 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_289
timestamp 1676037725
transform 1 0 27692 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_301
timestamp 1676037725
transform 1 0 28796 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_307
timestamp 1676037725
transform 1 0 29348 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_309
timestamp 1676037725
transform 1 0 29532 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_321
timestamp 1676037725
transform 1 0 30636 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_333
timestamp 1676037725
transform 1 0 31740 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_345
timestamp 1676037725
transform 1 0 32844 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_357
timestamp 1676037725
transform 1 0 33948 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_363
timestamp 1676037725
transform 1 0 34500 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_365
timestamp 1676037725
transform 1 0 34684 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_377
timestamp 1676037725
transform 1 0 35788 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_389
timestamp 1676037725
transform 1 0 36892 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_401
timestamp 1676037725
transform 1 0 37996 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_413
timestamp 1676037725
transform 1 0 39100 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_419
timestamp 1676037725
transform 1 0 39652 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_421
timestamp 1676037725
transform 1 0 39836 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_433
timestamp 1676037725
transform 1 0 40940 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_445
timestamp 1676037725
transform 1 0 42044 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_457
timestamp 1676037725
transform 1 0 43148 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_469
timestamp 1676037725
transform 1 0 44252 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_475
timestamp 1676037725
transform 1 0 44804 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_477
timestamp 1676037725
transform 1 0 44988 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_489
timestamp 1676037725
transform 1 0 46092 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_501
timestamp 1676037725
transform 1 0 47196 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_513
timestamp 1676037725
transform 1 0 48300 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_525
timestamp 1676037725
transform 1 0 49404 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_531
timestamp 1676037725
transform 1 0 49956 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_533
timestamp 1676037725
transform 1 0 50140 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_545
timestamp 1676037725
transform 1 0 51244 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_557
timestamp 1676037725
transform 1 0 52348 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_569
timestamp 1676037725
transform 1 0 53452 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_581
timestamp 1676037725
transform 1 0 54556 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_587
timestamp 1676037725
transform 1 0 55108 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_589
timestamp 1676037725
transform 1 0 55292 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_96_601
timestamp 1676037725
transform 1 0 56396 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_96_609
timestamp 1676037725
transform 1 0 57132 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_96_615
timestamp 1676037725
transform 1 0 57684 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_96_623
timestamp 1676037725
transform 1 0 58420 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_97_3
timestamp 1676037725
transform 1 0 1380 0 -1 55488
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_97_11
timestamp 1676037725
transform 1 0 2116 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_23
timestamp 1676037725
transform 1 0 3220 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_35
timestamp 1676037725
transform 1 0 4324 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_97_47
timestamp 1676037725
transform 1 0 5428 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_97_55
timestamp 1676037725
transform 1 0 6164 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_57
timestamp 1676037725
transform 1 0 6348 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_69
timestamp 1676037725
transform 1 0 7452 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_81
timestamp 1676037725
transform 1 0 8556 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_93
timestamp 1676037725
transform 1 0 9660 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_105
timestamp 1676037725
transform 1 0 10764 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_111
timestamp 1676037725
transform 1 0 11316 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_113
timestamp 1676037725
transform 1 0 11500 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_125
timestamp 1676037725
transform 1 0 12604 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_137
timestamp 1676037725
transform 1 0 13708 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_149
timestamp 1676037725
transform 1 0 14812 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_161
timestamp 1676037725
transform 1 0 15916 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_167
timestamp 1676037725
transform 1 0 16468 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_169
timestamp 1676037725
transform 1 0 16652 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_181
timestamp 1676037725
transform 1 0 17756 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_193
timestamp 1676037725
transform 1 0 18860 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_205
timestamp 1676037725
transform 1 0 19964 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_217
timestamp 1676037725
transform 1 0 21068 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_223
timestamp 1676037725
transform 1 0 21620 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_225
timestamp 1676037725
transform 1 0 21804 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_237
timestamp 1676037725
transform 1 0 22908 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_249
timestamp 1676037725
transform 1 0 24012 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_261
timestamp 1676037725
transform 1 0 25116 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_273
timestamp 1676037725
transform 1 0 26220 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_279
timestamp 1676037725
transform 1 0 26772 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_281
timestamp 1676037725
transform 1 0 26956 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_293
timestamp 1676037725
transform 1 0 28060 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_305
timestamp 1676037725
transform 1 0 29164 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_317
timestamp 1676037725
transform 1 0 30268 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_329
timestamp 1676037725
transform 1 0 31372 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_335
timestamp 1676037725
transform 1 0 31924 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_337
timestamp 1676037725
transform 1 0 32108 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_349
timestamp 1676037725
transform 1 0 33212 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_361
timestamp 1676037725
transform 1 0 34316 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_373
timestamp 1676037725
transform 1 0 35420 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_385
timestamp 1676037725
transform 1 0 36524 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_391
timestamp 1676037725
transform 1 0 37076 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_393
timestamp 1676037725
transform 1 0 37260 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_405
timestamp 1676037725
transform 1 0 38364 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_417
timestamp 1676037725
transform 1 0 39468 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_429
timestamp 1676037725
transform 1 0 40572 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_441
timestamp 1676037725
transform 1 0 41676 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_447
timestamp 1676037725
transform 1 0 42228 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_449
timestamp 1676037725
transform 1 0 42412 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_461
timestamp 1676037725
transform 1 0 43516 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_473
timestamp 1676037725
transform 1 0 44620 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_485
timestamp 1676037725
transform 1 0 45724 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_497
timestamp 1676037725
transform 1 0 46828 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_503
timestamp 1676037725
transform 1 0 47380 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_505
timestamp 1676037725
transform 1 0 47564 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_517
timestamp 1676037725
transform 1 0 48668 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_529
timestamp 1676037725
transform 1 0 49772 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_541
timestamp 1676037725
transform 1 0 50876 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_553
timestamp 1676037725
transform 1 0 51980 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_559
timestamp 1676037725
transform 1 0 52532 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_561
timestamp 1676037725
transform 1 0 52716 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_573
timestamp 1676037725
transform 1 0 53820 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_585
timestamp 1676037725
transform 1 0 54924 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_597
timestamp 1676037725
transform 1 0 56028 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_609
timestamp 1676037725
transform 1 0 57132 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_615
timestamp 1676037725
transform 1 0 57684 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_97_617
timestamp 1676037725
transform 1 0 57868 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_97_623
timestamp 1676037725
transform 1 0 58420 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_98_3
timestamp 1676037725
transform 1 0 1380 0 1 55488
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_98_11
timestamp 1676037725
transform 1 0 2116 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_98_23
timestamp 1676037725
transform 1 0 3220 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_98_27
timestamp 1676037725
transform 1 0 3588 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_29
timestamp 1676037725
transform 1 0 3772 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_41
timestamp 1676037725
transform 1 0 4876 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_53
timestamp 1676037725
transform 1 0 5980 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_65
timestamp 1676037725
transform 1 0 7084 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_77
timestamp 1676037725
transform 1 0 8188 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_83
timestamp 1676037725
transform 1 0 8740 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_85
timestamp 1676037725
transform 1 0 8924 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_97
timestamp 1676037725
transform 1 0 10028 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_109
timestamp 1676037725
transform 1 0 11132 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_121
timestamp 1676037725
transform 1 0 12236 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_133
timestamp 1676037725
transform 1 0 13340 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_139
timestamp 1676037725
transform 1 0 13892 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_141
timestamp 1676037725
transform 1 0 14076 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_153
timestamp 1676037725
transform 1 0 15180 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_165
timestamp 1676037725
transform 1 0 16284 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_177
timestamp 1676037725
transform 1 0 17388 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_189
timestamp 1676037725
transform 1 0 18492 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_195
timestamp 1676037725
transform 1 0 19044 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_197
timestamp 1676037725
transform 1 0 19228 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_209
timestamp 1676037725
transform 1 0 20332 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_221
timestamp 1676037725
transform 1 0 21436 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_233
timestamp 1676037725
transform 1 0 22540 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_245
timestamp 1676037725
transform 1 0 23644 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_251
timestamp 1676037725
transform 1 0 24196 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_253
timestamp 1676037725
transform 1 0 24380 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_265
timestamp 1676037725
transform 1 0 25484 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_277
timestamp 1676037725
transform 1 0 26588 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_289
timestamp 1676037725
transform 1 0 27692 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_301
timestamp 1676037725
transform 1 0 28796 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_307
timestamp 1676037725
transform 1 0 29348 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_309
timestamp 1676037725
transform 1 0 29532 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_321
timestamp 1676037725
transform 1 0 30636 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_333
timestamp 1676037725
transform 1 0 31740 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_345
timestamp 1676037725
transform 1 0 32844 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_357
timestamp 1676037725
transform 1 0 33948 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_363
timestamp 1676037725
transform 1 0 34500 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_365
timestamp 1676037725
transform 1 0 34684 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_377
timestamp 1676037725
transform 1 0 35788 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_389
timestamp 1676037725
transform 1 0 36892 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_401
timestamp 1676037725
transform 1 0 37996 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_413
timestamp 1676037725
transform 1 0 39100 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_419
timestamp 1676037725
transform 1 0 39652 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_421
timestamp 1676037725
transform 1 0 39836 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_433
timestamp 1676037725
transform 1 0 40940 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_445
timestamp 1676037725
transform 1 0 42044 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_457
timestamp 1676037725
transform 1 0 43148 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_469
timestamp 1676037725
transform 1 0 44252 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_475
timestamp 1676037725
transform 1 0 44804 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_477
timestamp 1676037725
transform 1 0 44988 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_489
timestamp 1676037725
transform 1 0 46092 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_501
timestamp 1676037725
transform 1 0 47196 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_513
timestamp 1676037725
transform 1 0 48300 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_525
timestamp 1676037725
transform 1 0 49404 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_531
timestamp 1676037725
transform 1 0 49956 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_533
timestamp 1676037725
transform 1 0 50140 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_545
timestamp 1676037725
transform 1 0 51244 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_557
timestamp 1676037725
transform 1 0 52348 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_569
timestamp 1676037725
transform 1 0 53452 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_581
timestamp 1676037725
transform 1 0 54556 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_587
timestamp 1676037725
transform 1 0 55108 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_589
timestamp 1676037725
transform 1 0 55292 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_98_601
timestamp 1676037725
transform 1 0 56396 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_98_609
timestamp 1676037725
transform 1 0 57132 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_98_615
timestamp 1676037725
transform 1 0 57684 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_98_623
timestamp 1676037725
transform 1 0 58420 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_99_3
timestamp 1676037725
transform 1 0 1380 0 -1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_99_11
timestamp 1676037725
transform 1 0 2116 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_23
timestamp 1676037725
transform 1 0 3220 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_35
timestamp 1676037725
transform 1 0 4324 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_99_47
timestamp 1676037725
transform 1 0 5428 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_99_55
timestamp 1676037725
transform 1 0 6164 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_57
timestamp 1676037725
transform 1 0 6348 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_69
timestamp 1676037725
transform 1 0 7452 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_81
timestamp 1676037725
transform 1 0 8556 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_93
timestamp 1676037725
transform 1 0 9660 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_105
timestamp 1676037725
transform 1 0 10764 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_111
timestamp 1676037725
transform 1 0 11316 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_113
timestamp 1676037725
transform 1 0 11500 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_125
timestamp 1676037725
transform 1 0 12604 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_137
timestamp 1676037725
transform 1 0 13708 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_149
timestamp 1676037725
transform 1 0 14812 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_161
timestamp 1676037725
transform 1 0 15916 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_167
timestamp 1676037725
transform 1 0 16468 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_169
timestamp 1676037725
transform 1 0 16652 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_181
timestamp 1676037725
transform 1 0 17756 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_193
timestamp 1676037725
transform 1 0 18860 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_205
timestamp 1676037725
transform 1 0 19964 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_217
timestamp 1676037725
transform 1 0 21068 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_223
timestamp 1676037725
transform 1 0 21620 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_225
timestamp 1676037725
transform 1 0 21804 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_237
timestamp 1676037725
transform 1 0 22908 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_249
timestamp 1676037725
transform 1 0 24012 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_261
timestamp 1676037725
transform 1 0 25116 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_273
timestamp 1676037725
transform 1 0 26220 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_279
timestamp 1676037725
transform 1 0 26772 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_281
timestamp 1676037725
transform 1 0 26956 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_293
timestamp 1676037725
transform 1 0 28060 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_305
timestamp 1676037725
transform 1 0 29164 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_317
timestamp 1676037725
transform 1 0 30268 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_329
timestamp 1676037725
transform 1 0 31372 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_335
timestamp 1676037725
transform 1 0 31924 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_337
timestamp 1676037725
transform 1 0 32108 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_349
timestamp 1676037725
transform 1 0 33212 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_361
timestamp 1676037725
transform 1 0 34316 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_373
timestamp 1676037725
transform 1 0 35420 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_385
timestamp 1676037725
transform 1 0 36524 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_391
timestamp 1676037725
transform 1 0 37076 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_393
timestamp 1676037725
transform 1 0 37260 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_405
timestamp 1676037725
transform 1 0 38364 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_417
timestamp 1676037725
transform 1 0 39468 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_429
timestamp 1676037725
transform 1 0 40572 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_441
timestamp 1676037725
transform 1 0 41676 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_447
timestamp 1676037725
transform 1 0 42228 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_449
timestamp 1676037725
transform 1 0 42412 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_461
timestamp 1676037725
transform 1 0 43516 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_473
timestamp 1676037725
transform 1 0 44620 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_485
timestamp 1676037725
transform 1 0 45724 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_497
timestamp 1676037725
transform 1 0 46828 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_503
timestamp 1676037725
transform 1 0 47380 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_505
timestamp 1676037725
transform 1 0 47564 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_517
timestamp 1676037725
transform 1 0 48668 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_529
timestamp 1676037725
transform 1 0 49772 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_541
timestamp 1676037725
transform 1 0 50876 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_553
timestamp 1676037725
transform 1 0 51980 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_559
timestamp 1676037725
transform 1 0 52532 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_561
timestamp 1676037725
transform 1 0 52716 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_573
timestamp 1676037725
transform 1 0 53820 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_99_585
timestamp 1676037725
transform 1 0 54924 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_99_593
timestamp 1676037725
transform 1 0 55660 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_598
timestamp 1676037725
transform 1 0 56120 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_606
timestamp 1676037725
transform 1 0 56856 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_99_614
timestamp 1676037725
transform 1 0 57592 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_99_617
timestamp 1676037725
transform 1 0 57868 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_99_623
timestamp 1676037725
transform 1 0 58420 0 -1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_100_3
timestamp 1676037725
transform 1 0 1380 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_15
timestamp 1676037725
transform 1 0 2484 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_100_27
timestamp 1676037725
transform 1 0 3588 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_29
timestamp 1676037725
transform 1 0 3772 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_41
timestamp 1676037725
transform 1 0 4876 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_53
timestamp 1676037725
transform 1 0 5980 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_65
timestamp 1676037725
transform 1 0 7084 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_77
timestamp 1676037725
transform 1 0 8188 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_83
timestamp 1676037725
transform 1 0 8740 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_85
timestamp 1676037725
transform 1 0 8924 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_97
timestamp 1676037725
transform 1 0 10028 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_109
timestamp 1676037725
transform 1 0 11132 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_121
timestamp 1676037725
transform 1 0 12236 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_133
timestamp 1676037725
transform 1 0 13340 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_139
timestamp 1676037725
transform 1 0 13892 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_141
timestamp 1676037725
transform 1 0 14076 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_153
timestamp 1676037725
transform 1 0 15180 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_165
timestamp 1676037725
transform 1 0 16284 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_177
timestamp 1676037725
transform 1 0 17388 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_189
timestamp 1676037725
transform 1 0 18492 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_195
timestamp 1676037725
transform 1 0 19044 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_197
timestamp 1676037725
transform 1 0 19228 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_209
timestamp 1676037725
transform 1 0 20332 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_221
timestamp 1676037725
transform 1 0 21436 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_233
timestamp 1676037725
transform 1 0 22540 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_245
timestamp 1676037725
transform 1 0 23644 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_251
timestamp 1676037725
transform 1 0 24196 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_253
timestamp 1676037725
transform 1 0 24380 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_265
timestamp 1676037725
transform 1 0 25484 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_277
timestamp 1676037725
transform 1 0 26588 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_289
timestamp 1676037725
transform 1 0 27692 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_301
timestamp 1676037725
transform 1 0 28796 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_307
timestamp 1676037725
transform 1 0 29348 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_309
timestamp 1676037725
transform 1 0 29532 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_321
timestamp 1676037725
transform 1 0 30636 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_333
timestamp 1676037725
transform 1 0 31740 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_345
timestamp 1676037725
transform 1 0 32844 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_357
timestamp 1676037725
transform 1 0 33948 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_363
timestamp 1676037725
transform 1 0 34500 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_365
timestamp 1676037725
transform 1 0 34684 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_377
timestamp 1676037725
transform 1 0 35788 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_389
timestamp 1676037725
transform 1 0 36892 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_401
timestamp 1676037725
transform 1 0 37996 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_413
timestamp 1676037725
transform 1 0 39100 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_419
timestamp 1676037725
transform 1 0 39652 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_421
timestamp 1676037725
transform 1 0 39836 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_433
timestamp 1676037725
transform 1 0 40940 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_445
timestamp 1676037725
transform 1 0 42044 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_457
timestamp 1676037725
transform 1 0 43148 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_469
timestamp 1676037725
transform 1 0 44252 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_475
timestamp 1676037725
transform 1 0 44804 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_477
timestamp 1676037725
transform 1 0 44988 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_489
timestamp 1676037725
transform 1 0 46092 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_501
timestamp 1676037725
transform 1 0 47196 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_513
timestamp 1676037725
transform 1 0 48300 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_525
timestamp 1676037725
transform 1 0 49404 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_531
timestamp 1676037725
transform 1 0 49956 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_533
timestamp 1676037725
transform 1 0 50140 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_545
timestamp 1676037725
transform 1 0 51244 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_557
timestamp 1676037725
transform 1 0 52348 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_569
timestamp 1676037725
transform 1 0 53452 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_581
timestamp 1676037725
transform 1 0 54556 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_587
timestamp 1676037725
transform 1 0 55108 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_100_589
timestamp 1676037725
transform 1 0 55292 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_100_601
timestamp 1676037725
transform 1 0 56396 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_611
timestamp 1676037725
transform 1 0 57316 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_621
timestamp 1676037725
transform 1 0 58236 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_3
timestamp 1676037725
transform 1 0 1380 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_101_11
timestamp 1676037725
transform 1 0 2116 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_101_17
timestamp 1676037725
transform 1 0 2668 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_101_25
timestamp 1676037725
transform 1 0 3404 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_101_29
timestamp 1676037725
transform 1 0 3772 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_101_35
timestamp 1676037725
transform 1 0 4324 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_101_45
timestamp 1676037725
transform 1 0 5244 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_101_53
timestamp 1676037725
transform 1 0 5980 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_101_57
timestamp 1676037725
transform 1 0 6348 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_101_63
timestamp 1676037725
transform 1 0 6900 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_101_73
timestamp 1676037725
transform 1 0 7820 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_101_81
timestamp 1676037725
transform 1 0 8556 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_101_85
timestamp 1676037725
transform 1 0 8924 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_101_91
timestamp 1676037725
transform 1 0 9476 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_101_101
timestamp 1676037725
transform 1 0 10396 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_101_109
timestamp 1676037725
transform 1 0 11132 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_101_113
timestamp 1676037725
transform 1 0 11500 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_101_119
timestamp 1676037725
transform 1 0 12052 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_101_131
timestamp 1676037725
transform 1 0 13156 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_101_139
timestamp 1676037725
transform 1 0 13892 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_101_141
timestamp 1676037725
transform 1 0 14076 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_149
timestamp 1676037725
transform 1 0 14812 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_157
timestamp 1676037725
transform 1 0 15548 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_101_165
timestamp 1676037725
transform 1 0 16284 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_101_169
timestamp 1676037725
transform 1 0 16652 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_101_175
timestamp 1676037725
transform 1 0 17204 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_101_185
timestamp 1676037725
transform 1 0 18124 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_101_193
timestamp 1676037725
transform 1 0 18860 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_101_197
timestamp 1676037725
transform 1 0 19228 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_101_203
timestamp 1676037725
transform 1 0 19780 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_101_213
timestamp 1676037725
transform 1 0 20700 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_101_221
timestamp 1676037725
transform 1 0 21436 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_101_225
timestamp 1676037725
transform 1 0 21804 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_101_231
timestamp 1676037725
transform 1 0 22356 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_101_243
timestamp 1676037725
transform 1 0 23460 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_101_251
timestamp 1676037725
transform 1 0 24196 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_101_253
timestamp 1676037725
transform 1 0 24380 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_101_259
timestamp 1676037725
transform 1 0 24932 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_101_269
timestamp 1676037725
transform 1 0 25852 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_101_277
timestamp 1676037725
transform 1 0 26588 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_101_281
timestamp 1676037725
transform 1 0 26956 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_101_287
timestamp 1676037725
transform 1 0 27508 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_101_297
timestamp 1676037725
transform 1 0 28428 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_101_305
timestamp 1676037725
transform 1 0 29164 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_101_309
timestamp 1676037725
transform 1 0 29532 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_101_315
timestamp 1676037725
transform 1 0 30084 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_101_325
timestamp 1676037725
transform 1 0 31004 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_101_333
timestamp 1676037725
transform 1 0 31740 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_101_337
timestamp 1676037725
transform 1 0 32108 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_101_343
timestamp 1676037725
transform 1 0 32660 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_101_353
timestamp 1676037725
transform 1 0 33580 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_101_361
timestamp 1676037725
transform 1 0 34316 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_101_365
timestamp 1676037725
transform 1 0 34684 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_101_371
timestamp 1676037725
transform 1 0 35236 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_101_381
timestamp 1676037725
transform 1 0 36156 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_101_389
timestamp 1676037725
transform 1 0 36892 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_101_393
timestamp 1676037725
transform 1 0 37260 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_101_399
timestamp 1676037725
transform 1 0 37812 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_101_409
timestamp 1676037725
transform 1 0 38732 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_101_417
timestamp 1676037725
transform 1 0 39468 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_101_421
timestamp 1676037725
transform 1 0 39836 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_101_427
timestamp 1676037725
transform 1 0 40388 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_101_437
timestamp 1676037725
transform 1 0 41308 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_101_445
timestamp 1676037725
transform 1 0 42044 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_101_449
timestamp 1676037725
transform 1 0 42412 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_101_455
timestamp 1676037725
transform 1 0 42964 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_101_465
timestamp 1676037725
transform 1 0 43884 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_101_473
timestamp 1676037725
transform 1 0 44620 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_101_477
timestamp 1676037725
transform 1 0 44988 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_101_483
timestamp 1676037725
transform 1 0 45540 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_101_493
timestamp 1676037725
transform 1 0 46460 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_101_501
timestamp 1676037725
transform 1 0 47196 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_101_505
timestamp 1676037725
transform 1 0 47564 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_101_511
timestamp 1676037725
transform 1 0 48116 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_101_521
timestamp 1676037725
transform 1 0 49036 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_101_529
timestamp 1676037725
transform 1 0 49772 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_101_533
timestamp 1676037725
transform 1 0 50140 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_101_539
timestamp 1676037725
transform 1 0 50692 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_101_549
timestamp 1676037725
transform 1 0 51612 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_101_557
timestamp 1676037725
transform 1 0 52348 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_101_561
timestamp 1676037725
transform 1 0 52716 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_101_567
timestamp 1676037725
transform 1 0 53268 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_101_579
timestamp 1676037725
transform 1 0 54372 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_101_587
timestamp 1676037725
transform 1 0 55108 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_101_589
timestamp 1676037725
transform 1 0 55292 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_595
timestamp 1676037725
transform 1 0 55844 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_599
timestamp 1676037725
transform 1 0 56212 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_604
timestamp 1676037725
transform 1 0 56672 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_614
timestamp 1676037725
transform 1 0 57592 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_617
timestamp 1676037725
transform 1 0 57868 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_623
timestamp 1676037725
transform 1 0 58420 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 58880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 58880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 58880 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 58880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 58880 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 58880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 58880 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 58880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 58880 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 58880 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 58880 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 58880 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 58880 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 58880 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 58880 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 58880 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1676037725
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1676037725
transform -1 0 58880 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1676037725
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1676037725
transform -1 0 58880 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1676037725
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1676037725
transform -1 0 58880 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1676037725
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1676037725
transform -1 0 58880 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1676037725
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1676037725
transform -1 0 58880 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1676037725
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1676037725
transform -1 0 58880 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1676037725
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1676037725
transform -1 0 58880 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1676037725
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1676037725
transform -1 0 58880 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1676037725
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1676037725
transform -1 0 58880 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1676037725
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1676037725
transform -1 0 58880 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1676037725
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1676037725
transform -1 0 58880 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1676037725
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1676037725
transform -1 0 58880 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1676037725
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1676037725
transform -1 0 58880 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1676037725
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1676037725
transform -1 0 58880 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1676037725
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1676037725
transform -1 0 58880 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1676037725
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1676037725
transform -1 0 58880 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1676037725
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1676037725
transform -1 0 58880 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1676037725
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1676037725
transform -1 0 58880 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1676037725
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1676037725
transform -1 0 58880 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1676037725
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1676037725
transform -1 0 58880 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1676037725
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1676037725
transform -1 0 58880 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1676037725
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1676037725
transform -1 0 58880 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1676037725
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1676037725
transform -1 0 58880 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1676037725
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1676037725
transform -1 0 58880 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1676037725
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1676037725
transform -1 0 58880 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1676037725
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1676037725
transform -1 0 58880 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1676037725
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1676037725
transform -1 0 58880 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1676037725
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1676037725
transform -1 0 58880 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1676037725
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1676037725
transform -1 0 58880 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1676037725
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1676037725
transform -1 0 58880 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1676037725
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1676037725
transform -1 0 58880 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1676037725
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1676037725
transform -1 0 58880 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1676037725
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1676037725
transform -1 0 58880 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1676037725
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1676037725
transform -1 0 58880 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1676037725
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1676037725
transform -1 0 58880 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1676037725
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1676037725
transform -1 0 58880 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1676037725
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1676037725
transform -1 0 58880 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1676037725
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1676037725
transform -1 0 58880 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1676037725
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1676037725
transform -1 0 58880 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1676037725
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1676037725
transform -1 0 58880 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1676037725
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1676037725
transform -1 0 58880 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1676037725
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1676037725
transform -1 0 58880 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1676037725
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1676037725
transform -1 0 58880 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1676037725
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1676037725
transform -1 0 58880 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1676037725
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1676037725
transform -1 0 58880 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1676037725
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1676037725
transform -1 0 58880 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1676037725
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1676037725
transform -1 0 58880 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1676037725
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1676037725
transform -1 0 58880 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1676037725
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1676037725
transform -1 0 58880 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1676037725
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1676037725
transform -1 0 58880 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1676037725
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1676037725
transform -1 0 58880 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1676037725
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1676037725
transform -1 0 58880 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1676037725
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1676037725
transform -1 0 58880 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1676037725
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1676037725
transform -1 0 58880 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1676037725
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1676037725
transform -1 0 58880 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1676037725
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1676037725
transform -1 0 58880 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1676037725
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1676037725
transform -1 0 58880 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1676037725
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1676037725
transform -1 0 58880 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1676037725
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1676037725
transform -1 0 58880 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1676037725
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1676037725
transform -1 0 58880 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1676037725
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1676037725
transform -1 0 58880 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1676037725
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1676037725
transform -1 0 58880 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1676037725
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1676037725
transform -1 0 58880 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1676037725
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1676037725
transform -1 0 58880 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1676037725
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1676037725
transform -1 0 58880 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1676037725
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1676037725
transform -1 0 58880 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1676037725
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1676037725
transform -1 0 58880 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1676037725
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1676037725
transform -1 0 58880 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1676037725
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1676037725
transform -1 0 58880 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1676037725
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1676037725
transform -1 0 58880 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1676037725
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1676037725
transform -1 0 58880 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1676037725
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1676037725
transform -1 0 58880 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1676037725
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1676037725
transform -1 0 58880 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1676037725
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1676037725
transform -1 0 58880 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1676037725
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1676037725
transform -1 0 58880 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1676037725
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1676037725
transform -1 0 58880 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1676037725
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1676037725
transform -1 0 58880 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1676037725
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1676037725
transform -1 0 58880 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1676037725
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1676037725
transform -1 0 58880 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1676037725
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1676037725
transform -1 0 58880 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1676037725
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1676037725
transform -1 0 58880 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 1676037725
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 1676037725
transform -1 0 58880 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 1676037725
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 1676037725
transform -1 0 58880 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 1676037725
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 1676037725
transform -1 0 58880 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 1676037725
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 1676037725
transform -1 0 58880 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 1676037725
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 1676037725
transform -1 0 58880 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1676037725
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1676037725
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1676037725
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1676037725
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1676037725
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1676037725
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1676037725
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1676037725
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1676037725
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1676037725
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1676037725
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1676037725
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1676037725
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1676037725
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1676037725
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1676037725
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1676037725
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1676037725
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1676037725
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1676037725
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1676037725
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1676037725
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1676037725
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1676037725
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1676037725
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1676037725
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1676037725
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1676037725
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1676037725
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1676037725
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1676037725
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1676037725
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1676037725
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1676037725
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1676037725
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1676037725
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1676037725
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1676037725
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1676037725
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1676037725
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1676037725
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1676037725
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1676037725
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1676037725
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1676037725
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1676037725
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1676037725
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1676037725
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1676037725
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1676037725
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1676037725
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1676037725
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1676037725
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1676037725
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1676037725
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1676037725
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1676037725
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1676037725
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1676037725
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1676037725
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1676037725
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1676037725
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1676037725
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1676037725
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1676037725
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1676037725
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1676037725
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1676037725
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1676037725
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1676037725
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1676037725
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1676037725
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1676037725
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1676037725
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1676037725
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1676037725
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1676037725
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1676037725
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1676037725
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1676037725
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1676037725
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1676037725
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1676037725
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1676037725
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1676037725
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1676037725
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1676037725
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1676037725
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1676037725
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1676037725
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1676037725
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1676037725
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1676037725
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1676037725
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1676037725
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1676037725
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1676037725
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1676037725
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1676037725
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1676037725
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1676037725
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1676037725
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1676037725
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1676037725
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1676037725
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1676037725
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1676037725
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1676037725
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1676037725
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1676037725
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1676037725
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1676037725
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1676037725
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1676037725
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1676037725
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1676037725
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1676037725
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1676037725
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1676037725
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1676037725
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1676037725
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1676037725
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1676037725
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1676037725
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1676037725
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1676037725
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1676037725
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1676037725
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1676037725
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1676037725
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1676037725
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1676037725
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1676037725
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1676037725
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1676037725
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1676037725
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1676037725
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1676037725
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1676037725
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1676037725
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1676037725
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1676037725
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1676037725
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1676037725
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1676037725
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1676037725
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1676037725
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1676037725
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1676037725
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1676037725
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1676037725
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1676037725
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1676037725
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1676037725
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1676037725
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1676037725
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1676037725
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1676037725
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1676037725
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1676037725
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1676037725
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1676037725
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1676037725
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1676037725
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1676037725
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1676037725
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1676037725
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1676037725
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1676037725
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1676037725
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1676037725
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1676037725
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1676037725
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1676037725
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1676037725
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1676037725
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1676037725
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1676037725
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1676037725
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1676037725
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1676037725
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1676037725
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1676037725
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1676037725
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1676037725
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1676037725
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1676037725
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1676037725
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1676037725
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1676037725
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1676037725
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1676037725
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1676037725
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1676037725
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1676037725
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1676037725
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1676037725
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1676037725
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1676037725
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1676037725
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1676037725
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1676037725
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1676037725
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1676037725
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1676037725
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1676037725
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1676037725
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1676037725
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1676037725
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1676037725
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1676037725
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1676037725
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1676037725
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1676037725
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1676037725
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1676037725
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1676037725
transform 1 0 57776 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1676037725
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1676037725
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1676037725
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1676037725
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1676037725
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1676037725
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1676037725
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1676037725
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1676037725
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1676037725
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1676037725
transform 1 0 55200 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1676037725
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1676037725
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1676037725
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1676037725
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1676037725
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1676037725
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1676037725
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1676037725
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1676037725
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1676037725
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1676037725
transform 1 0 57776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1676037725
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1676037725
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1676037725
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1676037725
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1676037725
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1676037725
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1676037725
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1676037725
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1676037725
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1676037725
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1676037725
transform 1 0 55200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1676037725
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1676037725
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1676037725
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1676037725
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1676037725
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1676037725
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1676037725
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1676037725
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1676037725
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1676037725
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1676037725
transform 1 0 57776 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1676037725
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1676037725
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1676037725
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1676037725
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1676037725
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1676037725
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1676037725
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1676037725
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1676037725
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1676037725
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1676037725
transform 1 0 55200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1676037725
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1676037725
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1676037725
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1676037725
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1676037725
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1676037725
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1676037725
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1676037725
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1676037725
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1676037725
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1676037725
transform 1 0 57776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1676037725
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1676037725
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1676037725
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1676037725
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1676037725
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1676037725
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1676037725
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1676037725
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1676037725
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1676037725
transform 1 0 50048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1676037725
transform 1 0 55200 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1676037725
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1676037725
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1676037725
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1676037725
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1676037725
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1676037725
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1676037725
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1676037725
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1676037725
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1676037725
transform 1 0 52624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1676037725
transform 1 0 57776 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1676037725
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1676037725
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1676037725
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1676037725
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1676037725
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1676037725
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1676037725
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1676037725
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1676037725
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1676037725
transform 1 0 50048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1676037725
transform 1 0 55200 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1676037725
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1676037725
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1676037725
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1676037725
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1676037725
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1676037725
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1676037725
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1676037725
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1676037725
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1676037725
transform 1 0 52624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1676037725
transform 1 0 57776 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1676037725
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1676037725
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1676037725
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1676037725
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1676037725
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1676037725
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1676037725
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1676037725
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1676037725
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1676037725
transform 1 0 50048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1676037725
transform 1 0 55200 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1676037725
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1676037725
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1676037725
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1676037725
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1676037725
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1676037725
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1676037725
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1676037725
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1676037725
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1676037725
transform 1 0 52624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1676037725
transform 1 0 57776 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1676037725
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1676037725
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1676037725
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1676037725
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1676037725
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1676037725
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1676037725
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1676037725
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1676037725
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1676037725
transform 1 0 50048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1676037725
transform 1 0 55200 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1676037725
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1676037725
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1676037725
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1676037725
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1676037725
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1676037725
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1676037725
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1676037725
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1676037725
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1676037725
transform 1 0 52624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1676037725
transform 1 0 57776 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1676037725
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1676037725
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1676037725
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1676037725
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1676037725
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1676037725
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1676037725
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1676037725
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1676037725
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1676037725
transform 1 0 50048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1676037725
transform 1 0 55200 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1676037725
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1676037725
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1676037725
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1676037725
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1676037725
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1676037725
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1676037725
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1676037725
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1676037725
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1676037725
transform 1 0 52624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1676037725
transform 1 0 57776 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1676037725
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1676037725
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1676037725
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1676037725
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1676037725
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1676037725
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1676037725
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1676037725
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1676037725
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1676037725
transform 1 0 50048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1676037725
transform 1 0 55200 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1676037725
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1676037725
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1676037725
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1676037725
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1676037725
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1676037725
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1676037725
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1676037725
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1676037725
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1676037725
transform 1 0 52624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1676037725
transform 1 0 57776 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1676037725
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1676037725
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1676037725
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1676037725
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1676037725
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1676037725
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1676037725
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1676037725
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1676037725
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1676037725
transform 1 0 50048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1676037725
transform 1 0 55200 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1676037725
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1676037725
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1676037725
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1676037725
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1676037725
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1676037725
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1676037725
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1676037725
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1676037725
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1676037725
transform 1 0 52624 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1676037725
transform 1 0 57776 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1676037725
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1676037725
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1676037725
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1676037725
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1676037725
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1676037725
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1676037725
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1676037725
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1676037725
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1676037725
transform 1 0 50048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1676037725
transform 1 0 55200 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1676037725
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1676037725
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1676037725
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1676037725
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1676037725
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1676037725
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1676037725
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1676037725
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1676037725
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1676037725
transform 1 0 52624 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1676037725
transform 1 0 57776 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1676037725
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1676037725
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1676037725
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1676037725
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1676037725
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1676037725
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1676037725
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1676037725
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1676037725
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1676037725
transform 1 0 50048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1676037725
transform 1 0 55200 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1676037725
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1676037725
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1676037725
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1676037725
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1676037725
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1676037725
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1676037725
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1676037725
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1676037725
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1676037725
transform 1 0 52624 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1676037725
transform 1 0 57776 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1676037725
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1676037725
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1676037725
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1676037725
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1676037725
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1676037725
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1676037725
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1676037725
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1676037725
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1676037725
transform 1 0 50048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1676037725
transform 1 0 55200 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1676037725
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1676037725
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1676037725
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1676037725
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1676037725
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1676037725
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1676037725
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1676037725
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1676037725
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1676037725
transform 1 0 52624 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1676037725
transform 1 0 57776 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1676037725
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1676037725
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1676037725
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1676037725
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1676037725
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1676037725
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1676037725
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1676037725
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1676037725
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1676037725
transform 1 0 50048 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1676037725
transform 1 0 55200 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1676037725
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1676037725
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1676037725
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1676037725
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1676037725
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1676037725
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1676037725
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1676037725
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1676037725
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1676037725
transform 1 0 52624 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1676037725
transform 1 0 57776 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1676037725
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1676037725
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1676037725
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1676037725
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1676037725
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1676037725
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1676037725
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1676037725
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1676037725
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1676037725
transform 1 0 50048 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1676037725
transform 1 0 55200 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1676037725
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1676037725
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1676037725
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1676037725
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1676037725
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1676037725
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1676037725
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1676037725
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1676037725
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1676037725
transform 1 0 52624 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1676037725
transform 1 0 57776 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1676037725
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1676037725
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1676037725
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1676037725
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1676037725
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1676037725
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1676037725
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1676037725
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1676037725
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1676037725
transform 1 0 50048 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1676037725
transform 1 0 55200 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1676037725
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1676037725
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1676037725
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1676037725
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1676037725
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1676037725
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1676037725
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1676037725
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1676037725
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1676037725
transform 1 0 52624 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1676037725
transform 1 0 57776 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1676037725
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1676037725
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1676037725
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1676037725
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1676037725
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1676037725
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1676037725
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1676037725
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1676037725
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1676037725
transform 1 0 50048 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1676037725
transform 1 0 55200 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1676037725
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1676037725
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1676037725
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1676037725
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1676037725
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1676037725
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1676037725
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1676037725
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1676037725
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1676037725
transform 1 0 52624 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1676037725
transform 1 0 57776 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1676037725
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1676037725
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1676037725
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1676037725
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1676037725
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1676037725
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1676037725
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1676037725
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1676037725
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1676037725
transform 1 0 50048 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1676037725
transform 1 0 55200 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1676037725
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1676037725
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1676037725
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1676037725
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1676037725
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1676037725
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1676037725
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1676037725
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1676037725
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1676037725
transform 1 0 52624 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1676037725
transform 1 0 57776 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1676037725
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1676037725
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1676037725
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1676037725
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1676037725
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1676037725
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1676037725
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1676037725
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1676037725
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1676037725
transform 1 0 50048 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1676037725
transform 1 0 55200 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1676037725
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1676037725
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1676037725
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1676037725
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1676037725
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1676037725
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1676037725
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1676037725
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1676037725
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1676037725
transform 1 0 52624 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1676037725
transform 1 0 57776 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1676037725
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1676037725
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1676037725
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1676037725
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1676037725
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1676037725
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1676037725
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1676037725
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1676037725
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1676037725
transform 1 0 50048 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1676037725
transform 1 0 55200 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1676037725
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1676037725
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1676037725
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1676037725
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1676037725
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1676037725
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1676037725
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1676037725
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1676037725
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1676037725
transform 1 0 52624 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1676037725
transform 1 0 57776 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1676037725
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1676037725
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1676037725
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1676037725
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1676037725
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1676037725
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1676037725
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1676037725
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1676037725
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1676037725
transform 1 0 50048 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1676037725
transform 1 0 55200 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1676037725
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1676037725
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1676037725
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1676037725
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1676037725
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1676037725
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1676037725
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1676037725
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1676037725
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1676037725
transform 1 0 52624 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1676037725
transform 1 0 57776 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1676037725
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1676037725
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1676037725
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1676037725
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1676037725
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1676037725
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1676037725
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1676037725
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1676037725
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1676037725
transform 1 0 50048 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1676037725
transform 1 0 55200 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1676037725
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1676037725
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1676037725
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1676037725
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1676037725
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1676037725
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1676037725
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1676037725
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1676037725
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1676037725
transform 1 0 52624 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1676037725
transform 1 0 57776 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1676037725
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1676037725
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1676037725
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1676037725
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1676037725
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1676037725
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1676037725
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1676037725
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1676037725
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1676037725
transform 1 0 50048 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1676037725
transform 1 0 55200 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1676037725
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1676037725
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1676037725
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1676037725
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1676037725
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1676037725
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1676037725
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1676037725
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1676037725
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1676037725
transform 1 0 52624 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1676037725
transform 1 0 57776 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1676037725
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1676037725
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1676037725
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1676037725
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1676037725
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_968
timestamp 1676037725
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_969
timestamp 1676037725
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_970
timestamp 1676037725
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_971
timestamp 1676037725
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_972
timestamp 1676037725
transform 1 0 50048 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_973
timestamp 1676037725
transform 1 0 55200 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_974
timestamp 1676037725
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_975
timestamp 1676037725
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_976
timestamp 1676037725
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_977
timestamp 1676037725
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_978
timestamp 1676037725
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_979
timestamp 1676037725
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_980
timestamp 1676037725
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_981
timestamp 1676037725
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_982
timestamp 1676037725
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_983
timestamp 1676037725
transform 1 0 52624 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_984
timestamp 1676037725
transform 1 0 57776 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_985
timestamp 1676037725
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_986
timestamp 1676037725
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_987
timestamp 1676037725
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_988
timestamp 1676037725
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_989
timestamp 1676037725
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_990
timestamp 1676037725
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_991
timestamp 1676037725
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_992
timestamp 1676037725
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_993
timestamp 1676037725
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_994
timestamp 1676037725
transform 1 0 50048 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_995
timestamp 1676037725
transform 1 0 55200 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_996
timestamp 1676037725
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_997
timestamp 1676037725
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_998
timestamp 1676037725
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_999
timestamp 1676037725
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1000
timestamp 1676037725
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1001
timestamp 1676037725
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1002
timestamp 1676037725
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1003
timestamp 1676037725
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1004
timestamp 1676037725
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1005
timestamp 1676037725
transform 1 0 52624 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1006
timestamp 1676037725
transform 1 0 57776 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1007
timestamp 1676037725
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1008
timestamp 1676037725
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1009
timestamp 1676037725
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1010
timestamp 1676037725
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1011
timestamp 1676037725
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1012
timestamp 1676037725
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1013
timestamp 1676037725
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1014
timestamp 1676037725
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1015
timestamp 1676037725
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1016
timestamp 1676037725
transform 1 0 50048 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1017
timestamp 1676037725
transform 1 0 55200 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1018
timestamp 1676037725
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1019
timestamp 1676037725
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1020
timestamp 1676037725
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1021
timestamp 1676037725
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1022
timestamp 1676037725
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1023
timestamp 1676037725
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1024
timestamp 1676037725
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1025
timestamp 1676037725
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1026
timestamp 1676037725
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1027
timestamp 1676037725
transform 1 0 52624 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1028
timestamp 1676037725
transform 1 0 57776 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1029
timestamp 1676037725
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1030
timestamp 1676037725
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1031
timestamp 1676037725
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1032
timestamp 1676037725
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1033
timestamp 1676037725
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1034
timestamp 1676037725
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1035
timestamp 1676037725
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1036
timestamp 1676037725
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1037
timestamp 1676037725
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1038
timestamp 1676037725
transform 1 0 50048 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1039
timestamp 1676037725
transform 1 0 55200 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1040
timestamp 1676037725
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1041
timestamp 1676037725
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1042
timestamp 1676037725
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1043
timestamp 1676037725
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1044
timestamp 1676037725
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1045
timestamp 1676037725
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1046
timestamp 1676037725
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1047
timestamp 1676037725
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1048
timestamp 1676037725
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1049
timestamp 1676037725
transform 1 0 52624 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1050
timestamp 1676037725
transform 1 0 57776 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1051
timestamp 1676037725
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1052
timestamp 1676037725
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1053
timestamp 1676037725
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1054
timestamp 1676037725
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1055
timestamp 1676037725
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1056
timestamp 1676037725
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1057
timestamp 1676037725
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1058
timestamp 1676037725
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1059
timestamp 1676037725
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1060
timestamp 1676037725
transform 1 0 50048 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1061
timestamp 1676037725
transform 1 0 55200 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1062
timestamp 1676037725
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1063
timestamp 1676037725
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1064
timestamp 1676037725
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1065
timestamp 1676037725
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1066
timestamp 1676037725
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1067
timestamp 1676037725
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1068
timestamp 1676037725
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1069
timestamp 1676037725
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1070
timestamp 1676037725
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1071
timestamp 1676037725
transform 1 0 52624 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1072
timestamp 1676037725
transform 1 0 57776 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1073
timestamp 1676037725
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1074
timestamp 1676037725
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1075
timestamp 1676037725
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1076
timestamp 1676037725
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1077
timestamp 1676037725
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1078
timestamp 1676037725
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1079
timestamp 1676037725
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1080
timestamp 1676037725
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1081
timestamp 1676037725
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1082
timestamp 1676037725
transform 1 0 50048 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1083
timestamp 1676037725
transform 1 0 55200 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1084
timestamp 1676037725
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1085
timestamp 1676037725
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1086
timestamp 1676037725
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1087
timestamp 1676037725
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1088
timestamp 1676037725
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1089
timestamp 1676037725
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1090
timestamp 1676037725
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1091
timestamp 1676037725
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1092
timestamp 1676037725
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1093
timestamp 1676037725
transform 1 0 52624 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1094
timestamp 1676037725
transform 1 0 57776 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1095
timestamp 1676037725
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1096
timestamp 1676037725
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1097
timestamp 1676037725
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1098
timestamp 1676037725
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1099
timestamp 1676037725
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1100
timestamp 1676037725
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1101
timestamp 1676037725
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1102
timestamp 1676037725
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1103
timestamp 1676037725
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1104
timestamp 1676037725
transform 1 0 50048 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1105
timestamp 1676037725
transform 1 0 55200 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1106
timestamp 1676037725
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1107
timestamp 1676037725
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1108
timestamp 1676037725
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1109
timestamp 1676037725
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1110
timestamp 1676037725
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1111
timestamp 1676037725
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1112
timestamp 1676037725
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1113
timestamp 1676037725
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1114
timestamp 1676037725
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1115
timestamp 1676037725
transform 1 0 52624 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1116
timestamp 1676037725
transform 1 0 57776 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1117
timestamp 1676037725
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1118
timestamp 1676037725
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1119
timestamp 1676037725
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1120
timestamp 1676037725
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1121
timestamp 1676037725
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1122
timestamp 1676037725
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1123
timestamp 1676037725
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1124
timestamp 1676037725
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1125
timestamp 1676037725
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1126
timestamp 1676037725
transform 1 0 50048 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1127
timestamp 1676037725
transform 1 0 55200 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1128
timestamp 1676037725
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1129
timestamp 1676037725
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1130
timestamp 1676037725
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1131
timestamp 1676037725
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1132
timestamp 1676037725
transform 1 0 26864 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1133
timestamp 1676037725
transform 1 0 32016 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1134
timestamp 1676037725
transform 1 0 37168 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1135
timestamp 1676037725
transform 1 0 42320 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1136
timestamp 1676037725
transform 1 0 47472 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1137
timestamp 1676037725
transform 1 0 52624 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1138
timestamp 1676037725
transform 1 0 57776 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1139
timestamp 1676037725
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1140
timestamp 1676037725
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1141
timestamp 1676037725
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1142
timestamp 1676037725
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1143
timestamp 1676037725
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1144
timestamp 1676037725
transform 1 0 29440 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1145
timestamp 1676037725
transform 1 0 34592 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1146
timestamp 1676037725
transform 1 0 39744 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1147
timestamp 1676037725
transform 1 0 44896 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1148
timestamp 1676037725
transform 1 0 50048 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1149
timestamp 1676037725
transform 1 0 55200 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1150
timestamp 1676037725
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1151
timestamp 1676037725
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1152
timestamp 1676037725
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1153
timestamp 1676037725
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1154
timestamp 1676037725
transform 1 0 26864 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1155
timestamp 1676037725
transform 1 0 32016 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1156
timestamp 1676037725
transform 1 0 37168 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1157
timestamp 1676037725
transform 1 0 42320 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1158
timestamp 1676037725
transform 1 0 47472 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1159
timestamp 1676037725
transform 1 0 52624 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1160
timestamp 1676037725
transform 1 0 57776 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1161
timestamp 1676037725
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1162
timestamp 1676037725
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1163
timestamp 1676037725
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1164
timestamp 1676037725
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1165
timestamp 1676037725
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1166
timestamp 1676037725
transform 1 0 29440 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1167
timestamp 1676037725
transform 1 0 34592 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1168
timestamp 1676037725
transform 1 0 39744 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1169
timestamp 1676037725
transform 1 0 44896 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1170
timestamp 1676037725
transform 1 0 50048 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1171
timestamp 1676037725
transform 1 0 55200 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1172
timestamp 1676037725
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1173
timestamp 1676037725
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1174
timestamp 1676037725
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1175
timestamp 1676037725
transform 1 0 21712 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1176
timestamp 1676037725
transform 1 0 26864 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1177
timestamp 1676037725
transform 1 0 32016 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1178
timestamp 1676037725
transform 1 0 37168 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1179
timestamp 1676037725
transform 1 0 42320 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1180
timestamp 1676037725
transform 1 0 47472 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1181
timestamp 1676037725
transform 1 0 52624 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1182
timestamp 1676037725
transform 1 0 57776 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1183
timestamp 1676037725
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1184
timestamp 1676037725
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1185
timestamp 1676037725
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1186
timestamp 1676037725
transform 1 0 19136 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1187
timestamp 1676037725
transform 1 0 24288 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1188
timestamp 1676037725
transform 1 0 29440 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1189
timestamp 1676037725
transform 1 0 34592 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1190
timestamp 1676037725
transform 1 0 39744 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1191
timestamp 1676037725
transform 1 0 44896 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1192
timestamp 1676037725
transform 1 0 50048 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1193
timestamp 1676037725
transform 1 0 55200 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1194
timestamp 1676037725
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1195
timestamp 1676037725
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1196
timestamp 1676037725
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1197
timestamp 1676037725
transform 1 0 21712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1198
timestamp 1676037725
transform 1 0 26864 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1199
timestamp 1676037725
transform 1 0 32016 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1200
timestamp 1676037725
transform 1 0 37168 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1201
timestamp 1676037725
transform 1 0 42320 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1202
timestamp 1676037725
transform 1 0 47472 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1203
timestamp 1676037725
transform 1 0 52624 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1204
timestamp 1676037725
transform 1 0 57776 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1205
timestamp 1676037725
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1206
timestamp 1676037725
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1207
timestamp 1676037725
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1208
timestamp 1676037725
transform 1 0 19136 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1209
timestamp 1676037725
transform 1 0 24288 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1210
timestamp 1676037725
transform 1 0 29440 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1211
timestamp 1676037725
transform 1 0 34592 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1212
timestamp 1676037725
transform 1 0 39744 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1213
timestamp 1676037725
transform 1 0 44896 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1214
timestamp 1676037725
transform 1 0 50048 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1215
timestamp 1676037725
transform 1 0 55200 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1216
timestamp 1676037725
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1217
timestamp 1676037725
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1218
timestamp 1676037725
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1219
timestamp 1676037725
transform 1 0 21712 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1220
timestamp 1676037725
transform 1 0 26864 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1221
timestamp 1676037725
transform 1 0 32016 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1222
timestamp 1676037725
transform 1 0 37168 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1223
timestamp 1676037725
transform 1 0 42320 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1224
timestamp 1676037725
transform 1 0 47472 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1225
timestamp 1676037725
transform 1 0 52624 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1226
timestamp 1676037725
transform 1 0 57776 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1227
timestamp 1676037725
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1228
timestamp 1676037725
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1229
timestamp 1676037725
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1230
timestamp 1676037725
transform 1 0 19136 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1231
timestamp 1676037725
transform 1 0 24288 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1232
timestamp 1676037725
transform 1 0 29440 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1233
timestamp 1676037725
transform 1 0 34592 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1234
timestamp 1676037725
transform 1 0 39744 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1235
timestamp 1676037725
transform 1 0 44896 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1236
timestamp 1676037725
transform 1 0 50048 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1237
timestamp 1676037725
transform 1 0 55200 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1238
timestamp 1676037725
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1239
timestamp 1676037725
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1240
timestamp 1676037725
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1241
timestamp 1676037725
transform 1 0 21712 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1242
timestamp 1676037725
transform 1 0 26864 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1243
timestamp 1676037725
transform 1 0 32016 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1244
timestamp 1676037725
transform 1 0 37168 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1245
timestamp 1676037725
transform 1 0 42320 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1246
timestamp 1676037725
transform 1 0 47472 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1247
timestamp 1676037725
transform 1 0 52624 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1248
timestamp 1676037725
transform 1 0 57776 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1249
timestamp 1676037725
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1250
timestamp 1676037725
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1251
timestamp 1676037725
transform 1 0 13984 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1252
timestamp 1676037725
transform 1 0 19136 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1253
timestamp 1676037725
transform 1 0 24288 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1254
timestamp 1676037725
transform 1 0 29440 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1255
timestamp 1676037725
transform 1 0 34592 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1256
timestamp 1676037725
transform 1 0 39744 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1257
timestamp 1676037725
transform 1 0 44896 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1258
timestamp 1676037725
transform 1 0 50048 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1259
timestamp 1676037725
transform 1 0 55200 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1260
timestamp 1676037725
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1261
timestamp 1676037725
transform 1 0 11408 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1262
timestamp 1676037725
transform 1 0 16560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1263
timestamp 1676037725
transform 1 0 21712 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1264
timestamp 1676037725
transform 1 0 26864 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1265
timestamp 1676037725
transform 1 0 32016 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1266
timestamp 1676037725
transform 1 0 37168 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1267
timestamp 1676037725
transform 1 0 42320 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1268
timestamp 1676037725
transform 1 0 47472 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1269
timestamp 1676037725
transform 1 0 52624 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1270
timestamp 1676037725
transform 1 0 57776 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1271
timestamp 1676037725
transform 1 0 3680 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1272
timestamp 1676037725
transform 1 0 8832 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1273
timestamp 1676037725
transform 1 0 13984 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1274
timestamp 1676037725
transform 1 0 19136 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1275
timestamp 1676037725
transform 1 0 24288 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1276
timestamp 1676037725
transform 1 0 29440 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1277
timestamp 1676037725
transform 1 0 34592 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1278
timestamp 1676037725
transform 1 0 39744 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1279
timestamp 1676037725
transform 1 0 44896 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1280
timestamp 1676037725
transform 1 0 50048 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1281
timestamp 1676037725
transform 1 0 55200 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1282
timestamp 1676037725
transform 1 0 6256 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1283
timestamp 1676037725
transform 1 0 11408 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1284
timestamp 1676037725
transform 1 0 16560 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1285
timestamp 1676037725
transform 1 0 21712 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1286
timestamp 1676037725
transform 1 0 26864 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1287
timestamp 1676037725
transform 1 0 32016 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1288
timestamp 1676037725
transform 1 0 37168 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1289
timestamp 1676037725
transform 1 0 42320 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1290
timestamp 1676037725
transform 1 0 47472 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1291
timestamp 1676037725
transform 1 0 52624 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1292
timestamp 1676037725
transform 1 0 57776 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1293
timestamp 1676037725
transform 1 0 3680 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1294
timestamp 1676037725
transform 1 0 8832 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1295
timestamp 1676037725
transform 1 0 13984 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1296
timestamp 1676037725
transform 1 0 19136 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1297
timestamp 1676037725
transform 1 0 24288 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1298
timestamp 1676037725
transform 1 0 29440 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1299
timestamp 1676037725
transform 1 0 34592 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1300
timestamp 1676037725
transform 1 0 39744 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1301
timestamp 1676037725
transform 1 0 44896 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1302
timestamp 1676037725
transform 1 0 50048 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1303
timestamp 1676037725
transform 1 0 55200 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1304
timestamp 1676037725
transform 1 0 6256 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1305
timestamp 1676037725
transform 1 0 11408 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1306
timestamp 1676037725
transform 1 0 16560 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1307
timestamp 1676037725
transform 1 0 21712 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1308
timestamp 1676037725
transform 1 0 26864 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1309
timestamp 1676037725
transform 1 0 32016 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1310
timestamp 1676037725
transform 1 0 37168 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1311
timestamp 1676037725
transform 1 0 42320 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1312
timestamp 1676037725
transform 1 0 47472 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1313
timestamp 1676037725
transform 1 0 52624 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1314
timestamp 1676037725
transform 1 0 57776 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1315
timestamp 1676037725
transform 1 0 3680 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1316
timestamp 1676037725
transform 1 0 8832 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1317
timestamp 1676037725
transform 1 0 13984 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1318
timestamp 1676037725
transform 1 0 19136 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1319
timestamp 1676037725
transform 1 0 24288 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1320
timestamp 1676037725
transform 1 0 29440 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1321
timestamp 1676037725
transform 1 0 34592 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1322
timestamp 1676037725
transform 1 0 39744 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1323
timestamp 1676037725
transform 1 0 44896 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1324
timestamp 1676037725
transform 1 0 50048 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1325
timestamp 1676037725
transform 1 0 55200 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1326
timestamp 1676037725
transform 1 0 3680 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1327
timestamp 1676037725
transform 1 0 6256 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1328
timestamp 1676037725
transform 1 0 8832 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1329
timestamp 1676037725
transform 1 0 11408 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1330
timestamp 1676037725
transform 1 0 13984 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1331
timestamp 1676037725
transform 1 0 16560 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1332
timestamp 1676037725
transform 1 0 19136 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1333
timestamp 1676037725
transform 1 0 21712 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1334
timestamp 1676037725
transform 1 0 24288 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1335
timestamp 1676037725
transform 1 0 26864 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1336
timestamp 1676037725
transform 1 0 29440 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1337
timestamp 1676037725
transform 1 0 32016 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1338
timestamp 1676037725
transform 1 0 34592 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1339
timestamp 1676037725
transform 1 0 37168 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1340
timestamp 1676037725
transform 1 0 39744 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1341
timestamp 1676037725
transform 1 0 42320 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1342
timestamp 1676037725
transform 1 0 44896 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1343
timestamp 1676037725
transform 1 0 47472 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1344
timestamp 1676037725
transform 1 0 50048 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1345
timestamp 1676037725
transform 1 0 52624 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1346
timestamp 1676037725
transform 1 0 55200 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1347
timestamp 1676037725
transform 1 0 57776 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  _0446_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 41492 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0447_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 37260 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0448_
timestamp 1676037725
transform 1 0 35604 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0449_
timestamp 1676037725
transform 1 0 29164 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0450_
timestamp 1676037725
transform 1 0 31556 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0451_
timestamp 1676037725
transform 1 0 37352 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0452_
timestamp 1676037725
transform 1 0 40112 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0453_
timestamp 1676037725
transform 1 0 43976 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0454_
timestamp 1676037725
transform 1 0 46644 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0455_
timestamp 1676037725
transform 1 0 48760 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0456_
timestamp 1676037725
transform 1 0 43424 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0457_
timestamp 1676037725
transform 1 0 26772 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_2  _0458_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25024 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__nor4b_4  _0459_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 22908 0 -1 28288
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_4  _0460_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9108 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2b_2  _0461_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21896 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nor4b_4  _0462_
timestamp 1676037725
transform 1 0 22908 0 -1 29376
box -38 -48 1786 592
use sky130_fd_sc_hd__nand2b_1  _0463_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15732 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_4  _0464_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 22632 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_2  _0465_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23920 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_4  _0466_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 22816 0 -1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2b_1  _0467_
timestamp 1676037725
transform 1 0 2484 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_4  _0468_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24748 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nand2b_1  _0469_
timestamp 1676037725
transform 1 0 24012 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nor4b_4  _0470_
timestamp 1676037725
transform 1 0 23000 0 -1 25024
box -38 -48 1786 592
use sky130_fd_sc_hd__nand2b_1  _0471_
timestamp 1676037725
transform 1 0 2484 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_4  _0472_
timestamp 1676037725
transform 1 0 22908 0 1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2b_1  _0473_
timestamp 1676037725
transform 1 0 2484 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_4  _0474_
timestamp 1676037725
transform 1 0 22908 0 1 28288
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2b_1  _0475_
timestamp 1676037725
transform 1 0 2484 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _0476_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25208 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or3_4  _0477_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 22816 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__nor3b_2  _0478_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24564 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__nor4b_2  _0479_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25024 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2b_2  _0480_
timestamp 1676037725
transform 1 0 21712 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_4  _0481_
timestamp 1676037725
transform 1 0 22908 0 1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2b_2  _0482_
timestamp 1676037725
transform 1 0 21896 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_4  _0483_
timestamp 1676037725
transform 1 0 22816 0 -1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2b_2  _0484_
timestamp 1676037725
transform 1 0 20884 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_4  _0485_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23184 0 -1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__nand2b_2  _0486_
timestamp 1676037725
transform 1 0 21988 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_1  _0487_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 22632 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__nand2b_1  _0488_
timestamp 1676037725
transform 1 0 2484 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0489_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25300 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _0490_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 38364 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0491_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25760 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0492_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 26128 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_4  _0493_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 26312 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _0494_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 29532 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0495_
timestamp 1676037725
transform 1 0 30268 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0496_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 26220 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _0497_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27140 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or3_4  _0498_
timestamp 1676037725
transform 1 0 27508 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__or2_2  _0499_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 31096 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_4  _0500_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10672 0 1 15232
box -38 -48 1326 592
use sky130_fd_sc_hd__a21o_2  _0501_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23644 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or3_4  _0502_
timestamp 1676037725
transform 1 0 24564 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _0503_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24012 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _0504_
timestamp 1676037725
transform 1 0 14812 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _0505_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24564 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_2  _0506_
timestamp 1676037725
transform 1 0 26128 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_4  _0507_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24656 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__nor4_4  _0508_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23184 0 -1 23936
box -38 -48 1602 592
use sky130_fd_sc_hd__a211o_1  _0509_
timestamp 1676037725
transform 1 0 34500 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _0510_
timestamp 1676037725
transform 1 0 33764 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or3_4  _0511_
timestamp 1676037725
transform 1 0 25852 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and2_4  _0512_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 31464 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0513_
timestamp 1676037725
transform 1 0 37444 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0514_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 29716 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0515_
timestamp 1676037725
transform 1 0 29716 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0516_
timestamp 1676037725
transform 1 0 37260 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or3_4  _0517_
timestamp 1676037725
transform 1 0 30084 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0518_
timestamp 1676037725
transform 1 0 37260 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0519_
timestamp 1676037725
transform 1 0 27692 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0520_
timestamp 1676037725
transform 1 0 27140 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0521_
timestamp 1676037725
transform 1 0 28152 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0522_
timestamp 1676037725
transform 1 0 27508 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or3_4  _0523_
timestamp 1676037725
transform 1 0 28152 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_2  _0524_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24840 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_4  _0525_
timestamp 1676037725
transform 1 0 29992 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _0526_
timestamp 1676037725
transform 1 0 31004 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0527_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 32016 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_2  _0528_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 30728 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_2  _0529_
timestamp 1676037725
transform 1 0 26404 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0530_
timestamp 1676037725
transform 1 0 33304 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or3_2  _0531_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 31372 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0532_
timestamp 1676037725
transform 1 0 47748 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0533_
timestamp 1676037725
transform 1 0 28428 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0534_
timestamp 1676037725
transform 1 0 28520 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0535_
timestamp 1676037725
transform 1 0 27876 0 -1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _0536_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 28612 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_2  _0537_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 31372 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0538_
timestamp 1676037725
transform 1 0 47564 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_2  _0539_
timestamp 1676037725
transform 1 0 47748 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_2  _0540_
timestamp 1676037725
transform 1 0 29716 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0541_
timestamp 1676037725
transform 1 0 16836 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_2  _0542_
timestamp 1676037725
transform 1 0 28244 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__or3_4  _0543_
timestamp 1676037725
transform 1 0 29716 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0544_
timestamp 1676037725
transform 1 0 41308 0 1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_2  _0545_
timestamp 1676037725
transform 1 0 42320 0 1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0546_
timestamp 1676037725
transform 1 0 2024 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0547_
timestamp 1676037725
transform 1 0 30176 0 1 48960
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0548_
timestamp 1676037725
transform 1 0 32108 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0549_
timestamp 1676037725
transform 1 0 30452 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0550_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 31280 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or2_4  _0551_
timestamp 1676037725
transform 1 0 31556 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0552_
timestamp 1676037725
transform 1 0 27600 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0553_
timestamp 1676037725
transform 1 0 2024 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_2  _0554_
timestamp 1676037725
transform 1 0 3312 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _0555_
timestamp 1676037725
transform 1 0 27876 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _0556_
timestamp 1676037725
transform 1 0 31004 0 1 47872
box -38 -48 866 592
use sky130_fd_sc_hd__or3_4  _0557_
timestamp 1676037725
transform 1 0 28980 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_4  _0558_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 48392 0 1 44608
box -38 -48 1326 592
use sky130_fd_sc_hd__a221o_4  _0559_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 47748 0 -1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__a22o_1  _0560_
timestamp 1676037725
transform 1 0 19872 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0561_
timestamp 1676037725
transform 1 0 27968 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0562_
timestamp 1676037725
transform 1 0 2024 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_2  _0563_
timestamp 1676037725
transform 1 0 2300 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__or3_4  _0564_
timestamp 1676037725
transform 1 0 28428 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0565_
timestamp 1676037725
transform 1 0 34868 0 1 47872
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_4  _0566_
timestamp 1676037725
transform 1 0 30268 0 -1 48960
box -38 -48 1602 592
use sky130_fd_sc_hd__a22o_1  _0567_
timestamp 1676037725
transform 1 0 2668 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_4  _0568_
timestamp 1676037725
transform 1 0 3128 0 -1 36992
box -38 -48 1602 592
use sky130_fd_sc_hd__a22o_1  _0569_
timestamp 1676037725
transform 1 0 30452 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__nor4_4  _0570_
timestamp 1676037725
transform 1 0 30176 0 1 35904
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _0571_
timestamp 1676037725
transform 1 0 21252 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _0572_
timestamp 1676037725
transform 1 0 3956 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0573_
timestamp 1676037725
transform 1 0 32660 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0574_
timestamp 1676037725
transform 1 0 35328 0 -1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_2  _0575_
timestamp 1676037725
transform 1 0 36432 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _0576_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 33856 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__nor4b_4  _0577_
timestamp 1676037725
transform 1 0 33120 0 -1 33728
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _0578_
timestamp 1676037725
transform 1 0 21988 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0579_
timestamp 1676037725
transform 1 0 34868 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_4  _0580_
timestamp 1676037725
transform 1 0 32292 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_2  _0581_
timestamp 1676037725
transform 1 0 4692 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0582_
timestamp 1676037725
transform 1 0 32476 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0583_
timestamp 1676037725
transform 1 0 36432 0 1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_2  _0584_
timestamp 1676037725
transform 1 0 36892 0 1 51136
box -38 -48 866 592
use sky130_fd_sc_hd__or4_4  _0585_
timestamp 1676037725
transform 1 0 33764 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0586_
timestamp 1676037725
transform 1 0 32660 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0587_
timestamp 1676037725
transform 1 0 32292 0 -1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0588_
timestamp 1676037725
transform 1 0 33028 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0589_
timestamp 1676037725
transform 1 0 31832 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0590_
timestamp 1676037725
transform 1 0 32292 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__or3_4  _0591_
timestamp 1676037725
transform 1 0 32844 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_4  _0592_
timestamp 1676037725
transform 1 0 41860 0 1 3264
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_2  _0593_
timestamp 1676037725
transform 1 0 7360 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0594_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 22080 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0595_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 22540 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a2111o_2  _0596_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 32200 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__a211oi_4  _0597_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 32936 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _0598_
timestamp 1676037725
transform 1 0 23828 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _0599_
timestamp 1676037725
transform 1 0 9108 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0600_
timestamp 1676037725
transform 1 0 30728 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0601_
timestamp 1676037725
transform 1 0 42596 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0602_
timestamp 1676037725
transform 1 0 40020 0 1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _0603_
timestamp 1676037725
transform 1 0 31188 0 1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0604_
timestamp 1676037725
transform 1 0 48392 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0605_
timestamp 1676037725
transform 1 0 9936 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _0606_
timestamp 1676037725
transform 1 0 41308 0 -1 47872
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _0607_
timestamp 1676037725
transform 1 0 42228 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0608_
timestamp 1676037725
transform 1 0 41492 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0609_
timestamp 1676037725
transform 1 0 42136 0 1 52224
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0610_
timestamp 1676037725
transform 1 0 42780 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_4  _0611_
timestamp 1676037725
transform 1 0 42596 0 -1 34816
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_2  _0612_
timestamp 1676037725
transform 1 0 49036 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a311o_1  _0613_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 26404 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _0614_
timestamp 1676037725
transform 1 0 43240 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _0615_
timestamp 1676037725
transform 1 0 26312 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_4  _0616_
timestamp 1676037725
transform 1 0 42596 0 -1 50048
box -38 -48 1326 592
use sky130_fd_sc_hd__a221o_2  _0617_
timestamp 1676037725
transform 1 0 43516 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_4  _0618_
timestamp 1676037725
transform 1 0 43332 0 -1 18496
box -38 -48 1326 592
use sky130_fd_sc_hd__a31o_2  _0619_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25024 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0620_
timestamp 1676037725
transform 1 0 47840 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0621_
timestamp 1676037725
transform 1 0 46000 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _0622_
timestamp 1676037725
transform 1 0 48208 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_4  _0623_
timestamp 1676037725
transform 1 0 47564 0 -1 51136
box -38 -48 1326 592
use sky130_fd_sc_hd__a221o_2  _0624_
timestamp 1676037725
transform 1 0 46920 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_4  _0625_
timestamp 1676037725
transform 1 0 47380 0 1 17408
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_2  _0626_
timestamp 1676037725
transform 1 0 46828 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _0627_
timestamp 1676037725
transform 1 0 47012 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_4  _0628_
timestamp 1676037725
transform 1 0 47196 0 1 33728
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_4  _0629_
timestamp 1676037725
transform 1 0 47748 0 -1 52224
box -38 -48 1326 592
use sky130_fd_sc_hd__a221o_2  _0630_
timestamp 1676037725
transform 1 0 48024 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_4  _0631_
timestamp 1676037725
transform 1 0 47748 0 -1 18496
box -38 -48 1326 592
use sky130_fd_sc_hd__a31o_2  _0632_
timestamp 1676037725
transform 1 0 25944 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0633_
timestamp 1676037725
transform 1 0 48944 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0634_
timestamp 1676037725
transform 1 0 47104 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _0635_
timestamp 1676037725
transform 1 0 47748 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_4  _0636_
timestamp 1676037725
transform 1 0 47380 0 1 52224
box -38 -48 1326 592
use sky130_fd_sc_hd__a221o_2  _0637_
timestamp 1676037725
transform 1 0 47932 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_4  _0638_
timestamp 1676037725
transform 1 0 47932 0 1 18496
box -38 -48 1326 592
use sky130_fd_sc_hd__a221o_1  _0639_
timestamp 1676037725
transform 1 0 49404 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_4  _0640_
timestamp 1676037725
transform 1 0 48116 0 1 3264
box -38 -48 1326 592
use sky130_fd_sc_hd__a211o_4  _0641_
timestamp 1676037725
transform 1 0 48300 0 1 50048
box -38 -48 1326 592
use sky130_fd_sc_hd__a221o_4  _0642_
timestamp 1676037725
transform 1 0 47932 0 1 51136
box -38 -48 1602 592
use sky130_fd_sc_hd__a22o_1  _0643_
timestamp 1676037725
transform 1 0 48208 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_4  _0644_
timestamp 1676037725
transform 1 0 48484 0 -1 11968
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_4  _0645_
timestamp 1676037725
transform 1 0 47748 0 -1 53312
box -38 -48 1326 592
use sky130_fd_sc_hd__a221o_2  _0646_
timestamp 1676037725
transform 1 0 47840 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_4  _0647_
timestamp 1676037725
transform 1 0 48116 0 -1 17408
box -38 -48 1326 592
use sky130_fd_sc_hd__a211o_4  _0648_
timestamp 1676037725
transform 1 0 23644 0 -1 20672
box -38 -48 1326 592
use sky130_fd_sc_hd__mux2_2  _0649_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25392 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _0650_
timestamp 1676037725
transform 1 0 24932 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0651_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11684 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _0652_
timestamp 1676037725
transform 1 0 22816 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0653_
timestamp 1676037725
transform 1 0 10672 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0654_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9660 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0655_
timestamp 1676037725
transform 1 0 9660 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0656_
timestamp 1676037725
transform 1 0 9752 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0657_
timestamp 1676037725
transform 1 0 11684 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _0658_
timestamp 1676037725
transform 1 0 26036 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0659_
timestamp 1676037725
transform 1 0 10580 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0660_
timestamp 1676037725
transform 1 0 10396 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0661_
timestamp 1676037725
transform 1 0 17388 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0662_
timestamp 1676037725
transform 1 0 17756 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0663_
timestamp 1676037725
transform 1 0 10672 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0664_
timestamp 1676037725
transform 1 0 10948 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0665_
timestamp 1676037725
transform 1 0 10028 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0666_
timestamp 1676037725
transform 1 0 10580 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0667_
timestamp 1676037725
transform 1 0 12972 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0668_
timestamp 1676037725
transform 1 0 12144 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0669_
timestamp 1676037725
transform 1 0 11776 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0670_
timestamp 1676037725
transform 1 0 12236 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0671_
timestamp 1676037725
transform 1 0 12052 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0672_
timestamp 1676037725
transform 1 0 12328 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0673_
timestamp 1676037725
transform 1 0 13340 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0674_
timestamp 1676037725
transform 1 0 12328 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0675_
timestamp 1676037725
transform 1 0 13340 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0676_
timestamp 1676037725
transform 1 0 14260 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0677_
timestamp 1676037725
transform 1 0 16744 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0678_
timestamp 1676037725
transform 1 0 17664 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0679_
timestamp 1676037725
transform 1 0 12420 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0680_
timestamp 1676037725
transform 1 0 13064 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0681_
timestamp 1676037725
transform 1 0 13064 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0682_
timestamp 1676037725
transform 1 0 13156 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0683_
timestamp 1676037725
transform 1 0 20700 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_4  _0684_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 35144 0 -1 6528
box -38 -48 1326 592
use sky130_fd_sc_hd__and2b_1  _0685_
timestamp 1676037725
transform 1 0 20424 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_4  _0686_
timestamp 1676037725
transform 1 0 37168 0 1 7616
box -38 -48 1326 592
use sky130_fd_sc_hd__and2b_1  _0687_
timestamp 1676037725
transform 1 0 20056 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_4  _0688_
timestamp 1676037725
transform 1 0 35512 0 1 7616
box -38 -48 1326 592
use sky130_fd_sc_hd__and2b_1  _0689_
timestamp 1676037725
transform 1 0 19504 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_4  _0690_
timestamp 1676037725
transform 1 0 35512 0 1 5440
box -38 -48 1326 592
use sky130_fd_sc_hd__and2b_2  _0691_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19964 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_4  _0692_
timestamp 1676037725
transform 1 0 35512 0 -1 8704
box -38 -48 1326 592
use sky130_fd_sc_hd__and2b_1  _0693_
timestamp 1676037725
transform 1 0 15824 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0694_
timestamp 1676037725
transform 1 0 14536 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_2  _0695_
timestamp 1676037725
transform 1 0 20332 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_4  _0696_
timestamp 1676037725
transform 1 0 37444 0 -1 7616
box -38 -48 1326 592
use sky130_fd_sc_hd__and2b_1  _0697_
timestamp 1676037725
transform 1 0 15088 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0698_
timestamp 1676037725
transform 1 0 15088 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_2  _0699_
timestamp 1676037725
transform 1 0 20240 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_4  _0700_
timestamp 1676037725
transform 1 0 35512 0 1 8704
box -38 -48 1326 592
use sky130_fd_sc_hd__and2b_2  _0701_
timestamp 1676037725
transform 1 0 20056 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_4  _0702_
timestamp 1676037725
transform 1 0 35512 0 -1 5440
box -38 -48 1326 592
use sky130_fd_sc_hd__and2b_1  _0703_
timestamp 1676037725
transform 1 0 15732 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0704_
timestamp 1676037725
transform 1 0 15548 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0705_
timestamp 1676037725
transform 1 0 19412 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _0706_
timestamp 1676037725
transform 1 0 20056 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _0707_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 57408 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _0708_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 57132 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and3_4  _0709_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 44804 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0710_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 37444 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0711_
timestamp 1676037725
transform 1 0 34316 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0712_
timestamp 1676037725
transform 1 0 43240 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0713_
timestamp 1676037725
transform 1 0 43056 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0714_
timestamp 1676037725
transform 1 0 38548 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0715_
timestamp 1676037725
transform 1 0 39100 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0716_
timestamp 1676037725
transform 1 0 35420 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0717_
timestamp 1676037725
transform 1 0 34684 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0718_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 54740 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0719_
timestamp 1676037725
transform 1 0 33212 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0720_
timestamp 1676037725
transform 1 0 27876 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0721_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 45080 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0722_
timestamp 1676037725
transform 1 0 44436 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0723_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 45172 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_2  _0724_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 46000 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0725_
timestamp 1676037725
transform 1 0 27692 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0726_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27692 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0727_
timestamp 1676037725
transform 1 0 32568 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0728_
timestamp 1676037725
transform 1 0 32476 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0729_
timestamp 1676037725
transform 1 0 31372 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0730_
timestamp 1676037725
transform 1 0 31648 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0731_
timestamp 1676037725
transform 1 0 27048 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0732_
timestamp 1676037725
transform 1 0 28336 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0733_
timestamp 1676037725
transform 1 0 30268 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0734_
timestamp 1676037725
transform 1 0 29716 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0735_
timestamp 1676037725
transform 1 0 32384 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0736_
timestamp 1676037725
transform 1 0 33396 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0737_
timestamp 1676037725
transform 1 0 28796 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0738_
timestamp 1676037725
transform 1 0 27876 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0739_
timestamp 1676037725
transform 1 0 31372 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0740_
timestamp 1676037725
transform 1 0 29716 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0741_
timestamp 1676037725
transform 1 0 28244 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0742_
timestamp 1676037725
transform 1 0 29072 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0743_
timestamp 1676037725
transform 1 0 33304 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0744_
timestamp 1676037725
transform 1 0 33672 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0745_
timestamp 1676037725
transform 1 0 38548 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0746_
timestamp 1676037725
transform 1 0 37536 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0747_
timestamp 1676037725
transform 1 0 41676 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0748_
timestamp 1676037725
transform 1 0 42596 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0749_
timestamp 1676037725
transform 1 0 43148 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0750_
timestamp 1676037725
transform 1 0 43976 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0751_
timestamp 1676037725
transform 1 0 43792 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0752_
timestamp 1676037725
transform 1 0 43976 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0753_
timestamp 1676037725
transform 1 0 42596 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0754_
timestamp 1676037725
transform 1 0 38364 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0755_
timestamp 1676037725
transform 1 0 40020 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0756_
timestamp 1676037725
transform 1 0 38640 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0757_
timestamp 1676037725
transform 1 0 34684 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0758_
timestamp 1676037725
transform 1 0 35420 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0759_
timestamp 1676037725
transform 1 0 37904 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0760_
timestamp 1676037725
transform 1 0 38732 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0761_
timestamp 1676037725
transform 1 0 44528 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0762_
timestamp 1676037725
transform 1 0 45172 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0763_
timestamp 1676037725
transform 1 0 42596 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0764_
timestamp 1676037725
transform 1 0 42872 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0765_
timestamp 1676037725
transform 1 0 40940 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0766_
timestamp 1676037725
transform 1 0 41308 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0767_
timestamp 1676037725
transform 1 0 41308 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0768_
timestamp 1676037725
transform 1 0 41584 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0769_
timestamp 1676037725
transform 1 0 44160 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0770_
timestamp 1676037725
transform 1 0 43608 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0771_
timestamp 1676037725
transform 1 0 41676 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0772_
timestamp 1676037725
transform 1 0 38824 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0773_
timestamp 1676037725
transform 1 0 56580 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0774_
timestamp 1676037725
transform 1 0 47656 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0775_
timestamp 1676037725
transform 1 0 25208 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0776_
timestamp 1676037725
transform 1 0 29808 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0777_
timestamp 1676037725
transform 1 0 27140 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0778_
timestamp 1676037725
transform 1 0 27140 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0779_
timestamp 1676037725
transform 1 0 24932 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0780_
timestamp 1676037725
transform 1 0 24840 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0781_
timestamp 1676037725
transform 1 0 25024 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0782_
timestamp 1676037725
transform 1 0 25300 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0783_
timestamp 1676037725
transform 1 0 27048 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0784_
timestamp 1676037725
transform 1 0 26220 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0785_
timestamp 1676037725
transform 1 0 38180 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0786_
timestamp 1676037725
transform 1 0 41492 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0787_
timestamp 1676037725
transform 1 0 42688 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0788_
timestamp 1676037725
transform 1 0 43516 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0789_
timestamp 1676037725
transform 1 0 37444 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0790_
timestamp 1676037725
transform 1 0 37444 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0791_
timestamp 1676037725
transform 1 0 35880 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0792_
timestamp 1676037725
transform 1 0 37444 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0793_
timestamp 1676037725
transform 1 0 45172 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0794_
timestamp 1676037725
transform 1 0 42596 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0795_
timestamp 1676037725
transform 1 0 40664 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0796_
timestamp 1676037725
transform 1 0 41216 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0797_
timestamp 1676037725
transform 1 0 42964 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0798_
timestamp 1676037725
transform 1 0 40020 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0799_
timestamp 1676037725
transform 1 0 46368 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0800_
timestamp 1676037725
transform 1 0 45356 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0801_
timestamp 1676037725
transform 1 0 46368 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0802_
timestamp 1676037725
transform 1 0 40480 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0803_
timestamp 1676037725
transform 1 0 22816 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0804_
timestamp 1676037725
transform 1 0 22724 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0805_
timestamp 1676037725
transform 1 0 22172 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0806_
timestamp 1676037725
transform 1 0 22264 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0807_
timestamp 1676037725
transform 1 0 23460 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0808_
timestamp 1676037725
transform 1 0 23276 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0809_
timestamp 1676037725
transform 1 0 23276 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0810_
timestamp 1676037725
transform 1 0 22908 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _0811_
timestamp 1676037725
transform 1 0 45172 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0812_
timestamp 1676037725
transform 1 0 46000 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0813_
timestamp 1676037725
transform 1 0 55108 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0814_
timestamp 1676037725
transform 1 0 28980 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0815_
timestamp 1676037725
transform 1 0 30912 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0816_
timestamp 1676037725
transform 1 0 30360 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0817_
timestamp 1676037725
transform 1 0 39744 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_2  _0818_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 38640 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0819_
timestamp 1676037725
transform 1 0 58052 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0820_
timestamp 1676037725
transform 1 0 56120 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0821_
timestamp 1676037725
transform 1 0 32292 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0822_
timestamp 1676037725
transform 1 0 30360 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0823_
timestamp 1676037725
transform 1 0 40388 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_2  _0824_
timestamp 1676037725
transform 1 0 40388 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0825_
timestamp 1676037725
transform 1 0 55568 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0826_
timestamp 1676037725
transform 1 0 56948 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0827_
timestamp 1676037725
transform 1 0 29992 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0828_
timestamp 1676037725
transform 1 0 30912 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0829_
timestamp 1676037725
transform 1 0 39100 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_2  _0830_
timestamp 1676037725
transform 1 0 39100 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0831_
timestamp 1676037725
transform 1 0 56304 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_2  _0832_
timestamp 1676037725
transform 1 0 30176 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _0833_
timestamp 1676037725
transform 1 0 44804 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0834_
timestamp 1676037725
transform 1 0 46000 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0835_
timestamp 1676037725
transform 1 0 47748 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0836_
timestamp 1676037725
transform 1 0 56396 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o31ai_4  _0837_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 29992 0 -1 30464
box -38 -48 1602 592
use sky130_fd_sc_hd__o221a_1  _0838_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 31004 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _0839_
timestamp 1676037725
transform 1 0 38824 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0840_
timestamp 1676037725
transform 1 0 56028 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0841_
timestamp 1676037725
transform 1 0 58052 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _0842_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 32292 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a221oi_4  _0843_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 31096 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__a211o_2  _0844_
timestamp 1676037725
transform 1 0 37996 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0845_
timestamp 1676037725
transform 1 0 56304 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a22oi_4  _0846_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 30360 0 1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__nor2_4  _0847_
timestamp 1676037725
transform 1 0 54188 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _0848_
timestamp 1676037725
transform 1 0 51520 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _0849_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 50324 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0850_
timestamp 1676037725
transform 1 0 49404 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _0851_
timestamp 1676037725
transform 1 0 30360 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0852_
timestamp 1676037725
transform 1 0 55568 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0853_
timestamp 1676037725
transform 1 0 56304 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0854_
timestamp 1676037725
transform 1 0 32476 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _0855_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 32292 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _0856_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 50232 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0857_
timestamp 1676037725
transform 1 0 49588 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0858_
timestamp 1676037725
transform 1 0 33028 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _0859_
timestamp 1676037725
transform 1 0 50416 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0860_
timestamp 1676037725
transform 1 0 50140 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _0861_
timestamp 1676037725
transform 1 0 33580 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _0862_
timestamp 1676037725
transform 1 0 34868 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0863_
timestamp 1676037725
transform 1 0 55936 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0864_
timestamp 1676037725
transform 1 0 56028 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a22oi_4  _0865_
timestamp 1676037725
transform 1 0 35420 0 -1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__o2bb2a_1  _0866_
timestamp 1676037725
transform 1 0 51704 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0867_
timestamp 1676037725
transform 1 0 51888 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _0868_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 33396 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0869_
timestamp 1676037725
transform 1 0 47104 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0870_
timestamp 1676037725
transform 1 0 47472 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0871_
timestamp 1676037725
transform 1 0 47748 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0872_
timestamp 1676037725
transform 1 0 29716 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0873_
timestamp 1676037725
transform 1 0 46920 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0874_
timestamp 1676037725
transform 1 0 46552 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0875_
timestamp 1676037725
transform 1 0 48944 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _0876_
timestamp 1676037725
transform 1 0 40020 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _0877_
timestamp 1676037725
transform 1 0 40940 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _0878_
timestamp 1676037725
transform 1 0 52900 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0879_
timestamp 1676037725
transform 1 0 51980 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_4  _0880_
timestamp 1676037725
transform 1 0 41216 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__o2bb2a_1  _0881_
timestamp 1676037725
transform 1 0 53820 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0882_
timestamp 1676037725
transform 1 0 52164 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0883_
timestamp 1676037725
transform 1 0 36616 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0884_
timestamp 1676037725
transform 1 0 48208 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0885_
timestamp 1676037725
transform 1 0 48484 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0886_
timestamp 1676037725
transform 1 0 43148 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__a22oi_1  _0887_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 55660 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0888_
timestamp 1676037725
transform 1 0 55752 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0889_
timestamp 1676037725
transform 1 0 47104 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0890_
timestamp 1676037725
transform 1 0 51060 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0891_
timestamp 1676037725
transform 1 0 51520 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0892_
timestamp 1676037725
transform 1 0 44988 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__a22oi_1  _0893_
timestamp 1676037725
transform 1 0 56672 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0894_
timestamp 1676037725
transform 1 0 56212 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0895_
timestamp 1676037725
transform 1 0 45540 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0896_
timestamp 1676037725
transform 1 0 53544 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0897_
timestamp 1676037725
transform 1 0 52900 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0898_
timestamp 1676037725
transform 1 0 49036 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_2  _0899_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 47656 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__o2bb2a_1  _0900_
timestamp 1676037725
transform 1 0 50324 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0901_
timestamp 1676037725
transform 1 0 50140 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0902_
timestamp 1676037725
transform 1 0 46184 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0903_
timestamp 1676037725
transform 1 0 57684 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0904_
timestamp 1676037725
transform 1 0 56120 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _0905_
timestamp 1676037725
transform 1 0 47748 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _0906_
timestamp 1676037725
transform 1 0 48944 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0907_
timestamp 1676037725
transform 1 0 48760 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0908_
timestamp 1676037725
transform 1 0 55752 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0909_
timestamp 1676037725
transform 1 0 55292 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0910_
timestamp 1676037725
transform 1 0 55660 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0911_
timestamp 1676037725
transform 1 0 56212 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0912_
timestamp 1676037725
transform 1 0 54648 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _0913_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 48392 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0914_
timestamp 1676037725
transform 1 0 53452 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _0915_
timestamp 1676037725
transform 1 0 55844 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0916_
timestamp 1676037725
transform 1 0 55844 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0917_
timestamp 1676037725
transform 1 0 21252 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0918_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20608 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0919_
timestamp 1676037725
transform 1 0 19780 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_2  _0920_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21988 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _0921_
timestamp 1676037725
transform 1 0 21160 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0922_
timestamp 1676037725
transform 1 0 19964 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0923_
timestamp 1676037725
transform 1 0 17848 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0924_
timestamp 1676037725
transform 1 0 18216 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0925_
timestamp 1676037725
transform 1 0 17572 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0926_
timestamp 1676037725
transform 1 0 17204 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and4_4  _0927_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 22264 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _0928_
timestamp 1676037725
transform 1 0 22080 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0929_
timestamp 1676037725
transform 1 0 23092 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _0930_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 28336 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0931_
timestamp 1676037725
transform 1 0 30728 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0932_
timestamp 1676037725
transform 1 0 30544 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0933_
timestamp 1676037725
transform 1 0 27968 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0934_
timestamp 1676037725
transform 1 0 30176 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0935_
timestamp 1676037725
transform 1 0 29716 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0936_
timestamp 1676037725
transform 1 0 32292 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0937_
timestamp 1676037725
transform 1 0 31372 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0938_
timestamp 1676037725
transform 1 0 31372 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0939_
timestamp 1676037725
transform 1 0 32292 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and4_2  _0940_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 31648 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0941_
timestamp 1676037725
transform 1 0 34500 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0942_
timestamp 1676037725
transform 1 0 31464 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _0943_
timestamp 1676037725
transform 1 0 35696 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0944_
timestamp 1676037725
transform 1 0 36708 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0945_
timestamp 1676037725
transform 1 0 35696 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0946_
timestamp 1676037725
transform 1 0 35696 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0947_
timestamp 1676037725
transform 1 0 36340 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0948_
timestamp 1676037725
transform 1 0 38916 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0949_
timestamp 1676037725
transform 1 0 37444 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0950_
timestamp 1676037725
transform 1 0 36524 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0951_
timestamp 1676037725
transform 1 0 37444 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0952_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 35788 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _0953_
timestamp 1676037725
transform 1 0 36340 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__and4_2  _0954_
timestamp 1676037725
transform 1 0 35236 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0955_
timestamp 1676037725
transform 1 0 37444 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0956_
timestamp 1676037725
transform 1 0 34132 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0957_
timestamp 1676037725
transform 1 0 27876 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0958_
timestamp 1676037725
transform 1 0 27140 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0959_
timestamp 1676037725
transform 1 0 26036 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and4_2  _0960_
timestamp 1676037725
transform 1 0 28520 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0961_
timestamp 1676037725
transform 1 0 28428 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0962_
timestamp 1676037725
transform 1 0 27784 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0963_
timestamp 1676037725
transform 1 0 30452 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0964_
timestamp 1676037725
transform 1 0 28704 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0965_
timestamp 1676037725
transform 1 0 29716 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0966_
timestamp 1676037725
transform 1 0 31004 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0967_
timestamp 1676037725
transform 1 0 30912 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0968_
timestamp 1676037725
transform 1 0 31004 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0969_
timestamp 1676037725
transform 1 0 32568 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0970_
timestamp 1676037725
transform 1 0 40020 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0971_
timestamp 1676037725
transform 1 0 39100 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0972_
timestamp 1676037725
transform 1 0 27876 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0973_
timestamp 1676037725
transform 1 0 36616 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0974_
timestamp 1676037725
transform 1 0 35788 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  _0975_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 35604 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _0976_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 42872 0 -1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0977_
timestamp 1676037725
transform 1 0 38180 0 -1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _0978_
timestamp 1676037725
transform 1 0 35144 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0979_
timestamp 1676037725
transform 1 0 27140 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0980_
timestamp 1676037725
transform 1 0 55568 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _0981_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27784 0 -1 5440
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _0982_
timestamp 1676037725
transform 1 0 32292 0 -1 5440
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _0983_
timestamp 1676037725
transform 1 0 32292 0 -1 4352
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _0984_
timestamp 1676037725
transform 1 0 27508 0 1 6528
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _0985_
timestamp 1676037725
transform 1 0 29992 0 -1 8704
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _0986_
timestamp 1676037725
transform 1 0 32660 0 -1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0987_
timestamp 1676037725
transform 1 0 28980 0 -1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _0988_
timestamp 1676037725
transform 1 0 29532 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0989_
timestamp 1676037725
transform 1 0 29716 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0990_
timestamp 1676037725
transform 1 0 33948 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0991_
timestamp 1676037725
transform 1 0 38088 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _0992_
timestamp 1676037725
transform 1 0 42228 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0993_
timestamp 1676037725
transform 1 0 45172 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _0994_
timestamp 1676037725
transform 1 0 44620 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0995_
timestamp 1676037725
transform 1 0 38180 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _0996_
timestamp 1676037725
transform 1 0 39744 0 -1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _0997_
timestamp 1676037725
transform 1 0 35512 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _0998_
timestamp 1676037725
transform 1 0 39100 0 -1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0999_
timestamp 1676037725
transform 1 0 45172 0 1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1000_
timestamp 1676037725
transform 1 0 43240 0 -1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1001_
timestamp 1676037725
transform 1 0 42596 0 -1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1002_
timestamp 1676037725
transform 1 0 42044 0 1 21760
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _1003_
timestamp 1676037725
transform 1 0 44068 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1004_
timestamp 1676037725
transform 1 0 38456 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1005_
timestamp 1676037725
transform 1 0 56856 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1006_
timestamp 1676037725
transform 1 0 24380 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1007_
timestamp 1676037725
transform 1 0 29164 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1008_
timestamp 1676037725
transform 1 0 25852 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1009_
timestamp 1676037725
transform 1 0 25392 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1010_
timestamp 1676037725
transform 1 0 24104 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1011_
timestamp 1676037725
transform 1 0 24104 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1012_
timestamp 1676037725
transform 1 0 24196 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1013_
timestamp 1676037725
transform 1 0 24564 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1014_
timestamp 1676037725
transform 1 0 25208 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1015_
timestamp 1676037725
transform 1 0 25208 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1016_
timestamp 1676037725
transform 1 0 37628 0 -1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1017_
timestamp 1676037725
transform 1 0 40572 0 -1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1018_
timestamp 1676037725
transform 1 0 41676 0 1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1019_
timestamp 1676037725
transform 1 0 42964 0 1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1020_
timestamp 1676037725
transform 1 0 36340 0 1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1021_
timestamp 1676037725
transform 1 0 36156 0 1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1022_
timestamp 1676037725
transform 1 0 34040 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1023_
timestamp 1676037725
transform 1 0 35512 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1024_
timestamp 1676037725
transform 1 0 44068 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1025_
timestamp 1676037725
transform 1 0 42596 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1026_
timestamp 1676037725
transform 1 0 40020 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1027_
timestamp 1676037725
transform 1 0 40664 0 1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1028_
timestamp 1676037725
transform 1 0 42596 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1029_
timestamp 1676037725
transform 1 0 38640 0 -1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1030_
timestamp 1676037725
transform 1 0 44528 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1031_
timestamp 1676037725
transform 1 0 45172 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1032_
timestamp 1676037725
transform 1 0 45540 0 1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1033_
timestamp 1676037725
transform 1 0 39928 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1034_
timestamp 1676037725
transform 1 0 23920 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1035_
timestamp 1676037725
transform 1 0 24564 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1036_
timestamp 1676037725
transform 1 0 24564 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1037_
timestamp 1676037725
transform 1 0 24104 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1038_
timestamp 1676037725
transform 1 0 56764 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1039_
timestamp 1676037725
transform 1 0 55752 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1040_
timestamp 1676037725
transform 1 0 56672 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1041_
timestamp 1676037725
transform 1 0 47472 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1042_
timestamp 1676037725
transform 1 0 56764 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1043_
timestamp 1676037725
transform 1 0 56764 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1044_
timestamp 1676037725
transform 1 0 50324 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1045_
timestamp 1676037725
transform 1 0 56764 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1046_
timestamp 1676037725
transform 1 0 50324 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1047_
timestamp 1676037725
transform 1 0 50048 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1048_
timestamp 1676037725
transform 1 0 56856 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1049_
timestamp 1676037725
transform 1 0 51796 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1050_
timestamp 1676037725
transform 1 0 47748 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1051_
timestamp 1676037725
transform 1 0 48300 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1052_
timestamp 1676037725
transform 1 0 51980 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1053_
timestamp 1676037725
transform 1 0 52900 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1054_
timestamp 1676037725
transform 1 0 48484 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1055_
timestamp 1676037725
transform 1 0 55752 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1056_
timestamp 1676037725
transform 1 0 51704 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1057_
timestamp 1676037725
transform 1 0 56856 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1058_
timestamp 1676037725
transform 1 0 52900 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1059_
timestamp 1676037725
transform 1 0 50048 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1060_
timestamp 1676037725
transform 1 0 56856 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1061_
timestamp 1676037725
transform 1 0 48392 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1062_
timestamp 1676037725
transform 1 0 55844 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1063_
timestamp 1676037725
transform 1 0 56764 0 1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1064_
timestamp 1676037725
transform 1 0 54188 0 -1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1065_
timestamp 1676037725
transform 1 0 56120 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _1066_
timestamp 1676037725
transform 1 0 21620 0 1 18496
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1067_
timestamp 1676037725
transform 1 0 20056 0 1 16320
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1068_
timestamp 1676037725
transform 1 0 19596 0 -1 16320
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1069_
timestamp 1676037725
transform 1 0 17020 0 -1 16320
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1070_
timestamp 1676037725
transform 1 0 17204 0 1 16320
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1071_
timestamp 1676037725
transform 1 0 22172 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1072_
timestamp 1676037725
transform 1 0 28704 0 -1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1073_
timestamp 1676037725
transform 1 0 28704 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1074_
timestamp 1676037725
transform 1 0 29716 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1075_
timestamp 1676037725
transform 1 0 31832 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1076_
timestamp 1676037725
transform 1 0 32660 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1077_
timestamp 1676037725
transform 1 0 32844 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1078_
timestamp 1676037725
transform 1 0 33488 0 -1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1079_
timestamp 1676037725
transform 1 0 32936 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1080_
timestamp 1676037725
transform 1 0 33212 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1081_
timestamp 1676037725
transform 1 0 33304 0 -1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1082_
timestamp 1676037725
transform 1 0 34868 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1083_
timestamp 1676037725
transform 1 0 26312 0 1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1084_
timestamp 1676037725
transform 1 0 25944 0 1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1085_
timestamp 1676037725
transform 1 0 27876 0 -1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1086_
timestamp 1676037725
transform 1 0 29716 0 1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1087_
timestamp 1676037725
transform 1 0 29992 0 -1 20672
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _1088_
timestamp 1676037725
transform 1 0 31648 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1089_
timestamp 1676037725
transform 1 0 33028 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1090_
timestamp 1676037725
transform 1 0 39100 0 -1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1091_
timestamp 1676037725
transform 1 0 27140 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1092_
timestamp 1676037725
transform 1 0 36248 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_2  _1113_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 28888 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1114_
timestamp 1676037725
transform 1 0 30912 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1115_
timestamp 1676037725
transform 1 0 32752 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1116_
timestamp 1676037725
transform 1 0 33488 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1117_
timestamp 1676037725
transform 1 0 36524 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1118_
timestamp 1676037725
transform 1 0 40020 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1119_
timestamp 1676037725
transform 1 0 34500 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1120_
timestamp 1676037725
transform 1 0 40756 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1121_
timestamp 1676037725
transform 1 0 34040 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1122_
timestamp 1676037725
transform 1 0 38088 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1123_
timestamp 1676037725
transform 1 0 35052 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1124_
timestamp 1676037725
transform 1 0 40940 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1125_
timestamp 1676037725
transform 1 0 40388 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1126_
timestamp 1676037725
transform 1 0 38364 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 41768 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_wb_clk_i
timestamp 1676037725
transform 1 0 28612 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_wb_clk_i
timestamp 1676037725
transform 1 0 33764 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_wb_clk_i
timestamp 1676037725
transform 1 0 31188 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_wb_clk_i
timestamp 1676037725
transform 1 0 33764 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_wb_clk_i
timestamp 1676037725
transform 1 0 46828 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_wb_clk_i
timestamp 1676037725
transform 1 0 49404 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_wb_clk_i
timestamp 1676037725
transform 1 0 44160 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_wb_clk_i
timestamp 1676037725
transform 1 0 49404 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_4  fanout400 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 55844 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout401 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 44160 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout402
timestamp 1676037725
transform 1 0 43792 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout403
timestamp 1676037725
transform 1 0 50692 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout404
timestamp 1676037725
transform 1 0 50784 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout405
timestamp 1676037725
transform 1 0 51612 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout406
timestamp 1676037725
transform 1 0 46460 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout407 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 36248 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout408
timestamp 1676037725
transform 1 0 46368 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  fanout409 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 42780 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout410
timestamp 1676037725
transform 1 0 45908 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout411
timestamp 1676037725
transform 1 0 45172 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout412
timestamp 1676037725
transform 1 0 46092 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout413
timestamp 1676037725
transform 1 0 45172 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  fanout414 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 44712 0 -1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_16  fanout415
timestamp 1676037725
transform 1 0 29716 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_4  fanout416
timestamp 1676037725
transform 1 0 33856 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout417
timestamp 1676037725
transform 1 0 37444 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout419
timestamp 1676037725
transform 1 0 27784 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout420
timestamp 1676037725
transform 1 0 42136 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout421
timestamp 1676037725
transform 1 0 27140 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout422
timestamp 1676037725
transform 1 0 28060 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout423
timestamp 1676037725
transform 1 0 39284 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout424
timestamp 1676037725
transform 1 0 24196 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout425
timestamp 1676037725
transform 1 0 21988 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout426
timestamp 1676037725
transform 1 0 37444 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  fanout427
timestamp 1676037725
transform 1 0 38548 0 1 3264
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  fanout428
timestamp 1676037725
transform 1 0 37628 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout429
timestamp 1676037725
transform 1 0 29532 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout430
timestamp 1676037725
transform 1 0 29716 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  fanout431 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  fanout432
timestamp 1676037725
transform 1 0 38548 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout433
timestamp 1676037725
transform 1 0 28980 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout434
timestamp 1676037725
transform 1 0 27876 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_16  fanout435
timestamp 1676037725
transform 1 0 19688 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_12  fanout436 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 29440 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_8  fanout437
timestamp 1676037725
transform 1 0 23000 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_16  fanout438
timestamp 1676037725
transform 1 0 28704 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_4  fanout439
timestamp 1676037725
transform 1 0 2116 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_16  fanout440
timestamp 1676037725
transform 1 0 22356 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_6  fanout441
timestamp 1676037725
transform 1 0 41308 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout442
timestamp 1676037725
transform 1 0 33028 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout443
timestamp 1676037725
transform 1 0 13156 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout444
timestamp 1676037725
transform 1 0 11592 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout445
timestamp 1676037725
transform 1 0 15272 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout446
timestamp 1676037725
transform 1 0 12604 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout447
timestamp 1676037725
transform 1 0 23368 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout448
timestamp 1676037725
transform 1 0 23368 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout449
timestamp 1676037725
transform 1 0 37444 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout450
timestamp 1676037725
transform 1 0 37444 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout451
timestamp 1676037725
transform 1 0 27140 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout452
timestamp 1676037725
transform 1 0 24380 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout453
timestamp 1676037725
transform 1 0 24564 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout454
timestamp 1676037725
transform 1 0 23644 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  fanout455
timestamp 1676037725
transform 1 0 25300 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  fanout456
timestamp 1676037725
transform 1 0 23276 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout457
timestamp 1676037725
transform 1 0 23000 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout458
timestamp 1676037725
transform 1 0 23828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout459
timestamp 1676037725
transform 1 0 24564 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout460
timestamp 1676037725
transform 1 0 25668 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout461
timestamp 1676037725
transform 1 0 22724 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout462
timestamp 1676037725
transform 1 0 25116 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  fanout463
timestamp 1676037725
transform 1 0 23736 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout464
timestamp 1676037725
transform 1 0 23276 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  fanout465
timestamp 1676037725
transform 1 0 34868 0 1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_2  fanout466
timestamp 1676037725
transform 1 0 40204 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout467
timestamp 1676037725
transform 1 0 37168 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout468
timestamp 1676037725
transform 1 0 44896 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout469
timestamp 1676037725
transform 1 0 46092 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  fanout470
timestamp 1676037725
transform 1 0 43056 0 1 5440
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_6  fanout471
timestamp 1676037725
transform 1 0 32292 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  fanout472
timestamp 1676037725
transform 1 0 46000 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  fanout473
timestamp 1676037725
transform 1 0 44068 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout474
timestamp 1676037725
transform 1 0 31464 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout475
timestamp 1676037725
transform 1 0 56580 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout476
timestamp 1676037725
transform 1 0 56120 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout477
timestamp 1676037725
transform 1 0 55936 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout478
timestamp 1676037725
transform 1 0 58052 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  fanout479
timestamp 1676037725
transform 1 0 55936 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  hold1
timestamp 1676037725
transform 1 0 41400 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold2
timestamp 1676037725
transform 1 0 37444 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold3
timestamp 1676037725
transform 1 0 38180 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold4
timestamp 1676037725
transform 1 0 25208 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold5
timestamp 1676037725
transform 1 0 35880 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold6
timestamp 1676037725
transform 1 0 29716 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold7
timestamp 1676037725
transform 1 0 35236 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold8
timestamp 1676037725
transform 1 0 27600 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold9
timestamp 1676037725
transform 1 0 28888 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold10
timestamp 1676037725
transform 1 0 28704 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold11
timestamp 1676037725
transform 1 0 37812 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold12
timestamp 1676037725
transform 1 0 30268 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold13
timestamp 1676037725
transform 1 0 27140 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold14
timestamp 1676037725
transform 1 0 21988 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold15
timestamp 1676037725
transform 1 0 25116 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold16
timestamp 1676037725
transform 1 0 21160 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold17
timestamp 1676037725
transform 1 0 40020 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold18
timestamp 1676037725
transform 1 0 37444 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold19
timestamp 1676037725
transform 1 0 33212 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold20
timestamp 1676037725
transform 1 0 24564 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold21
timestamp 1676037725
transform 1 0 16468 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold22
timestamp 1676037725
transform 1 0 32292 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold23
timestamp 1676037725
transform 1 0 30452 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold24
timestamp 1676037725
transform 1 0 29900 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold25
timestamp 1676037725
transform 1 0 40848 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold26
timestamp 1676037725
transform 1 0 40020 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold27
timestamp 1676037725
transform 1 0 34040 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold28
timestamp 1676037725
transform 1 0 37444 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold29
timestamp 1676037725
transform 1 0 37444 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold30
timestamp 1676037725
transform 1 0 36708 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold31
timestamp 1676037725
transform 1 0 37444 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold32
timestamp 1676037725
transform 1 0 33120 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold33
timestamp 1676037725
transform 1 0 32384 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold34
timestamp 1676037725
transform 1 0 34040 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold35
timestamp 1676037725
transform 1 0 33672 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold36
timestamp 1676037725
transform 1 0 32108 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold37
timestamp 1676037725
transform 1 0 40112 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold38
timestamp 1676037725
transform 1 0 36708 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold39
timestamp 1676037725
transform 1 0 34868 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold40
timestamp 1676037725
transform 1 0 30084 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold41
timestamp 1676037725
transform 1 0 29440 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold42
timestamp 1676037725
transform 1 0 30636 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold43
timestamp 1676037725
transform 1 0 41584 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold44
timestamp 1676037725
transform 1 0 34960 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold45
timestamp 1676037725
transform 1 0 45908 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold46
timestamp 1676037725
transform 1 0 37444 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold47
timestamp 1676037725
transform 1 0 38456 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold48
timestamp 1676037725
transform 1 0 39192 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold49
timestamp 1676037725
transform 1 0 28244 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold50
timestamp 1676037725
transform 1 0 27968 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold51
timestamp 1676037725
transform 1 0 27048 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold52
timestamp 1676037725
transform 1 0 21068 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold53
timestamp 1676037725
transform 1 0 20240 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold54
timestamp 1676037725
transform 1 0 27508 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold55
timestamp 1676037725
transform 1 0 23460 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold56
timestamp 1676037725
transform 1 0 22908 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold57
timestamp 1676037725
transform 1 0 39100 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold58
timestamp 1676037725
transform 1 0 32016 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold59
timestamp 1676037725
transform 1 0 32752 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold60
timestamp 1676037725
transform 1 0 22540 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold61
timestamp 1676037725
transform 1 0 18308 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold62
timestamp 1676037725
transform 1 0 17480 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold63
timestamp 1676037725
transform 1 0 29624 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold64
timestamp 1676037725
transform 1 0 28428 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold65
timestamp 1676037725
transform 1 0 29716 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold66
timestamp 1676037725
transform 1 0 30452 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold67
timestamp 1676037725
transform 1 0 40204 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold68
timestamp 1676037725
transform 1 0 33948 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold69
timestamp 1676037725
transform 1 0 30268 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold70
timestamp 1676037725
transform 1 0 31004 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold71
timestamp 1676037725
transform 1 0 43332 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold72
timestamp 1676037725
transform 1 0 32292 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold73
timestamp 1676037725
transform 1 0 26220 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold74
timestamp 1676037725
transform 1 0 26312 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold75
timestamp 1676037725
transform 1 0 43424 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold76
timestamp 1676037725
transform 1 0 39192 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold77
timestamp 1676037725
transform 1 0 35972 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold78
timestamp 1676037725
transform 1 0 36708 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold79
timestamp 1676037725
transform 1 0 40940 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold80
timestamp 1676037725
transform 1 0 33488 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold81
timestamp 1676037725
transform 1 0 28888 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold82
timestamp 1676037725
transform 1 0 29532 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold83
timestamp 1676037725
transform 1 0 40020 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold84
timestamp 1676037725
transform 1 0 31740 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold85
timestamp 1676037725
transform 1 0 26312 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold86
timestamp 1676037725
transform 1 0 26864 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold87
timestamp 1676037725
transform 1 0 30820 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold88
timestamp 1676037725
transform 1 0 23644 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold89
timestamp 1676037725
transform 1 0 20792 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold90
timestamp 1676037725
transform 1 0 20516 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold91
timestamp 1676037725
transform 1 0 40112 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold92
timestamp 1676037725
transform 1 0 41676 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold93
timestamp 1676037725
transform 1 0 37168 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold94
timestamp 1676037725
transform 1 0 35052 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold95
timestamp 1676037725
transform 1 0 26404 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold96
timestamp 1676037725
transform 1 0 23184 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold97
timestamp 1676037725
transform 1 0 20424 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold98
timestamp 1676037725
transform 1 0 21988 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold99
timestamp 1676037725
transform 1 0 28060 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold100
timestamp 1676037725
transform 1 0 21160 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold101
timestamp 1676037725
transform 1 0 16008 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold102
timestamp 1676037725
transform 1 0 17572 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold103
timestamp 1676037725
transform 1 0 36616 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold104
timestamp 1676037725
transform 1 0 38180 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold105
timestamp 1676037725
transform 1 0 37444 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold106
timestamp 1676037725
transform 1 0 36524 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold107
timestamp 1676037725
transform 1 0 35788 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold108
timestamp 1676037725
transform 1 0 36524 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold109
timestamp 1676037725
transform 1 0 40296 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold110
timestamp 1676037725
transform 1 0 40756 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold111
timestamp 1676037725
transform 1 0 38364 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold112
timestamp 1676037725
transform 1 0 34868 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold113
timestamp 1676037725
transform 1 0 33580 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold114
timestamp 1676037725
transform 1 0 33488 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold115
timestamp 1676037725
transform 1 0 39376 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold116
timestamp 1676037725
transform 1 0 35420 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold117
timestamp 1676037725
transform 1 0 33856 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold118
timestamp 1676037725
transform 1 0 32292 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold119
timestamp 1676037725
transform 1 0 42596 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold120
timestamp 1676037725
transform 1 0 40020 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold121
timestamp 1676037725
transform 1 0 38916 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold122
timestamp 1676037725
transform 1 0 36616 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold123
timestamp 1676037725
transform 1 0 34684 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold124
timestamp 1676037725
transform 1 0 30820 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold125
timestamp 1676037725
transform 1 0 28152 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold126
timestamp 1676037725
transform 1 0 28888 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold127
timestamp 1676037725
transform 1 0 31556 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold128
timestamp 1676037725
transform 1 0 31096 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold129
timestamp 1676037725
transform 1 0 28888 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold130
timestamp 1676037725
transform 1 0 34868 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold131
timestamp 1676037725
transform 1 0 34408 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold132
timestamp 1676037725
transform 1 0 32752 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold133
timestamp 1676037725
transform 1 0 31464 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold134
timestamp 1676037725
transform 1 0 41032 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold135
timestamp 1676037725
transform 1 0 38456 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold136
timestamp 1676037725
transform 1 0 38180 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold137
timestamp 1676037725
transform 1 0 33304 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold138
timestamp 1676037725
transform 1 0 44344 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold139
timestamp 1676037725
transform 1 0 40848 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold140
timestamp 1676037725
transform 1 0 40756 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold141
timestamp 1676037725
transform 1 0 26312 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold142
timestamp 1676037725
transform 1 0 21068 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold143
timestamp 1676037725
transform 1 0 18400 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold144
timestamp 1676037725
transform 1 0 40756 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold145
timestamp 1676037725
transform 1 0 32568 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold146
timestamp 1676037725
transform 1 0 27140 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold147
timestamp 1676037725
transform 1 0 42596 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold148
timestamp 1676037725
transform 1 0 35052 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold149
timestamp 1676037725
transform 1 0 30268 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold150
timestamp 1676037725
transform 1 0 29256 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold151
timestamp 1676037725
transform 1 0 25944 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold152
timestamp 1676037725
transform 1 0 20976 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold153
timestamp 1676037725
transform 1 0 28888 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold154
timestamp 1676037725
transform 1 0 25024 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold155
timestamp 1676037725
transform 1 0 42688 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold156
timestamp 1676037725
transform 1 0 45172 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold157
timestamp 1676037725
transform 1 0 40020 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1676037725
transform 1 0 44252 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input2
timestamp 1676037725
transform 1 0 41584 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input3
timestamp 1676037725
transform 1 0 42596 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 1676037725
transform 1 0 42688 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1676037725
transform 1 0 45908 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input6
timestamp 1676037725
transform 1 0 44068 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1676037725
transform 1 0 45172 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1676037725
transform 1 0 44804 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1676037725
transform 1 0 45172 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 1676037725
transform 1 0 46644 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input11
timestamp 1676037725
transform 1 0 49956 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input12
timestamp 1676037725
transform 1 0 43332 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1676037725
transform 1 0 45540 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1676037725
transform 1 0 45908 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input15
timestamp 1676037725
transform 1 0 46644 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1676037725
transform 1 0 46276 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp 1676037725
transform 1 0 46184 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input18
timestamp 1676037725
transform 1 0 45724 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 1676037725
transform 1 0 46460 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input20
timestamp 1676037725
transform 1 0 43700 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input21
timestamp 1676037725
transform 1 0 40020 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input22
timestamp 1676037725
transform 1 0 44436 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input23
timestamp 1676037725
transform 1 0 41032 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input24
timestamp 1676037725
transform 1 0 41952 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input25
timestamp 1676037725
transform 1 0 45172 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input26
timestamp 1676037725
transform 1 0 41032 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input27
timestamp 1676037725
transform 1 0 41768 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input28
timestamp 1676037725
transform 1 0 2300 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input29
timestamp 1676037725
transform 1 0 1564 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input30
timestamp 1676037725
transform 1 0 1564 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input31
timestamp 1676037725
transform 1 0 1564 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input32
timestamp 1676037725
transform 1 0 1564 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input33
timestamp 1676037725
transform 1 0 2300 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input34
timestamp 1676037725
transform 1 0 1564 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input35
timestamp 1676037725
transform 1 0 1564 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input36
timestamp 1676037725
transform 1 0 46276 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input37
timestamp 1676037725
transform 1 0 52900 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input38
timestamp 1676037725
transform 1 0 50324 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input39
timestamp 1676037725
transform 1 0 50416 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input40
timestamp 1676037725
transform 1 0 51060 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input41
timestamp 1676037725
transform 1 0 51796 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input42
timestamp 1676037725
transform 1 0 54372 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input43
timestamp 1676037725
transform 1 0 51152 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input44
timestamp 1676037725
transform 1 0 53636 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input45
timestamp 1676037725
transform 1 0 51888 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input46
timestamp 1676037725
transform 1 0 52532 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input47
timestamp 1676037725
transform 1 0 47196 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input48
timestamp 1676037725
transform 1 0 55108 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input49
timestamp 1676037725
transform 1 0 53268 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 1676037725
transform 1 0 52900 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input51
timestamp 1676037725
transform 1 0 55844 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input52
timestamp 1676037725
transform 1 0 58052 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input53
timestamp 1676037725
transform 1 0 54004 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input54
timestamp 1676037725
transform 1 0 55476 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input55
timestamp 1676037725
transform 1 0 50692 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input56
timestamp 1676037725
transform 1 0 51428 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input57
timestamp 1676037725
transform 1 0 52900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input58
timestamp 1676037725
transform 1 0 50324 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input59
timestamp 1676037725
transform 1 0 49128 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input60
timestamp 1676037725
transform 1 0 49680 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input61
timestamp 1676037725
transform 1 0 49036 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input62
timestamp 1676037725
transform 1 0 51428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input63
timestamp 1676037725
transform 1 0 24564 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input64
timestamp 1676037725
transform 1 0 37444 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input65
timestamp 1676037725
transform 1 0 38364 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input66
timestamp 1676037725
transform 1 0 40020 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input67
timestamp 1676037725
transform 1 0 40940 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input68
timestamp 1676037725
transform 1 0 42596 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input69
timestamp 1676037725
transform 1 0 43516 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input70
timestamp 1676037725
transform 1 0 45172 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input71
timestamp 1676037725
transform 1 0 46092 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input72
timestamp 1676037725
transform 1 0 47748 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input73
timestamp 1676037725
transform 1 0 48668 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input74
timestamp 1676037725
transform 1 0 25484 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input75
timestamp 1676037725
transform 1 0 50324 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input76
timestamp 1676037725
transform 1 0 51244 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input77
timestamp 1676037725
transform 1 0 52900 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input78
timestamp 1676037725
transform 1 0 53820 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input79
timestamp 1676037725
transform 1 0 55476 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input80
timestamp 1676037725
transform 1 0 56304 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input81
timestamp 1676037725
transform 1 0 57684 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input82
timestamp 1676037725
transform 1 0 27140 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input83
timestamp 1676037725
transform 1 0 28060 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input84
timestamp 1676037725
transform 1 0 29716 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input85
timestamp 1676037725
transform 1 0 30636 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input86
timestamp 1676037725
transform 1 0 32292 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input87
timestamp 1676037725
transform 1 0 33212 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input88
timestamp 1676037725
transform 1 0 34868 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input89
timestamp 1676037725
transform 1 0 35788 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input90
timestamp 1676037725
transform 1 0 1564 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input91
timestamp 1676037725
transform 1 0 1564 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input92
timestamp 1676037725
transform 1 0 1564 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input93
timestamp 1676037725
transform 1 0 1564 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input94
timestamp 1676037725
transform 1 0 1564 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input95
timestamp 1676037725
transform 1 0 1564 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input96
timestamp 1676037725
transform 1 0 1564 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input97
timestamp 1676037725
transform 1 0 1564 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input98
timestamp 1676037725
transform 1 0 1564 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input99
timestamp 1676037725
transform 1 0 1564 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input100
timestamp 1676037725
transform 1 0 1564 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input101
timestamp 1676037725
transform 1 0 1564 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input102
timestamp 1676037725
transform 1 0 1564 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input103
timestamp 1676037725
transform 1 0 1564 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input104
timestamp 1676037725
transform 1 0 1564 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input105
timestamp 1676037725
transform 1 0 1564 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input106
timestamp 1676037725
transform 1 0 1564 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input107
timestamp 1676037725
transform 1 0 1564 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input108
timestamp 1676037725
transform 1 0 1564 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input109
timestamp 1676037725
transform 1 0 1564 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input110
timestamp 1676037725
transform 1 0 1564 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input111
timestamp 1676037725
transform 1 0 1564 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input112
timestamp 1676037725
transform 1 0 1564 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input113
timestamp 1676037725
transform 1 0 1564 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input114
timestamp 1676037725
transform 1 0 1564 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input115
timestamp 1676037725
transform 1 0 1564 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input116
timestamp 1676037725
transform 1 0 1564 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input117
timestamp 1676037725
transform 1 0 1564 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input118
timestamp 1676037725
transform 1 0 58052 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input119
timestamp 1676037725
transform 1 0 57224 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input120
timestamp 1676037725
transform 1 0 58052 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input121
timestamp 1676037725
transform 1 0 57868 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input122
timestamp 1676037725
transform 1 0 58052 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input123
timestamp 1676037725
transform 1 0 58052 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input124
timestamp 1676037725
transform 1 0 58052 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input125
timestamp 1676037725
transform 1 0 58052 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input126
timestamp 1676037725
transform 1 0 57316 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input127
timestamp 1676037725
transform 1 0 58052 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input128
timestamp 1676037725
transform 1 0 58052 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input129
timestamp 1676037725
transform 1 0 57132 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input130
timestamp 1676037725
transform 1 0 57224 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input131
timestamp 1676037725
transform 1 0 58052 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input132
timestamp 1676037725
transform 1 0 56028 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input133
timestamp 1676037725
transform 1 0 57316 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input134
timestamp 1676037725
transform 1 0 56488 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input135
timestamp 1676037725
transform 1 0 57040 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input136
timestamp 1676037725
transform 1 0 55752 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input137
timestamp 1676037725
transform 1 0 57868 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input138
timestamp 1676037725
transform 1 0 57868 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input139
timestamp 1676037725
transform 1 0 58052 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input140
timestamp 1676037725
transform 1 0 58052 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input141
timestamp 1676037725
transform 1 0 58052 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input142
timestamp 1676037725
transform 1 0 58052 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input143
timestamp 1676037725
transform 1 0 58052 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input144
timestamp 1676037725
transform 1 0 57316 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input145
timestamp 1676037725
transform 1 0 58052 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input146
timestamp 1676037725
transform 1 0 58052 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input147
timestamp 1676037725
transform 1 0 57224 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input148
timestamp 1676037725
transform 1 0 57868 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input149
timestamp 1676037725
transform 1 0 58052 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input150
timestamp 1676037725
transform 1 0 58052 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input151
timestamp 1676037725
transform 1 0 58052 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input152
timestamp 1676037725
transform 1 0 57132 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input153
timestamp 1676037725
transform 1 0 57868 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input154
timestamp 1676037725
transform 1 0 58052 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input155
timestamp 1676037725
transform 1 0 57868 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input156
timestamp 1676037725
transform 1 0 58052 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input157
timestamp 1676037725
transform 1 0 12604 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input158
timestamp 1676037725
transform 1 0 14260 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input159
timestamp 1676037725
transform 1 0 15180 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input160
timestamp 1676037725
transform 1 0 16836 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input161
timestamp 1676037725
transform 1 0 17756 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input162
timestamp 1676037725
transform 1 0 19412 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input163
timestamp 1676037725
transform 1 0 20332 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input164
timestamp 1676037725
transform 1 0 21988 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input165
timestamp 1676037725
transform 1 0 1564 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input166
timestamp 1676037725
transform 1 0 2300 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input167
timestamp 1676037725
transform 1 0 1564 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input168
timestamp 1676037725
transform 1 0 1564 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input169
timestamp 1676037725
transform 1 0 1564 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input170
timestamp 1676037725
transform 1 0 1564 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input171
timestamp 1676037725
transform 1 0 1564 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input172
timestamp 1676037725
transform 1 0 1564 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input173
timestamp 1676037725
transform 1 0 1564 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input174
timestamp 1676037725
transform 1 0 2300 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input175
timestamp 1676037725
transform 1 0 3956 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input176
timestamp 1676037725
transform 1 0 4876 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input177
timestamp 1676037725
transform 1 0 6532 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input178
timestamp 1676037725
transform 1 0 7452 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input179
timestamp 1676037725
transform 1 0 9108 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input180
timestamp 1676037725
transform 1 0 10028 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input181
timestamp 1676037725
transform 1 0 11684 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input182
timestamp 1676037725
transform 1 0 41676 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input183
timestamp 1676037725
transform 1 0 43516 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input184
timestamp 1676037725
transform 1 0 38824 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input185
timestamp 1676037725
transform 1 0 42596 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input186
timestamp 1676037725
transform 1 0 1564 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input187
timestamp 1676037725
transform 1 0 1564 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input188
timestamp 1676037725
transform 1 0 1564 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input189
timestamp 1676037725
transform 1 0 1564 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input190
timestamp 1676037725
transform 1 0 1564 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input191
timestamp 1676037725
transform 1 0 1564 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input192
timestamp 1676037725
transform 1 0 1564 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input193
timestamp 1676037725
transform 1 0 1564 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input194
timestamp 1676037725
transform 1 0 54004 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input195
timestamp 1676037725
transform 1 0 5704 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input196
timestamp 1676037725
transform 1 0 8280 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input197
timestamp 1676037725
transform 1 0 9016 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input198
timestamp 1676037725
transform 1 0 7452 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input199
timestamp 1676037725
transform 1 0 6808 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input200
timestamp 1676037725
transform 1 0 8188 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input201
timestamp 1676037725
transform 1 0 7544 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input202
timestamp 1676037725
transform 1 0 10396 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input203
timestamp 1676037725
transform 1 0 8924 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input204
timestamp 1676037725
transform 1 0 8280 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input205
timestamp 1676037725
transform 1 0 10856 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input206
timestamp 1676037725
transform 1 0 11500 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input207
timestamp 1676037725
transform 1 0 9384 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input208
timestamp 1676037725
transform 1 0 10120 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input209
timestamp 1676037725
transform 1 0 10856 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input210
timestamp 1676037725
transform 1 0 10856 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input211
timestamp 1676037725
transform 1 0 12696 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input212
timestamp 1676037725
transform 1 0 11960 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input213
timestamp 1676037725
transform 1 0 13432 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input214
timestamp 1676037725
transform 1 0 12880 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input215
timestamp 1676037725
transform 1 0 12696 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input216
timestamp 1676037725
transform 1 0 14260 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input217
timestamp 1676037725
transform 1 0 13616 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input218
timestamp 1676037725
transform 1 0 13432 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input219
timestamp 1676037725
transform 1 0 14352 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input220
timestamp 1676037725
transform 1 0 15088 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input221
timestamp 1676037725
transform 1 0 15640 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input222
timestamp 1676037725
transform 1 0 15088 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input223
timestamp 1676037725
transform 1 0 15824 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input224
timestamp 1676037725
transform 1 0 5704 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input225
timestamp 1676037725
transform 1 0 6808 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input226
timestamp 1676037725
transform 1 0 6716 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input227
timestamp 1676037725
transform 1 0 8188 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input228
timestamp 1676037725
transform 1 0 7544 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input229
timestamp 1676037725
transform 1 0 41216 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input230
timestamp 1676037725
transform 1 0 58052 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input231
timestamp 1676037725
transform 1 0 22908 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input232
timestamp 1676037725
transform 1 0 1564 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input233
timestamp 1676037725
transform 1 0 56764 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input234
timestamp 1676037725
transform 1 0 1564 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input235
timestamp 1676037725
transform 1 0 55200 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input236
timestamp 1676037725
transform 1 0 58052 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input237
timestamp 1676037725
transform 1 0 58052 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input238
timestamp 1676037725
transform 1 0 57868 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input239
timestamp 1676037725
transform 1 0 56212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input240
timestamp 1676037725
transform 1 0 58052 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input241
timestamp 1676037725
transform 1 0 58052 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input242
timestamp 1676037725
transform 1 0 58052 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input243
timestamp 1676037725
transform 1 0 58052 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input244
timestamp 1676037725
transform 1 0 58052 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input245
timestamp 1676037725
transform 1 0 58052 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input246
timestamp 1676037725
transform 1 0 58052 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input247
timestamp 1676037725
transform 1 0 58052 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input248
timestamp 1676037725
transform 1 0 58052 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input249
timestamp 1676037725
transform 1 0 58052 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input250
timestamp 1676037725
transform 1 0 58052 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input251
timestamp 1676037725
transform 1 0 58052 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input252
timestamp 1676037725
transform 1 0 58052 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input253
timestamp 1676037725
transform 1 0 58052 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input254
timestamp 1676037725
transform 1 0 58052 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input255
timestamp 1676037725
transform 1 0 58052 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input256
timestamp 1676037725
transform 1 0 58052 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input257
timestamp 1676037725
transform 1 0 58052 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input258
timestamp 1676037725
transform 1 0 58052 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input259
timestamp 1676037725
transform 1 0 58052 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input260
timestamp 1676037725
transform 1 0 55752 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input261
timestamp 1676037725
transform 1 0 58052 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input262
timestamp 1676037725
transform 1 0 58052 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input263
timestamp 1676037725
transform 1 0 56948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input264
timestamp 1676037725
transform 1 0 58052 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input265
timestamp 1676037725
transform 1 0 58052 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input266
timestamp 1676037725
transform 1 0 58052 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input267
timestamp 1676037725
transform 1 0 58052 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input268
timestamp 1676037725
transform 1 0 55384 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input269
timestamp 1676037725
transform 1 0 54464 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  max_cap418
timestamp 1676037725
transform 1 0 24196 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  multiplexer_480 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 26404 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_481
timestamp 1676037725
transform 1 0 26404 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_482
timestamp 1676037725
transform 1 0 27048 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_483
timestamp 1676037725
transform 1 0 24380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_484
timestamp 1676037725
transform 1 0 14260 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_485
timestamp 1676037725
transform 1 0 18308 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_486
timestamp 1676037725
transform 1 0 18400 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_487
timestamp 1676037725
transform 1 0 16836 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_488
timestamp 1676037725
transform 1 0 16836 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_489
timestamp 1676037725
transform 1 0 19412 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_490
timestamp 1676037725
transform 1 0 58144 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_491
timestamp 1676037725
transform 1 0 58144 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_492
timestamp 1676037725
transform 1 0 58144 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_493
timestamp 1676037725
transform 1 0 58144 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_494
timestamp 1676037725
transform 1 0 28796 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_495
timestamp 1676037725
transform 1 0 28520 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_496
timestamp 1676037725
transform 1 0 28244 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_497
timestamp 1676037725
transform 1 0 28060 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_498
timestamp 1676037725
transform 1 0 28612 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_499
timestamp 1676037725
transform 1 0 29256 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output270
timestamp 1676037725
transform 1 0 2484 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  output271
timestamp 1676037725
transform 1 0 1564 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output272
timestamp 1676037725
transform 1 0 1564 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output273
timestamp 1676037725
transform 1 0 1564 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output274
timestamp 1676037725
transform 1 0 1564 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output275
timestamp 1676037725
transform 1 0 1564 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output276
timestamp 1676037725
transform 1 0 1564 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output277
timestamp 1676037725
transform 1 0 1564 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output278
timestamp 1676037725
transform 1 0 1564 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output279
timestamp 1676037725
transform 1 0 1564 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output280
timestamp 1676037725
transform 1 0 1564 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output281
timestamp 1676037725
transform 1 0 1564 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output282
timestamp 1676037725
transform 1 0 1564 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output283
timestamp 1676037725
transform 1 0 1564 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output284
timestamp 1676037725
transform 1 0 1564 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output285
timestamp 1676037725
transform 1 0 1564 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output286
timestamp 1676037725
transform 1 0 1564 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output287
timestamp 1676037725
transform 1 0 1564 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output288
timestamp 1676037725
transform 1 0 1564 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output289
timestamp 1676037725
transform 1 0 1564 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output290
timestamp 1676037725
transform 1 0 1564 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output291
timestamp 1676037725
transform 1 0 1564 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output292
timestamp 1676037725
transform 1 0 1564 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output293
timestamp 1676037725
transform 1 0 1564 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output294
timestamp 1676037725
transform 1 0 1564 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output295
timestamp 1676037725
transform 1 0 1564 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output296
timestamp 1676037725
transform 1 0 1564 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output297
timestamp 1676037725
transform 1 0 1564 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output298
timestamp 1676037725
transform 1 0 1564 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output299
timestamp 1676037725
transform 1 0 27140 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output300
timestamp 1676037725
transform 1 0 28704 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output301
timestamp 1676037725
transform 1 0 29900 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output302
timestamp 1676037725
transform 1 0 30176 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output303
timestamp 1676037725
transform 1 0 30820 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output304
timestamp 1676037725
transform 1 0 31096 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output305
timestamp 1676037725
transform 1 0 32292 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output306
timestamp 1676037725
transform 1 0 32292 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output307
timestamp 1676037725
transform 1 0 33212 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output308
timestamp 1676037725
transform 1 0 33212 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output309
timestamp 1676037725
transform 1 0 32936 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output310
timestamp 1676037725
transform 1 0 34132 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output311
timestamp 1676037725
transform 1 0 34868 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output312
timestamp 1676037725
transform 1 0 33856 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output313
timestamp 1676037725
transform 1 0 35052 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output314
timestamp 1676037725
transform 1 0 35788 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output315
timestamp 1676037725
transform 1 0 34868 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output316
timestamp 1676037725
transform 1 0 35972 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output317
timestamp 1676037725
transform 1 0 34684 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output318
timestamp 1676037725
transform 1 0 37444 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output319
timestamp 1676037725
transform 1 0 35604 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output320
timestamp 1676037725
transform 1 0 37444 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output321
timestamp 1676037725
transform 1 0 38364 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output322
timestamp 1676037725
transform 1 0 37444 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output323
timestamp 1676037725
transform 1 0 39468 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output324
timestamp 1676037725
transform 1 0 40020 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output325
timestamp 1676037725
transform 1 0 38364 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output326
timestamp 1676037725
transform 1 0 37812 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output327
timestamp 1676037725
transform 1 0 14904 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output328
timestamp 1676037725
transform 1 0 15824 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output329
timestamp 1676037725
transform 1 0 19780 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output330
timestamp 1676037725
transform 1 0 17480 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output331
timestamp 1676037725
transform 1 0 19412 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output332
timestamp 1676037725
transform 1 0 18400 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output333
timestamp 1676037725
transform 1 0 19136 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output334
timestamp 1676037725
transform 1 0 20332 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output335
timestamp 1676037725
transform 1 0 20976 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output336
timestamp 1676037725
transform 1 0 17480 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output337
timestamp 1676037725
transform 1 0 15824 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output338
timestamp 1676037725
transform 1 0 18400 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output339
timestamp 1676037725
transform 1 0 19412 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output340
timestamp 1676037725
transform 1 0 18400 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output341
timestamp 1676037725
transform 1 0 19320 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output342
timestamp 1676037725
transform 1 0 21068 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output343
timestamp 1676037725
transform 1 0 20056 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output344
timestamp 1676037725
transform 1 0 21896 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output345
timestamp 1676037725
transform 1 0 22448 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output346
timestamp 1676037725
transform 1 0 20976 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output347
timestamp 1676037725
transform 1 0 22540 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output348
timestamp 1676037725
transform 1 0 16560 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output349
timestamp 1676037725
transform 1 0 24288 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output350
timestamp 1676037725
transform 1 0 22632 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output351
timestamp 1676037725
transform 1 0 23460 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output352
timestamp 1676037725
transform 1 0 23552 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output353
timestamp 1676037725
transform 1 0 24932 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output354
timestamp 1676037725
transform 1 0 25208 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output355
timestamp 1676037725
transform 1 0 27140 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output356
timestamp 1676037725
transform 1 0 26128 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output357
timestamp 1676037725
transform 1 0 17296 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output358
timestamp 1676037725
transform 1 0 17480 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output359
timestamp 1676037725
transform 1 0 1564 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output360
timestamp 1676037725
transform 1 0 1564 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output361
timestamp 1676037725
transform 1 0 1564 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output362
timestamp 1676037725
transform 1 0 1564 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output363
timestamp 1676037725
transform 1 0 1564 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output364
timestamp 1676037725
transform 1 0 1564 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output365
timestamp 1676037725
transform 1 0 1564 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output366
timestamp 1676037725
transform 1 0 1564 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output367
timestamp 1676037725
transform 1 0 1564 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output368
timestamp 1676037725
transform 1 0 1564 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output369
timestamp 1676037725
transform 1 0 1564 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output370
timestamp 1676037725
transform 1 0 1564 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output371
timestamp 1676037725
transform 1 0 57040 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output372
timestamp 1676037725
transform 1 0 56120 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output373
timestamp 1676037725
transform 1 0 57040 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output374
timestamp 1676037725
transform 1 0 56948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output375
timestamp 1676037725
transform 1 0 57868 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output376
timestamp 1676037725
transform 1 0 57868 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output377
timestamp 1676037725
transform 1 0 56948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output378
timestamp 1676037725
transform 1 0 57868 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output379
timestamp 1676037725
transform 1 0 57868 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output380
timestamp 1676037725
transform 1 0 57868 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output381
timestamp 1676037725
transform 1 0 57868 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output382
timestamp 1676037725
transform 1 0 57868 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output383
timestamp 1676037725
transform 1 0 57040 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output384
timestamp 1676037725
transform 1 0 57868 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output385
timestamp 1676037725
transform 1 0 57868 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output386
timestamp 1676037725
transform 1 0 56948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output387
timestamp 1676037725
transform 1 0 57868 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output388
timestamp 1676037725
transform 1 0 57868 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output389
timestamp 1676037725
transform 1 0 57868 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output390
timestamp 1676037725
transform 1 0 57868 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output391
timestamp 1676037725
transform 1 0 57868 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output392
timestamp 1676037725
transform 1 0 57040 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output393
timestamp 1676037725
transform 1 0 57868 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output394
timestamp 1676037725
transform 1 0 57040 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output395
timestamp 1676037725
transform 1 0 57040 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output396
timestamp 1676037725
transform 1 0 57868 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output397
timestamp 1676037725
transform 1 0 57040 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output398
timestamp 1676037725
transform 1 0 57868 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output399
timestamp 1676037725
transform 1 0 57868 0 1 15232
box -38 -48 590 592
<< labels >>
flabel metal3 s 0 19320 800 19440 0 FreeSans 480 0 0 0 design_clk_o
port 0 nsew signal tristate
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 dsi_all[0]
port 1 nsew signal tristate
flabel metal3 s 0 9528 800 9648 0 FreeSans 480 0 0 0 dsi_all[10]
port 2 nsew signal tristate
flabel metal3 s 0 10072 800 10192 0 FreeSans 480 0 0 0 dsi_all[11]
port 3 nsew signal tristate
flabel metal3 s 0 10616 800 10736 0 FreeSans 480 0 0 0 dsi_all[12]
port 4 nsew signal tristate
flabel metal3 s 0 11160 800 11280 0 FreeSans 480 0 0 0 dsi_all[13]
port 5 nsew signal tristate
flabel metal3 s 0 11704 800 11824 0 FreeSans 480 0 0 0 dsi_all[14]
port 6 nsew signal tristate
flabel metal3 s 0 12248 800 12368 0 FreeSans 480 0 0 0 dsi_all[15]
port 7 nsew signal tristate
flabel metal3 s 0 12792 800 12912 0 FreeSans 480 0 0 0 dsi_all[16]
port 8 nsew signal tristate
flabel metal3 s 0 13336 800 13456 0 FreeSans 480 0 0 0 dsi_all[17]
port 9 nsew signal tristate
flabel metal3 s 0 13880 800 14000 0 FreeSans 480 0 0 0 dsi_all[18]
port 10 nsew signal tristate
flabel metal3 s 0 14424 800 14544 0 FreeSans 480 0 0 0 dsi_all[19]
port 11 nsew signal tristate
flabel metal3 s 0 4632 800 4752 0 FreeSans 480 0 0 0 dsi_all[1]
port 12 nsew signal tristate
flabel metal3 s 0 14968 800 15088 0 FreeSans 480 0 0 0 dsi_all[20]
port 13 nsew signal tristate
flabel metal3 s 0 15512 800 15632 0 FreeSans 480 0 0 0 dsi_all[21]
port 14 nsew signal tristate
flabel metal3 s 0 16056 800 16176 0 FreeSans 480 0 0 0 dsi_all[22]
port 15 nsew signal tristate
flabel metal3 s 0 16600 800 16720 0 FreeSans 480 0 0 0 dsi_all[23]
port 16 nsew signal tristate
flabel metal3 s 0 17144 800 17264 0 FreeSans 480 0 0 0 dsi_all[24]
port 17 nsew signal tristate
flabel metal3 s 0 17688 800 17808 0 FreeSans 480 0 0 0 dsi_all[25]
port 18 nsew signal tristate
flabel metal3 s 0 18232 800 18352 0 FreeSans 480 0 0 0 dsi_all[26]
port 19 nsew signal tristate
flabel metal3 s 0 18776 800 18896 0 FreeSans 480 0 0 0 dsi_all[27]
port 20 nsew signal tristate
flabel metal3 s 0 5176 800 5296 0 FreeSans 480 0 0 0 dsi_all[2]
port 21 nsew signal tristate
flabel metal3 s 0 5720 800 5840 0 FreeSans 480 0 0 0 dsi_all[3]
port 22 nsew signal tristate
flabel metal3 s 0 6264 800 6384 0 FreeSans 480 0 0 0 dsi_all[4]
port 23 nsew signal tristate
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 dsi_all[5]
port 24 nsew signal tristate
flabel metal3 s 0 7352 800 7472 0 FreeSans 480 0 0 0 dsi_all[6]
port 25 nsew signal tristate
flabel metal3 s 0 7896 800 8016 0 FreeSans 480 0 0 0 dsi_all[7]
port 26 nsew signal tristate
flabel metal3 s 0 8440 800 8560 0 FreeSans 480 0 0 0 dsi_all[8]
port 27 nsew signal tristate
flabel metal3 s 0 8984 800 9104 0 FreeSans 480 0 0 0 dsi_all[9]
port 28 nsew signal tristate
flabel metal2 s 38750 0 38806 800 0 FreeSans 224 90 0 0 dso_6502[0]
port 29 nsew signal input
flabel metal2 s 41510 0 41566 800 0 FreeSans 224 90 0 0 dso_6502[10]
port 30 nsew signal input
flabel metal2 s 41786 0 41842 800 0 FreeSans 224 90 0 0 dso_6502[11]
port 31 nsew signal input
flabel metal2 s 42062 0 42118 800 0 FreeSans 224 90 0 0 dso_6502[12]
port 32 nsew signal input
flabel metal2 s 42338 0 42394 800 0 FreeSans 224 90 0 0 dso_6502[13]
port 33 nsew signal input
flabel metal2 s 42614 0 42670 800 0 FreeSans 224 90 0 0 dso_6502[14]
port 34 nsew signal input
flabel metal2 s 42890 0 42946 800 0 FreeSans 224 90 0 0 dso_6502[15]
port 35 nsew signal input
flabel metal2 s 43166 0 43222 800 0 FreeSans 224 90 0 0 dso_6502[16]
port 36 nsew signal input
flabel metal2 s 43442 0 43498 800 0 FreeSans 224 90 0 0 dso_6502[17]
port 37 nsew signal input
flabel metal2 s 43718 0 43774 800 0 FreeSans 224 90 0 0 dso_6502[18]
port 38 nsew signal input
flabel metal2 s 43994 0 44050 800 0 FreeSans 224 90 0 0 dso_6502[19]
port 39 nsew signal input
flabel metal2 s 39026 0 39082 800 0 FreeSans 224 90 0 0 dso_6502[1]
port 40 nsew signal input
flabel metal2 s 44270 0 44326 800 0 FreeSans 224 90 0 0 dso_6502[20]
port 41 nsew signal input
flabel metal2 s 44546 0 44602 800 0 FreeSans 224 90 0 0 dso_6502[21]
port 42 nsew signal input
flabel metal2 s 44822 0 44878 800 0 FreeSans 224 90 0 0 dso_6502[22]
port 43 nsew signal input
flabel metal2 s 45098 0 45154 800 0 FreeSans 224 90 0 0 dso_6502[23]
port 44 nsew signal input
flabel metal2 s 45374 0 45430 800 0 FreeSans 224 90 0 0 dso_6502[24]
port 45 nsew signal input
flabel metal2 s 45650 0 45706 800 0 FreeSans 224 90 0 0 dso_6502[25]
port 46 nsew signal input
flabel metal2 s 45926 0 45982 800 0 FreeSans 224 90 0 0 dso_6502[26]
port 47 nsew signal input
flabel metal2 s 39302 0 39358 800 0 FreeSans 224 90 0 0 dso_6502[2]
port 48 nsew signal input
flabel metal2 s 39578 0 39634 800 0 FreeSans 224 90 0 0 dso_6502[3]
port 49 nsew signal input
flabel metal2 s 39854 0 39910 800 0 FreeSans 224 90 0 0 dso_6502[4]
port 50 nsew signal input
flabel metal2 s 40130 0 40186 800 0 FreeSans 224 90 0 0 dso_6502[5]
port 51 nsew signal input
flabel metal2 s 40406 0 40462 800 0 FreeSans 224 90 0 0 dso_6502[6]
port 52 nsew signal input
flabel metal2 s 40682 0 40738 800 0 FreeSans 224 90 0 0 dso_6502[7]
port 53 nsew signal input
flabel metal2 s 40958 0 41014 800 0 FreeSans 224 90 0 0 dso_6502[8]
port 54 nsew signal input
flabel metal2 s 41234 0 41290 800 0 FreeSans 224 90 0 0 dso_6502[9]
port 55 nsew signal input
flabel metal3 s 0 26392 800 26512 0 FreeSans 480 0 0 0 dso_LCD[0]
port 56 nsew signal input
flabel metal3 s 0 26936 800 27056 0 FreeSans 480 0 0 0 dso_LCD[1]
port 57 nsew signal input
flabel metal3 s 0 27480 800 27600 0 FreeSans 480 0 0 0 dso_LCD[2]
port 58 nsew signal input
flabel metal3 s 0 28024 800 28144 0 FreeSans 480 0 0 0 dso_LCD[3]
port 59 nsew signal input
flabel metal3 s 0 28568 800 28688 0 FreeSans 480 0 0 0 dso_LCD[4]
port 60 nsew signal input
flabel metal3 s 0 29112 800 29232 0 FreeSans 480 0 0 0 dso_LCD[5]
port 61 nsew signal input
flabel metal3 s 0 29656 800 29776 0 FreeSans 480 0 0 0 dso_LCD[6]
port 62 nsew signal input
flabel metal3 s 0 30200 800 30320 0 FreeSans 480 0 0 0 dso_LCD[7]
port 63 nsew signal input
flabel metal2 s 46202 0 46258 800 0 FreeSans 224 90 0 0 dso_as1802[0]
port 64 nsew signal input
flabel metal2 s 48962 0 49018 800 0 FreeSans 224 90 0 0 dso_as1802[10]
port 65 nsew signal input
flabel metal2 s 49238 0 49294 800 0 FreeSans 224 90 0 0 dso_as1802[11]
port 66 nsew signal input
flabel metal2 s 49514 0 49570 800 0 FreeSans 224 90 0 0 dso_as1802[12]
port 67 nsew signal input
flabel metal2 s 49790 0 49846 800 0 FreeSans 224 90 0 0 dso_as1802[13]
port 68 nsew signal input
flabel metal2 s 50066 0 50122 800 0 FreeSans 224 90 0 0 dso_as1802[14]
port 69 nsew signal input
flabel metal2 s 50342 0 50398 800 0 FreeSans 224 90 0 0 dso_as1802[15]
port 70 nsew signal input
flabel metal2 s 50618 0 50674 800 0 FreeSans 224 90 0 0 dso_as1802[16]
port 71 nsew signal input
flabel metal2 s 50894 0 50950 800 0 FreeSans 224 90 0 0 dso_as1802[17]
port 72 nsew signal input
flabel metal2 s 51170 0 51226 800 0 FreeSans 224 90 0 0 dso_as1802[18]
port 73 nsew signal input
flabel metal2 s 51446 0 51502 800 0 FreeSans 224 90 0 0 dso_as1802[19]
port 74 nsew signal input
flabel metal2 s 46478 0 46534 800 0 FreeSans 224 90 0 0 dso_as1802[1]
port 75 nsew signal input
flabel metal2 s 51722 0 51778 800 0 FreeSans 224 90 0 0 dso_as1802[20]
port 76 nsew signal input
flabel metal2 s 51998 0 52054 800 0 FreeSans 224 90 0 0 dso_as1802[21]
port 77 nsew signal input
flabel metal2 s 52274 0 52330 800 0 FreeSans 224 90 0 0 dso_as1802[22]
port 78 nsew signal input
flabel metal2 s 52550 0 52606 800 0 FreeSans 224 90 0 0 dso_as1802[23]
port 79 nsew signal input
flabel metal2 s 52826 0 52882 800 0 FreeSans 224 90 0 0 dso_as1802[24]
port 80 nsew signal input
flabel metal2 s 53102 0 53158 800 0 FreeSans 224 90 0 0 dso_as1802[25]
port 81 nsew signal input
flabel metal2 s 53378 0 53434 800 0 FreeSans 224 90 0 0 dso_as1802[26]
port 82 nsew signal input
flabel metal2 s 46754 0 46810 800 0 FreeSans 224 90 0 0 dso_as1802[2]
port 83 nsew signal input
flabel metal2 s 47030 0 47086 800 0 FreeSans 224 90 0 0 dso_as1802[3]
port 84 nsew signal input
flabel metal2 s 47306 0 47362 800 0 FreeSans 224 90 0 0 dso_as1802[4]
port 85 nsew signal input
flabel metal2 s 47582 0 47638 800 0 FreeSans 224 90 0 0 dso_as1802[5]
port 86 nsew signal input
flabel metal2 s 47858 0 47914 800 0 FreeSans 224 90 0 0 dso_as1802[6]
port 87 nsew signal input
flabel metal2 s 48134 0 48190 800 0 FreeSans 224 90 0 0 dso_as1802[7]
port 88 nsew signal input
flabel metal2 s 48410 0 48466 800 0 FreeSans 224 90 0 0 dso_as1802[8]
port 89 nsew signal input
flabel metal2 s 48686 0 48742 800 0 FreeSans 224 90 0 0 dso_as1802[9]
port 90 nsew signal input
flabel metal2 s 24122 59200 24178 60000 0 FreeSans 224 90 0 0 dso_as2650[0]
port 91 nsew signal input
flabel metal2 s 37002 59200 37058 60000 0 FreeSans 224 90 0 0 dso_as2650[10]
port 92 nsew signal input
flabel metal2 s 38290 59200 38346 60000 0 FreeSans 224 90 0 0 dso_as2650[11]
port 93 nsew signal input
flabel metal2 s 39578 59200 39634 60000 0 FreeSans 224 90 0 0 dso_as2650[12]
port 94 nsew signal input
flabel metal2 s 40866 59200 40922 60000 0 FreeSans 224 90 0 0 dso_as2650[13]
port 95 nsew signal input
flabel metal2 s 42154 59200 42210 60000 0 FreeSans 224 90 0 0 dso_as2650[14]
port 96 nsew signal input
flabel metal2 s 43442 59200 43498 60000 0 FreeSans 224 90 0 0 dso_as2650[15]
port 97 nsew signal input
flabel metal2 s 44730 59200 44786 60000 0 FreeSans 224 90 0 0 dso_as2650[16]
port 98 nsew signal input
flabel metal2 s 46018 59200 46074 60000 0 FreeSans 224 90 0 0 dso_as2650[17]
port 99 nsew signal input
flabel metal2 s 47306 59200 47362 60000 0 FreeSans 224 90 0 0 dso_as2650[18]
port 100 nsew signal input
flabel metal2 s 48594 59200 48650 60000 0 FreeSans 224 90 0 0 dso_as2650[19]
port 101 nsew signal input
flabel metal2 s 25410 59200 25466 60000 0 FreeSans 224 90 0 0 dso_as2650[1]
port 102 nsew signal input
flabel metal2 s 49882 59200 49938 60000 0 FreeSans 224 90 0 0 dso_as2650[20]
port 103 nsew signal input
flabel metal2 s 51170 59200 51226 60000 0 FreeSans 224 90 0 0 dso_as2650[21]
port 104 nsew signal input
flabel metal2 s 52458 59200 52514 60000 0 FreeSans 224 90 0 0 dso_as2650[22]
port 105 nsew signal input
flabel metal2 s 53746 59200 53802 60000 0 FreeSans 224 90 0 0 dso_as2650[23]
port 106 nsew signal input
flabel metal2 s 55034 59200 55090 60000 0 FreeSans 224 90 0 0 dso_as2650[24]
port 107 nsew signal input
flabel metal2 s 56322 59200 56378 60000 0 FreeSans 224 90 0 0 dso_as2650[25]
port 108 nsew signal input
flabel metal2 s 57610 59200 57666 60000 0 FreeSans 224 90 0 0 dso_as2650[26]
port 109 nsew signal input
flabel metal2 s 26698 59200 26754 60000 0 FreeSans 224 90 0 0 dso_as2650[2]
port 110 nsew signal input
flabel metal2 s 27986 59200 28042 60000 0 FreeSans 224 90 0 0 dso_as2650[3]
port 111 nsew signal input
flabel metal2 s 29274 59200 29330 60000 0 FreeSans 224 90 0 0 dso_as2650[4]
port 112 nsew signal input
flabel metal2 s 30562 59200 30618 60000 0 FreeSans 224 90 0 0 dso_as2650[5]
port 113 nsew signal input
flabel metal2 s 31850 59200 31906 60000 0 FreeSans 224 90 0 0 dso_as2650[6]
port 114 nsew signal input
flabel metal2 s 33138 59200 33194 60000 0 FreeSans 224 90 0 0 dso_as2650[7]
port 115 nsew signal input
flabel metal2 s 34426 59200 34482 60000 0 FreeSans 224 90 0 0 dso_as2650[8]
port 116 nsew signal input
flabel metal2 s 35714 59200 35770 60000 0 FreeSans 224 90 0 0 dso_as2650[9]
port 117 nsew signal input
flabel metal3 s 0 40536 800 40656 0 FreeSans 480 0 0 0 dso_as512512512[0]
port 118 nsew signal input
flabel metal3 s 0 45976 800 46096 0 FreeSans 480 0 0 0 dso_as512512512[10]
port 119 nsew signal input
flabel metal3 s 0 46520 800 46640 0 FreeSans 480 0 0 0 dso_as512512512[11]
port 120 nsew signal input
flabel metal3 s 0 47064 800 47184 0 FreeSans 480 0 0 0 dso_as512512512[12]
port 121 nsew signal input
flabel metal3 s 0 47608 800 47728 0 FreeSans 480 0 0 0 dso_as512512512[13]
port 122 nsew signal input
flabel metal3 s 0 48152 800 48272 0 FreeSans 480 0 0 0 dso_as512512512[14]
port 123 nsew signal input
flabel metal3 s 0 48696 800 48816 0 FreeSans 480 0 0 0 dso_as512512512[15]
port 124 nsew signal input
flabel metal3 s 0 49240 800 49360 0 FreeSans 480 0 0 0 dso_as512512512[16]
port 125 nsew signal input
flabel metal3 s 0 49784 800 49904 0 FreeSans 480 0 0 0 dso_as512512512[17]
port 126 nsew signal input
flabel metal3 s 0 50328 800 50448 0 FreeSans 480 0 0 0 dso_as512512512[18]
port 127 nsew signal input
flabel metal3 s 0 50872 800 50992 0 FreeSans 480 0 0 0 dso_as512512512[19]
port 128 nsew signal input
flabel metal3 s 0 41080 800 41200 0 FreeSans 480 0 0 0 dso_as512512512[1]
port 129 nsew signal input
flabel metal3 s 0 51416 800 51536 0 FreeSans 480 0 0 0 dso_as512512512[20]
port 130 nsew signal input
flabel metal3 s 0 51960 800 52080 0 FreeSans 480 0 0 0 dso_as512512512[21]
port 131 nsew signal input
flabel metal3 s 0 52504 800 52624 0 FreeSans 480 0 0 0 dso_as512512512[22]
port 132 nsew signal input
flabel metal3 s 0 53048 800 53168 0 FreeSans 480 0 0 0 dso_as512512512[23]
port 133 nsew signal input
flabel metal3 s 0 53592 800 53712 0 FreeSans 480 0 0 0 dso_as512512512[24]
port 134 nsew signal input
flabel metal3 s 0 54136 800 54256 0 FreeSans 480 0 0 0 dso_as512512512[25]
port 135 nsew signal input
flabel metal3 s 0 54680 800 54800 0 FreeSans 480 0 0 0 dso_as512512512[26]
port 136 nsew signal input
flabel metal3 s 0 55224 800 55344 0 FreeSans 480 0 0 0 dso_as512512512[27]
port 137 nsew signal input
flabel metal3 s 0 41624 800 41744 0 FreeSans 480 0 0 0 dso_as512512512[2]
port 138 nsew signal input
flabel metal3 s 0 42168 800 42288 0 FreeSans 480 0 0 0 dso_as512512512[3]
port 139 nsew signal input
flabel metal3 s 0 42712 800 42832 0 FreeSans 480 0 0 0 dso_as512512512[4]
port 140 nsew signal input
flabel metal3 s 0 43256 800 43376 0 FreeSans 480 0 0 0 dso_as512512512[5]
port 141 nsew signal input
flabel metal3 s 0 43800 800 43920 0 FreeSans 480 0 0 0 dso_as512512512[6]
port 142 nsew signal input
flabel metal3 s 0 44344 800 44464 0 FreeSans 480 0 0 0 dso_as512512512[7]
port 143 nsew signal input
flabel metal3 s 0 44888 800 45008 0 FreeSans 480 0 0 0 dso_as512512512[8]
port 144 nsew signal input
flabel metal3 s 0 45432 800 45552 0 FreeSans 480 0 0 0 dso_as512512512[9]
port 145 nsew signal input
flabel metal3 s 59200 47608 60000 47728 0 FreeSans 480 0 0 0 dso_as5401[0]
port 146 nsew signal input
flabel metal3 s 59200 51688 60000 51808 0 FreeSans 480 0 0 0 dso_as5401[10]
port 147 nsew signal input
flabel metal3 s 59200 52096 60000 52216 0 FreeSans 480 0 0 0 dso_as5401[11]
port 148 nsew signal input
flabel metal3 s 59200 52504 60000 52624 0 FreeSans 480 0 0 0 dso_as5401[12]
port 149 nsew signal input
flabel metal3 s 59200 52912 60000 53032 0 FreeSans 480 0 0 0 dso_as5401[13]
port 150 nsew signal input
flabel metal3 s 59200 53320 60000 53440 0 FreeSans 480 0 0 0 dso_as5401[14]
port 151 nsew signal input
flabel metal3 s 59200 53728 60000 53848 0 FreeSans 480 0 0 0 dso_as5401[15]
port 152 nsew signal input
flabel metal3 s 59200 54136 60000 54256 0 FreeSans 480 0 0 0 dso_as5401[16]
port 153 nsew signal input
flabel metal3 s 59200 54544 60000 54664 0 FreeSans 480 0 0 0 dso_as5401[17]
port 154 nsew signal input
flabel metal3 s 59200 54952 60000 55072 0 FreeSans 480 0 0 0 dso_as5401[18]
port 155 nsew signal input
flabel metal3 s 59200 55360 60000 55480 0 FreeSans 480 0 0 0 dso_as5401[19]
port 156 nsew signal input
flabel metal3 s 59200 48016 60000 48136 0 FreeSans 480 0 0 0 dso_as5401[1]
port 157 nsew signal input
flabel metal3 s 59200 55768 60000 55888 0 FreeSans 480 0 0 0 dso_as5401[20]
port 158 nsew signal input
flabel metal3 s 59200 56176 60000 56296 0 FreeSans 480 0 0 0 dso_as5401[21]
port 159 nsew signal input
flabel metal3 s 59200 56584 60000 56704 0 FreeSans 480 0 0 0 dso_as5401[22]
port 160 nsew signal input
flabel metal3 s 59200 56992 60000 57112 0 FreeSans 480 0 0 0 dso_as5401[23]
port 161 nsew signal input
flabel metal3 s 59200 57400 60000 57520 0 FreeSans 480 0 0 0 dso_as5401[24]
port 162 nsew signal input
flabel metal3 s 59200 57808 60000 57928 0 FreeSans 480 0 0 0 dso_as5401[25]
port 163 nsew signal input
flabel metal3 s 59200 58216 60000 58336 0 FreeSans 480 0 0 0 dso_as5401[26]
port 164 nsew signal input
flabel metal3 s 59200 48424 60000 48544 0 FreeSans 480 0 0 0 dso_as5401[2]
port 165 nsew signal input
flabel metal3 s 59200 48832 60000 48952 0 FreeSans 480 0 0 0 dso_as5401[3]
port 166 nsew signal input
flabel metal3 s 59200 49240 60000 49360 0 FreeSans 480 0 0 0 dso_as5401[4]
port 167 nsew signal input
flabel metal3 s 59200 49648 60000 49768 0 FreeSans 480 0 0 0 dso_as5401[5]
port 168 nsew signal input
flabel metal3 s 59200 50056 60000 50176 0 FreeSans 480 0 0 0 dso_as5401[6]
port 169 nsew signal input
flabel metal3 s 59200 50464 60000 50584 0 FreeSans 480 0 0 0 dso_as5401[7]
port 170 nsew signal input
flabel metal3 s 59200 50872 60000 50992 0 FreeSans 480 0 0 0 dso_as5401[8]
port 171 nsew signal input
flabel metal3 s 59200 51280 60000 51400 0 FreeSans 480 0 0 0 dso_as5401[9]
port 172 nsew signal input
flabel metal3 s 59200 42712 60000 42832 0 FreeSans 480 0 0 0 dso_counter[0]
port 173 nsew signal input
flabel metal3 s 59200 46792 60000 46912 0 FreeSans 480 0 0 0 dso_counter[10]
port 174 nsew signal input
flabel metal3 s 59200 47200 60000 47320 0 FreeSans 480 0 0 0 dso_counter[11]
port 175 nsew signal input
flabel metal3 s 59200 43120 60000 43240 0 FreeSans 480 0 0 0 dso_counter[1]
port 176 nsew signal input
flabel metal3 s 59200 43528 60000 43648 0 FreeSans 480 0 0 0 dso_counter[2]
port 177 nsew signal input
flabel metal3 s 59200 43936 60000 44056 0 FreeSans 480 0 0 0 dso_counter[3]
port 178 nsew signal input
flabel metal3 s 59200 44344 60000 44464 0 FreeSans 480 0 0 0 dso_counter[4]
port 179 nsew signal input
flabel metal3 s 59200 44752 60000 44872 0 FreeSans 480 0 0 0 dso_counter[5]
port 180 nsew signal input
flabel metal3 s 59200 45160 60000 45280 0 FreeSans 480 0 0 0 dso_counter[6]
port 181 nsew signal input
flabel metal3 s 59200 45568 60000 45688 0 FreeSans 480 0 0 0 dso_counter[7]
port 182 nsew signal input
flabel metal3 s 59200 45976 60000 46096 0 FreeSans 480 0 0 0 dso_counter[8]
port 183 nsew signal input
flabel metal3 s 59200 46384 60000 46504 0 FreeSans 480 0 0 0 dso_counter[9]
port 184 nsew signal input
flabel metal2 s 12530 59200 12586 60000 0 FreeSans 224 90 0 0 dso_diceroll[0]
port 185 nsew signal input
flabel metal2 s 13818 59200 13874 60000 0 FreeSans 224 90 0 0 dso_diceroll[1]
port 186 nsew signal input
flabel metal2 s 15106 59200 15162 60000 0 FreeSans 224 90 0 0 dso_diceroll[2]
port 187 nsew signal input
flabel metal2 s 16394 59200 16450 60000 0 FreeSans 224 90 0 0 dso_diceroll[3]
port 188 nsew signal input
flabel metal2 s 17682 59200 17738 60000 0 FreeSans 224 90 0 0 dso_diceroll[4]
port 189 nsew signal input
flabel metal2 s 18970 59200 19026 60000 0 FreeSans 224 90 0 0 dso_diceroll[5]
port 190 nsew signal input
flabel metal2 s 20258 59200 20314 60000 0 FreeSans 224 90 0 0 dso_diceroll[6]
port 191 nsew signal input
flabel metal2 s 21546 59200 21602 60000 0 FreeSans 224 90 0 0 dso_diceroll[7]
port 192 nsew signal input
flabel metal3 s 0 30744 800 30864 0 FreeSans 480 0 0 0 dso_mc14500[0]
port 193 nsew signal input
flabel metal3 s 0 31288 800 31408 0 FreeSans 480 0 0 0 dso_mc14500[1]
port 194 nsew signal input
flabel metal3 s 0 31832 800 31952 0 FreeSans 480 0 0 0 dso_mc14500[2]
port 195 nsew signal input
flabel metal3 s 0 32376 800 32496 0 FreeSans 480 0 0 0 dso_mc14500[3]
port 196 nsew signal input
flabel metal3 s 0 32920 800 33040 0 FreeSans 480 0 0 0 dso_mc14500[4]
port 197 nsew signal input
flabel metal3 s 0 33464 800 33584 0 FreeSans 480 0 0 0 dso_mc14500[5]
port 198 nsew signal input
flabel metal3 s 0 34008 800 34128 0 FreeSans 480 0 0 0 dso_mc14500[6]
port 199 nsew signal input
flabel metal3 s 0 34552 800 34672 0 FreeSans 480 0 0 0 dso_mc14500[7]
port 200 nsew signal input
flabel metal3 s 0 35096 800 35216 0 FreeSans 480 0 0 0 dso_mc14500[8]
port 201 nsew signal input
flabel metal2 s 2226 59200 2282 60000 0 FreeSans 224 90 0 0 dso_multiplier[0]
port 202 nsew signal input
flabel metal2 s 3514 59200 3570 60000 0 FreeSans 224 90 0 0 dso_multiplier[1]
port 203 nsew signal input
flabel metal2 s 4802 59200 4858 60000 0 FreeSans 224 90 0 0 dso_multiplier[2]
port 204 nsew signal input
flabel metal2 s 6090 59200 6146 60000 0 FreeSans 224 90 0 0 dso_multiplier[3]
port 205 nsew signal input
flabel metal2 s 7378 59200 7434 60000 0 FreeSans 224 90 0 0 dso_multiplier[4]
port 206 nsew signal input
flabel metal2 s 8666 59200 8722 60000 0 FreeSans 224 90 0 0 dso_multiplier[5]
port 207 nsew signal input
flabel metal2 s 9954 59200 10010 60000 0 FreeSans 224 90 0 0 dso_multiplier[6]
port 208 nsew signal input
flabel metal2 s 11242 59200 11298 60000 0 FreeSans 224 90 0 0 dso_multiplier[7]
port 209 nsew signal input
flabel metal2 s 37370 0 37426 800 0 FreeSans 224 90 0 0 dso_posit[0]
port 210 nsew signal input
flabel metal2 s 37646 0 37702 800 0 FreeSans 224 90 0 0 dso_posit[1]
port 211 nsew signal input
flabel metal2 s 37922 0 37978 800 0 FreeSans 224 90 0 0 dso_posit[2]
port 212 nsew signal input
flabel metal2 s 38198 0 38254 800 0 FreeSans 224 90 0 0 dso_posit[3]
port 213 nsew signal input
flabel metal3 s 0 36184 800 36304 0 FreeSans 480 0 0 0 dso_tbb1143[0]
port 214 nsew signal input
flabel metal3 s 0 36728 800 36848 0 FreeSans 480 0 0 0 dso_tbb1143[1]
port 215 nsew signal input
flabel metal3 s 0 37272 800 37392 0 FreeSans 480 0 0 0 dso_tbb1143[2]
port 216 nsew signal input
flabel metal3 s 0 37816 800 37936 0 FreeSans 480 0 0 0 dso_tbb1143[3]
port 217 nsew signal input
flabel metal3 s 0 38360 800 38480 0 FreeSans 480 0 0 0 dso_tbb1143[4]
port 218 nsew signal input
flabel metal3 s 0 38904 800 39024 0 FreeSans 480 0 0 0 dso_tbb1143[5]
port 219 nsew signal input
flabel metal3 s 0 39448 800 39568 0 FreeSans 480 0 0 0 dso_tbb1143[6]
port 220 nsew signal input
flabel metal3 s 0 39992 800 40112 0 FreeSans 480 0 0 0 dso_tbb1143[7]
port 221 nsew signal input
flabel metal2 s 53930 0 53986 800 0 FreeSans 224 90 0 0 dso_tune
port 222 nsew signal input
flabel metal2 s 5906 0 5962 800 0 FreeSans 224 90 0 0 io_in[0]
port 223 nsew signal input
flabel metal2 s 8666 0 8722 800 0 FreeSans 224 90 0 0 io_in[10]
port 224 nsew signal input
flabel metal2 s 8942 0 8998 800 0 FreeSans 224 90 0 0 io_in[11]
port 225 nsew signal input
flabel metal2 s 9218 0 9274 800 0 FreeSans 224 90 0 0 io_in[12]
port 226 nsew signal input
flabel metal2 s 9494 0 9550 800 0 FreeSans 224 90 0 0 io_in[13]
port 227 nsew signal input
flabel metal2 s 9770 0 9826 800 0 FreeSans 224 90 0 0 io_in[14]
port 228 nsew signal input
flabel metal2 s 10046 0 10102 800 0 FreeSans 224 90 0 0 io_in[15]
port 229 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 io_in[16]
port 230 nsew signal input
flabel metal2 s 10598 0 10654 800 0 FreeSans 224 90 0 0 io_in[17]
port 231 nsew signal input
flabel metal2 s 10874 0 10930 800 0 FreeSans 224 90 0 0 io_in[18]
port 232 nsew signal input
flabel metal2 s 11150 0 11206 800 0 FreeSans 224 90 0 0 io_in[19]
port 233 nsew signal input
flabel metal2 s 6182 0 6238 800 0 FreeSans 224 90 0 0 io_in[1]
port 234 nsew signal input
flabel metal2 s 11426 0 11482 800 0 FreeSans 224 90 0 0 io_in[20]
port 235 nsew signal input
flabel metal2 s 11702 0 11758 800 0 FreeSans 224 90 0 0 io_in[21]
port 236 nsew signal input
flabel metal2 s 11978 0 12034 800 0 FreeSans 224 90 0 0 io_in[22]
port 237 nsew signal input
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 io_in[23]
port 238 nsew signal input
flabel metal2 s 12530 0 12586 800 0 FreeSans 224 90 0 0 io_in[24]
port 239 nsew signal input
flabel metal2 s 12806 0 12862 800 0 FreeSans 224 90 0 0 io_in[25]
port 240 nsew signal input
flabel metal2 s 13082 0 13138 800 0 FreeSans 224 90 0 0 io_in[26]
port 241 nsew signal input
flabel metal2 s 13358 0 13414 800 0 FreeSans 224 90 0 0 io_in[27]
port 242 nsew signal input
flabel metal2 s 13634 0 13690 800 0 FreeSans 224 90 0 0 io_in[28]
port 243 nsew signal input
flabel metal2 s 13910 0 13966 800 0 FreeSans 224 90 0 0 io_in[29]
port 244 nsew signal input
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 io_in[2]
port 245 nsew signal input
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 io_in[30]
port 246 nsew signal input
flabel metal2 s 14462 0 14518 800 0 FreeSans 224 90 0 0 io_in[31]
port 247 nsew signal input
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 io_in[32]
port 248 nsew signal input
flabel metal2 s 15014 0 15070 800 0 FreeSans 224 90 0 0 io_in[33]
port 249 nsew signal input
flabel metal2 s 15290 0 15346 800 0 FreeSans 224 90 0 0 io_in[34]
port 250 nsew signal input
flabel metal2 s 15566 0 15622 800 0 FreeSans 224 90 0 0 io_in[35]
port 251 nsew signal input
flabel metal2 s 15842 0 15898 800 0 FreeSans 224 90 0 0 io_in[36]
port 252 nsew signal input
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 io_in[37]
port 253 nsew signal input
flabel metal2 s 6734 0 6790 800 0 FreeSans 224 90 0 0 io_in[3]
port 254 nsew signal input
flabel metal2 s 7010 0 7066 800 0 FreeSans 224 90 0 0 io_in[4]
port 255 nsew signal input
flabel metal2 s 7286 0 7342 800 0 FreeSans 224 90 0 0 io_in[5]
port 256 nsew signal input
flabel metal2 s 7562 0 7618 800 0 FreeSans 224 90 0 0 io_in[6]
port 257 nsew signal input
flabel metal2 s 7838 0 7894 800 0 FreeSans 224 90 0 0 io_in[7]
port 258 nsew signal input
flabel metal2 s 8114 0 8170 800 0 FreeSans 224 90 0 0 io_in[8]
port 259 nsew signal input
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 io_in[9]
port 260 nsew signal input
flabel metal2 s 26882 0 26938 800 0 FreeSans 224 90 0 0 io_oeb[0]
port 261 nsew signal tristate
flabel metal2 s 29642 0 29698 800 0 FreeSans 224 90 0 0 io_oeb[10]
port 262 nsew signal tristate
flabel metal2 s 29918 0 29974 800 0 FreeSans 224 90 0 0 io_oeb[11]
port 263 nsew signal tristate
flabel metal2 s 30194 0 30250 800 0 FreeSans 224 90 0 0 io_oeb[12]
port 264 nsew signal tristate
flabel metal2 s 30470 0 30526 800 0 FreeSans 224 90 0 0 io_oeb[13]
port 265 nsew signal tristate
flabel metal2 s 30746 0 30802 800 0 FreeSans 224 90 0 0 io_oeb[14]
port 266 nsew signal tristate
flabel metal2 s 31022 0 31078 800 0 FreeSans 224 90 0 0 io_oeb[15]
port 267 nsew signal tristate
flabel metal2 s 31298 0 31354 800 0 FreeSans 224 90 0 0 io_oeb[16]
port 268 nsew signal tristate
flabel metal2 s 31574 0 31630 800 0 FreeSans 224 90 0 0 io_oeb[17]
port 269 nsew signal tristate
flabel metal2 s 31850 0 31906 800 0 FreeSans 224 90 0 0 io_oeb[18]
port 270 nsew signal tristate
flabel metal2 s 32126 0 32182 800 0 FreeSans 224 90 0 0 io_oeb[19]
port 271 nsew signal tristate
flabel metal2 s 27158 0 27214 800 0 FreeSans 224 90 0 0 io_oeb[1]
port 272 nsew signal tristate
flabel metal2 s 32402 0 32458 800 0 FreeSans 224 90 0 0 io_oeb[20]
port 273 nsew signal tristate
flabel metal2 s 32678 0 32734 800 0 FreeSans 224 90 0 0 io_oeb[21]
port 274 nsew signal tristate
flabel metal2 s 32954 0 33010 800 0 FreeSans 224 90 0 0 io_oeb[22]
port 275 nsew signal tristate
flabel metal2 s 33230 0 33286 800 0 FreeSans 224 90 0 0 io_oeb[23]
port 276 nsew signal tristate
flabel metal2 s 33506 0 33562 800 0 FreeSans 224 90 0 0 io_oeb[24]
port 277 nsew signal tristate
flabel metal2 s 33782 0 33838 800 0 FreeSans 224 90 0 0 io_oeb[25]
port 278 nsew signal tristate
flabel metal2 s 34058 0 34114 800 0 FreeSans 224 90 0 0 io_oeb[26]
port 279 nsew signal tristate
flabel metal2 s 34334 0 34390 800 0 FreeSans 224 90 0 0 io_oeb[27]
port 280 nsew signal tristate
flabel metal2 s 34610 0 34666 800 0 FreeSans 224 90 0 0 io_oeb[28]
port 281 nsew signal tristate
flabel metal2 s 34886 0 34942 800 0 FreeSans 224 90 0 0 io_oeb[29]
port 282 nsew signal tristate
flabel metal2 s 27434 0 27490 800 0 FreeSans 224 90 0 0 io_oeb[2]
port 283 nsew signal tristate
flabel metal2 s 35162 0 35218 800 0 FreeSans 224 90 0 0 io_oeb[30]
port 284 nsew signal tristate
flabel metal2 s 35438 0 35494 800 0 FreeSans 224 90 0 0 io_oeb[31]
port 285 nsew signal tristate
flabel metal2 s 35714 0 35770 800 0 FreeSans 224 90 0 0 io_oeb[32]
port 286 nsew signal tristate
flabel metal2 s 35990 0 36046 800 0 FreeSans 224 90 0 0 io_oeb[33]
port 287 nsew signal tristate
flabel metal2 s 36266 0 36322 800 0 FreeSans 224 90 0 0 io_oeb[34]
port 288 nsew signal tristate
flabel metal2 s 36542 0 36598 800 0 FreeSans 224 90 0 0 io_oeb[35]
port 289 nsew signal tristate
flabel metal2 s 36818 0 36874 800 0 FreeSans 224 90 0 0 io_oeb[36]
port 290 nsew signal tristate
flabel metal2 s 37094 0 37150 800 0 FreeSans 224 90 0 0 io_oeb[37]
port 291 nsew signal tristate
flabel metal2 s 27710 0 27766 800 0 FreeSans 224 90 0 0 io_oeb[3]
port 292 nsew signal tristate
flabel metal2 s 27986 0 28042 800 0 FreeSans 224 90 0 0 io_oeb[4]
port 293 nsew signal tristate
flabel metal2 s 28262 0 28318 800 0 FreeSans 224 90 0 0 io_oeb[5]
port 294 nsew signal tristate
flabel metal2 s 28538 0 28594 800 0 FreeSans 224 90 0 0 io_oeb[6]
port 295 nsew signal tristate
flabel metal2 s 28814 0 28870 800 0 FreeSans 224 90 0 0 io_oeb[7]
port 296 nsew signal tristate
flabel metal2 s 29090 0 29146 800 0 FreeSans 224 90 0 0 io_oeb[8]
port 297 nsew signal tristate
flabel metal2 s 29366 0 29422 800 0 FreeSans 224 90 0 0 io_oeb[9]
port 298 nsew signal tristate
flabel metal2 s 16394 0 16450 800 0 FreeSans 224 90 0 0 io_out[0]
port 299 nsew signal tristate
flabel metal2 s 19154 0 19210 800 0 FreeSans 224 90 0 0 io_out[10]
port 300 nsew signal tristate
flabel metal2 s 19430 0 19486 800 0 FreeSans 224 90 0 0 io_out[11]
port 301 nsew signal tristate
flabel metal2 s 19706 0 19762 800 0 FreeSans 224 90 0 0 io_out[12]
port 302 nsew signal tristate
flabel metal2 s 19982 0 20038 800 0 FreeSans 224 90 0 0 io_out[13]
port 303 nsew signal tristate
flabel metal2 s 20258 0 20314 800 0 FreeSans 224 90 0 0 io_out[14]
port 304 nsew signal tristate
flabel metal2 s 20534 0 20590 800 0 FreeSans 224 90 0 0 io_out[15]
port 305 nsew signal tristate
flabel metal2 s 20810 0 20866 800 0 FreeSans 224 90 0 0 io_out[16]
port 306 nsew signal tristate
flabel metal2 s 21086 0 21142 800 0 FreeSans 224 90 0 0 io_out[17]
port 307 nsew signal tristate
flabel metal2 s 21362 0 21418 800 0 FreeSans 224 90 0 0 io_out[18]
port 308 nsew signal tristate
flabel metal2 s 21638 0 21694 800 0 FreeSans 224 90 0 0 io_out[19]
port 309 nsew signal tristate
flabel metal2 s 16670 0 16726 800 0 FreeSans 224 90 0 0 io_out[1]
port 310 nsew signal tristate
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 io_out[20]
port 311 nsew signal tristate
flabel metal2 s 22190 0 22246 800 0 FreeSans 224 90 0 0 io_out[21]
port 312 nsew signal tristate
flabel metal2 s 22466 0 22522 800 0 FreeSans 224 90 0 0 io_out[22]
port 313 nsew signal tristate
flabel metal2 s 22742 0 22798 800 0 FreeSans 224 90 0 0 io_out[23]
port 314 nsew signal tristate
flabel metal2 s 23018 0 23074 800 0 FreeSans 224 90 0 0 io_out[24]
port 315 nsew signal tristate
flabel metal2 s 23294 0 23350 800 0 FreeSans 224 90 0 0 io_out[25]
port 316 nsew signal tristate
flabel metal2 s 23570 0 23626 800 0 FreeSans 224 90 0 0 io_out[26]
port 317 nsew signal tristate
flabel metal2 s 23846 0 23902 800 0 FreeSans 224 90 0 0 io_out[27]
port 318 nsew signal tristate
flabel metal2 s 24122 0 24178 800 0 FreeSans 224 90 0 0 io_out[28]
port 319 nsew signal tristate
flabel metal2 s 24398 0 24454 800 0 FreeSans 224 90 0 0 io_out[29]
port 320 nsew signal tristate
flabel metal2 s 16946 0 17002 800 0 FreeSans 224 90 0 0 io_out[2]
port 321 nsew signal tristate
flabel metal2 s 24674 0 24730 800 0 FreeSans 224 90 0 0 io_out[30]
port 322 nsew signal tristate
flabel metal2 s 24950 0 25006 800 0 FreeSans 224 90 0 0 io_out[31]
port 323 nsew signal tristate
flabel metal2 s 25226 0 25282 800 0 FreeSans 224 90 0 0 io_out[32]
port 324 nsew signal tristate
flabel metal2 s 25502 0 25558 800 0 FreeSans 224 90 0 0 io_out[33]
port 325 nsew signal tristate
flabel metal2 s 25778 0 25834 800 0 FreeSans 224 90 0 0 io_out[34]
port 326 nsew signal tristate
flabel metal2 s 26054 0 26110 800 0 FreeSans 224 90 0 0 io_out[35]
port 327 nsew signal tristate
flabel metal2 s 26330 0 26386 800 0 FreeSans 224 90 0 0 io_out[36]
port 328 nsew signal tristate
flabel metal2 s 26606 0 26662 800 0 FreeSans 224 90 0 0 io_out[37]
port 329 nsew signal tristate
flabel metal2 s 17222 0 17278 800 0 FreeSans 224 90 0 0 io_out[3]
port 330 nsew signal tristate
flabel metal2 s 17498 0 17554 800 0 FreeSans 224 90 0 0 io_out[4]
port 331 nsew signal tristate
flabel metal2 s 17774 0 17830 800 0 FreeSans 224 90 0 0 io_out[5]
port 332 nsew signal tristate
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 io_out[6]
port 333 nsew signal tristate
flabel metal2 s 18326 0 18382 800 0 FreeSans 224 90 0 0 io_out[7]
port 334 nsew signal tristate
flabel metal2 s 18602 0 18658 800 0 FreeSans 224 90 0 0 io_out[8]
port 335 nsew signal tristate
flabel metal2 s 18878 0 18934 800 0 FreeSans 224 90 0 0 io_out[9]
port 336 nsew signal tristate
flabel metal2 s 38474 0 38530 800 0 FreeSans 224 90 0 0 oeb_6502
port 337 nsew signal input
flabel metal2 s 53654 0 53710 800 0 FreeSans 224 90 0 0 oeb_as1802
port 338 nsew signal input
flabel metal2 s 22834 59200 22890 60000 0 FreeSans 224 90 0 0 oeb_as2650
port 339 nsew signal input
flabel metal3 s 0 55768 800 55888 0 FreeSans 480 0 0 0 oeb_as512512512
port 340 nsew signal input
flabel metal3 s 59200 58624 60000 58744 0 FreeSans 480 0 0 0 oeb_as5401
port 341 nsew signal input
flabel metal3 s 0 35640 800 35760 0 FreeSans 480 0 0 0 oeb_mc14500
port 342 nsew signal input
flabel metal3 s 0 19864 800 19984 0 FreeSans 480 0 0 0 rst_6502
port 343 nsew signal tristate
flabel metal3 s 0 20408 800 20528 0 FreeSans 480 0 0 0 rst_LCD
port 344 nsew signal tristate
flabel metal3 s 0 20952 800 21072 0 FreeSans 480 0 0 0 rst_as1802
port 345 nsew signal tristate
flabel metal3 s 0 21496 800 21616 0 FreeSans 480 0 0 0 rst_as2650
port 346 nsew signal tristate
flabel metal3 s 0 22584 800 22704 0 FreeSans 480 0 0 0 rst_as512512512
port 347 nsew signal tristate
flabel metal3 s 0 22040 800 22160 0 FreeSans 480 0 0 0 rst_as5401
port 348 nsew signal tristate
flabel metal3 s 0 23128 800 23248 0 FreeSans 480 0 0 0 rst_counter
port 349 nsew signal tristate
flabel metal3 s 0 23672 800 23792 0 FreeSans 480 0 0 0 rst_diceroll
port 350 nsew signal tristate
flabel metal3 s 0 24216 800 24336 0 FreeSans 480 0 0 0 rst_mc14500
port 351 nsew signal tristate
flabel metal3 s 0 24760 800 24880 0 FreeSans 480 0 0 0 rst_posit
port 352 nsew signal tristate
flabel metal3 s 0 25304 800 25424 0 FreeSans 480 0 0 0 rst_tbb1143
port 353 nsew signal tristate
flabel metal3 s 0 25848 800 25968 0 FreeSans 480 0 0 0 rst_tune
port 354 nsew signal tristate
flabel metal4 s 4208 2128 4528 57712 0 FreeSans 1920 90 0 0 vccd1
port 355 nsew power bidirectional
flabel metal4 s 34928 2128 35248 57712 0 FreeSans 1920 90 0 0 vccd1
port 355 nsew power bidirectional
flabel metal4 s 19568 2128 19888 57712 0 FreeSans 1920 90 0 0 vssd1
port 356 nsew ground bidirectional
flabel metal4 s 50288 2128 50608 57712 0 FreeSans 1920 90 0 0 vssd1
port 356 nsew ground bidirectional
flabel metal3 s 59200 1096 60000 1216 0 FreeSans 480 0 0 0 wb_clk_i
port 357 nsew signal input
flabel metal3 s 59200 1504 60000 1624 0 FreeSans 480 0 0 0 wb_rst_i
port 358 nsew signal input
flabel metal3 s 59200 1912 60000 2032 0 FreeSans 480 0 0 0 wbs_ack_o
port 359 nsew signal tristate
flabel metal3 s 59200 3544 60000 3664 0 FreeSans 480 0 0 0 wbs_adr_i[0]
port 360 nsew signal input
flabel metal3 s 59200 15784 60000 15904 0 FreeSans 480 0 0 0 wbs_adr_i[10]
port 361 nsew signal input
flabel metal3 s 59200 17008 60000 17128 0 FreeSans 480 0 0 0 wbs_adr_i[11]
port 362 nsew signal input
flabel metal3 s 59200 18232 60000 18352 0 FreeSans 480 0 0 0 wbs_adr_i[12]
port 363 nsew signal input
flabel metal3 s 59200 19456 60000 19576 0 FreeSans 480 0 0 0 wbs_adr_i[13]
port 364 nsew signal input
flabel metal3 s 59200 20680 60000 20800 0 FreeSans 480 0 0 0 wbs_adr_i[14]
port 365 nsew signal input
flabel metal3 s 59200 21904 60000 22024 0 FreeSans 480 0 0 0 wbs_adr_i[15]
port 366 nsew signal input
flabel metal3 s 59200 23128 60000 23248 0 FreeSans 480 0 0 0 wbs_adr_i[16]
port 367 nsew signal input
flabel metal3 s 59200 24352 60000 24472 0 FreeSans 480 0 0 0 wbs_adr_i[17]
port 368 nsew signal input
flabel metal3 s 59200 25576 60000 25696 0 FreeSans 480 0 0 0 wbs_adr_i[18]
port 369 nsew signal input
flabel metal3 s 59200 26800 60000 26920 0 FreeSans 480 0 0 0 wbs_adr_i[19]
port 370 nsew signal input
flabel metal3 s 59200 4768 60000 4888 0 FreeSans 480 0 0 0 wbs_adr_i[1]
port 371 nsew signal input
flabel metal3 s 59200 28024 60000 28144 0 FreeSans 480 0 0 0 wbs_adr_i[20]
port 372 nsew signal input
flabel metal3 s 59200 29248 60000 29368 0 FreeSans 480 0 0 0 wbs_adr_i[21]
port 373 nsew signal input
flabel metal3 s 59200 30472 60000 30592 0 FreeSans 480 0 0 0 wbs_adr_i[22]
port 374 nsew signal input
flabel metal3 s 59200 31696 60000 31816 0 FreeSans 480 0 0 0 wbs_adr_i[23]
port 375 nsew signal input
flabel metal3 s 59200 32920 60000 33040 0 FreeSans 480 0 0 0 wbs_adr_i[24]
port 376 nsew signal input
flabel metal3 s 59200 34144 60000 34264 0 FreeSans 480 0 0 0 wbs_adr_i[25]
port 377 nsew signal input
flabel metal3 s 59200 35368 60000 35488 0 FreeSans 480 0 0 0 wbs_adr_i[26]
port 378 nsew signal input
flabel metal3 s 59200 36592 60000 36712 0 FreeSans 480 0 0 0 wbs_adr_i[27]
port 379 nsew signal input
flabel metal3 s 59200 37816 60000 37936 0 FreeSans 480 0 0 0 wbs_adr_i[28]
port 380 nsew signal input
flabel metal3 s 59200 39040 60000 39160 0 FreeSans 480 0 0 0 wbs_adr_i[29]
port 381 nsew signal input
flabel metal3 s 59200 5992 60000 6112 0 FreeSans 480 0 0 0 wbs_adr_i[2]
port 382 nsew signal input
flabel metal3 s 59200 40264 60000 40384 0 FreeSans 480 0 0 0 wbs_adr_i[30]
port 383 nsew signal input
flabel metal3 s 59200 41488 60000 41608 0 FreeSans 480 0 0 0 wbs_adr_i[31]
port 384 nsew signal input
flabel metal3 s 59200 7216 60000 7336 0 FreeSans 480 0 0 0 wbs_adr_i[3]
port 385 nsew signal input
flabel metal3 s 59200 8440 60000 8560 0 FreeSans 480 0 0 0 wbs_adr_i[4]
port 386 nsew signal input
flabel metal3 s 59200 9664 60000 9784 0 FreeSans 480 0 0 0 wbs_adr_i[5]
port 387 nsew signal input
flabel metal3 s 59200 10888 60000 11008 0 FreeSans 480 0 0 0 wbs_adr_i[6]
port 388 nsew signal input
flabel metal3 s 59200 12112 60000 12232 0 FreeSans 480 0 0 0 wbs_adr_i[7]
port 389 nsew signal input
flabel metal3 s 59200 13336 60000 13456 0 FreeSans 480 0 0 0 wbs_adr_i[8]
port 390 nsew signal input
flabel metal3 s 59200 14560 60000 14680 0 FreeSans 480 0 0 0 wbs_adr_i[9]
port 391 nsew signal input
flabel metal3 s 59200 2320 60000 2440 0 FreeSans 480 0 0 0 wbs_cyc_i
port 392 nsew signal input
flabel metal3 s 59200 3952 60000 4072 0 FreeSans 480 0 0 0 wbs_dat_i[0]
port 393 nsew signal input
flabel metal3 s 59200 16192 60000 16312 0 FreeSans 480 0 0 0 wbs_dat_i[10]
port 394 nsew signal input
flabel metal3 s 59200 17416 60000 17536 0 FreeSans 480 0 0 0 wbs_dat_i[11]
port 395 nsew signal input
flabel metal3 s 59200 18640 60000 18760 0 FreeSans 480 0 0 0 wbs_dat_i[12]
port 396 nsew signal input
flabel metal3 s 59200 19864 60000 19984 0 FreeSans 480 0 0 0 wbs_dat_i[13]
port 397 nsew signal input
flabel metal3 s 59200 21088 60000 21208 0 FreeSans 480 0 0 0 wbs_dat_i[14]
port 398 nsew signal input
flabel metal3 s 59200 22312 60000 22432 0 FreeSans 480 0 0 0 wbs_dat_i[15]
port 399 nsew signal input
flabel metal3 s 59200 23536 60000 23656 0 FreeSans 480 0 0 0 wbs_dat_i[16]
port 400 nsew signal input
flabel metal3 s 59200 24760 60000 24880 0 FreeSans 480 0 0 0 wbs_dat_i[17]
port 401 nsew signal input
flabel metal3 s 59200 25984 60000 26104 0 FreeSans 480 0 0 0 wbs_dat_i[18]
port 402 nsew signal input
flabel metal3 s 59200 27208 60000 27328 0 FreeSans 480 0 0 0 wbs_dat_i[19]
port 403 nsew signal input
flabel metal3 s 59200 5176 60000 5296 0 FreeSans 480 0 0 0 wbs_dat_i[1]
port 404 nsew signal input
flabel metal3 s 59200 28432 60000 28552 0 FreeSans 480 0 0 0 wbs_dat_i[20]
port 405 nsew signal input
flabel metal3 s 59200 29656 60000 29776 0 FreeSans 480 0 0 0 wbs_dat_i[21]
port 406 nsew signal input
flabel metal3 s 59200 30880 60000 31000 0 FreeSans 480 0 0 0 wbs_dat_i[22]
port 407 nsew signal input
flabel metal3 s 59200 32104 60000 32224 0 FreeSans 480 0 0 0 wbs_dat_i[23]
port 408 nsew signal input
flabel metal3 s 59200 33328 60000 33448 0 FreeSans 480 0 0 0 wbs_dat_i[24]
port 409 nsew signal input
flabel metal3 s 59200 34552 60000 34672 0 FreeSans 480 0 0 0 wbs_dat_i[25]
port 410 nsew signal input
flabel metal3 s 59200 35776 60000 35896 0 FreeSans 480 0 0 0 wbs_dat_i[26]
port 411 nsew signal input
flabel metal3 s 59200 37000 60000 37120 0 FreeSans 480 0 0 0 wbs_dat_i[27]
port 412 nsew signal input
flabel metal3 s 59200 38224 60000 38344 0 FreeSans 480 0 0 0 wbs_dat_i[28]
port 413 nsew signal input
flabel metal3 s 59200 39448 60000 39568 0 FreeSans 480 0 0 0 wbs_dat_i[29]
port 414 nsew signal input
flabel metal3 s 59200 6400 60000 6520 0 FreeSans 480 0 0 0 wbs_dat_i[2]
port 415 nsew signal input
flabel metal3 s 59200 40672 60000 40792 0 FreeSans 480 0 0 0 wbs_dat_i[30]
port 416 nsew signal input
flabel metal3 s 59200 41896 60000 42016 0 FreeSans 480 0 0 0 wbs_dat_i[31]
port 417 nsew signal input
flabel metal3 s 59200 7624 60000 7744 0 FreeSans 480 0 0 0 wbs_dat_i[3]
port 418 nsew signal input
flabel metal3 s 59200 8848 60000 8968 0 FreeSans 480 0 0 0 wbs_dat_i[4]
port 419 nsew signal input
flabel metal3 s 59200 10072 60000 10192 0 FreeSans 480 0 0 0 wbs_dat_i[5]
port 420 nsew signal input
flabel metal3 s 59200 11296 60000 11416 0 FreeSans 480 0 0 0 wbs_dat_i[6]
port 421 nsew signal input
flabel metal3 s 59200 12520 60000 12640 0 FreeSans 480 0 0 0 wbs_dat_i[7]
port 422 nsew signal input
flabel metal3 s 59200 13744 60000 13864 0 FreeSans 480 0 0 0 wbs_dat_i[8]
port 423 nsew signal input
flabel metal3 s 59200 14968 60000 15088 0 FreeSans 480 0 0 0 wbs_dat_i[9]
port 424 nsew signal input
flabel metal3 s 59200 4360 60000 4480 0 FreeSans 480 0 0 0 wbs_dat_o[0]
port 425 nsew signal tristate
flabel metal3 s 59200 16600 60000 16720 0 FreeSans 480 0 0 0 wbs_dat_o[10]
port 426 nsew signal tristate
flabel metal3 s 59200 17824 60000 17944 0 FreeSans 480 0 0 0 wbs_dat_o[11]
port 427 nsew signal tristate
flabel metal3 s 59200 19048 60000 19168 0 FreeSans 480 0 0 0 wbs_dat_o[12]
port 428 nsew signal tristate
flabel metal3 s 59200 20272 60000 20392 0 FreeSans 480 0 0 0 wbs_dat_o[13]
port 429 nsew signal tristate
flabel metal3 s 59200 21496 60000 21616 0 FreeSans 480 0 0 0 wbs_dat_o[14]
port 430 nsew signal tristate
flabel metal3 s 59200 22720 60000 22840 0 FreeSans 480 0 0 0 wbs_dat_o[15]
port 431 nsew signal tristate
flabel metal3 s 59200 23944 60000 24064 0 FreeSans 480 0 0 0 wbs_dat_o[16]
port 432 nsew signal tristate
flabel metal3 s 59200 25168 60000 25288 0 FreeSans 480 0 0 0 wbs_dat_o[17]
port 433 nsew signal tristate
flabel metal3 s 59200 26392 60000 26512 0 FreeSans 480 0 0 0 wbs_dat_o[18]
port 434 nsew signal tristate
flabel metal3 s 59200 27616 60000 27736 0 FreeSans 480 0 0 0 wbs_dat_o[19]
port 435 nsew signal tristate
flabel metal3 s 59200 5584 60000 5704 0 FreeSans 480 0 0 0 wbs_dat_o[1]
port 436 nsew signal tristate
flabel metal3 s 59200 28840 60000 28960 0 FreeSans 480 0 0 0 wbs_dat_o[20]
port 437 nsew signal tristate
flabel metal3 s 59200 30064 60000 30184 0 FreeSans 480 0 0 0 wbs_dat_o[21]
port 438 nsew signal tristate
flabel metal3 s 59200 31288 60000 31408 0 FreeSans 480 0 0 0 wbs_dat_o[22]
port 439 nsew signal tristate
flabel metal3 s 59200 32512 60000 32632 0 FreeSans 480 0 0 0 wbs_dat_o[23]
port 440 nsew signal tristate
flabel metal3 s 59200 33736 60000 33856 0 FreeSans 480 0 0 0 wbs_dat_o[24]
port 441 nsew signal tristate
flabel metal3 s 59200 34960 60000 35080 0 FreeSans 480 0 0 0 wbs_dat_o[25]
port 442 nsew signal tristate
flabel metal3 s 59200 36184 60000 36304 0 FreeSans 480 0 0 0 wbs_dat_o[26]
port 443 nsew signal tristate
flabel metal3 s 59200 37408 60000 37528 0 FreeSans 480 0 0 0 wbs_dat_o[27]
port 444 nsew signal tristate
flabel metal3 s 59200 38632 60000 38752 0 FreeSans 480 0 0 0 wbs_dat_o[28]
port 445 nsew signal tristate
flabel metal3 s 59200 39856 60000 39976 0 FreeSans 480 0 0 0 wbs_dat_o[29]
port 446 nsew signal tristate
flabel metal3 s 59200 6808 60000 6928 0 FreeSans 480 0 0 0 wbs_dat_o[2]
port 447 nsew signal tristate
flabel metal3 s 59200 41080 60000 41200 0 FreeSans 480 0 0 0 wbs_dat_o[30]
port 448 nsew signal tristate
flabel metal3 s 59200 42304 60000 42424 0 FreeSans 480 0 0 0 wbs_dat_o[31]
port 449 nsew signal tristate
flabel metal3 s 59200 8032 60000 8152 0 FreeSans 480 0 0 0 wbs_dat_o[3]
port 450 nsew signal tristate
flabel metal3 s 59200 9256 60000 9376 0 FreeSans 480 0 0 0 wbs_dat_o[4]
port 451 nsew signal tristate
flabel metal3 s 59200 10480 60000 10600 0 FreeSans 480 0 0 0 wbs_dat_o[5]
port 452 nsew signal tristate
flabel metal3 s 59200 11704 60000 11824 0 FreeSans 480 0 0 0 wbs_dat_o[6]
port 453 nsew signal tristate
flabel metal3 s 59200 12928 60000 13048 0 FreeSans 480 0 0 0 wbs_dat_o[7]
port 454 nsew signal tristate
flabel metal3 s 59200 14152 60000 14272 0 FreeSans 480 0 0 0 wbs_dat_o[8]
port 455 nsew signal tristate
flabel metal3 s 59200 15376 60000 15496 0 FreeSans 480 0 0 0 wbs_dat_o[9]
port 456 nsew signal tristate
flabel metal3 s 59200 2728 60000 2848 0 FreeSans 480 0 0 0 wbs_stb_i
port 457 nsew signal input
flabel metal3 s 59200 3136 60000 3256 0 FreeSans 480 0 0 0 wbs_we_i
port 458 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 60000 60000
<< end >>
