magic
tech sky130B
magscale 1 2
timestamp 1680267177
<< obsli1 >>
rect 1104 2159 58880 61489
<< obsm1 >>
rect 842 1300 59234 61520
<< metal2 >>
rect 846 63200 902 64000
rect 1582 63200 1638 64000
rect 2318 63200 2374 64000
rect 3054 63200 3110 64000
rect 3790 63200 3846 64000
rect 4526 63200 4582 64000
rect 5262 63200 5318 64000
rect 5998 63200 6054 64000
rect 6734 63200 6790 64000
rect 7470 63200 7526 64000
rect 8206 63200 8262 64000
rect 8942 63200 8998 64000
rect 9678 63200 9734 64000
rect 10414 63200 10470 64000
rect 11150 63200 11206 64000
rect 11886 63200 11942 64000
rect 12622 63200 12678 64000
rect 13358 63200 13414 64000
rect 14094 63200 14150 64000
rect 14830 63200 14886 64000
rect 15566 63200 15622 64000
rect 16302 63200 16358 64000
rect 17038 63200 17094 64000
rect 17774 63200 17830 64000
rect 18510 63200 18566 64000
rect 19246 63200 19302 64000
rect 19982 63200 20038 64000
rect 20718 63200 20774 64000
rect 21454 63200 21510 64000
rect 22190 63200 22246 64000
rect 22926 63200 22982 64000
rect 23662 63200 23718 64000
rect 24398 63200 24454 64000
rect 25134 63200 25190 64000
rect 25870 63200 25926 64000
rect 26606 63200 26662 64000
rect 27342 63200 27398 64000
rect 28078 63200 28134 64000
rect 28814 63200 28870 64000
rect 29550 63200 29606 64000
rect 30286 63200 30342 64000
rect 31022 63200 31078 64000
rect 31758 63200 31814 64000
rect 32494 63200 32550 64000
rect 33230 63200 33286 64000
rect 33966 63200 34022 64000
rect 34702 63200 34758 64000
rect 35438 63200 35494 64000
rect 36174 63200 36230 64000
rect 36910 63200 36966 64000
rect 37646 63200 37702 64000
rect 38382 63200 38438 64000
rect 39118 63200 39174 64000
rect 39854 63200 39910 64000
rect 40590 63200 40646 64000
rect 41326 63200 41382 64000
rect 42062 63200 42118 64000
rect 42798 63200 42854 64000
rect 43534 63200 43590 64000
rect 44270 63200 44326 64000
rect 45006 63200 45062 64000
rect 45742 63200 45798 64000
rect 46478 63200 46534 64000
rect 47214 63200 47270 64000
rect 47950 63200 48006 64000
rect 48686 63200 48742 64000
rect 49422 63200 49478 64000
rect 50158 63200 50214 64000
rect 50894 63200 50950 64000
rect 51630 63200 51686 64000
rect 52366 63200 52422 64000
rect 53102 63200 53158 64000
rect 53838 63200 53894 64000
rect 54574 63200 54630 64000
rect 55310 63200 55366 64000
rect 56046 63200 56102 64000
rect 56782 63200 56838 64000
rect 57518 63200 57574 64000
rect 58254 63200 58310 64000
rect 58990 63200 59046 64000
rect 5906 0 5962 800
rect 6182 0 6238 800
rect 6458 0 6514 800
rect 6734 0 6790 800
rect 7010 0 7066 800
rect 7286 0 7342 800
rect 7562 0 7618 800
rect 7838 0 7894 800
rect 8114 0 8170 800
rect 8390 0 8446 800
rect 8666 0 8722 800
rect 8942 0 8998 800
rect 9218 0 9274 800
rect 9494 0 9550 800
rect 9770 0 9826 800
rect 10046 0 10102 800
rect 10322 0 10378 800
rect 10598 0 10654 800
rect 10874 0 10930 800
rect 11150 0 11206 800
rect 11426 0 11482 800
rect 11702 0 11758 800
rect 11978 0 12034 800
rect 12254 0 12310 800
rect 12530 0 12586 800
rect 12806 0 12862 800
rect 13082 0 13138 800
rect 13358 0 13414 800
rect 13634 0 13690 800
rect 13910 0 13966 800
rect 14186 0 14242 800
rect 14462 0 14518 800
rect 14738 0 14794 800
rect 15014 0 15070 800
rect 15290 0 15346 800
rect 15566 0 15622 800
rect 15842 0 15898 800
rect 16118 0 16174 800
rect 16394 0 16450 800
rect 16670 0 16726 800
rect 16946 0 17002 800
rect 17222 0 17278 800
rect 17498 0 17554 800
rect 17774 0 17830 800
rect 18050 0 18106 800
rect 18326 0 18382 800
rect 18602 0 18658 800
rect 18878 0 18934 800
rect 19154 0 19210 800
rect 19430 0 19486 800
rect 19706 0 19762 800
rect 19982 0 20038 800
rect 20258 0 20314 800
rect 20534 0 20590 800
rect 20810 0 20866 800
rect 21086 0 21142 800
rect 21362 0 21418 800
rect 21638 0 21694 800
rect 21914 0 21970 800
rect 22190 0 22246 800
rect 22466 0 22522 800
rect 22742 0 22798 800
rect 23018 0 23074 800
rect 23294 0 23350 800
rect 23570 0 23626 800
rect 23846 0 23902 800
rect 24122 0 24178 800
rect 24398 0 24454 800
rect 24674 0 24730 800
rect 24950 0 25006 800
rect 25226 0 25282 800
rect 25502 0 25558 800
rect 25778 0 25834 800
rect 26054 0 26110 800
rect 26330 0 26386 800
rect 26606 0 26662 800
rect 26882 0 26938 800
rect 27158 0 27214 800
rect 27434 0 27490 800
rect 27710 0 27766 800
rect 27986 0 28042 800
rect 28262 0 28318 800
rect 28538 0 28594 800
rect 28814 0 28870 800
rect 29090 0 29146 800
rect 29366 0 29422 800
rect 29642 0 29698 800
rect 29918 0 29974 800
rect 30194 0 30250 800
rect 30470 0 30526 800
rect 30746 0 30802 800
rect 31022 0 31078 800
rect 31298 0 31354 800
rect 31574 0 31630 800
rect 31850 0 31906 800
rect 32126 0 32182 800
rect 32402 0 32458 800
rect 32678 0 32734 800
rect 32954 0 33010 800
rect 33230 0 33286 800
rect 33506 0 33562 800
rect 33782 0 33838 800
rect 34058 0 34114 800
rect 34334 0 34390 800
rect 34610 0 34666 800
rect 34886 0 34942 800
rect 35162 0 35218 800
rect 35438 0 35494 800
rect 35714 0 35770 800
rect 35990 0 36046 800
rect 36266 0 36322 800
rect 36542 0 36598 800
rect 36818 0 36874 800
rect 37094 0 37150 800
rect 37370 0 37426 800
rect 37646 0 37702 800
rect 37922 0 37978 800
rect 38198 0 38254 800
rect 38474 0 38530 800
rect 38750 0 38806 800
rect 39026 0 39082 800
rect 39302 0 39358 800
rect 39578 0 39634 800
rect 39854 0 39910 800
rect 40130 0 40186 800
rect 40406 0 40462 800
rect 40682 0 40738 800
rect 40958 0 41014 800
rect 41234 0 41290 800
rect 41510 0 41566 800
rect 41786 0 41842 800
rect 42062 0 42118 800
rect 42338 0 42394 800
rect 42614 0 42670 800
rect 42890 0 42946 800
rect 43166 0 43222 800
rect 43442 0 43498 800
rect 43718 0 43774 800
rect 43994 0 44050 800
rect 44270 0 44326 800
rect 44546 0 44602 800
rect 44822 0 44878 800
rect 45098 0 45154 800
rect 45374 0 45430 800
rect 45650 0 45706 800
rect 45926 0 45982 800
rect 46202 0 46258 800
rect 46478 0 46534 800
rect 46754 0 46810 800
rect 47030 0 47086 800
rect 47306 0 47362 800
rect 47582 0 47638 800
rect 47858 0 47914 800
rect 48134 0 48190 800
rect 48410 0 48466 800
rect 48686 0 48742 800
rect 48962 0 49018 800
rect 49238 0 49294 800
rect 49514 0 49570 800
rect 49790 0 49846 800
rect 50066 0 50122 800
rect 50342 0 50398 800
rect 50618 0 50674 800
rect 50894 0 50950 800
rect 51170 0 51226 800
rect 51446 0 51502 800
rect 51722 0 51778 800
rect 51998 0 52054 800
rect 52274 0 52330 800
rect 52550 0 52606 800
rect 52826 0 52882 800
rect 53102 0 53158 800
rect 53378 0 53434 800
rect 53654 0 53710 800
rect 53930 0 53986 800
<< obsm2 >>
rect 958 63144 1526 63322
rect 1694 63144 2262 63322
rect 2430 63144 2998 63322
rect 3166 63144 3734 63322
rect 3902 63144 4470 63322
rect 4638 63144 5206 63322
rect 5374 63144 5942 63322
rect 6110 63144 6678 63322
rect 6846 63144 7414 63322
rect 7582 63144 8150 63322
rect 8318 63144 8886 63322
rect 9054 63144 9622 63322
rect 9790 63144 10358 63322
rect 10526 63144 11094 63322
rect 11262 63144 11830 63322
rect 11998 63144 12566 63322
rect 12734 63144 13302 63322
rect 13470 63144 14038 63322
rect 14206 63144 14774 63322
rect 14942 63144 15510 63322
rect 15678 63144 16246 63322
rect 16414 63144 16982 63322
rect 17150 63144 17718 63322
rect 17886 63144 18454 63322
rect 18622 63144 19190 63322
rect 19358 63144 19926 63322
rect 20094 63144 20662 63322
rect 20830 63144 21398 63322
rect 21566 63144 22134 63322
rect 22302 63144 22870 63322
rect 23038 63144 23606 63322
rect 23774 63144 24342 63322
rect 24510 63144 25078 63322
rect 25246 63144 25814 63322
rect 25982 63144 26550 63322
rect 26718 63144 27286 63322
rect 27454 63144 28022 63322
rect 28190 63144 28758 63322
rect 28926 63144 29494 63322
rect 29662 63144 30230 63322
rect 30398 63144 30966 63322
rect 31134 63144 31702 63322
rect 31870 63144 32438 63322
rect 32606 63144 33174 63322
rect 33342 63144 33910 63322
rect 34078 63144 34646 63322
rect 34814 63144 35382 63322
rect 35550 63144 36118 63322
rect 36286 63144 36854 63322
rect 37022 63144 37590 63322
rect 37758 63144 38326 63322
rect 38494 63144 39062 63322
rect 39230 63144 39798 63322
rect 39966 63144 40534 63322
rect 40702 63144 41270 63322
rect 41438 63144 42006 63322
rect 42174 63144 42742 63322
rect 42910 63144 43478 63322
rect 43646 63144 44214 63322
rect 44382 63144 44950 63322
rect 45118 63144 45686 63322
rect 45854 63144 46422 63322
rect 46590 63144 47158 63322
rect 47326 63144 47894 63322
rect 48062 63144 48630 63322
rect 48798 63144 49366 63322
rect 49534 63144 50102 63322
rect 50270 63144 50838 63322
rect 51006 63144 51574 63322
rect 51742 63144 52310 63322
rect 52478 63144 53046 63322
rect 53214 63144 53782 63322
rect 53950 63144 54518 63322
rect 54686 63144 55254 63322
rect 55422 63144 55990 63322
rect 56158 63144 56726 63322
rect 56894 63144 57462 63322
rect 57630 63144 58198 63322
rect 58366 63144 58934 63322
rect 59102 63144 59228 63322
rect 848 856 59228 63144
rect 848 800 5850 856
rect 6018 800 6126 856
rect 6294 800 6402 856
rect 6570 800 6678 856
rect 6846 800 6954 856
rect 7122 800 7230 856
rect 7398 800 7506 856
rect 7674 800 7782 856
rect 7950 800 8058 856
rect 8226 800 8334 856
rect 8502 800 8610 856
rect 8778 800 8886 856
rect 9054 800 9162 856
rect 9330 800 9438 856
rect 9606 800 9714 856
rect 9882 800 9990 856
rect 10158 800 10266 856
rect 10434 800 10542 856
rect 10710 800 10818 856
rect 10986 800 11094 856
rect 11262 800 11370 856
rect 11538 800 11646 856
rect 11814 800 11922 856
rect 12090 800 12198 856
rect 12366 800 12474 856
rect 12642 800 12750 856
rect 12918 800 13026 856
rect 13194 800 13302 856
rect 13470 800 13578 856
rect 13746 800 13854 856
rect 14022 800 14130 856
rect 14298 800 14406 856
rect 14574 800 14682 856
rect 14850 800 14958 856
rect 15126 800 15234 856
rect 15402 800 15510 856
rect 15678 800 15786 856
rect 15954 800 16062 856
rect 16230 800 16338 856
rect 16506 800 16614 856
rect 16782 800 16890 856
rect 17058 800 17166 856
rect 17334 800 17442 856
rect 17610 800 17718 856
rect 17886 800 17994 856
rect 18162 800 18270 856
rect 18438 800 18546 856
rect 18714 800 18822 856
rect 18990 800 19098 856
rect 19266 800 19374 856
rect 19542 800 19650 856
rect 19818 800 19926 856
rect 20094 800 20202 856
rect 20370 800 20478 856
rect 20646 800 20754 856
rect 20922 800 21030 856
rect 21198 800 21306 856
rect 21474 800 21582 856
rect 21750 800 21858 856
rect 22026 800 22134 856
rect 22302 800 22410 856
rect 22578 800 22686 856
rect 22854 800 22962 856
rect 23130 800 23238 856
rect 23406 800 23514 856
rect 23682 800 23790 856
rect 23958 800 24066 856
rect 24234 800 24342 856
rect 24510 800 24618 856
rect 24786 800 24894 856
rect 25062 800 25170 856
rect 25338 800 25446 856
rect 25614 800 25722 856
rect 25890 800 25998 856
rect 26166 800 26274 856
rect 26442 800 26550 856
rect 26718 800 26826 856
rect 26994 800 27102 856
rect 27270 800 27378 856
rect 27546 800 27654 856
rect 27822 800 27930 856
rect 28098 800 28206 856
rect 28374 800 28482 856
rect 28650 800 28758 856
rect 28926 800 29034 856
rect 29202 800 29310 856
rect 29478 800 29586 856
rect 29754 800 29862 856
rect 30030 800 30138 856
rect 30306 800 30414 856
rect 30582 800 30690 856
rect 30858 800 30966 856
rect 31134 800 31242 856
rect 31410 800 31518 856
rect 31686 800 31794 856
rect 31962 800 32070 856
rect 32238 800 32346 856
rect 32514 800 32622 856
rect 32790 800 32898 856
rect 33066 800 33174 856
rect 33342 800 33450 856
rect 33618 800 33726 856
rect 33894 800 34002 856
rect 34170 800 34278 856
rect 34446 800 34554 856
rect 34722 800 34830 856
rect 34998 800 35106 856
rect 35274 800 35382 856
rect 35550 800 35658 856
rect 35826 800 35934 856
rect 36102 800 36210 856
rect 36378 800 36486 856
rect 36654 800 36762 856
rect 36930 800 37038 856
rect 37206 800 37314 856
rect 37482 800 37590 856
rect 37758 800 37866 856
rect 38034 800 38142 856
rect 38310 800 38418 856
rect 38586 800 38694 856
rect 38862 800 38970 856
rect 39138 800 39246 856
rect 39414 800 39522 856
rect 39690 800 39798 856
rect 39966 800 40074 856
rect 40242 800 40350 856
rect 40518 800 40626 856
rect 40794 800 40902 856
rect 41070 800 41178 856
rect 41346 800 41454 856
rect 41622 800 41730 856
rect 41898 800 42006 856
rect 42174 800 42282 856
rect 42450 800 42558 856
rect 42726 800 42834 856
rect 43002 800 43110 856
rect 43278 800 43386 856
rect 43554 800 43662 856
rect 43830 800 43938 856
rect 44106 800 44214 856
rect 44382 800 44490 856
rect 44658 800 44766 856
rect 44934 800 45042 856
rect 45210 800 45318 856
rect 45486 800 45594 856
rect 45762 800 45870 856
rect 46038 800 46146 856
rect 46314 800 46422 856
rect 46590 800 46698 856
rect 46866 800 46974 856
rect 47142 800 47250 856
rect 47418 800 47526 856
rect 47694 800 47802 856
rect 47970 800 48078 856
rect 48246 800 48354 856
rect 48522 800 48630 856
rect 48798 800 48906 856
rect 49074 800 49182 856
rect 49350 800 49458 856
rect 49626 800 49734 856
rect 49902 800 50010 856
rect 50178 800 50286 856
rect 50454 800 50562 856
rect 50730 800 50838 856
rect 51006 800 51114 856
rect 51282 800 51390 856
rect 51558 800 51666 856
rect 51834 800 51942 856
rect 52110 800 52218 856
rect 52386 800 52494 856
rect 52662 800 52770 856
rect 52938 800 53046 856
rect 53214 800 53322 856
rect 53490 800 53598 856
rect 53766 800 53874 856
rect 54042 800 59228 856
<< metal3 >>
rect 59200 62568 60000 62688
rect 59200 62024 60000 62144
rect 0 61480 800 61600
rect 59200 61480 60000 61600
rect 0 60800 800 60920
rect 59200 60936 60000 61056
rect 59200 60392 60000 60512
rect 0 60120 800 60240
rect 59200 59848 60000 59968
rect 0 59440 800 59560
rect 59200 59304 60000 59424
rect 0 58760 800 58880
rect 59200 58760 60000 58880
rect 0 58080 800 58200
rect 59200 58216 60000 58336
rect 59200 57672 60000 57792
rect 0 57400 800 57520
rect 59200 57128 60000 57248
rect 0 56720 800 56840
rect 59200 56584 60000 56704
rect 0 56040 800 56160
rect 59200 56040 60000 56160
rect 0 55360 800 55480
rect 59200 55496 60000 55616
rect 59200 54952 60000 55072
rect 0 54680 800 54800
rect 59200 54408 60000 54528
rect 0 54000 800 54120
rect 59200 53864 60000 53984
rect 0 53320 800 53440
rect 59200 53320 60000 53440
rect 0 52640 800 52760
rect 59200 52776 60000 52896
rect 59200 52232 60000 52352
rect 0 51960 800 52080
rect 59200 51688 60000 51808
rect 0 51280 800 51400
rect 59200 51144 60000 51264
rect 0 50600 800 50720
rect 59200 50600 60000 50720
rect 0 49920 800 50040
rect 59200 50056 60000 50176
rect 59200 49512 60000 49632
rect 0 49240 800 49360
rect 59200 48968 60000 49088
rect 0 48560 800 48680
rect 59200 48424 60000 48544
rect 0 47880 800 48000
rect 59200 47880 60000 48000
rect 0 47200 800 47320
rect 59200 47336 60000 47456
rect 59200 46792 60000 46912
rect 0 46520 800 46640
rect 59200 46248 60000 46368
rect 0 45840 800 45960
rect 59200 45704 60000 45824
rect 0 45160 800 45280
rect 59200 45160 60000 45280
rect 0 44480 800 44600
rect 59200 44616 60000 44736
rect 59200 44072 60000 44192
rect 0 43800 800 43920
rect 59200 43528 60000 43648
rect 0 43120 800 43240
rect 59200 42984 60000 43104
rect 0 42440 800 42560
rect 59200 42440 60000 42560
rect 0 41760 800 41880
rect 59200 41896 60000 42016
rect 59200 41352 60000 41472
rect 0 41080 800 41200
rect 59200 40808 60000 40928
rect 0 40400 800 40520
rect 59200 40264 60000 40384
rect 0 39720 800 39840
rect 59200 39720 60000 39840
rect 0 39040 800 39160
rect 59200 39176 60000 39296
rect 59200 38632 60000 38752
rect 0 38360 800 38480
rect 59200 38088 60000 38208
rect 0 37680 800 37800
rect 59200 37544 60000 37664
rect 0 37000 800 37120
rect 59200 37000 60000 37120
rect 0 36320 800 36440
rect 59200 36456 60000 36576
rect 59200 35912 60000 36032
rect 0 35640 800 35760
rect 59200 35368 60000 35488
rect 0 34960 800 35080
rect 59200 34824 60000 34944
rect 0 34280 800 34400
rect 59200 34280 60000 34400
rect 0 33600 800 33720
rect 59200 33736 60000 33856
rect 59200 33192 60000 33312
rect 0 32920 800 33040
rect 59200 32648 60000 32768
rect 0 32240 800 32360
rect 59200 32104 60000 32224
rect 0 31560 800 31680
rect 59200 31560 60000 31680
rect 0 30880 800 31000
rect 59200 31016 60000 31136
rect 59200 30472 60000 30592
rect 0 30200 800 30320
rect 59200 29928 60000 30048
rect 0 29520 800 29640
rect 59200 29384 60000 29504
rect 0 28840 800 28960
rect 59200 28840 60000 28960
rect 0 28160 800 28280
rect 59200 28296 60000 28416
rect 59200 27752 60000 27872
rect 0 27480 800 27600
rect 59200 27208 60000 27328
rect 0 26800 800 26920
rect 59200 26664 60000 26784
rect 0 26120 800 26240
rect 59200 26120 60000 26240
rect 0 25440 800 25560
rect 59200 25576 60000 25696
rect 59200 25032 60000 25152
rect 0 24760 800 24880
rect 59200 24488 60000 24608
rect 0 24080 800 24200
rect 59200 23944 60000 24064
rect 0 23400 800 23520
rect 59200 23400 60000 23520
rect 0 22720 800 22840
rect 59200 22856 60000 22976
rect 59200 22312 60000 22432
rect 0 22040 800 22160
rect 59200 21768 60000 21888
rect 0 21360 800 21480
rect 59200 21224 60000 21344
rect 0 20680 800 20800
rect 59200 20680 60000 20800
rect 0 20000 800 20120
rect 59200 20136 60000 20256
rect 59200 19592 60000 19712
rect 0 19320 800 19440
rect 59200 19048 60000 19168
rect 0 18640 800 18760
rect 59200 18504 60000 18624
rect 0 17960 800 18080
rect 59200 17960 60000 18080
rect 0 17280 800 17400
rect 59200 17416 60000 17536
rect 59200 16872 60000 16992
rect 0 16600 800 16720
rect 59200 16328 60000 16448
rect 0 15920 800 16040
rect 59200 15784 60000 15904
rect 0 15240 800 15360
rect 59200 15240 60000 15360
rect 0 14560 800 14680
rect 59200 14696 60000 14816
rect 59200 14152 60000 14272
rect 0 13880 800 14000
rect 59200 13608 60000 13728
rect 0 13200 800 13320
rect 59200 13064 60000 13184
rect 0 12520 800 12640
rect 59200 12520 60000 12640
rect 0 11840 800 11960
rect 59200 11976 60000 12096
rect 59200 11432 60000 11552
rect 0 11160 800 11280
rect 59200 10888 60000 11008
rect 0 10480 800 10600
rect 59200 10344 60000 10464
rect 0 9800 800 9920
rect 59200 9800 60000 9920
rect 0 9120 800 9240
rect 59200 9256 60000 9376
rect 59200 8712 60000 8832
rect 0 8440 800 8560
rect 59200 8168 60000 8288
rect 0 7760 800 7880
rect 59200 7624 60000 7744
rect 0 7080 800 7200
rect 59200 7080 60000 7200
rect 0 6400 800 6520
rect 59200 6536 60000 6656
rect 59200 5992 60000 6112
rect 0 5720 800 5840
rect 59200 5448 60000 5568
rect 0 5040 800 5160
rect 59200 4904 60000 5024
rect 0 4360 800 4480
rect 59200 4360 60000 4480
rect 0 3680 800 3800
rect 59200 3816 60000 3936
rect 59200 3272 60000 3392
rect 0 3000 800 3120
rect 59200 2728 60000 2848
rect 0 2320 800 2440
rect 59200 2184 60000 2304
rect 59200 1640 60000 1760
rect 59200 1096 60000 1216
<< obsm3 >>
rect 800 62488 59120 62661
rect 800 62224 59200 62488
rect 800 61944 59120 62224
rect 800 61680 59200 61944
rect 880 61400 59120 61680
rect 800 61136 59200 61400
rect 800 61000 59120 61136
rect 880 60856 59120 61000
rect 880 60720 59200 60856
rect 800 60592 59200 60720
rect 800 60320 59120 60592
rect 880 60312 59120 60320
rect 880 60048 59200 60312
rect 880 60040 59120 60048
rect 800 59768 59120 60040
rect 800 59640 59200 59768
rect 880 59504 59200 59640
rect 880 59360 59120 59504
rect 800 59224 59120 59360
rect 800 58960 59200 59224
rect 880 58680 59120 58960
rect 800 58416 59200 58680
rect 800 58280 59120 58416
rect 880 58136 59120 58280
rect 880 58000 59200 58136
rect 800 57872 59200 58000
rect 800 57600 59120 57872
rect 880 57592 59120 57600
rect 880 57328 59200 57592
rect 880 57320 59120 57328
rect 800 57048 59120 57320
rect 800 56920 59200 57048
rect 880 56784 59200 56920
rect 880 56640 59120 56784
rect 800 56504 59120 56640
rect 800 56240 59200 56504
rect 880 55960 59120 56240
rect 800 55696 59200 55960
rect 800 55560 59120 55696
rect 880 55416 59120 55560
rect 880 55280 59200 55416
rect 800 55152 59200 55280
rect 800 54880 59120 55152
rect 880 54872 59120 54880
rect 880 54608 59200 54872
rect 880 54600 59120 54608
rect 800 54328 59120 54600
rect 800 54200 59200 54328
rect 880 54064 59200 54200
rect 880 53920 59120 54064
rect 800 53784 59120 53920
rect 800 53520 59200 53784
rect 880 53240 59120 53520
rect 800 52976 59200 53240
rect 800 52840 59120 52976
rect 880 52696 59120 52840
rect 880 52560 59200 52696
rect 800 52432 59200 52560
rect 800 52160 59120 52432
rect 880 52152 59120 52160
rect 880 51888 59200 52152
rect 880 51880 59120 51888
rect 800 51608 59120 51880
rect 800 51480 59200 51608
rect 880 51344 59200 51480
rect 880 51200 59120 51344
rect 800 51064 59120 51200
rect 800 50800 59200 51064
rect 880 50520 59120 50800
rect 800 50256 59200 50520
rect 800 50120 59120 50256
rect 880 49976 59120 50120
rect 880 49840 59200 49976
rect 800 49712 59200 49840
rect 800 49440 59120 49712
rect 880 49432 59120 49440
rect 880 49168 59200 49432
rect 880 49160 59120 49168
rect 800 48888 59120 49160
rect 800 48760 59200 48888
rect 880 48624 59200 48760
rect 880 48480 59120 48624
rect 800 48344 59120 48480
rect 800 48080 59200 48344
rect 880 47800 59120 48080
rect 800 47536 59200 47800
rect 800 47400 59120 47536
rect 880 47256 59120 47400
rect 880 47120 59200 47256
rect 800 46992 59200 47120
rect 800 46720 59120 46992
rect 880 46712 59120 46720
rect 880 46448 59200 46712
rect 880 46440 59120 46448
rect 800 46168 59120 46440
rect 800 46040 59200 46168
rect 880 45904 59200 46040
rect 880 45760 59120 45904
rect 800 45624 59120 45760
rect 800 45360 59200 45624
rect 880 45080 59120 45360
rect 800 44816 59200 45080
rect 800 44680 59120 44816
rect 880 44536 59120 44680
rect 880 44400 59200 44536
rect 800 44272 59200 44400
rect 800 44000 59120 44272
rect 880 43992 59120 44000
rect 880 43728 59200 43992
rect 880 43720 59120 43728
rect 800 43448 59120 43720
rect 800 43320 59200 43448
rect 880 43184 59200 43320
rect 880 43040 59120 43184
rect 800 42904 59120 43040
rect 800 42640 59200 42904
rect 880 42360 59120 42640
rect 800 42096 59200 42360
rect 800 41960 59120 42096
rect 880 41816 59120 41960
rect 880 41680 59200 41816
rect 800 41552 59200 41680
rect 800 41280 59120 41552
rect 880 41272 59120 41280
rect 880 41008 59200 41272
rect 880 41000 59120 41008
rect 800 40728 59120 41000
rect 800 40600 59200 40728
rect 880 40464 59200 40600
rect 880 40320 59120 40464
rect 800 40184 59120 40320
rect 800 39920 59200 40184
rect 880 39640 59120 39920
rect 800 39376 59200 39640
rect 800 39240 59120 39376
rect 880 39096 59120 39240
rect 880 38960 59200 39096
rect 800 38832 59200 38960
rect 800 38560 59120 38832
rect 880 38552 59120 38560
rect 880 38288 59200 38552
rect 880 38280 59120 38288
rect 800 38008 59120 38280
rect 800 37880 59200 38008
rect 880 37744 59200 37880
rect 880 37600 59120 37744
rect 800 37464 59120 37600
rect 800 37200 59200 37464
rect 880 36920 59120 37200
rect 800 36656 59200 36920
rect 800 36520 59120 36656
rect 880 36376 59120 36520
rect 880 36240 59200 36376
rect 800 36112 59200 36240
rect 800 35840 59120 36112
rect 880 35832 59120 35840
rect 880 35568 59200 35832
rect 880 35560 59120 35568
rect 800 35288 59120 35560
rect 800 35160 59200 35288
rect 880 35024 59200 35160
rect 880 34880 59120 35024
rect 800 34744 59120 34880
rect 800 34480 59200 34744
rect 880 34200 59120 34480
rect 800 33936 59200 34200
rect 800 33800 59120 33936
rect 880 33656 59120 33800
rect 880 33520 59200 33656
rect 800 33392 59200 33520
rect 800 33120 59120 33392
rect 880 33112 59120 33120
rect 880 32848 59200 33112
rect 880 32840 59120 32848
rect 800 32568 59120 32840
rect 800 32440 59200 32568
rect 880 32304 59200 32440
rect 880 32160 59120 32304
rect 800 32024 59120 32160
rect 800 31760 59200 32024
rect 880 31480 59120 31760
rect 800 31216 59200 31480
rect 800 31080 59120 31216
rect 880 30936 59120 31080
rect 880 30800 59200 30936
rect 800 30672 59200 30800
rect 800 30400 59120 30672
rect 880 30392 59120 30400
rect 880 30128 59200 30392
rect 880 30120 59120 30128
rect 800 29848 59120 30120
rect 800 29720 59200 29848
rect 880 29584 59200 29720
rect 880 29440 59120 29584
rect 800 29304 59120 29440
rect 800 29040 59200 29304
rect 880 28760 59120 29040
rect 800 28496 59200 28760
rect 800 28360 59120 28496
rect 880 28216 59120 28360
rect 880 28080 59200 28216
rect 800 27952 59200 28080
rect 800 27680 59120 27952
rect 880 27672 59120 27680
rect 880 27408 59200 27672
rect 880 27400 59120 27408
rect 800 27128 59120 27400
rect 800 27000 59200 27128
rect 880 26864 59200 27000
rect 880 26720 59120 26864
rect 800 26584 59120 26720
rect 800 26320 59200 26584
rect 880 26040 59120 26320
rect 800 25776 59200 26040
rect 800 25640 59120 25776
rect 880 25496 59120 25640
rect 880 25360 59200 25496
rect 800 25232 59200 25360
rect 800 24960 59120 25232
rect 880 24952 59120 24960
rect 880 24688 59200 24952
rect 880 24680 59120 24688
rect 800 24408 59120 24680
rect 800 24280 59200 24408
rect 880 24144 59200 24280
rect 880 24000 59120 24144
rect 800 23864 59120 24000
rect 800 23600 59200 23864
rect 880 23320 59120 23600
rect 800 23056 59200 23320
rect 800 22920 59120 23056
rect 880 22776 59120 22920
rect 880 22640 59200 22776
rect 800 22512 59200 22640
rect 800 22240 59120 22512
rect 880 22232 59120 22240
rect 880 21968 59200 22232
rect 880 21960 59120 21968
rect 800 21688 59120 21960
rect 800 21560 59200 21688
rect 880 21424 59200 21560
rect 880 21280 59120 21424
rect 800 21144 59120 21280
rect 800 20880 59200 21144
rect 880 20600 59120 20880
rect 800 20336 59200 20600
rect 800 20200 59120 20336
rect 880 20056 59120 20200
rect 880 19920 59200 20056
rect 800 19792 59200 19920
rect 800 19520 59120 19792
rect 880 19512 59120 19520
rect 880 19248 59200 19512
rect 880 19240 59120 19248
rect 800 18968 59120 19240
rect 800 18840 59200 18968
rect 880 18704 59200 18840
rect 880 18560 59120 18704
rect 800 18424 59120 18560
rect 800 18160 59200 18424
rect 880 17880 59120 18160
rect 800 17616 59200 17880
rect 800 17480 59120 17616
rect 880 17336 59120 17480
rect 880 17200 59200 17336
rect 800 17072 59200 17200
rect 800 16800 59120 17072
rect 880 16792 59120 16800
rect 880 16528 59200 16792
rect 880 16520 59120 16528
rect 800 16248 59120 16520
rect 800 16120 59200 16248
rect 880 15984 59200 16120
rect 880 15840 59120 15984
rect 800 15704 59120 15840
rect 800 15440 59200 15704
rect 880 15160 59120 15440
rect 800 14896 59200 15160
rect 800 14760 59120 14896
rect 880 14616 59120 14760
rect 880 14480 59200 14616
rect 800 14352 59200 14480
rect 800 14080 59120 14352
rect 880 14072 59120 14080
rect 880 13808 59200 14072
rect 880 13800 59120 13808
rect 800 13528 59120 13800
rect 800 13400 59200 13528
rect 880 13264 59200 13400
rect 880 13120 59120 13264
rect 800 12984 59120 13120
rect 800 12720 59200 12984
rect 880 12440 59120 12720
rect 800 12176 59200 12440
rect 800 12040 59120 12176
rect 880 11896 59120 12040
rect 880 11760 59200 11896
rect 800 11632 59200 11760
rect 800 11360 59120 11632
rect 880 11352 59120 11360
rect 880 11088 59200 11352
rect 880 11080 59120 11088
rect 800 10808 59120 11080
rect 800 10680 59200 10808
rect 880 10544 59200 10680
rect 880 10400 59120 10544
rect 800 10264 59120 10400
rect 800 10000 59200 10264
rect 880 9720 59120 10000
rect 800 9456 59200 9720
rect 800 9320 59120 9456
rect 880 9176 59120 9320
rect 880 9040 59200 9176
rect 800 8912 59200 9040
rect 800 8640 59120 8912
rect 880 8632 59120 8640
rect 880 8368 59200 8632
rect 880 8360 59120 8368
rect 800 8088 59120 8360
rect 800 7960 59200 8088
rect 880 7824 59200 7960
rect 880 7680 59120 7824
rect 800 7544 59120 7680
rect 800 7280 59200 7544
rect 880 7000 59120 7280
rect 800 6736 59200 7000
rect 800 6600 59120 6736
rect 880 6456 59120 6600
rect 880 6320 59200 6456
rect 800 6192 59200 6320
rect 800 5920 59120 6192
rect 880 5912 59120 5920
rect 880 5648 59200 5912
rect 880 5640 59120 5648
rect 800 5368 59120 5640
rect 800 5240 59200 5368
rect 880 5104 59200 5240
rect 880 4960 59120 5104
rect 800 4824 59120 4960
rect 800 4560 59200 4824
rect 880 4280 59120 4560
rect 800 4016 59200 4280
rect 800 3880 59120 4016
rect 880 3736 59120 3880
rect 880 3600 59200 3736
rect 800 3472 59200 3600
rect 800 3200 59120 3472
rect 880 3192 59120 3200
rect 880 2928 59200 3192
rect 880 2920 59120 2928
rect 800 2648 59120 2920
rect 800 2520 59200 2648
rect 880 2384 59200 2520
rect 880 2240 59120 2384
rect 800 2104 59120 2240
rect 800 1840 59200 2104
rect 800 1560 59120 1840
rect 800 1296 59200 1560
rect 800 1123 59120 1296
<< metal4 >>
rect 4208 2128 4528 61520
rect 19568 2128 19888 61520
rect 34928 2128 35248 61520
rect 50288 2128 50608 61520
<< obsm4 >>
rect 18275 2347 19488 61165
rect 19968 2347 34848 61165
rect 35328 2347 40973 61165
<< labels >>
rlabel metal3 s 0 21360 800 21480 6 design_clk_o
port 1 nsew signal output
rlabel metal3 s 0 2320 800 2440 6 dsi_all[0]
port 2 nsew signal output
rlabel metal3 s 0 9120 800 9240 6 dsi_all[10]
port 3 nsew signal output
rlabel metal3 s 0 9800 800 9920 6 dsi_all[11]
port 4 nsew signal output
rlabel metal3 s 0 10480 800 10600 6 dsi_all[12]
port 5 nsew signal output
rlabel metal3 s 0 11160 800 11280 6 dsi_all[13]
port 6 nsew signal output
rlabel metal3 s 0 11840 800 11960 6 dsi_all[14]
port 7 nsew signal output
rlabel metal3 s 0 12520 800 12640 6 dsi_all[15]
port 8 nsew signal output
rlabel metal3 s 0 13200 800 13320 6 dsi_all[16]
port 9 nsew signal output
rlabel metal3 s 0 13880 800 14000 6 dsi_all[17]
port 10 nsew signal output
rlabel metal3 s 0 14560 800 14680 6 dsi_all[18]
port 11 nsew signal output
rlabel metal3 s 0 15240 800 15360 6 dsi_all[19]
port 12 nsew signal output
rlabel metal3 s 0 3000 800 3120 6 dsi_all[1]
port 13 nsew signal output
rlabel metal3 s 0 15920 800 16040 6 dsi_all[20]
port 14 nsew signal output
rlabel metal3 s 0 16600 800 16720 6 dsi_all[21]
port 15 nsew signal output
rlabel metal3 s 0 17280 800 17400 6 dsi_all[22]
port 16 nsew signal output
rlabel metal3 s 0 17960 800 18080 6 dsi_all[23]
port 17 nsew signal output
rlabel metal3 s 0 18640 800 18760 6 dsi_all[24]
port 18 nsew signal output
rlabel metal3 s 0 19320 800 19440 6 dsi_all[25]
port 19 nsew signal output
rlabel metal3 s 0 20000 800 20120 6 dsi_all[26]
port 20 nsew signal output
rlabel metal3 s 0 20680 800 20800 6 dsi_all[27]
port 21 nsew signal output
rlabel metal3 s 0 3680 800 3800 6 dsi_all[2]
port 22 nsew signal output
rlabel metal3 s 0 4360 800 4480 6 dsi_all[3]
port 23 nsew signal output
rlabel metal3 s 0 5040 800 5160 6 dsi_all[4]
port 24 nsew signal output
rlabel metal3 s 0 5720 800 5840 6 dsi_all[5]
port 25 nsew signal output
rlabel metal3 s 0 6400 800 6520 6 dsi_all[6]
port 26 nsew signal output
rlabel metal3 s 0 7080 800 7200 6 dsi_all[7]
port 27 nsew signal output
rlabel metal3 s 0 7760 800 7880 6 dsi_all[8]
port 28 nsew signal output
rlabel metal3 s 0 8440 800 8560 6 dsi_all[9]
port 29 nsew signal output
rlabel metal2 s 38750 0 38806 800 6 dso_6502[0]
port 30 nsew signal input
rlabel metal2 s 41510 0 41566 800 6 dso_6502[10]
port 31 nsew signal input
rlabel metal2 s 41786 0 41842 800 6 dso_6502[11]
port 32 nsew signal input
rlabel metal2 s 42062 0 42118 800 6 dso_6502[12]
port 33 nsew signal input
rlabel metal2 s 42338 0 42394 800 6 dso_6502[13]
port 34 nsew signal input
rlabel metal2 s 42614 0 42670 800 6 dso_6502[14]
port 35 nsew signal input
rlabel metal2 s 42890 0 42946 800 6 dso_6502[15]
port 36 nsew signal input
rlabel metal2 s 43166 0 43222 800 6 dso_6502[16]
port 37 nsew signal input
rlabel metal2 s 43442 0 43498 800 6 dso_6502[17]
port 38 nsew signal input
rlabel metal2 s 43718 0 43774 800 6 dso_6502[18]
port 39 nsew signal input
rlabel metal2 s 43994 0 44050 800 6 dso_6502[19]
port 40 nsew signal input
rlabel metal2 s 39026 0 39082 800 6 dso_6502[1]
port 41 nsew signal input
rlabel metal2 s 44270 0 44326 800 6 dso_6502[20]
port 42 nsew signal input
rlabel metal2 s 44546 0 44602 800 6 dso_6502[21]
port 43 nsew signal input
rlabel metal2 s 44822 0 44878 800 6 dso_6502[22]
port 44 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 dso_6502[23]
port 45 nsew signal input
rlabel metal2 s 45374 0 45430 800 6 dso_6502[24]
port 46 nsew signal input
rlabel metal2 s 45650 0 45706 800 6 dso_6502[25]
port 47 nsew signal input
rlabel metal2 s 45926 0 45982 800 6 dso_6502[26]
port 48 nsew signal input
rlabel metal2 s 39302 0 39358 800 6 dso_6502[2]
port 49 nsew signal input
rlabel metal2 s 39578 0 39634 800 6 dso_6502[3]
port 50 nsew signal input
rlabel metal2 s 39854 0 39910 800 6 dso_6502[4]
port 51 nsew signal input
rlabel metal2 s 40130 0 40186 800 6 dso_6502[5]
port 52 nsew signal input
rlabel metal2 s 40406 0 40462 800 6 dso_6502[6]
port 53 nsew signal input
rlabel metal2 s 40682 0 40738 800 6 dso_6502[7]
port 54 nsew signal input
rlabel metal2 s 40958 0 41014 800 6 dso_6502[8]
port 55 nsew signal input
rlabel metal2 s 41234 0 41290 800 6 dso_6502[9]
port 56 nsew signal input
rlabel metal2 s 53838 63200 53894 64000 6 dso_LCD[0]
port 57 nsew signal input
rlabel metal2 s 54574 63200 54630 64000 6 dso_LCD[1]
port 58 nsew signal input
rlabel metal2 s 55310 63200 55366 64000 6 dso_LCD[2]
port 59 nsew signal input
rlabel metal2 s 56046 63200 56102 64000 6 dso_LCD[3]
port 60 nsew signal input
rlabel metal2 s 56782 63200 56838 64000 6 dso_LCD[4]
port 61 nsew signal input
rlabel metal2 s 57518 63200 57574 64000 6 dso_LCD[5]
port 62 nsew signal input
rlabel metal2 s 58254 63200 58310 64000 6 dso_LCD[6]
port 63 nsew signal input
rlabel metal2 s 58990 63200 59046 64000 6 dso_LCD[7]
port 64 nsew signal input
rlabel metal2 s 46202 0 46258 800 6 dso_as1802[0]
port 65 nsew signal input
rlabel metal2 s 48962 0 49018 800 6 dso_as1802[10]
port 66 nsew signal input
rlabel metal2 s 49238 0 49294 800 6 dso_as1802[11]
port 67 nsew signal input
rlabel metal2 s 49514 0 49570 800 6 dso_as1802[12]
port 68 nsew signal input
rlabel metal2 s 49790 0 49846 800 6 dso_as1802[13]
port 69 nsew signal input
rlabel metal2 s 50066 0 50122 800 6 dso_as1802[14]
port 70 nsew signal input
rlabel metal2 s 50342 0 50398 800 6 dso_as1802[15]
port 71 nsew signal input
rlabel metal2 s 50618 0 50674 800 6 dso_as1802[16]
port 72 nsew signal input
rlabel metal2 s 50894 0 50950 800 6 dso_as1802[17]
port 73 nsew signal input
rlabel metal2 s 51170 0 51226 800 6 dso_as1802[18]
port 74 nsew signal input
rlabel metal2 s 51446 0 51502 800 6 dso_as1802[19]
port 75 nsew signal input
rlabel metal2 s 46478 0 46534 800 6 dso_as1802[1]
port 76 nsew signal input
rlabel metal2 s 51722 0 51778 800 6 dso_as1802[20]
port 77 nsew signal input
rlabel metal2 s 51998 0 52054 800 6 dso_as1802[21]
port 78 nsew signal input
rlabel metal2 s 52274 0 52330 800 6 dso_as1802[22]
port 79 nsew signal input
rlabel metal2 s 52550 0 52606 800 6 dso_as1802[23]
port 80 nsew signal input
rlabel metal2 s 52826 0 52882 800 6 dso_as1802[24]
port 81 nsew signal input
rlabel metal2 s 53102 0 53158 800 6 dso_as1802[25]
port 82 nsew signal input
rlabel metal2 s 53378 0 53434 800 6 dso_as1802[26]
port 83 nsew signal input
rlabel metal2 s 46754 0 46810 800 6 dso_as1802[2]
port 84 nsew signal input
rlabel metal2 s 47030 0 47086 800 6 dso_as1802[3]
port 85 nsew signal input
rlabel metal2 s 47306 0 47362 800 6 dso_as1802[4]
port 86 nsew signal input
rlabel metal2 s 47582 0 47638 800 6 dso_as1802[5]
port 87 nsew signal input
rlabel metal2 s 47858 0 47914 800 6 dso_as1802[6]
port 88 nsew signal input
rlabel metal2 s 48134 0 48190 800 6 dso_as1802[7]
port 89 nsew signal input
rlabel metal2 s 48410 0 48466 800 6 dso_as1802[8]
port 90 nsew signal input
rlabel metal2 s 48686 0 48742 800 6 dso_as1802[9]
port 91 nsew signal input
rlabel metal2 s 13358 63200 13414 64000 6 dso_as2650[0]
port 92 nsew signal input
rlabel metal2 s 20718 63200 20774 64000 6 dso_as2650[10]
port 93 nsew signal input
rlabel metal2 s 21454 63200 21510 64000 6 dso_as2650[11]
port 94 nsew signal input
rlabel metal2 s 22190 63200 22246 64000 6 dso_as2650[12]
port 95 nsew signal input
rlabel metal2 s 22926 63200 22982 64000 6 dso_as2650[13]
port 96 nsew signal input
rlabel metal2 s 23662 63200 23718 64000 6 dso_as2650[14]
port 97 nsew signal input
rlabel metal2 s 24398 63200 24454 64000 6 dso_as2650[15]
port 98 nsew signal input
rlabel metal2 s 25134 63200 25190 64000 6 dso_as2650[16]
port 99 nsew signal input
rlabel metal2 s 25870 63200 25926 64000 6 dso_as2650[17]
port 100 nsew signal input
rlabel metal2 s 26606 63200 26662 64000 6 dso_as2650[18]
port 101 nsew signal input
rlabel metal2 s 27342 63200 27398 64000 6 dso_as2650[19]
port 102 nsew signal input
rlabel metal2 s 14094 63200 14150 64000 6 dso_as2650[1]
port 103 nsew signal input
rlabel metal2 s 28078 63200 28134 64000 6 dso_as2650[20]
port 104 nsew signal input
rlabel metal2 s 28814 63200 28870 64000 6 dso_as2650[21]
port 105 nsew signal input
rlabel metal2 s 29550 63200 29606 64000 6 dso_as2650[22]
port 106 nsew signal input
rlabel metal2 s 30286 63200 30342 64000 6 dso_as2650[23]
port 107 nsew signal input
rlabel metal2 s 31022 63200 31078 64000 6 dso_as2650[24]
port 108 nsew signal input
rlabel metal2 s 31758 63200 31814 64000 6 dso_as2650[25]
port 109 nsew signal input
rlabel metal2 s 32494 63200 32550 64000 6 dso_as2650[26]
port 110 nsew signal input
rlabel metal2 s 14830 63200 14886 64000 6 dso_as2650[2]
port 111 nsew signal input
rlabel metal2 s 15566 63200 15622 64000 6 dso_as2650[3]
port 112 nsew signal input
rlabel metal2 s 16302 63200 16358 64000 6 dso_as2650[4]
port 113 nsew signal input
rlabel metal2 s 17038 63200 17094 64000 6 dso_as2650[5]
port 114 nsew signal input
rlabel metal2 s 17774 63200 17830 64000 6 dso_as2650[6]
port 115 nsew signal input
rlabel metal2 s 18510 63200 18566 64000 6 dso_as2650[7]
port 116 nsew signal input
rlabel metal2 s 19246 63200 19302 64000 6 dso_as2650[8]
port 117 nsew signal input
rlabel metal2 s 19982 63200 20038 64000 6 dso_as2650[9]
port 118 nsew signal input
rlabel metal3 s 0 42440 800 42560 6 dso_as512512512[0]
port 119 nsew signal input
rlabel metal3 s 0 49240 800 49360 6 dso_as512512512[10]
port 120 nsew signal input
rlabel metal3 s 0 49920 800 50040 6 dso_as512512512[11]
port 121 nsew signal input
rlabel metal3 s 0 50600 800 50720 6 dso_as512512512[12]
port 122 nsew signal input
rlabel metal3 s 0 51280 800 51400 6 dso_as512512512[13]
port 123 nsew signal input
rlabel metal3 s 0 51960 800 52080 6 dso_as512512512[14]
port 124 nsew signal input
rlabel metal3 s 0 52640 800 52760 6 dso_as512512512[15]
port 125 nsew signal input
rlabel metal3 s 0 53320 800 53440 6 dso_as512512512[16]
port 126 nsew signal input
rlabel metal3 s 0 54000 800 54120 6 dso_as512512512[17]
port 127 nsew signal input
rlabel metal3 s 0 54680 800 54800 6 dso_as512512512[18]
port 128 nsew signal input
rlabel metal3 s 0 55360 800 55480 6 dso_as512512512[19]
port 129 nsew signal input
rlabel metal3 s 0 43120 800 43240 6 dso_as512512512[1]
port 130 nsew signal input
rlabel metal3 s 0 56040 800 56160 6 dso_as512512512[20]
port 131 nsew signal input
rlabel metal3 s 0 56720 800 56840 6 dso_as512512512[21]
port 132 nsew signal input
rlabel metal3 s 0 57400 800 57520 6 dso_as512512512[22]
port 133 nsew signal input
rlabel metal3 s 0 58080 800 58200 6 dso_as512512512[23]
port 134 nsew signal input
rlabel metal3 s 0 58760 800 58880 6 dso_as512512512[24]
port 135 nsew signal input
rlabel metal3 s 0 59440 800 59560 6 dso_as512512512[25]
port 136 nsew signal input
rlabel metal3 s 0 60120 800 60240 6 dso_as512512512[26]
port 137 nsew signal input
rlabel metal3 s 0 60800 800 60920 6 dso_as512512512[27]
port 138 nsew signal input
rlabel metal3 s 0 43800 800 43920 6 dso_as512512512[2]
port 139 nsew signal input
rlabel metal3 s 0 44480 800 44600 6 dso_as512512512[3]
port 140 nsew signal input
rlabel metal3 s 0 45160 800 45280 6 dso_as512512512[4]
port 141 nsew signal input
rlabel metal3 s 0 45840 800 45960 6 dso_as512512512[5]
port 142 nsew signal input
rlabel metal3 s 0 46520 800 46640 6 dso_as512512512[6]
port 143 nsew signal input
rlabel metal3 s 0 47200 800 47320 6 dso_as512512512[7]
port 144 nsew signal input
rlabel metal3 s 0 47880 800 48000 6 dso_as512512512[8]
port 145 nsew signal input
rlabel metal3 s 0 48560 800 48680 6 dso_as512512512[9]
port 146 nsew signal input
rlabel metal2 s 33230 63200 33286 64000 6 dso_as5401[0]
port 147 nsew signal input
rlabel metal2 s 40590 63200 40646 64000 6 dso_as5401[10]
port 148 nsew signal input
rlabel metal2 s 41326 63200 41382 64000 6 dso_as5401[11]
port 149 nsew signal input
rlabel metal2 s 42062 63200 42118 64000 6 dso_as5401[12]
port 150 nsew signal input
rlabel metal2 s 42798 63200 42854 64000 6 dso_as5401[13]
port 151 nsew signal input
rlabel metal2 s 43534 63200 43590 64000 6 dso_as5401[14]
port 152 nsew signal input
rlabel metal2 s 44270 63200 44326 64000 6 dso_as5401[15]
port 153 nsew signal input
rlabel metal2 s 45006 63200 45062 64000 6 dso_as5401[16]
port 154 nsew signal input
rlabel metal2 s 45742 63200 45798 64000 6 dso_as5401[17]
port 155 nsew signal input
rlabel metal2 s 46478 63200 46534 64000 6 dso_as5401[18]
port 156 nsew signal input
rlabel metal2 s 47214 63200 47270 64000 6 dso_as5401[19]
port 157 nsew signal input
rlabel metal2 s 33966 63200 34022 64000 6 dso_as5401[1]
port 158 nsew signal input
rlabel metal2 s 47950 63200 48006 64000 6 dso_as5401[20]
port 159 nsew signal input
rlabel metal2 s 48686 63200 48742 64000 6 dso_as5401[21]
port 160 nsew signal input
rlabel metal2 s 49422 63200 49478 64000 6 dso_as5401[22]
port 161 nsew signal input
rlabel metal2 s 50158 63200 50214 64000 6 dso_as5401[23]
port 162 nsew signal input
rlabel metal2 s 50894 63200 50950 64000 6 dso_as5401[24]
port 163 nsew signal input
rlabel metal2 s 51630 63200 51686 64000 6 dso_as5401[25]
port 164 nsew signal input
rlabel metal2 s 52366 63200 52422 64000 6 dso_as5401[26]
port 165 nsew signal input
rlabel metal2 s 34702 63200 34758 64000 6 dso_as5401[2]
port 166 nsew signal input
rlabel metal2 s 35438 63200 35494 64000 6 dso_as5401[3]
port 167 nsew signal input
rlabel metal2 s 36174 63200 36230 64000 6 dso_as5401[4]
port 168 nsew signal input
rlabel metal2 s 36910 63200 36966 64000 6 dso_as5401[5]
port 169 nsew signal input
rlabel metal2 s 37646 63200 37702 64000 6 dso_as5401[6]
port 170 nsew signal input
rlabel metal2 s 38382 63200 38438 64000 6 dso_as5401[7]
port 171 nsew signal input
rlabel metal2 s 39118 63200 39174 64000 6 dso_as5401[8]
port 172 nsew signal input
rlabel metal2 s 39854 63200 39910 64000 6 dso_as5401[9]
port 173 nsew signal input
rlabel metal3 s 59200 56584 60000 56704 6 dso_counter[0]
port 174 nsew signal input
rlabel metal3 s 59200 62024 60000 62144 6 dso_counter[10]
port 175 nsew signal input
rlabel metal3 s 59200 62568 60000 62688 6 dso_counter[11]
port 176 nsew signal input
rlabel metal3 s 59200 57128 60000 57248 6 dso_counter[1]
port 177 nsew signal input
rlabel metal3 s 59200 57672 60000 57792 6 dso_counter[2]
port 178 nsew signal input
rlabel metal3 s 59200 58216 60000 58336 6 dso_counter[3]
port 179 nsew signal input
rlabel metal3 s 59200 58760 60000 58880 6 dso_counter[4]
port 180 nsew signal input
rlabel metal3 s 59200 59304 60000 59424 6 dso_counter[5]
port 181 nsew signal input
rlabel metal3 s 59200 59848 60000 59968 6 dso_counter[6]
port 182 nsew signal input
rlabel metal3 s 59200 60392 60000 60512 6 dso_counter[7]
port 183 nsew signal input
rlabel metal3 s 59200 60936 60000 61056 6 dso_counter[8]
port 184 nsew signal input
rlabel metal3 s 59200 61480 60000 61600 6 dso_counter[9]
port 185 nsew signal input
rlabel metal2 s 6734 63200 6790 64000 6 dso_diceroll[0]
port 186 nsew signal input
rlabel metal2 s 7470 63200 7526 64000 6 dso_diceroll[1]
port 187 nsew signal input
rlabel metal2 s 8206 63200 8262 64000 6 dso_diceroll[2]
port 188 nsew signal input
rlabel metal2 s 8942 63200 8998 64000 6 dso_diceroll[3]
port 189 nsew signal input
rlabel metal2 s 9678 63200 9734 64000 6 dso_diceroll[4]
port 190 nsew signal input
rlabel metal2 s 10414 63200 10470 64000 6 dso_diceroll[5]
port 191 nsew signal input
rlabel metal2 s 11150 63200 11206 64000 6 dso_diceroll[6]
port 192 nsew signal input
rlabel metal2 s 11886 63200 11942 64000 6 dso_diceroll[7]
port 193 nsew signal input
rlabel metal3 s 0 30200 800 30320 6 dso_mc14500[0]
port 194 nsew signal input
rlabel metal3 s 0 30880 800 31000 6 dso_mc14500[1]
port 195 nsew signal input
rlabel metal3 s 0 31560 800 31680 6 dso_mc14500[2]
port 196 nsew signal input
rlabel metal3 s 0 32240 800 32360 6 dso_mc14500[3]
port 197 nsew signal input
rlabel metal3 s 0 32920 800 33040 6 dso_mc14500[4]
port 198 nsew signal input
rlabel metal3 s 0 33600 800 33720 6 dso_mc14500[5]
port 199 nsew signal input
rlabel metal3 s 0 34280 800 34400 6 dso_mc14500[6]
port 200 nsew signal input
rlabel metal3 s 0 34960 800 35080 6 dso_mc14500[7]
port 201 nsew signal input
rlabel metal3 s 0 35640 800 35760 6 dso_mc14500[8]
port 202 nsew signal input
rlabel metal2 s 846 63200 902 64000 6 dso_multiplier[0]
port 203 nsew signal input
rlabel metal2 s 1582 63200 1638 64000 6 dso_multiplier[1]
port 204 nsew signal input
rlabel metal2 s 2318 63200 2374 64000 6 dso_multiplier[2]
port 205 nsew signal input
rlabel metal2 s 3054 63200 3110 64000 6 dso_multiplier[3]
port 206 nsew signal input
rlabel metal2 s 3790 63200 3846 64000 6 dso_multiplier[4]
port 207 nsew signal input
rlabel metal2 s 4526 63200 4582 64000 6 dso_multiplier[5]
port 208 nsew signal input
rlabel metal2 s 5262 63200 5318 64000 6 dso_multiplier[6]
port 209 nsew signal input
rlabel metal2 s 5998 63200 6054 64000 6 dso_multiplier[7]
port 210 nsew signal input
rlabel metal2 s 37370 0 37426 800 6 dso_posit[0]
port 211 nsew signal input
rlabel metal2 s 37646 0 37702 800 6 dso_posit[1]
port 212 nsew signal input
rlabel metal2 s 37922 0 37978 800 6 dso_posit[2]
port 213 nsew signal input
rlabel metal2 s 38198 0 38254 800 6 dso_posit[3]
port 214 nsew signal input
rlabel metal3 s 0 37000 800 37120 6 dso_tbb1143[0]
port 215 nsew signal input
rlabel metal3 s 0 37680 800 37800 6 dso_tbb1143[1]
port 216 nsew signal input
rlabel metal3 s 0 38360 800 38480 6 dso_tbb1143[2]
port 217 nsew signal input
rlabel metal3 s 0 39040 800 39160 6 dso_tbb1143[3]
port 218 nsew signal input
rlabel metal3 s 0 39720 800 39840 6 dso_tbb1143[4]
port 219 nsew signal input
rlabel metal3 s 0 40400 800 40520 6 dso_tbb1143[5]
port 220 nsew signal input
rlabel metal3 s 0 41080 800 41200 6 dso_tbb1143[6]
port 221 nsew signal input
rlabel metal3 s 0 41760 800 41880 6 dso_tbb1143[7]
port 222 nsew signal input
rlabel metal2 s 53930 0 53986 800 6 dso_tune
port 223 nsew signal input
rlabel metal2 s 5906 0 5962 800 6 io_in[0]
port 224 nsew signal input
rlabel metal2 s 8666 0 8722 800 6 io_in[10]
port 225 nsew signal input
rlabel metal2 s 8942 0 8998 800 6 io_in[11]
port 226 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 io_in[12]
port 227 nsew signal input
rlabel metal2 s 9494 0 9550 800 6 io_in[13]
port 228 nsew signal input
rlabel metal2 s 9770 0 9826 800 6 io_in[14]
port 229 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 io_in[15]
port 230 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 io_in[16]
port 231 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 io_in[17]
port 232 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 io_in[18]
port 233 nsew signal input
rlabel metal2 s 11150 0 11206 800 6 io_in[19]
port 234 nsew signal input
rlabel metal2 s 6182 0 6238 800 6 io_in[1]
port 235 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 io_in[20]
port 236 nsew signal input
rlabel metal2 s 11702 0 11758 800 6 io_in[21]
port 237 nsew signal input
rlabel metal2 s 11978 0 12034 800 6 io_in[22]
port 238 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 io_in[23]
port 239 nsew signal input
rlabel metal2 s 12530 0 12586 800 6 io_in[24]
port 240 nsew signal input
rlabel metal2 s 12806 0 12862 800 6 io_in[25]
port 241 nsew signal input
rlabel metal2 s 13082 0 13138 800 6 io_in[26]
port 242 nsew signal input
rlabel metal2 s 13358 0 13414 800 6 io_in[27]
port 243 nsew signal input
rlabel metal2 s 13634 0 13690 800 6 io_in[28]
port 244 nsew signal input
rlabel metal2 s 13910 0 13966 800 6 io_in[29]
port 245 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 io_in[2]
port 246 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 io_in[30]
port 247 nsew signal input
rlabel metal2 s 14462 0 14518 800 6 io_in[31]
port 248 nsew signal input
rlabel metal2 s 14738 0 14794 800 6 io_in[32]
port 249 nsew signal input
rlabel metal2 s 15014 0 15070 800 6 io_in[33]
port 250 nsew signal input
rlabel metal2 s 15290 0 15346 800 6 io_in[34]
port 251 nsew signal input
rlabel metal2 s 15566 0 15622 800 6 io_in[35]
port 252 nsew signal input
rlabel metal2 s 15842 0 15898 800 6 io_in[36]
port 253 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 io_in[37]
port 254 nsew signal input
rlabel metal2 s 6734 0 6790 800 6 io_in[3]
port 255 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 io_in[4]
port 256 nsew signal input
rlabel metal2 s 7286 0 7342 800 6 io_in[5]
port 257 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 io_in[6]
port 258 nsew signal input
rlabel metal2 s 7838 0 7894 800 6 io_in[7]
port 259 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 io_in[8]
port 260 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 io_in[9]
port 261 nsew signal input
rlabel metal2 s 26882 0 26938 800 6 io_oeb[0]
port 262 nsew signal output
rlabel metal2 s 29642 0 29698 800 6 io_oeb[10]
port 263 nsew signal output
rlabel metal2 s 29918 0 29974 800 6 io_oeb[11]
port 264 nsew signal output
rlabel metal2 s 30194 0 30250 800 6 io_oeb[12]
port 265 nsew signal output
rlabel metal2 s 30470 0 30526 800 6 io_oeb[13]
port 266 nsew signal output
rlabel metal2 s 30746 0 30802 800 6 io_oeb[14]
port 267 nsew signal output
rlabel metal2 s 31022 0 31078 800 6 io_oeb[15]
port 268 nsew signal output
rlabel metal2 s 31298 0 31354 800 6 io_oeb[16]
port 269 nsew signal output
rlabel metal2 s 31574 0 31630 800 6 io_oeb[17]
port 270 nsew signal output
rlabel metal2 s 31850 0 31906 800 6 io_oeb[18]
port 271 nsew signal output
rlabel metal2 s 32126 0 32182 800 6 io_oeb[19]
port 272 nsew signal output
rlabel metal2 s 27158 0 27214 800 6 io_oeb[1]
port 273 nsew signal output
rlabel metal2 s 32402 0 32458 800 6 io_oeb[20]
port 274 nsew signal output
rlabel metal2 s 32678 0 32734 800 6 io_oeb[21]
port 275 nsew signal output
rlabel metal2 s 32954 0 33010 800 6 io_oeb[22]
port 276 nsew signal output
rlabel metal2 s 33230 0 33286 800 6 io_oeb[23]
port 277 nsew signal output
rlabel metal2 s 33506 0 33562 800 6 io_oeb[24]
port 278 nsew signal output
rlabel metal2 s 33782 0 33838 800 6 io_oeb[25]
port 279 nsew signal output
rlabel metal2 s 34058 0 34114 800 6 io_oeb[26]
port 280 nsew signal output
rlabel metal2 s 34334 0 34390 800 6 io_oeb[27]
port 281 nsew signal output
rlabel metal2 s 34610 0 34666 800 6 io_oeb[28]
port 282 nsew signal output
rlabel metal2 s 34886 0 34942 800 6 io_oeb[29]
port 283 nsew signal output
rlabel metal2 s 27434 0 27490 800 6 io_oeb[2]
port 284 nsew signal output
rlabel metal2 s 35162 0 35218 800 6 io_oeb[30]
port 285 nsew signal output
rlabel metal2 s 35438 0 35494 800 6 io_oeb[31]
port 286 nsew signal output
rlabel metal2 s 35714 0 35770 800 6 io_oeb[32]
port 287 nsew signal output
rlabel metal2 s 35990 0 36046 800 6 io_oeb[33]
port 288 nsew signal output
rlabel metal2 s 36266 0 36322 800 6 io_oeb[34]
port 289 nsew signal output
rlabel metal2 s 36542 0 36598 800 6 io_oeb[35]
port 290 nsew signal output
rlabel metal2 s 36818 0 36874 800 6 io_oeb[36]
port 291 nsew signal output
rlabel metal2 s 37094 0 37150 800 6 io_oeb[37]
port 292 nsew signal output
rlabel metal2 s 27710 0 27766 800 6 io_oeb[3]
port 293 nsew signal output
rlabel metal2 s 27986 0 28042 800 6 io_oeb[4]
port 294 nsew signal output
rlabel metal2 s 28262 0 28318 800 6 io_oeb[5]
port 295 nsew signal output
rlabel metal2 s 28538 0 28594 800 6 io_oeb[6]
port 296 nsew signal output
rlabel metal2 s 28814 0 28870 800 6 io_oeb[7]
port 297 nsew signal output
rlabel metal2 s 29090 0 29146 800 6 io_oeb[8]
port 298 nsew signal output
rlabel metal2 s 29366 0 29422 800 6 io_oeb[9]
port 299 nsew signal output
rlabel metal2 s 16394 0 16450 800 6 io_out[0]
port 300 nsew signal output
rlabel metal2 s 19154 0 19210 800 6 io_out[10]
port 301 nsew signal output
rlabel metal2 s 19430 0 19486 800 6 io_out[11]
port 302 nsew signal output
rlabel metal2 s 19706 0 19762 800 6 io_out[12]
port 303 nsew signal output
rlabel metal2 s 19982 0 20038 800 6 io_out[13]
port 304 nsew signal output
rlabel metal2 s 20258 0 20314 800 6 io_out[14]
port 305 nsew signal output
rlabel metal2 s 20534 0 20590 800 6 io_out[15]
port 306 nsew signal output
rlabel metal2 s 20810 0 20866 800 6 io_out[16]
port 307 nsew signal output
rlabel metal2 s 21086 0 21142 800 6 io_out[17]
port 308 nsew signal output
rlabel metal2 s 21362 0 21418 800 6 io_out[18]
port 309 nsew signal output
rlabel metal2 s 21638 0 21694 800 6 io_out[19]
port 310 nsew signal output
rlabel metal2 s 16670 0 16726 800 6 io_out[1]
port 311 nsew signal output
rlabel metal2 s 21914 0 21970 800 6 io_out[20]
port 312 nsew signal output
rlabel metal2 s 22190 0 22246 800 6 io_out[21]
port 313 nsew signal output
rlabel metal2 s 22466 0 22522 800 6 io_out[22]
port 314 nsew signal output
rlabel metal2 s 22742 0 22798 800 6 io_out[23]
port 315 nsew signal output
rlabel metal2 s 23018 0 23074 800 6 io_out[24]
port 316 nsew signal output
rlabel metal2 s 23294 0 23350 800 6 io_out[25]
port 317 nsew signal output
rlabel metal2 s 23570 0 23626 800 6 io_out[26]
port 318 nsew signal output
rlabel metal2 s 23846 0 23902 800 6 io_out[27]
port 319 nsew signal output
rlabel metal2 s 24122 0 24178 800 6 io_out[28]
port 320 nsew signal output
rlabel metal2 s 24398 0 24454 800 6 io_out[29]
port 321 nsew signal output
rlabel metal2 s 16946 0 17002 800 6 io_out[2]
port 322 nsew signal output
rlabel metal2 s 24674 0 24730 800 6 io_out[30]
port 323 nsew signal output
rlabel metal2 s 24950 0 25006 800 6 io_out[31]
port 324 nsew signal output
rlabel metal2 s 25226 0 25282 800 6 io_out[32]
port 325 nsew signal output
rlabel metal2 s 25502 0 25558 800 6 io_out[33]
port 326 nsew signal output
rlabel metal2 s 25778 0 25834 800 6 io_out[34]
port 327 nsew signal output
rlabel metal2 s 26054 0 26110 800 6 io_out[35]
port 328 nsew signal output
rlabel metal2 s 26330 0 26386 800 6 io_out[36]
port 329 nsew signal output
rlabel metal2 s 26606 0 26662 800 6 io_out[37]
port 330 nsew signal output
rlabel metal2 s 17222 0 17278 800 6 io_out[3]
port 331 nsew signal output
rlabel metal2 s 17498 0 17554 800 6 io_out[4]
port 332 nsew signal output
rlabel metal2 s 17774 0 17830 800 6 io_out[5]
port 333 nsew signal output
rlabel metal2 s 18050 0 18106 800 6 io_out[6]
port 334 nsew signal output
rlabel metal2 s 18326 0 18382 800 6 io_out[7]
port 335 nsew signal output
rlabel metal2 s 18602 0 18658 800 6 io_out[8]
port 336 nsew signal output
rlabel metal2 s 18878 0 18934 800 6 io_out[9]
port 337 nsew signal output
rlabel metal2 s 38474 0 38530 800 6 oeb_6502
port 338 nsew signal input
rlabel metal2 s 53654 0 53710 800 6 oeb_as1802
port 339 nsew signal input
rlabel metal2 s 12622 63200 12678 64000 6 oeb_as2650
port 340 nsew signal input
rlabel metal3 s 0 61480 800 61600 6 oeb_as512512512
port 341 nsew signal input
rlabel metal2 s 53102 63200 53158 64000 6 oeb_as5401
port 342 nsew signal input
rlabel metal3 s 0 36320 800 36440 6 oeb_mc14500
port 343 nsew signal input
rlabel metal3 s 0 22040 800 22160 6 rst_6502
port 344 nsew signal output
rlabel metal3 s 0 22720 800 22840 6 rst_LCD
port 345 nsew signal output
rlabel metal3 s 0 23400 800 23520 6 rst_as1802
port 346 nsew signal output
rlabel metal3 s 0 24080 800 24200 6 rst_as2650
port 347 nsew signal output
rlabel metal3 s 0 25440 800 25560 6 rst_as512512512
port 348 nsew signal output
rlabel metal3 s 0 24760 800 24880 6 rst_as5401
port 349 nsew signal output
rlabel metal3 s 0 26120 800 26240 6 rst_counter
port 350 nsew signal output
rlabel metal3 s 0 26800 800 26920 6 rst_diceroll
port 351 nsew signal output
rlabel metal3 s 0 27480 800 27600 6 rst_mc14500
port 352 nsew signal output
rlabel metal3 s 0 28160 800 28280 6 rst_posit
port 353 nsew signal output
rlabel metal3 s 0 28840 800 28960 6 rst_tbb1143
port 354 nsew signal output
rlabel metal3 s 0 29520 800 29640 6 rst_tune
port 355 nsew signal output
rlabel metal4 s 4208 2128 4528 61520 6 vccd1
port 356 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 61520 6 vccd1
port 356 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 61520 6 vssd1
port 357 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 61520 6 vssd1
port 357 nsew ground bidirectional
rlabel metal3 s 59200 1096 60000 1216 6 wb_clk_i
port 358 nsew signal input
rlabel metal3 s 59200 1640 60000 1760 6 wb_rst_i
port 359 nsew signal input
rlabel metal3 s 59200 2184 60000 2304 6 wbs_ack_o
port 360 nsew signal output
rlabel metal3 s 59200 4360 60000 4480 6 wbs_adr_i[0]
port 361 nsew signal input
rlabel metal3 s 59200 20680 60000 20800 6 wbs_adr_i[10]
port 362 nsew signal input
rlabel metal3 s 59200 22312 60000 22432 6 wbs_adr_i[11]
port 363 nsew signal input
rlabel metal3 s 59200 23944 60000 24064 6 wbs_adr_i[12]
port 364 nsew signal input
rlabel metal3 s 59200 25576 60000 25696 6 wbs_adr_i[13]
port 365 nsew signal input
rlabel metal3 s 59200 27208 60000 27328 6 wbs_adr_i[14]
port 366 nsew signal input
rlabel metal3 s 59200 28840 60000 28960 6 wbs_adr_i[15]
port 367 nsew signal input
rlabel metal3 s 59200 30472 60000 30592 6 wbs_adr_i[16]
port 368 nsew signal input
rlabel metal3 s 59200 32104 60000 32224 6 wbs_adr_i[17]
port 369 nsew signal input
rlabel metal3 s 59200 33736 60000 33856 6 wbs_adr_i[18]
port 370 nsew signal input
rlabel metal3 s 59200 35368 60000 35488 6 wbs_adr_i[19]
port 371 nsew signal input
rlabel metal3 s 59200 5992 60000 6112 6 wbs_adr_i[1]
port 372 nsew signal input
rlabel metal3 s 59200 37000 60000 37120 6 wbs_adr_i[20]
port 373 nsew signal input
rlabel metal3 s 59200 38632 60000 38752 6 wbs_adr_i[21]
port 374 nsew signal input
rlabel metal3 s 59200 40264 60000 40384 6 wbs_adr_i[22]
port 375 nsew signal input
rlabel metal3 s 59200 41896 60000 42016 6 wbs_adr_i[23]
port 376 nsew signal input
rlabel metal3 s 59200 43528 60000 43648 6 wbs_adr_i[24]
port 377 nsew signal input
rlabel metal3 s 59200 45160 60000 45280 6 wbs_adr_i[25]
port 378 nsew signal input
rlabel metal3 s 59200 46792 60000 46912 6 wbs_adr_i[26]
port 379 nsew signal input
rlabel metal3 s 59200 48424 60000 48544 6 wbs_adr_i[27]
port 380 nsew signal input
rlabel metal3 s 59200 50056 60000 50176 6 wbs_adr_i[28]
port 381 nsew signal input
rlabel metal3 s 59200 51688 60000 51808 6 wbs_adr_i[29]
port 382 nsew signal input
rlabel metal3 s 59200 7624 60000 7744 6 wbs_adr_i[2]
port 383 nsew signal input
rlabel metal3 s 59200 53320 60000 53440 6 wbs_adr_i[30]
port 384 nsew signal input
rlabel metal3 s 59200 54952 60000 55072 6 wbs_adr_i[31]
port 385 nsew signal input
rlabel metal3 s 59200 9256 60000 9376 6 wbs_adr_i[3]
port 386 nsew signal input
rlabel metal3 s 59200 10888 60000 11008 6 wbs_adr_i[4]
port 387 nsew signal input
rlabel metal3 s 59200 12520 60000 12640 6 wbs_adr_i[5]
port 388 nsew signal input
rlabel metal3 s 59200 14152 60000 14272 6 wbs_adr_i[6]
port 389 nsew signal input
rlabel metal3 s 59200 15784 60000 15904 6 wbs_adr_i[7]
port 390 nsew signal input
rlabel metal3 s 59200 17416 60000 17536 6 wbs_adr_i[8]
port 391 nsew signal input
rlabel metal3 s 59200 19048 60000 19168 6 wbs_adr_i[9]
port 392 nsew signal input
rlabel metal3 s 59200 2728 60000 2848 6 wbs_cyc_i
port 393 nsew signal input
rlabel metal3 s 59200 4904 60000 5024 6 wbs_dat_i[0]
port 394 nsew signal input
rlabel metal3 s 59200 21224 60000 21344 6 wbs_dat_i[10]
port 395 nsew signal input
rlabel metal3 s 59200 22856 60000 22976 6 wbs_dat_i[11]
port 396 nsew signal input
rlabel metal3 s 59200 24488 60000 24608 6 wbs_dat_i[12]
port 397 nsew signal input
rlabel metal3 s 59200 26120 60000 26240 6 wbs_dat_i[13]
port 398 nsew signal input
rlabel metal3 s 59200 27752 60000 27872 6 wbs_dat_i[14]
port 399 nsew signal input
rlabel metal3 s 59200 29384 60000 29504 6 wbs_dat_i[15]
port 400 nsew signal input
rlabel metal3 s 59200 31016 60000 31136 6 wbs_dat_i[16]
port 401 nsew signal input
rlabel metal3 s 59200 32648 60000 32768 6 wbs_dat_i[17]
port 402 nsew signal input
rlabel metal3 s 59200 34280 60000 34400 6 wbs_dat_i[18]
port 403 nsew signal input
rlabel metal3 s 59200 35912 60000 36032 6 wbs_dat_i[19]
port 404 nsew signal input
rlabel metal3 s 59200 6536 60000 6656 6 wbs_dat_i[1]
port 405 nsew signal input
rlabel metal3 s 59200 37544 60000 37664 6 wbs_dat_i[20]
port 406 nsew signal input
rlabel metal3 s 59200 39176 60000 39296 6 wbs_dat_i[21]
port 407 nsew signal input
rlabel metal3 s 59200 40808 60000 40928 6 wbs_dat_i[22]
port 408 nsew signal input
rlabel metal3 s 59200 42440 60000 42560 6 wbs_dat_i[23]
port 409 nsew signal input
rlabel metal3 s 59200 44072 60000 44192 6 wbs_dat_i[24]
port 410 nsew signal input
rlabel metal3 s 59200 45704 60000 45824 6 wbs_dat_i[25]
port 411 nsew signal input
rlabel metal3 s 59200 47336 60000 47456 6 wbs_dat_i[26]
port 412 nsew signal input
rlabel metal3 s 59200 48968 60000 49088 6 wbs_dat_i[27]
port 413 nsew signal input
rlabel metal3 s 59200 50600 60000 50720 6 wbs_dat_i[28]
port 414 nsew signal input
rlabel metal3 s 59200 52232 60000 52352 6 wbs_dat_i[29]
port 415 nsew signal input
rlabel metal3 s 59200 8168 60000 8288 6 wbs_dat_i[2]
port 416 nsew signal input
rlabel metal3 s 59200 53864 60000 53984 6 wbs_dat_i[30]
port 417 nsew signal input
rlabel metal3 s 59200 55496 60000 55616 6 wbs_dat_i[31]
port 418 nsew signal input
rlabel metal3 s 59200 9800 60000 9920 6 wbs_dat_i[3]
port 419 nsew signal input
rlabel metal3 s 59200 11432 60000 11552 6 wbs_dat_i[4]
port 420 nsew signal input
rlabel metal3 s 59200 13064 60000 13184 6 wbs_dat_i[5]
port 421 nsew signal input
rlabel metal3 s 59200 14696 60000 14816 6 wbs_dat_i[6]
port 422 nsew signal input
rlabel metal3 s 59200 16328 60000 16448 6 wbs_dat_i[7]
port 423 nsew signal input
rlabel metal3 s 59200 17960 60000 18080 6 wbs_dat_i[8]
port 424 nsew signal input
rlabel metal3 s 59200 19592 60000 19712 6 wbs_dat_i[9]
port 425 nsew signal input
rlabel metal3 s 59200 5448 60000 5568 6 wbs_dat_o[0]
port 426 nsew signal output
rlabel metal3 s 59200 21768 60000 21888 6 wbs_dat_o[10]
port 427 nsew signal output
rlabel metal3 s 59200 23400 60000 23520 6 wbs_dat_o[11]
port 428 nsew signal output
rlabel metal3 s 59200 25032 60000 25152 6 wbs_dat_o[12]
port 429 nsew signal output
rlabel metal3 s 59200 26664 60000 26784 6 wbs_dat_o[13]
port 430 nsew signal output
rlabel metal3 s 59200 28296 60000 28416 6 wbs_dat_o[14]
port 431 nsew signal output
rlabel metal3 s 59200 29928 60000 30048 6 wbs_dat_o[15]
port 432 nsew signal output
rlabel metal3 s 59200 31560 60000 31680 6 wbs_dat_o[16]
port 433 nsew signal output
rlabel metal3 s 59200 33192 60000 33312 6 wbs_dat_o[17]
port 434 nsew signal output
rlabel metal3 s 59200 34824 60000 34944 6 wbs_dat_o[18]
port 435 nsew signal output
rlabel metal3 s 59200 36456 60000 36576 6 wbs_dat_o[19]
port 436 nsew signal output
rlabel metal3 s 59200 7080 60000 7200 6 wbs_dat_o[1]
port 437 nsew signal output
rlabel metal3 s 59200 38088 60000 38208 6 wbs_dat_o[20]
port 438 nsew signal output
rlabel metal3 s 59200 39720 60000 39840 6 wbs_dat_o[21]
port 439 nsew signal output
rlabel metal3 s 59200 41352 60000 41472 6 wbs_dat_o[22]
port 440 nsew signal output
rlabel metal3 s 59200 42984 60000 43104 6 wbs_dat_o[23]
port 441 nsew signal output
rlabel metal3 s 59200 44616 60000 44736 6 wbs_dat_o[24]
port 442 nsew signal output
rlabel metal3 s 59200 46248 60000 46368 6 wbs_dat_o[25]
port 443 nsew signal output
rlabel metal3 s 59200 47880 60000 48000 6 wbs_dat_o[26]
port 444 nsew signal output
rlabel metal3 s 59200 49512 60000 49632 6 wbs_dat_o[27]
port 445 nsew signal output
rlabel metal3 s 59200 51144 60000 51264 6 wbs_dat_o[28]
port 446 nsew signal output
rlabel metal3 s 59200 52776 60000 52896 6 wbs_dat_o[29]
port 447 nsew signal output
rlabel metal3 s 59200 8712 60000 8832 6 wbs_dat_o[2]
port 448 nsew signal output
rlabel metal3 s 59200 54408 60000 54528 6 wbs_dat_o[30]
port 449 nsew signal output
rlabel metal3 s 59200 56040 60000 56160 6 wbs_dat_o[31]
port 450 nsew signal output
rlabel metal3 s 59200 10344 60000 10464 6 wbs_dat_o[3]
port 451 nsew signal output
rlabel metal3 s 59200 11976 60000 12096 6 wbs_dat_o[4]
port 452 nsew signal output
rlabel metal3 s 59200 13608 60000 13728 6 wbs_dat_o[5]
port 453 nsew signal output
rlabel metal3 s 59200 15240 60000 15360 6 wbs_dat_o[6]
port 454 nsew signal output
rlabel metal3 s 59200 16872 60000 16992 6 wbs_dat_o[7]
port 455 nsew signal output
rlabel metal3 s 59200 18504 60000 18624 6 wbs_dat_o[8]
port 456 nsew signal output
rlabel metal3 s 59200 20136 60000 20256 6 wbs_dat_o[9]
port 457 nsew signal output
rlabel metal3 s 59200 3272 60000 3392 6 wbs_stb_i
port 458 nsew signal input
rlabel metal3 s 59200 3816 60000 3936 6 wbs_we_i
port 459 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 60000 64000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 4594530
string GDS_FILE /run/media/tholin/e6042058-84c8-448b-be8a-b40bc065b34b/TMBoC/openlane/Multiplexer/runs/23_03_31_14_46/results/signoff/multiplexer.magic.gds
string GDS_START 687750
<< end >>

