VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_as512512512
  CLASS BLOCK ;
  FOREIGN wrapped_as512512512 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1700.000 BY 3200.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 1517.120 1700.000 1517.720 ;
    END
  END clk
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 29.960 1700.000 30.560 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 580.760 1700.000 581.360 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 635.840 1700.000 636.440 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 690.920 1700.000 691.520 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 746.000 1700.000 746.600 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 801.080 1700.000 801.680 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 856.160 1700.000 856.760 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 911.240 1700.000 911.840 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 966.320 1700.000 966.920 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 1021.400 1700.000 1022.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 1076.480 1700.000 1077.080 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 85.040 1700.000 85.640 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 1131.560 1700.000 1132.160 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 1186.640 1700.000 1187.240 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 1241.720 1700.000 1242.320 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 1296.800 1700.000 1297.400 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 1351.880 1700.000 1352.480 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 1406.960 1700.000 1407.560 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 1462.040 1700.000 1462.640 ;
    END
  END io_in[26]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 140.120 1700.000 140.720 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 195.200 1700.000 195.800 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 250.280 1700.000 250.880 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 305.360 1700.000 305.960 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 360.440 1700.000 361.040 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 415.520 1700.000 416.120 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 470.600 1700.000 471.200 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 525.680 1700.000 526.280 ;
    END
  END io_in[9]
  PIN io_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 3169.520 1700.000 3170.120 ;
    END
  END io_oeb
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 1627.280 1700.000 1627.880 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 2178.080 1700.000 2178.680 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 2233.160 1700.000 2233.760 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 2288.240 1700.000 2288.840 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 2343.320 1700.000 2343.920 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 2398.400 1700.000 2399.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 2453.480 1700.000 2454.080 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 2508.560 1700.000 2509.160 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 2563.640 1700.000 2564.240 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 2618.720 1700.000 2619.320 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 2673.800 1700.000 2674.400 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 1682.360 1700.000 1682.960 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 2728.880 1700.000 2729.480 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 2783.960 1700.000 2784.560 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 2839.040 1700.000 2839.640 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 2894.120 1700.000 2894.720 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 2949.200 1700.000 2949.800 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 3004.280 1700.000 3004.880 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 3059.360 1700.000 3059.960 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 3114.440 1700.000 3115.040 ;
    END
  END io_out[27]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 1737.440 1700.000 1738.040 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 1792.520 1700.000 1793.120 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 1847.600 1700.000 1848.200 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 1902.680 1700.000 1903.280 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 1957.760 1700.000 1958.360 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 2012.840 1700.000 2013.440 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 2067.920 1700.000 2068.520 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 2123.000 1700.000 2123.600 ;
    END
  END io_out[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 1572.200 1700.000 1572.800 ;
    END
  END rst
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 10.640 1558.640 3188.080 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1633.840 10.640 1635.440 3188.080 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 3183.705 1694.370 3186.535 ;
        RECT 5.330 3178.265 1694.370 3181.095 ;
        RECT 5.330 3172.825 1694.370 3175.655 ;
        RECT 5.330 3167.385 1694.370 3170.215 ;
        RECT 5.330 3161.945 1694.370 3164.775 ;
        RECT 5.330 3156.505 1694.370 3159.335 ;
        RECT 5.330 3151.065 1694.370 3153.895 ;
        RECT 5.330 3145.625 1694.370 3148.455 ;
        RECT 5.330 3140.185 1694.370 3143.015 ;
        RECT 5.330 3134.745 1694.370 3137.575 ;
        RECT 5.330 3129.305 1694.370 3132.135 ;
        RECT 5.330 3123.865 1694.370 3126.695 ;
        RECT 5.330 3118.425 1694.370 3121.255 ;
        RECT 5.330 3112.985 1694.370 3115.815 ;
        RECT 5.330 3107.545 1694.370 3110.375 ;
        RECT 5.330 3102.105 1694.370 3104.935 ;
        RECT 5.330 3096.665 1694.370 3099.495 ;
        RECT 5.330 3091.225 1694.370 3094.055 ;
        RECT 5.330 3085.785 1694.370 3088.615 ;
        RECT 5.330 3080.345 1694.370 3083.175 ;
        RECT 5.330 3074.905 1694.370 3077.735 ;
        RECT 5.330 3069.465 1694.370 3072.295 ;
        RECT 5.330 3064.025 1694.370 3066.855 ;
        RECT 5.330 3058.585 1694.370 3061.415 ;
        RECT 5.330 3053.145 1694.370 3055.975 ;
        RECT 5.330 3047.705 1694.370 3050.535 ;
        RECT 5.330 3042.265 1694.370 3045.095 ;
        RECT 5.330 3036.825 1694.370 3039.655 ;
        RECT 5.330 3031.385 1694.370 3034.215 ;
        RECT 5.330 3025.945 1694.370 3028.775 ;
        RECT 5.330 3020.505 1694.370 3023.335 ;
        RECT 5.330 3015.065 1694.370 3017.895 ;
        RECT 5.330 3009.625 1694.370 3012.455 ;
        RECT 5.330 3004.185 1694.370 3007.015 ;
        RECT 5.330 2998.745 1694.370 3001.575 ;
        RECT 5.330 2993.305 1694.370 2996.135 ;
        RECT 5.330 2987.865 1694.370 2990.695 ;
        RECT 5.330 2982.425 1694.370 2985.255 ;
        RECT 5.330 2976.985 1694.370 2979.815 ;
        RECT 5.330 2971.545 1694.370 2974.375 ;
        RECT 5.330 2966.105 1694.370 2968.935 ;
        RECT 5.330 2960.665 1694.370 2963.495 ;
        RECT 5.330 2955.225 1694.370 2958.055 ;
        RECT 5.330 2949.785 1694.370 2952.615 ;
        RECT 5.330 2944.345 1694.370 2947.175 ;
        RECT 5.330 2938.905 1694.370 2941.735 ;
        RECT 5.330 2933.465 1694.370 2936.295 ;
        RECT 5.330 2928.025 1694.370 2930.855 ;
        RECT 5.330 2922.585 1694.370 2925.415 ;
        RECT 5.330 2917.145 1694.370 2919.975 ;
        RECT 5.330 2911.705 1694.370 2914.535 ;
        RECT 5.330 2906.265 1694.370 2909.095 ;
        RECT 5.330 2900.825 1694.370 2903.655 ;
        RECT 5.330 2895.385 1694.370 2898.215 ;
        RECT 5.330 2889.945 1694.370 2892.775 ;
        RECT 5.330 2884.505 1694.370 2887.335 ;
        RECT 5.330 2879.065 1694.370 2881.895 ;
        RECT 5.330 2873.625 1694.370 2876.455 ;
        RECT 5.330 2868.185 1694.370 2871.015 ;
        RECT 5.330 2862.745 1694.370 2865.575 ;
        RECT 5.330 2857.305 1694.370 2860.135 ;
        RECT 5.330 2851.865 1694.370 2854.695 ;
        RECT 5.330 2846.425 1694.370 2849.255 ;
        RECT 5.330 2840.985 1694.370 2843.815 ;
        RECT 5.330 2835.545 1694.370 2838.375 ;
        RECT 5.330 2830.105 1694.370 2832.935 ;
        RECT 5.330 2824.665 1694.370 2827.495 ;
        RECT 5.330 2819.225 1694.370 2822.055 ;
        RECT 5.330 2813.785 1694.370 2816.615 ;
        RECT 5.330 2808.345 1694.370 2811.175 ;
        RECT 5.330 2802.905 1694.370 2805.735 ;
        RECT 5.330 2797.465 1694.370 2800.295 ;
        RECT 5.330 2792.025 1694.370 2794.855 ;
        RECT 5.330 2786.585 1694.370 2789.415 ;
        RECT 5.330 2781.145 1694.370 2783.975 ;
        RECT 5.330 2775.705 1694.370 2778.535 ;
        RECT 5.330 2770.265 1694.370 2773.095 ;
        RECT 5.330 2764.825 1694.370 2767.655 ;
        RECT 5.330 2759.385 1694.370 2762.215 ;
        RECT 5.330 2753.945 1694.370 2756.775 ;
        RECT 5.330 2748.505 1694.370 2751.335 ;
        RECT 5.330 2743.065 1694.370 2745.895 ;
        RECT 5.330 2737.625 1694.370 2740.455 ;
        RECT 5.330 2732.185 1694.370 2735.015 ;
        RECT 5.330 2726.745 1694.370 2729.575 ;
        RECT 5.330 2721.305 1694.370 2724.135 ;
        RECT 5.330 2715.865 1694.370 2718.695 ;
        RECT 5.330 2710.425 1694.370 2713.255 ;
        RECT 5.330 2704.985 1694.370 2707.815 ;
        RECT 5.330 2699.545 1694.370 2702.375 ;
        RECT 5.330 2694.105 1694.370 2696.935 ;
        RECT 5.330 2688.665 1694.370 2691.495 ;
        RECT 5.330 2683.225 1694.370 2686.055 ;
        RECT 5.330 2677.785 1694.370 2680.615 ;
        RECT 5.330 2672.345 1694.370 2675.175 ;
        RECT 5.330 2666.905 1694.370 2669.735 ;
        RECT 5.330 2661.465 1694.370 2664.295 ;
        RECT 5.330 2656.025 1694.370 2658.855 ;
        RECT 5.330 2650.585 1694.370 2653.415 ;
        RECT 5.330 2645.145 1694.370 2647.975 ;
        RECT 5.330 2639.705 1694.370 2642.535 ;
        RECT 5.330 2634.265 1694.370 2637.095 ;
        RECT 5.330 2628.825 1694.370 2631.655 ;
        RECT 5.330 2623.385 1694.370 2626.215 ;
        RECT 5.330 2617.945 1694.370 2620.775 ;
        RECT 5.330 2612.505 1694.370 2615.335 ;
        RECT 5.330 2607.065 1694.370 2609.895 ;
        RECT 5.330 2601.625 1694.370 2604.455 ;
        RECT 5.330 2596.185 1694.370 2599.015 ;
        RECT 5.330 2590.745 1694.370 2593.575 ;
        RECT 5.330 2585.305 1694.370 2588.135 ;
        RECT 5.330 2579.865 1694.370 2582.695 ;
        RECT 5.330 2574.425 1694.370 2577.255 ;
        RECT 5.330 2568.985 1694.370 2571.815 ;
        RECT 5.330 2563.545 1694.370 2566.375 ;
        RECT 5.330 2558.105 1694.370 2560.935 ;
        RECT 5.330 2552.665 1694.370 2555.495 ;
        RECT 5.330 2547.225 1694.370 2550.055 ;
        RECT 5.330 2541.785 1694.370 2544.615 ;
        RECT 5.330 2536.345 1694.370 2539.175 ;
        RECT 5.330 2530.905 1694.370 2533.735 ;
        RECT 5.330 2525.465 1694.370 2528.295 ;
        RECT 5.330 2520.025 1694.370 2522.855 ;
        RECT 5.330 2514.585 1694.370 2517.415 ;
        RECT 5.330 2509.145 1694.370 2511.975 ;
        RECT 5.330 2503.705 1694.370 2506.535 ;
        RECT 5.330 2498.265 1694.370 2501.095 ;
        RECT 5.330 2492.825 1694.370 2495.655 ;
        RECT 5.330 2487.385 1694.370 2490.215 ;
        RECT 5.330 2481.945 1694.370 2484.775 ;
        RECT 5.330 2476.505 1694.370 2479.335 ;
        RECT 5.330 2471.065 1694.370 2473.895 ;
        RECT 5.330 2465.625 1694.370 2468.455 ;
        RECT 5.330 2460.185 1694.370 2463.015 ;
        RECT 5.330 2454.745 1694.370 2457.575 ;
        RECT 5.330 2449.305 1694.370 2452.135 ;
        RECT 5.330 2443.865 1694.370 2446.695 ;
        RECT 5.330 2438.425 1694.370 2441.255 ;
        RECT 5.330 2432.985 1694.370 2435.815 ;
        RECT 5.330 2427.545 1694.370 2430.375 ;
        RECT 5.330 2422.105 1694.370 2424.935 ;
        RECT 5.330 2416.665 1694.370 2419.495 ;
        RECT 5.330 2411.225 1694.370 2414.055 ;
        RECT 5.330 2405.785 1694.370 2408.615 ;
        RECT 5.330 2400.345 1694.370 2403.175 ;
        RECT 5.330 2394.905 1694.370 2397.735 ;
        RECT 5.330 2389.465 1694.370 2392.295 ;
        RECT 5.330 2384.025 1694.370 2386.855 ;
        RECT 5.330 2378.585 1694.370 2381.415 ;
        RECT 5.330 2373.145 1694.370 2375.975 ;
        RECT 5.330 2367.705 1694.370 2370.535 ;
        RECT 5.330 2362.265 1694.370 2365.095 ;
        RECT 5.330 2356.825 1694.370 2359.655 ;
        RECT 5.330 2351.385 1694.370 2354.215 ;
        RECT 5.330 2345.945 1694.370 2348.775 ;
        RECT 5.330 2340.505 1694.370 2343.335 ;
        RECT 5.330 2335.065 1694.370 2337.895 ;
        RECT 5.330 2329.625 1694.370 2332.455 ;
        RECT 5.330 2324.185 1694.370 2327.015 ;
        RECT 5.330 2318.745 1694.370 2321.575 ;
        RECT 5.330 2313.305 1694.370 2316.135 ;
        RECT 5.330 2307.865 1694.370 2310.695 ;
        RECT 5.330 2302.425 1694.370 2305.255 ;
        RECT 5.330 2296.985 1694.370 2299.815 ;
        RECT 5.330 2291.545 1694.370 2294.375 ;
        RECT 5.330 2286.105 1694.370 2288.935 ;
        RECT 5.330 2280.665 1694.370 2283.495 ;
        RECT 5.330 2275.225 1694.370 2278.055 ;
        RECT 5.330 2269.785 1694.370 2272.615 ;
        RECT 5.330 2264.345 1694.370 2267.175 ;
        RECT 5.330 2258.905 1694.370 2261.735 ;
        RECT 5.330 2253.465 1694.370 2256.295 ;
        RECT 5.330 2248.025 1694.370 2250.855 ;
        RECT 5.330 2242.585 1694.370 2245.415 ;
        RECT 5.330 2237.145 1694.370 2239.975 ;
        RECT 5.330 2231.705 1694.370 2234.535 ;
        RECT 5.330 2226.265 1694.370 2229.095 ;
        RECT 5.330 2220.825 1694.370 2223.655 ;
        RECT 5.330 2215.385 1694.370 2218.215 ;
        RECT 5.330 2209.945 1694.370 2212.775 ;
        RECT 5.330 2204.505 1694.370 2207.335 ;
        RECT 5.330 2199.065 1694.370 2201.895 ;
        RECT 5.330 2193.625 1694.370 2196.455 ;
        RECT 5.330 2188.185 1694.370 2191.015 ;
        RECT 5.330 2182.745 1694.370 2185.575 ;
        RECT 5.330 2177.305 1694.370 2180.135 ;
        RECT 5.330 2171.865 1694.370 2174.695 ;
        RECT 5.330 2166.425 1694.370 2169.255 ;
        RECT 5.330 2160.985 1694.370 2163.815 ;
        RECT 5.330 2155.545 1694.370 2158.375 ;
        RECT 5.330 2150.105 1694.370 2152.935 ;
        RECT 5.330 2144.665 1694.370 2147.495 ;
        RECT 5.330 2139.225 1694.370 2142.055 ;
        RECT 5.330 2133.785 1694.370 2136.615 ;
        RECT 5.330 2128.345 1694.370 2131.175 ;
        RECT 5.330 2122.905 1694.370 2125.735 ;
        RECT 5.330 2117.465 1694.370 2120.295 ;
        RECT 5.330 2112.025 1694.370 2114.855 ;
        RECT 5.330 2106.585 1694.370 2109.415 ;
        RECT 5.330 2101.145 1694.370 2103.975 ;
        RECT 5.330 2095.705 1694.370 2098.535 ;
        RECT 5.330 2090.265 1694.370 2093.095 ;
        RECT 5.330 2084.825 1694.370 2087.655 ;
        RECT 5.330 2079.385 1694.370 2082.215 ;
        RECT 5.330 2073.945 1694.370 2076.775 ;
        RECT 5.330 2068.505 1694.370 2071.335 ;
        RECT 5.330 2063.065 1694.370 2065.895 ;
        RECT 5.330 2057.625 1694.370 2060.455 ;
        RECT 5.330 2052.185 1694.370 2055.015 ;
        RECT 5.330 2046.745 1694.370 2049.575 ;
        RECT 5.330 2041.305 1694.370 2044.135 ;
        RECT 5.330 2035.865 1694.370 2038.695 ;
        RECT 5.330 2030.425 1694.370 2033.255 ;
        RECT 5.330 2024.985 1694.370 2027.815 ;
        RECT 5.330 2019.545 1694.370 2022.375 ;
        RECT 5.330 2014.105 1694.370 2016.935 ;
        RECT 5.330 2008.665 1694.370 2011.495 ;
        RECT 5.330 2003.225 1694.370 2006.055 ;
        RECT 5.330 1997.785 1694.370 2000.615 ;
        RECT 5.330 1992.345 1694.370 1995.175 ;
        RECT 5.330 1986.905 1694.370 1989.735 ;
        RECT 5.330 1981.465 1694.370 1984.295 ;
        RECT 5.330 1976.025 1694.370 1978.855 ;
        RECT 5.330 1970.585 1694.370 1973.415 ;
        RECT 5.330 1965.145 1694.370 1967.975 ;
        RECT 5.330 1959.705 1694.370 1962.535 ;
        RECT 5.330 1954.265 1694.370 1957.095 ;
        RECT 5.330 1948.825 1694.370 1951.655 ;
        RECT 5.330 1943.385 1694.370 1946.215 ;
        RECT 5.330 1937.945 1694.370 1940.775 ;
        RECT 5.330 1932.505 1694.370 1935.335 ;
        RECT 5.330 1927.065 1694.370 1929.895 ;
        RECT 5.330 1921.625 1694.370 1924.455 ;
        RECT 5.330 1916.185 1694.370 1919.015 ;
        RECT 5.330 1910.745 1694.370 1913.575 ;
        RECT 5.330 1905.305 1694.370 1908.135 ;
        RECT 5.330 1899.865 1694.370 1902.695 ;
        RECT 5.330 1894.425 1694.370 1897.255 ;
        RECT 5.330 1888.985 1694.370 1891.815 ;
        RECT 5.330 1883.545 1694.370 1886.375 ;
        RECT 5.330 1878.105 1694.370 1880.935 ;
        RECT 5.330 1872.665 1694.370 1875.495 ;
        RECT 5.330 1867.225 1694.370 1870.055 ;
        RECT 5.330 1861.785 1694.370 1864.615 ;
        RECT 5.330 1856.345 1694.370 1859.175 ;
        RECT 5.330 1850.905 1694.370 1853.735 ;
        RECT 5.330 1845.465 1694.370 1848.295 ;
        RECT 5.330 1840.025 1694.370 1842.855 ;
        RECT 5.330 1834.585 1694.370 1837.415 ;
        RECT 5.330 1829.145 1694.370 1831.975 ;
        RECT 5.330 1823.705 1694.370 1826.535 ;
        RECT 5.330 1818.265 1694.370 1821.095 ;
        RECT 5.330 1812.825 1694.370 1815.655 ;
        RECT 5.330 1807.385 1694.370 1810.215 ;
        RECT 5.330 1801.945 1694.370 1804.775 ;
        RECT 5.330 1796.505 1694.370 1799.335 ;
        RECT 5.330 1791.065 1694.370 1793.895 ;
        RECT 5.330 1785.625 1694.370 1788.455 ;
        RECT 5.330 1780.185 1694.370 1783.015 ;
        RECT 5.330 1774.745 1694.370 1777.575 ;
        RECT 5.330 1769.305 1694.370 1772.135 ;
        RECT 5.330 1763.865 1694.370 1766.695 ;
        RECT 5.330 1758.425 1694.370 1761.255 ;
        RECT 5.330 1752.985 1694.370 1755.815 ;
        RECT 5.330 1747.545 1694.370 1750.375 ;
        RECT 5.330 1742.105 1694.370 1744.935 ;
        RECT 5.330 1736.665 1694.370 1739.495 ;
        RECT 5.330 1731.225 1694.370 1734.055 ;
        RECT 5.330 1725.785 1694.370 1728.615 ;
        RECT 5.330 1720.345 1694.370 1723.175 ;
        RECT 5.330 1714.905 1694.370 1717.735 ;
        RECT 5.330 1709.465 1694.370 1712.295 ;
        RECT 5.330 1704.025 1694.370 1706.855 ;
        RECT 5.330 1698.585 1694.370 1701.415 ;
        RECT 5.330 1693.145 1694.370 1695.975 ;
        RECT 5.330 1687.705 1694.370 1690.535 ;
        RECT 5.330 1682.265 1694.370 1685.095 ;
        RECT 5.330 1676.825 1694.370 1679.655 ;
        RECT 5.330 1671.385 1694.370 1674.215 ;
        RECT 5.330 1665.945 1694.370 1668.775 ;
        RECT 5.330 1660.505 1694.370 1663.335 ;
        RECT 5.330 1655.065 1694.370 1657.895 ;
        RECT 5.330 1649.625 1694.370 1652.455 ;
        RECT 5.330 1644.185 1694.370 1647.015 ;
        RECT 5.330 1638.745 1694.370 1641.575 ;
        RECT 5.330 1633.305 1694.370 1636.135 ;
        RECT 5.330 1627.865 1694.370 1630.695 ;
        RECT 5.330 1622.425 1694.370 1625.255 ;
        RECT 5.330 1616.985 1694.370 1619.815 ;
        RECT 5.330 1611.545 1694.370 1614.375 ;
        RECT 5.330 1606.105 1694.370 1608.935 ;
        RECT 5.330 1600.665 1694.370 1603.495 ;
        RECT 5.330 1595.225 1694.370 1598.055 ;
        RECT 5.330 1589.785 1694.370 1592.615 ;
        RECT 5.330 1584.345 1694.370 1587.175 ;
        RECT 5.330 1578.905 1694.370 1581.735 ;
        RECT 5.330 1573.465 1694.370 1576.295 ;
        RECT 5.330 1568.025 1694.370 1570.855 ;
        RECT 5.330 1562.585 1694.370 1565.415 ;
        RECT 5.330 1557.145 1694.370 1559.975 ;
        RECT 5.330 1551.705 1694.370 1554.535 ;
        RECT 5.330 1546.265 1694.370 1549.095 ;
        RECT 5.330 1540.825 1694.370 1543.655 ;
        RECT 5.330 1535.385 1694.370 1538.215 ;
        RECT 5.330 1529.945 1694.370 1532.775 ;
        RECT 5.330 1524.505 1694.370 1527.335 ;
        RECT 5.330 1519.065 1694.370 1521.895 ;
        RECT 5.330 1513.625 1694.370 1516.455 ;
        RECT 5.330 1508.185 1694.370 1511.015 ;
        RECT 5.330 1502.745 1694.370 1505.575 ;
        RECT 5.330 1497.305 1694.370 1500.135 ;
        RECT 5.330 1491.865 1694.370 1494.695 ;
        RECT 5.330 1486.425 1694.370 1489.255 ;
        RECT 5.330 1480.985 1694.370 1483.815 ;
        RECT 5.330 1475.545 1694.370 1478.375 ;
        RECT 5.330 1470.105 1694.370 1472.935 ;
        RECT 5.330 1464.665 1694.370 1467.495 ;
        RECT 5.330 1459.225 1694.370 1462.055 ;
        RECT 5.330 1453.785 1694.370 1456.615 ;
        RECT 5.330 1448.345 1694.370 1451.175 ;
        RECT 5.330 1442.905 1694.370 1445.735 ;
        RECT 5.330 1437.465 1694.370 1440.295 ;
        RECT 5.330 1432.025 1694.370 1434.855 ;
        RECT 5.330 1426.585 1694.370 1429.415 ;
        RECT 5.330 1421.145 1694.370 1423.975 ;
        RECT 5.330 1415.705 1694.370 1418.535 ;
        RECT 5.330 1410.265 1694.370 1413.095 ;
        RECT 5.330 1404.825 1694.370 1407.655 ;
        RECT 5.330 1399.385 1694.370 1402.215 ;
        RECT 5.330 1393.945 1694.370 1396.775 ;
        RECT 5.330 1388.505 1694.370 1391.335 ;
        RECT 5.330 1383.065 1694.370 1385.895 ;
        RECT 5.330 1377.625 1694.370 1380.455 ;
        RECT 5.330 1372.185 1694.370 1375.015 ;
        RECT 5.330 1366.745 1694.370 1369.575 ;
        RECT 5.330 1361.305 1694.370 1364.135 ;
        RECT 5.330 1355.865 1694.370 1358.695 ;
        RECT 5.330 1350.425 1694.370 1353.255 ;
        RECT 5.330 1344.985 1694.370 1347.815 ;
        RECT 5.330 1339.545 1694.370 1342.375 ;
        RECT 5.330 1334.105 1694.370 1336.935 ;
        RECT 5.330 1328.665 1694.370 1331.495 ;
        RECT 5.330 1323.225 1694.370 1326.055 ;
        RECT 5.330 1317.785 1694.370 1320.615 ;
        RECT 5.330 1312.345 1694.370 1315.175 ;
        RECT 5.330 1306.905 1694.370 1309.735 ;
        RECT 5.330 1301.465 1694.370 1304.295 ;
        RECT 5.330 1296.025 1694.370 1298.855 ;
        RECT 5.330 1290.585 1694.370 1293.415 ;
        RECT 5.330 1285.145 1694.370 1287.975 ;
        RECT 5.330 1279.705 1694.370 1282.535 ;
        RECT 5.330 1274.265 1694.370 1277.095 ;
        RECT 5.330 1268.825 1694.370 1271.655 ;
        RECT 5.330 1263.385 1694.370 1266.215 ;
        RECT 5.330 1257.945 1694.370 1260.775 ;
        RECT 5.330 1252.505 1694.370 1255.335 ;
        RECT 5.330 1247.065 1694.370 1249.895 ;
        RECT 5.330 1241.625 1694.370 1244.455 ;
        RECT 5.330 1236.185 1694.370 1239.015 ;
        RECT 5.330 1230.745 1694.370 1233.575 ;
        RECT 5.330 1225.305 1694.370 1228.135 ;
        RECT 5.330 1219.865 1694.370 1222.695 ;
        RECT 5.330 1214.425 1694.370 1217.255 ;
        RECT 5.330 1208.985 1694.370 1211.815 ;
        RECT 5.330 1203.545 1694.370 1206.375 ;
        RECT 5.330 1198.105 1694.370 1200.935 ;
        RECT 5.330 1192.665 1694.370 1195.495 ;
        RECT 5.330 1187.225 1694.370 1190.055 ;
        RECT 5.330 1181.785 1694.370 1184.615 ;
        RECT 5.330 1176.345 1694.370 1179.175 ;
        RECT 5.330 1170.905 1694.370 1173.735 ;
        RECT 5.330 1165.465 1694.370 1168.295 ;
        RECT 5.330 1160.025 1694.370 1162.855 ;
        RECT 5.330 1154.585 1694.370 1157.415 ;
        RECT 5.330 1149.145 1694.370 1151.975 ;
        RECT 5.330 1143.705 1694.370 1146.535 ;
        RECT 5.330 1138.265 1694.370 1141.095 ;
        RECT 5.330 1132.825 1694.370 1135.655 ;
        RECT 5.330 1127.385 1694.370 1130.215 ;
        RECT 5.330 1121.945 1694.370 1124.775 ;
        RECT 5.330 1116.505 1694.370 1119.335 ;
        RECT 5.330 1111.065 1694.370 1113.895 ;
        RECT 5.330 1105.625 1694.370 1108.455 ;
        RECT 5.330 1100.185 1694.370 1103.015 ;
        RECT 5.330 1094.745 1694.370 1097.575 ;
        RECT 5.330 1089.305 1694.370 1092.135 ;
        RECT 5.330 1083.865 1694.370 1086.695 ;
        RECT 5.330 1078.425 1694.370 1081.255 ;
        RECT 5.330 1072.985 1694.370 1075.815 ;
        RECT 5.330 1067.545 1694.370 1070.375 ;
        RECT 5.330 1062.105 1694.370 1064.935 ;
        RECT 5.330 1056.665 1694.370 1059.495 ;
        RECT 5.330 1051.225 1694.370 1054.055 ;
        RECT 5.330 1045.785 1694.370 1048.615 ;
        RECT 5.330 1040.345 1694.370 1043.175 ;
        RECT 5.330 1034.905 1694.370 1037.735 ;
        RECT 5.330 1029.465 1694.370 1032.295 ;
        RECT 5.330 1024.025 1694.370 1026.855 ;
        RECT 5.330 1018.585 1694.370 1021.415 ;
        RECT 5.330 1013.145 1694.370 1015.975 ;
        RECT 5.330 1007.705 1694.370 1010.535 ;
        RECT 5.330 1002.265 1694.370 1005.095 ;
        RECT 5.330 996.825 1694.370 999.655 ;
        RECT 5.330 991.385 1694.370 994.215 ;
        RECT 5.330 985.945 1694.370 988.775 ;
        RECT 5.330 980.505 1694.370 983.335 ;
        RECT 5.330 975.065 1694.370 977.895 ;
        RECT 5.330 969.625 1694.370 972.455 ;
        RECT 5.330 964.185 1694.370 967.015 ;
        RECT 5.330 958.745 1694.370 961.575 ;
        RECT 5.330 953.305 1694.370 956.135 ;
        RECT 5.330 947.865 1694.370 950.695 ;
        RECT 5.330 942.425 1694.370 945.255 ;
        RECT 5.330 936.985 1694.370 939.815 ;
        RECT 5.330 931.545 1694.370 934.375 ;
        RECT 5.330 926.105 1694.370 928.935 ;
        RECT 5.330 920.665 1694.370 923.495 ;
        RECT 5.330 915.225 1694.370 918.055 ;
        RECT 5.330 909.785 1694.370 912.615 ;
        RECT 5.330 904.345 1694.370 907.175 ;
        RECT 5.330 898.905 1694.370 901.735 ;
        RECT 5.330 893.465 1694.370 896.295 ;
        RECT 5.330 888.025 1694.370 890.855 ;
        RECT 5.330 882.585 1694.370 885.415 ;
        RECT 5.330 877.145 1694.370 879.975 ;
        RECT 5.330 871.705 1694.370 874.535 ;
        RECT 5.330 866.265 1694.370 869.095 ;
        RECT 5.330 860.825 1694.370 863.655 ;
        RECT 5.330 855.385 1694.370 858.215 ;
        RECT 5.330 849.945 1694.370 852.775 ;
        RECT 5.330 844.505 1694.370 847.335 ;
        RECT 5.330 839.065 1694.370 841.895 ;
        RECT 5.330 833.625 1694.370 836.455 ;
        RECT 5.330 828.185 1694.370 831.015 ;
        RECT 5.330 822.745 1694.370 825.575 ;
        RECT 5.330 817.305 1694.370 820.135 ;
        RECT 5.330 811.865 1694.370 814.695 ;
        RECT 5.330 806.425 1694.370 809.255 ;
        RECT 5.330 800.985 1694.370 803.815 ;
        RECT 5.330 795.545 1694.370 798.375 ;
        RECT 5.330 790.105 1694.370 792.935 ;
        RECT 5.330 784.665 1694.370 787.495 ;
        RECT 5.330 779.225 1694.370 782.055 ;
        RECT 5.330 773.785 1694.370 776.615 ;
        RECT 5.330 768.345 1694.370 771.175 ;
        RECT 5.330 762.905 1694.370 765.735 ;
        RECT 5.330 757.465 1694.370 760.295 ;
        RECT 5.330 752.025 1694.370 754.855 ;
        RECT 5.330 746.585 1694.370 749.415 ;
        RECT 5.330 741.145 1694.370 743.975 ;
        RECT 5.330 735.705 1694.370 738.535 ;
        RECT 5.330 730.265 1694.370 733.095 ;
        RECT 5.330 724.825 1694.370 727.655 ;
        RECT 5.330 719.385 1694.370 722.215 ;
        RECT 5.330 713.945 1694.370 716.775 ;
        RECT 5.330 708.505 1694.370 711.335 ;
        RECT 5.330 703.065 1694.370 705.895 ;
        RECT 5.330 697.625 1694.370 700.455 ;
        RECT 5.330 692.185 1694.370 695.015 ;
        RECT 5.330 686.745 1694.370 689.575 ;
        RECT 5.330 681.305 1694.370 684.135 ;
        RECT 5.330 675.865 1694.370 678.695 ;
        RECT 5.330 670.425 1694.370 673.255 ;
        RECT 5.330 664.985 1694.370 667.815 ;
        RECT 5.330 659.545 1694.370 662.375 ;
        RECT 5.330 654.105 1694.370 656.935 ;
        RECT 5.330 648.665 1694.370 651.495 ;
        RECT 5.330 643.225 1694.370 646.055 ;
        RECT 5.330 637.785 1694.370 640.615 ;
        RECT 5.330 632.345 1694.370 635.175 ;
        RECT 5.330 626.905 1694.370 629.735 ;
        RECT 5.330 621.465 1694.370 624.295 ;
        RECT 5.330 616.025 1694.370 618.855 ;
        RECT 5.330 610.585 1694.370 613.415 ;
        RECT 5.330 605.145 1694.370 607.975 ;
        RECT 5.330 599.705 1694.370 602.535 ;
        RECT 5.330 594.265 1694.370 597.095 ;
        RECT 5.330 588.825 1694.370 591.655 ;
        RECT 5.330 583.385 1694.370 586.215 ;
        RECT 5.330 577.945 1694.370 580.775 ;
        RECT 5.330 572.505 1694.370 575.335 ;
        RECT 5.330 567.065 1694.370 569.895 ;
        RECT 5.330 561.625 1694.370 564.455 ;
        RECT 5.330 556.185 1694.370 559.015 ;
        RECT 5.330 550.745 1694.370 553.575 ;
        RECT 5.330 545.305 1694.370 548.135 ;
        RECT 5.330 539.865 1694.370 542.695 ;
        RECT 5.330 534.425 1694.370 537.255 ;
        RECT 5.330 528.985 1694.370 531.815 ;
        RECT 5.330 523.545 1694.370 526.375 ;
        RECT 5.330 518.105 1694.370 520.935 ;
        RECT 5.330 512.665 1694.370 515.495 ;
        RECT 5.330 507.225 1694.370 510.055 ;
        RECT 5.330 501.785 1694.370 504.615 ;
        RECT 5.330 496.345 1694.370 499.175 ;
        RECT 5.330 490.905 1694.370 493.735 ;
        RECT 5.330 485.465 1694.370 488.295 ;
        RECT 5.330 480.025 1694.370 482.855 ;
        RECT 5.330 474.585 1694.370 477.415 ;
        RECT 5.330 469.145 1694.370 471.975 ;
        RECT 5.330 463.705 1694.370 466.535 ;
        RECT 5.330 458.265 1694.370 461.095 ;
        RECT 5.330 452.825 1694.370 455.655 ;
        RECT 5.330 447.385 1694.370 450.215 ;
        RECT 5.330 441.945 1694.370 444.775 ;
        RECT 5.330 436.505 1694.370 439.335 ;
        RECT 5.330 431.065 1694.370 433.895 ;
        RECT 5.330 425.625 1694.370 428.455 ;
        RECT 5.330 420.185 1694.370 423.015 ;
        RECT 5.330 414.745 1694.370 417.575 ;
        RECT 5.330 409.305 1694.370 412.135 ;
        RECT 5.330 403.865 1694.370 406.695 ;
        RECT 5.330 398.425 1694.370 401.255 ;
        RECT 5.330 392.985 1694.370 395.815 ;
        RECT 5.330 387.545 1694.370 390.375 ;
        RECT 5.330 382.105 1694.370 384.935 ;
        RECT 5.330 376.665 1694.370 379.495 ;
        RECT 5.330 371.225 1694.370 374.055 ;
        RECT 5.330 365.785 1694.370 368.615 ;
        RECT 5.330 360.345 1694.370 363.175 ;
        RECT 5.330 354.905 1694.370 357.735 ;
        RECT 5.330 349.465 1694.370 352.295 ;
        RECT 5.330 344.025 1694.370 346.855 ;
        RECT 5.330 338.585 1694.370 341.415 ;
        RECT 5.330 333.145 1694.370 335.975 ;
        RECT 5.330 327.705 1694.370 330.535 ;
        RECT 5.330 322.265 1694.370 325.095 ;
        RECT 5.330 316.825 1694.370 319.655 ;
        RECT 5.330 311.385 1694.370 314.215 ;
        RECT 5.330 305.945 1694.370 308.775 ;
        RECT 5.330 300.505 1694.370 303.335 ;
        RECT 5.330 295.065 1694.370 297.895 ;
        RECT 5.330 289.625 1694.370 292.455 ;
        RECT 5.330 284.185 1694.370 287.015 ;
        RECT 5.330 278.745 1694.370 281.575 ;
        RECT 5.330 273.305 1694.370 276.135 ;
        RECT 5.330 267.865 1694.370 270.695 ;
        RECT 5.330 262.425 1694.370 265.255 ;
        RECT 5.330 256.985 1694.370 259.815 ;
        RECT 5.330 251.545 1694.370 254.375 ;
        RECT 5.330 246.105 1694.370 248.935 ;
        RECT 5.330 240.665 1694.370 243.495 ;
        RECT 5.330 235.225 1694.370 238.055 ;
        RECT 5.330 229.785 1694.370 232.615 ;
        RECT 5.330 224.345 1694.370 227.175 ;
        RECT 5.330 218.905 1694.370 221.735 ;
        RECT 5.330 213.465 1694.370 216.295 ;
        RECT 5.330 208.025 1694.370 210.855 ;
        RECT 5.330 202.585 1694.370 205.415 ;
        RECT 5.330 197.145 1694.370 199.975 ;
        RECT 5.330 191.705 1694.370 194.535 ;
        RECT 5.330 186.265 1694.370 189.095 ;
        RECT 5.330 180.825 1694.370 183.655 ;
        RECT 5.330 175.385 1694.370 178.215 ;
        RECT 5.330 169.945 1694.370 172.775 ;
        RECT 5.330 164.505 1694.370 167.335 ;
        RECT 5.330 159.065 1694.370 161.895 ;
        RECT 5.330 153.625 1694.370 156.455 ;
        RECT 5.330 148.185 1694.370 151.015 ;
        RECT 5.330 142.745 1694.370 145.575 ;
        RECT 5.330 137.305 1694.370 140.135 ;
        RECT 5.330 131.865 1694.370 134.695 ;
        RECT 5.330 126.425 1694.370 129.255 ;
        RECT 5.330 120.985 1694.370 123.815 ;
        RECT 5.330 115.545 1694.370 118.375 ;
        RECT 5.330 110.105 1694.370 112.935 ;
        RECT 5.330 104.665 1694.370 107.495 ;
        RECT 5.330 99.225 1694.370 102.055 ;
        RECT 5.330 93.785 1694.370 96.615 ;
        RECT 5.330 88.345 1694.370 91.175 ;
        RECT 5.330 82.905 1694.370 85.735 ;
        RECT 5.330 77.465 1694.370 80.295 ;
        RECT 5.330 72.025 1694.370 74.855 ;
        RECT 5.330 66.585 1694.370 69.415 ;
        RECT 5.330 61.145 1694.370 63.975 ;
        RECT 5.330 55.705 1694.370 58.535 ;
        RECT 5.330 50.265 1694.370 53.095 ;
        RECT 5.330 44.825 1694.370 47.655 ;
        RECT 5.330 39.385 1694.370 42.215 ;
        RECT 5.330 33.945 1694.370 36.775 ;
        RECT 5.330 28.505 1694.370 31.335 ;
        RECT 5.330 23.065 1694.370 25.895 ;
        RECT 5.330 17.625 1694.370 20.455 ;
        RECT 5.330 12.185 1694.370 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 1694.180 3187.925 ;
      LAYER met1 ;
        RECT 5.520 10.640 1696.870 3188.080 ;
      LAYER met2 ;
        RECT 7.920 10.695 1696.840 3188.025 ;
      LAYER met3 ;
        RECT 21.050 3170.520 1696.000 3188.005 ;
        RECT 21.050 3169.120 1695.600 3170.520 ;
        RECT 21.050 3115.440 1696.000 3169.120 ;
        RECT 21.050 3114.040 1695.600 3115.440 ;
        RECT 21.050 3060.360 1696.000 3114.040 ;
        RECT 21.050 3058.960 1695.600 3060.360 ;
        RECT 21.050 3005.280 1696.000 3058.960 ;
        RECT 21.050 3003.880 1695.600 3005.280 ;
        RECT 21.050 2950.200 1696.000 3003.880 ;
        RECT 21.050 2948.800 1695.600 2950.200 ;
        RECT 21.050 2895.120 1696.000 2948.800 ;
        RECT 21.050 2893.720 1695.600 2895.120 ;
        RECT 21.050 2840.040 1696.000 2893.720 ;
        RECT 21.050 2838.640 1695.600 2840.040 ;
        RECT 21.050 2784.960 1696.000 2838.640 ;
        RECT 21.050 2783.560 1695.600 2784.960 ;
        RECT 21.050 2729.880 1696.000 2783.560 ;
        RECT 21.050 2728.480 1695.600 2729.880 ;
        RECT 21.050 2674.800 1696.000 2728.480 ;
        RECT 21.050 2673.400 1695.600 2674.800 ;
        RECT 21.050 2619.720 1696.000 2673.400 ;
        RECT 21.050 2618.320 1695.600 2619.720 ;
        RECT 21.050 2564.640 1696.000 2618.320 ;
        RECT 21.050 2563.240 1695.600 2564.640 ;
        RECT 21.050 2509.560 1696.000 2563.240 ;
        RECT 21.050 2508.160 1695.600 2509.560 ;
        RECT 21.050 2454.480 1696.000 2508.160 ;
        RECT 21.050 2453.080 1695.600 2454.480 ;
        RECT 21.050 2399.400 1696.000 2453.080 ;
        RECT 21.050 2398.000 1695.600 2399.400 ;
        RECT 21.050 2344.320 1696.000 2398.000 ;
        RECT 21.050 2342.920 1695.600 2344.320 ;
        RECT 21.050 2289.240 1696.000 2342.920 ;
        RECT 21.050 2287.840 1695.600 2289.240 ;
        RECT 21.050 2234.160 1696.000 2287.840 ;
        RECT 21.050 2232.760 1695.600 2234.160 ;
        RECT 21.050 2179.080 1696.000 2232.760 ;
        RECT 21.050 2177.680 1695.600 2179.080 ;
        RECT 21.050 2124.000 1696.000 2177.680 ;
        RECT 21.050 2122.600 1695.600 2124.000 ;
        RECT 21.050 2068.920 1696.000 2122.600 ;
        RECT 21.050 2067.520 1695.600 2068.920 ;
        RECT 21.050 2013.840 1696.000 2067.520 ;
        RECT 21.050 2012.440 1695.600 2013.840 ;
        RECT 21.050 1958.760 1696.000 2012.440 ;
        RECT 21.050 1957.360 1695.600 1958.760 ;
        RECT 21.050 1903.680 1696.000 1957.360 ;
        RECT 21.050 1902.280 1695.600 1903.680 ;
        RECT 21.050 1848.600 1696.000 1902.280 ;
        RECT 21.050 1847.200 1695.600 1848.600 ;
        RECT 21.050 1793.520 1696.000 1847.200 ;
        RECT 21.050 1792.120 1695.600 1793.520 ;
        RECT 21.050 1738.440 1696.000 1792.120 ;
        RECT 21.050 1737.040 1695.600 1738.440 ;
        RECT 21.050 1683.360 1696.000 1737.040 ;
        RECT 21.050 1681.960 1695.600 1683.360 ;
        RECT 21.050 1628.280 1696.000 1681.960 ;
        RECT 21.050 1626.880 1695.600 1628.280 ;
        RECT 21.050 1573.200 1696.000 1626.880 ;
        RECT 21.050 1571.800 1695.600 1573.200 ;
        RECT 21.050 1518.120 1696.000 1571.800 ;
        RECT 21.050 1516.720 1695.600 1518.120 ;
        RECT 21.050 1463.040 1696.000 1516.720 ;
        RECT 21.050 1461.640 1695.600 1463.040 ;
        RECT 21.050 1407.960 1696.000 1461.640 ;
        RECT 21.050 1406.560 1695.600 1407.960 ;
        RECT 21.050 1352.880 1696.000 1406.560 ;
        RECT 21.050 1351.480 1695.600 1352.880 ;
        RECT 21.050 1297.800 1696.000 1351.480 ;
        RECT 21.050 1296.400 1695.600 1297.800 ;
        RECT 21.050 1242.720 1696.000 1296.400 ;
        RECT 21.050 1241.320 1695.600 1242.720 ;
        RECT 21.050 1187.640 1696.000 1241.320 ;
        RECT 21.050 1186.240 1695.600 1187.640 ;
        RECT 21.050 1132.560 1696.000 1186.240 ;
        RECT 21.050 1131.160 1695.600 1132.560 ;
        RECT 21.050 1077.480 1696.000 1131.160 ;
        RECT 21.050 1076.080 1695.600 1077.480 ;
        RECT 21.050 1022.400 1696.000 1076.080 ;
        RECT 21.050 1021.000 1695.600 1022.400 ;
        RECT 21.050 967.320 1696.000 1021.000 ;
        RECT 21.050 965.920 1695.600 967.320 ;
        RECT 21.050 912.240 1696.000 965.920 ;
        RECT 21.050 910.840 1695.600 912.240 ;
        RECT 21.050 857.160 1696.000 910.840 ;
        RECT 21.050 855.760 1695.600 857.160 ;
        RECT 21.050 802.080 1696.000 855.760 ;
        RECT 21.050 800.680 1695.600 802.080 ;
        RECT 21.050 747.000 1696.000 800.680 ;
        RECT 21.050 745.600 1695.600 747.000 ;
        RECT 21.050 691.920 1696.000 745.600 ;
        RECT 21.050 690.520 1695.600 691.920 ;
        RECT 21.050 636.840 1696.000 690.520 ;
        RECT 21.050 635.440 1695.600 636.840 ;
        RECT 21.050 581.760 1696.000 635.440 ;
        RECT 21.050 580.360 1695.600 581.760 ;
        RECT 21.050 526.680 1696.000 580.360 ;
        RECT 21.050 525.280 1695.600 526.680 ;
        RECT 21.050 471.600 1696.000 525.280 ;
        RECT 21.050 470.200 1695.600 471.600 ;
        RECT 21.050 416.520 1696.000 470.200 ;
        RECT 21.050 415.120 1695.600 416.520 ;
        RECT 21.050 361.440 1696.000 415.120 ;
        RECT 21.050 360.040 1695.600 361.440 ;
        RECT 21.050 306.360 1696.000 360.040 ;
        RECT 21.050 304.960 1695.600 306.360 ;
        RECT 21.050 251.280 1696.000 304.960 ;
        RECT 21.050 249.880 1695.600 251.280 ;
        RECT 21.050 196.200 1696.000 249.880 ;
        RECT 21.050 194.800 1695.600 196.200 ;
        RECT 21.050 141.120 1696.000 194.800 ;
        RECT 21.050 139.720 1695.600 141.120 ;
        RECT 21.050 86.040 1696.000 139.720 ;
        RECT 21.050 84.640 1695.600 86.040 ;
        RECT 21.050 30.960 1696.000 84.640 ;
        RECT 21.050 29.560 1695.600 30.960 ;
        RECT 21.050 10.715 1696.000 29.560 ;
      LAYER met4 ;
        RECT 61.015 32.135 97.440 3136.665 ;
        RECT 99.840 32.135 174.240 3136.665 ;
        RECT 176.640 32.135 251.040 3136.665 ;
        RECT 253.440 32.135 327.840 3136.665 ;
        RECT 330.240 32.135 404.640 3136.665 ;
        RECT 407.040 32.135 481.440 3136.665 ;
        RECT 483.840 32.135 558.240 3136.665 ;
        RECT 560.640 32.135 635.040 3136.665 ;
        RECT 637.440 32.135 711.840 3136.665 ;
        RECT 714.240 32.135 788.640 3136.665 ;
        RECT 791.040 32.135 865.440 3136.665 ;
        RECT 867.840 32.135 942.240 3136.665 ;
        RECT 944.640 32.135 1019.040 3136.665 ;
        RECT 1021.440 32.135 1095.840 3136.665 ;
        RECT 1098.240 32.135 1172.640 3136.665 ;
        RECT 1175.040 32.135 1249.440 3136.665 ;
        RECT 1251.840 32.135 1326.240 3136.665 ;
        RECT 1328.640 32.135 1403.040 3136.665 ;
        RECT 1405.440 32.135 1479.840 3136.665 ;
        RECT 1482.240 32.135 1556.640 3136.665 ;
        RECT 1559.040 32.135 1633.440 3136.665 ;
        RECT 1635.840 32.135 1684.225 3136.665 ;
  END
END wrapped_as512512512
END LIBRARY

