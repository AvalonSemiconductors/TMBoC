* NGSPICE file created from posit_unit.ext - technology: sky130B

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_2 abstract view
.subckt sky130_fd_sc_hd__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_1 abstract view
.subckt sky130_fd_sc_hd__nor2b_1 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_2 abstract view
.subckt sky130_fd_sc_hd__nor4b_2 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_2 abstract view
.subckt sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_4 abstract view
.subckt sky130_fd_sc_hd__a2111oi_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_1 abstract view
.subckt sky130_fd_sc_hd__o32ai_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

.subckt posit_unit clk io_in[0] io_in[1] io_in[2] io_out[0] io_out[1] io_out[2] io_out[3]
+ rst vccd1 vssd1
XFILLER_100_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4935__A _4045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7963_ _3120_ _3146_ _3065_ vssd1 vssd1 vccd1 vccd1 _3147_ sky130_fd_sc_hd__mux2_1
XFILLER_39_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6914_ _1929_ _1938_ vssd1 vssd1 vccd1 vccd1 _1993_ sky130_fd_sc_hd__xnor2_1
XFILLER_54_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7894_ _3040_ vssd1 vssd1 vccd1 vccd1 _3071_ sky130_fd_sc_hd__clkinv_2
X_6845_ _1904_ _1910_ vssd1 vssd1 vccd1 vccd1 _1917_ sky130_fd_sc_hd__and2b_1
XFILLER_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6776_ _1801_ _1828_ vssd1 vssd1 vccd1 vccd1 _1841_ sky130_fd_sc_hd__xnor2_1
XFILLER_50_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5727_ _3866_ _0706_ _0703_ vssd1 vssd1 vccd1 vccd1 _0707_ sky130_fd_sc_hd__a21o_1
X_8515_ clknet_3_3__leaf_clk _0001_ vssd1 vssd1 vccd1 vccd1 cmd\[6\] sky130_fd_sc_hd__dfxtp_4
X_8446_ _3654_ vssd1 vssd1 vccd1 vccd1 _3655_ sky130_fd_sc_hd__buf_4
X_5658_ _3923_ _0628_ _0629_ _0630_ vssd1 vssd1 vccd1 vccd1 _0631_ sky130_fd_sc_hd__a31o_2
X_4609_ _3763_ _3702_ vssd1 vssd1 vccd1 vccd1 _3764_ sky130_fd_sc_hd__or2_1
X_8377_ _3547_ _3556_ _1319_ vssd1 vssd1 vccd1 vccd1 _3589_ sky130_fd_sc_hd__o21ai_1
X_5589_ _0533_ _0541_ _0480_ vssd1 vssd1 vccd1 vccd1 _0562_ sky130_fd_sc_hd__mux2_1
X_7328_ _2403_ _2404_ vssd1 vssd1 vccd1 vccd1 _2448_ sky130_fd_sc_hd__xor2_1
XFILLER_117_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7259_ _2371_ vssd1 vssd1 vccd1 vccd1 _2372_ sky130_fd_sc_hd__inv_2
XFILLER_104_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6136__A1 _0627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5895__B1 _3832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5111__A2 _0082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4960_ _4096_ _4114_ vssd1 vssd1 vccd1 vccd1 _4115_ sky130_fd_sc_hd__xnor2_1
X_4891_ _4045_ _3986_ vssd1 vssd1 vccd1 vccd1 _4046_ sky130_fd_sc_hd__nand2_1
X_6630_ _1677_ _1678_ vssd1 vssd1 vccd1 vccd1 _1680_ sky130_fd_sc_hd__or2_1
X_6561_ _1595_ _1597_ _1602_ vssd1 vssd1 vccd1 vccd1 _1604_ sky130_fd_sc_hd__or3_1
X_5512_ _0250_ _0325_ vssd1 vssd1 vccd1 vccd1 _0485_ sky130_fd_sc_hd__xor2_1
XFILLER_9_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8300_ _3481_ _3505_ _3499_ vssd1 vssd1 vccd1 vccd1 _3507_ sky130_fd_sc_hd__or3_1
XFILLER_118_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6492_ _1526_ _1527_ vssd1 vssd1 vccd1 vccd1 _1529_ sky130_fd_sc_hd__and2b_1
XFILLER_118_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8231_ _3427_ _3433_ _0600_ vssd1 vssd1 vccd1 vccd1 _3434_ sky130_fd_sc_hd__a21oi_1
X_5443_ _0415_ vssd1 vssd1 vccd1 vccd1 _0416_ sky130_fd_sc_hd__inv_2
X_8162_ _0570_ vssd1 vssd1 vccd1 vccd1 _3361_ sky130_fd_sc_hd__clkinv_2
X_5374_ _1781_ vssd1 vssd1 vccd1 vccd1 _0347_ sky130_fd_sc_hd__inv_2
XFILLER_99_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7113_ _2207_ _2211_ vssd1 vssd1 vccd1 vccd1 _2212_ sky130_fd_sc_hd__nand2_1
XFILLER_87_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4325_ posit_add.in2\[7\] posit_add.in2\[5\] posit_add.in2\[4\] posit_add.in2\[6\]
+ vssd1 vssd1 vccd1 vccd1 _1363_ sky130_fd_sc_hd__or4_1
XFILLER_113_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8093_ _2486_ _2614_ _3286_ vssd1 vssd1 vccd1 vccd1 _3287_ sky130_fd_sc_hd__o21a_1
XFILLER_101_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7044_ _1454_ _1531_ _1537_ _2086_ vssd1 vssd1 vccd1 vccd1 _2136_ sky130_fd_sc_hd__or4_1
XFILLER_95_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6850__A2 _1531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7946_ _3126_ _3127_ _3038_ _3089_ vssd1 vssd1 vccd1 vccd1 _3128_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_42_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7877_ _2923_ _2932_ _2971_ vssd1 vssd1 vccd1 vccd1 _3052_ sky130_fd_sc_hd__mux2_1
X_6828_ _1761_ _1897_ vssd1 vssd1 vccd1 vccd1 _1898_ sky130_fd_sc_hd__nand2_1
XFILLER_50_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6759_ _1804_ _1821_ vssd1 vssd1 vccd1 vccd1 _1822_ sky130_fd_sc_hd__xor2_1
XFILLER_109_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8429_ _0679_ _3639_ vssd1 vssd1 vccd1 vccd1 _3641_ sky130_fd_sc_hd__nor2_1
XFILLER_2_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4741__C _3838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6949__B _1538_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7306__B1 _2335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5090_ _4243_ _4244_ vssd1 vssd1 vccd1 vccd1 _4245_ sky130_fd_sc_hd__and2_1
XFILLER_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4843__A1 _3881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5992_ _0984_ _0987_ _0985_ vssd1 vssd1 vccd1 vccd1 _0989_ sky130_fd_sc_hd__o21a_1
XFILLER_92_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7800_ _2898_ _2901_ _2894_ vssd1 vssd1 vccd1 vccd1 _2967_ sky130_fd_sc_hd__o21a_1
XFILLER_25_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4943_ _4072_ _4088_ vssd1 vssd1 vccd1 vccd1 _4098_ sky130_fd_sc_hd__and2_1
XFILLER_17_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7731_ _2842_ _2890_ vssd1 vssd1 vccd1 vccd1 _2891_ sky130_fd_sc_hd__or2b_1
X_7662_ _2788_ _2789_ vssd1 vssd1 vccd1 vccd1 _2816_ sky130_fd_sc_hd__nor2_1
XFILLER_32_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6613_ _1301_ _1300_ vssd1 vssd1 vccd1 vccd1 _1662_ sky130_fd_sc_hd__and2_1
X_4874_ _3890_ _3913_ vssd1 vssd1 vccd1 vccd1 _4029_ sky130_fd_sc_hd__and2b_1
XFILLER_60_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7593_ _0113_ _4153_ _2721_ vssd1 vssd1 vccd1 vccd1 _2740_ sky130_fd_sc_hd__mux2_2
X_6544_ _1468_ _1471_ vssd1 vssd1 vccd1 vccd1 _1586_ sky130_fd_sc_hd__nand2_1
X_6475_ _1509_ vssd1 vssd1 vccd1 vccd1 _1510_ sky130_fd_sc_hd__buf_4
XFILLER_118_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8214_ _2491_ _2611_ vssd1 vssd1 vccd1 vccd1 _3416_ sky130_fd_sc_hd__nor2_4
X_5426_ _3328_ _1781_ vssd1 vssd1 vccd1 vccd1 _0399_ sky130_fd_sc_hd__nand2_2
XANTENNA__4379__B _1946_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8145_ _3166_ _3336_ _3342_ vssd1 vssd1 vccd1 vccd1 _3343_ sky130_fd_sc_hd__o21a_1
X_5357_ _0328_ _0329_ vssd1 vssd1 vccd1 vccd1 _0330_ sky130_fd_sc_hd__and2b_1
XFILLER_101_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5288_ _4163_ _4162_ vssd1 vssd1 vccd1 vccd1 _0261_ sky130_fd_sc_hd__and2b_1
X_4308_ _0701_ vssd1 vssd1 vccd1 vccd1 _1177_ sky130_fd_sc_hd__buf_4
X_8076_ _0600_ _3268_ vssd1 vssd1 vccd1 vccd1 _3269_ sky130_fd_sc_hd__nor2_1
X_7027_ _2116_ _2080_ vssd1 vssd1 vccd1 vccd1 _2117_ sky130_fd_sc_hd__xor2_1
XFILLER_87_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5003__B _3930_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7929_ _2899_ _2906_ _2971_ vssd1 vssd1 vccd1 vccd1 _3109_ sky130_fd_sc_hd__mux2_1
XANTENNA__6115__A _4017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8264__B2 _0600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5250__A1 _3988_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5864__A _3815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4590_ _3339_ _3349_ _2936_ _3360_ vssd1 vssd1 vccd1 vccd1 _3745_ sky130_fd_sc_hd__o211a_1
X_6260_ _1261_ _1272_ vssd1 vssd1 vccd1 vccd1 _1273_ sky130_fd_sc_hd__xnor2_1
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6191_ _0779_ _0992_ vssd1 vssd1 vccd1 vccd1 _1198_ sky130_fd_sc_hd__nor2_1
X_5211_ _4017_ _3930_ vssd1 vssd1 vccd1 vccd1 _0184_ sky130_fd_sc_hd__nor2_2
XFILLER_69_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5142_ _0104_ _0110_ vssd1 vssd1 vccd1 vccd1 _0115_ sky130_fd_sc_hd__xor2_1
XFILLER_111_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5073_ _3827_ vssd1 vssd1 vccd1 vccd1 _4228_ sky130_fd_sc_hd__buf_4
XFILLER_56_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5975_ _0968_ _0969_ _0970_ vssd1 vssd1 vccd1 vccd1 _0971_ sky130_fd_sc_hd__and3_1
XFILLER_80_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4926_ _4058_ _4059_ vssd1 vssd1 vccd1 vccd1 _4081_ sky130_fd_sc_hd__xor2_1
XFILLER_21_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7714_ _2796_ _2798_ _2800_ vssd1 vssd1 vccd1 vccd1 _2873_ sky130_fd_sc_hd__a21o_1
XFILLER_40_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4857_ _3929_ _3931_ vssd1 vssd1 vccd1 vccd1 _4012_ sky130_fd_sc_hd__and2_1
X_7645_ _2676_ _2731_ _2732_ vssd1 vssd1 vccd1 vccd1 _2797_ sky130_fd_sc_hd__and3_1
XFILLER_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7576_ _2713_ vssd1 vssd1 vccd1 vccd1 _2721_ sky130_fd_sc_hd__buf_4
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6527_ _0080_ _1510_ vssd1 vssd1 vccd1 vccd1 _1567_ sky130_fd_sc_hd__nor2_2
X_4788_ _3722_ _3754_ vssd1 vssd1 vccd1 vccd1 _3943_ sky130_fd_sc_hd__and2_1
XFILLER_119_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8494__A1 in_reg\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6458_ _1469_ _1470_ vssd1 vssd1 vccd1 vccd1 _1491_ sky130_fd_sc_hd__xnor2_1
X_6389_ _4217_ _1414_ vssd1 vssd1 vccd1 vccd1 _1415_ sky130_fd_sc_hd__nand2_1
X_5409_ _2309_ _0359_ _0381_ vssd1 vssd1 vccd1 vccd1 _0382_ sky130_fd_sc_hd__o21a_1
X_8128_ _3166_ _3323_ vssd1 vssd1 vccd1 vccd1 _3324_ sky130_fd_sc_hd__or2_1
XFILLER_114_391 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8059_ _2348_ _2522_ _3204_ vssd1 vssd1 vccd1 vccd1 _3250_ sky130_fd_sc_hd__o21ai_1
XFILLER_18_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7883__B _2941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4747__B _3868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5578__B _0548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5760_ _0732_ _0738_ _3762_ vssd1 vssd1 vccd1 vccd1 _0742_ sky130_fd_sc_hd__a21o_1
XFILLER_62_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_581 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4711_ _3865_ vssd1 vssd1 vccd1 vccd1 _3866_ sky130_fd_sc_hd__clkbuf_4
X_5691_ _0616_ _0609_ _3814_ vssd1 vssd1 vccd1 vccd1 _0667_ sky130_fd_sc_hd__a21o_1
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4642_ _3781_ _3790_ _3796_ vssd1 vssd1 vccd1 vccd1 _3797_ sky130_fd_sc_hd__a21bo_1
X_7430_ _2451_ _2436_ _2514_ _2541_ _2559_ vssd1 vssd1 vccd1 vccd1 _2560_ sky130_fd_sc_hd__o41a_1
XFILLER_116_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4573_ _3704_ _3727_ vssd1 vssd1 vccd1 vccd1 _3728_ sky130_fd_sc_hd__nand2_2
X_7361_ _2481_ _2483_ vssd1 vssd1 vccd1 vccd1 _2484_ sky130_fd_sc_hd__or2_1
XFILLER_116_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6312_ _1306_ _1310_ _1323_ _1329_ vssd1 vssd1 vccd1 vccd1 _1331_ sky130_fd_sc_hd__a211o_1
X_7292_ _2379_ _2396_ _2407_ vssd1 vssd1 vccd1 vccd1 _2409_ sky130_fd_sc_hd__or3_1
X_6243_ _1251_ _1252_ vssd1 vssd1 vccd1 vccd1 _1255_ sky130_fd_sc_hd__nor2_1
X_6174_ _1031_ _1179_ vssd1 vssd1 vccd1 vccd1 _1180_ sky130_fd_sc_hd__nor2_1
XFILLER_111_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5125_ _0095_ _0097_ vssd1 vssd1 vccd1 vccd1 _0098_ sky130_fd_sc_hd__nor2_1
X_5056_ _4210_ _3615_ vssd1 vssd1 vccd1 vccd1 _4211_ sky130_fd_sc_hd__or2_1
XFILLER_38_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4673__A _3735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_662 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8400__A1 _2993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5958_ _0948_ _0952_ vssd1 vssd1 vccd1 vccd1 _0953_ sky130_fd_sc_hd__and2b_1
XFILLER_53_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4909_ _4049_ _4063_ vssd1 vssd1 vccd1 vccd1 _4064_ sky130_fd_sc_hd__and2b_1
XFILLER_40_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5889_ _0864_ _0865_ _0879_ _0876_ vssd1 vssd1 vccd1 vccd1 _0880_ sky130_fd_sc_hd__a211o_1
X_7628_ _2736_ _2777_ _2748_ vssd1 vssd1 vccd1 vccd1 _2778_ sky130_fd_sc_hd__mux2_1
XFILLER_119_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7559_ _0465_ _2696_ _2697_ _2701_ vssd1 vssd1 vccd1 vccd1 _2702_ sky130_fd_sc_hd__a211oi_4
XFILLER_107_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8467__A1 posit_add.in1\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6930_ _1408_ _1409_ _3804_ vssd1 vssd1 vccd1 vccd1 _2010_ sky130_fd_sc_hd__and3_1
XFILLER_47_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4493__A _2969_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6861_ _0303_ _1718_ _1930_ vssd1 vssd1 vccd1 vccd1 _1934_ sky130_fd_sc_hd__o21ai_1
XANTENNA__8394__B1 _2621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5812_ _3763_ _3815_ _0627_ _0634_ vssd1 vssd1 vccd1 vccd1 _0798_ sky130_fd_sc_hd__or4b_1
X_6792_ _1775_ _1777_ vssd1 vssd1 vccd1 vccd1 _1859_ sky130_fd_sc_hd__xnor2_1
X_5743_ _0720_ _0721_ _0724_ vssd1 vssd1 vccd1 vccd1 _0725_ sky130_fd_sc_hd__nand3_1
X_8531_ clknet_3_5__leaf_clk _0017_ vssd1 vssd1 vccd1 vccd1 in_reg\[14\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__4404__C1 _1858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8412__B cmd\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5674_ _0616_ _0648_ _3865_ vssd1 vssd1 vccd1 vccd1 _0649_ sky130_fd_sc_hd__a21oi_1
X_8462_ _3664_ vssd1 vssd1 vccd1 vccd1 _0050_ sky130_fd_sc_hd__clkbuf_1
X_7413_ _2239_ _2240_ vssd1 vssd1 vccd1 vccd1 _2542_ sky130_fd_sc_hd__and2b_1
X_4625_ _3756_ _3779_ vssd1 vssd1 vccd1 vccd1 _3780_ sky130_fd_sc_hd__xnor2_1
X_8393_ _3585_ _3602_ _3605_ vssd1 vssd1 vccd1 vccd1 _3606_ sky130_fd_sc_hd__a21oi_1
XANTENNA__8449__A1 posit_add.in1\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4556_ _2485_ _1737_ vssd1 vssd1 vccd1 vccd1 _3711_ sky130_fd_sc_hd__nand2_1
XANTENNA__7743__S _1297_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7344_ _2425_ _2426_ _2427_ _2465_ vssd1 vssd1 vccd1 vccd1 _2466_ sky130_fd_sc_hd__a31o_1
XFILLER_116_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7044__A _1454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4487_ _2804_ _3002_ _3134_ vssd1 vssd1 vccd1 vccd1 _3145_ sky130_fd_sc_hd__a21o_1
X_7275_ _2365_ _2389_ vssd1 vssd1 vccd1 vccd1 _2390_ sky130_fd_sc_hd__xor2_1
X_6226_ _0795_ _1164_ _1234_ vssd1 vssd1 vccd1 vccd1 _1236_ sky130_fd_sc_hd__a21oi_1
XANTENNA__4387__B _1803_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6157_ _1160_ _1159_ _1161_ vssd1 vssd1 vccd1 vccd1 _1162_ sky130_fd_sc_hd__nand3_1
XFILLER_112_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5683__A1 _3762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5108_ _0080_ _3925_ _4251_ _4254_ vssd1 vssd1 vccd1 vccd1 _0081_ sky130_fd_sc_hd__o31a_1
X_6088_ _1079_ _1081_ _1088_ vssd1 vssd1 vccd1 vccd1 _1089_ sky130_fd_sc_hd__a21bo_1
XFILLER_85_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5039_ _4170_ _4193_ vssd1 vssd1 vccd1 vccd1 _4194_ sky130_fd_sc_hd__xnor2_1
XFILLER_72_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5665__C _3770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6777__B _1718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7129__A _1531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4410_ _2012_ _2276_ _2287_ _1550_ vssd1 vssd1 vccd1 vccd1 _2298_ sky130_fd_sc_hd__a211oi_2
XFILLER_8_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7351__A1 _1428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5390_ _0357_ _1748_ _0361_ _0362_ vssd1 vssd1 vccd1 vccd1 _0363_ sky130_fd_sc_hd__a31o_2
XFILLER_99_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4341_ posit_add.in2\[13\] _1528_ vssd1 vssd1 vccd1 vccd1 _1539_ sky130_fd_sc_hd__xnor2_4
XFILLER_113_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7060_ _2134_ _2142_ vssd1 vssd1 vccd1 vccd1 _2153_ sky130_fd_sc_hd__xor2_1
X_4272_ net1 _0786_ vssd1 vssd1 vccd1 vccd1 _0797_ sky130_fd_sc_hd__nand2_1
X_6011_ _4017_ _0773_ _0992_ vssd1 vssd1 vccd1 vccd1 _1008_ sky130_fd_sc_hd__or3_2
XFILLER_39_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4935__B _4089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6208__A _1164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7962_ _3130_ _3139_ _2999_ vssd1 vssd1 vccd1 vccd1 _3146_ sky130_fd_sc_hd__mux2_1
XFILLER_27_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6913_ _1987_ _1989_ _1991_ vssd1 vssd1 vccd1 vccd1 _1992_ sky130_fd_sc_hd__a21bo_1
X_7893_ _3069_ _3052_ _2954_ vssd1 vssd1 vccd1 vccd1 _3070_ sky130_fd_sc_hd__mux2_1
XFILLER_35_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6844_ _1912_ _1915_ vssd1 vssd1 vccd1 vccd1 _1916_ sky130_fd_sc_hd__xnor2_1
XFILLER_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6775_ _1838_ _1839_ vssd1 vssd1 vccd1 vccd1 _1840_ sky130_fd_sc_hd__and2_1
XFILLER_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5726_ _0705_ vssd1 vssd1 vccd1 vccd1 _0706_ sky130_fd_sc_hd__clkbuf_4
X_8514_ clknet_3_0__leaf_clk _0000_ vssd1 vssd1 vccd1 vccd1 cmd\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_22_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8445_ _3653_ vssd1 vssd1 vccd1 vccd1 _3654_ sky130_fd_sc_hd__clkbuf_4
XFILLER_108_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5782__A _0113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6878__A _1428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5657_ _3761_ _3813_ _0604_ _3717_ _3699_ vssd1 vssd1 vccd1 vccd1 _0630_ sky130_fd_sc_hd__o311a_1
X_4608_ _3762_ vssd1 vssd1 vccd1 vccd1 _3763_ sky130_fd_sc_hd__clkbuf_4
X_8376_ _3555_ _3587_ vssd1 vssd1 vccd1 vccd1 _3588_ sky130_fd_sc_hd__xor2_1
X_5588_ _0559_ _0560_ _0535_ vssd1 vssd1 vccd1 vccd1 _0561_ sky130_fd_sc_hd__mux2_1
XFILLER_104_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4539_ _1385_ _1726_ vssd1 vssd1 vccd1 vccd1 _3678_ sky130_fd_sc_hd__nor2_4
X_7327_ _2443_ _2446_ _2410_ vssd1 vssd1 vccd1 vccd1 _2447_ sky130_fd_sc_hd__mux2_1
X_7258_ _2352_ _2355_ _2357_ vssd1 vssd1 vccd1 vccd1 _2371_ sky130_fd_sc_hd__a21oi_1
X_6209_ _1208_ _1210_ vssd1 vssd1 vccd1 vccd1 _1217_ sky130_fd_sc_hd__and2b_1
X_7189_ _2269_ _2294_ vssd1 vssd1 vccd1 vccd1 _2295_ sky130_fd_sc_hd__nand2_1
XFILLER_93_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_6__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_6__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_60_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5895__B2 _0722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5895__A1 _3892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5867__A _2529_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4890_ _4044_ vssd1 vssd1 vccd1 vccd1 _4045_ sky130_fd_sc_hd__buf_4
XANTENNA__4771__A _3925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6895__A1_N _1665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6560_ _1595_ _1597_ _1602_ vssd1 vssd1 vccd1 vccd1 _1603_ sky130_fd_sc_hd__o21ai_1
X_5511_ _0482_ _0483_ _0338_ vssd1 vssd1 vccd1 vccd1 _0484_ sky130_fd_sc_hd__mux2_1
X_6491_ _1505_ _1525_ vssd1 vssd1 vccd1 vccd1 _1527_ sky130_fd_sc_hd__nand2_1
XFILLER_8_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8230_ _3431_ _3432_ vssd1 vssd1 vccd1 vccd1 _3433_ sky130_fd_sc_hd__nand2_1
X_5442_ _0413_ _0414_ vssd1 vssd1 vccd1 vccd1 _0415_ sky130_fd_sc_hd__or2_1
X_8161_ _3336_ _3342_ vssd1 vssd1 vccd1 vccd1 _3359_ sky130_fd_sc_hd__nand2_1
X_5373_ _0342_ _0345_ vssd1 vssd1 vccd1 vccd1 _0346_ sky130_fd_sc_hd__nor2_1
X_7112_ _2160_ _2209_ vssd1 vssd1 vccd1 vccd1 _2211_ sky130_fd_sc_hd__and2_1
XANTENNA__5107__A _4228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4324_ _1341_ vssd1 vssd1 vccd1 vccd1 _1352_ sky130_fd_sc_hd__buf_2
X_8092_ _2392_ _2486_ vssd1 vssd1 vccd1 vccd1 _3286_ sky130_fd_sc_hd__nand2_2
XFILLER_113_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7043_ _1456_ _1537_ _2063_ vssd1 vssd1 vccd1 vccd1 _2135_ sky130_fd_sc_hd__o21ai_1
XANTENNA__5638__A1 _3762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4946__A _3828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7322__A _2416_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6880__B _1782_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7945_ _2901_ _3034_ _3109_ _3044_ _2941_ vssd1 vssd1 vccd1 vccd1 _3127_ sky130_fd_sc_hd__a221o_1
X_7876_ _3043_ _3050_ _2999_ vssd1 vssd1 vccd1 vccd1 _3051_ sky130_fd_sc_hd__mux2_1
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6827_ _1746_ _1752_ _1760_ vssd1 vssd1 vccd1 vccd1 _1897_ sky130_fd_sc_hd__nand3_1
XFILLER_23_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6758_ _1805_ _1820_ _1818_ vssd1 vssd1 vccd1 vccd1 _1821_ sky130_fd_sc_hd__a21oi_1
XFILLER_10_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5709_ _0604_ _0607_ vssd1 vssd1 vccd1 vccd1 _0687_ sky130_fd_sc_hd__and2_2
XANTENNA__8512__A0 _1275_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6689_ _1738_ _1744_ vssd1 vssd1 vccd1 vccd1 _1745_ sky130_fd_sc_hd__xnor2_1
XANTENNA__7315__A1 _1456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6401__A _4037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8428_ _3639_ _3640_ vssd1 vssd1 vccd1 vccd1 _0037_ sky130_fd_sc_hd__nor2_1
XFILLER_105_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5877__A1 _3776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8359_ _3502_ _3528_ _3568_ vssd1 vssd1 vccd1 vccd1 _3570_ sky130_fd_sc_hd__a21oi_1
XANTENNA__5017__A _3893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7306__A1 _1676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4843__A2 _3883_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7242__B1 _2352_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5991_ _0882_ _0853_ vssd1 vssd1 vccd1 vccd1 _0987_ sky130_fd_sc_hd__and2b_1
XFILLER_92_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4942_ _2540_ _3930_ vssd1 vssd1 vccd1 vccd1 _4097_ sky130_fd_sc_hd__nor2_1
XFILLER_17_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7730_ _2843_ _2889_ vssd1 vssd1 vccd1 vccd1 _2890_ sky130_fd_sc_hd__xor2_1
X_7661_ _2801_ _2812_ _2813_ vssd1 vssd1 vccd1 vccd1 _2814_ sky130_fd_sc_hd__o21a_1
XFILLER_32_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4873_ _4011_ _4027_ vssd1 vssd1 vccd1 vccd1 _4028_ sky130_fd_sc_hd__xnor2_2
X_6612_ _1420_ _1510_ vssd1 vssd1 vccd1 vccd1 _1661_ sky130_fd_sc_hd__nor2_1
XFILLER_60_593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7592_ _2729_ _2737_ vssd1 vssd1 vccd1 vccd1 _2739_ sky130_fd_sc_hd__nand2_1
XFILLER_32_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6543_ _1496_ _1502_ _1503_ _1450_ vssd1 vssd1 vccd1 vccd1 _1585_ sky130_fd_sc_hd__a2bb2o_1
X_6474_ _1157_ _1508_ vssd1 vssd1 vccd1 vccd1 _1509_ sky130_fd_sc_hd__xnor2_2
XANTENNA__6221__A _0702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8213_ _3322_ _3355_ _3408_ _3323_ vssd1 vssd1 vccd1 vccd1 _3415_ sky130_fd_sc_hd__or4bb_1
X_5425_ _0397_ vssd1 vssd1 vccd1 vccd1 _0398_ sky130_fd_sc_hd__inv_2
XANTENNA__7751__S _1297_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5356_ _0133_ _0163_ vssd1 vssd1 vccd1 vccd1 _0329_ sky130_fd_sc_hd__xor2_1
X_8144_ _3340_ _3341_ vssd1 vssd1 vccd1 vccd1 _3342_ sky130_fd_sc_hd__nand2_1
XFILLER_101_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4307_ _1156_ vssd1 vssd1 vccd1 vccd1 _0018_ sky130_fd_sc_hd__clkbuf_1
X_5287_ _0257_ _0259_ vssd1 vssd1 vccd1 vccd1 _0260_ sky130_fd_sc_hd__xnor2_1
XANTENNA__4676__A _3690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8075_ _3166_ _3257_ _3267_ vssd1 vssd1 vccd1 vccd1 _3268_ sky130_fd_sc_hd__o21a_1
XFILLER_101_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7026_ _4217_ _2079_ vssd1 vssd1 vccd1 vccd1 _2116_ sky130_fd_sc_hd__nand2_1
XFILLER_87_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4598__A1 _2969_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7928_ _3094_ _3107_ _2998_ vssd1 vssd1 vccd1 vccd1 _3108_ sky130_fd_sc_hd__mux2_1
XFILLER_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7859_ _2999_ _3021_ _3030_ _3031_ vssd1 vssd1 vccd1 vccd1 _3032_ sky130_fd_sc_hd__o211a_1
XFILLER_51_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6009__C _0773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5210__A _3701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5210_ _3701_ _3817_ vssd1 vssd1 vccd1 vccd1 _0183_ sky130_fd_sc_hd__nor2_1
XANTENNA__7571__S _2652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6190_ _0773_ _1095_ vssd1 vssd1 vccd1 vccd1 _1197_ sky130_fd_sc_hd__nor2_1
XFILLER_97_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5710__B1 _3762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5141_ _0113_ _4217_ vssd1 vssd1 vccd1 vccd1 _0114_ sky130_fd_sc_hd__nand2_1
X_5072_ _4216_ _4226_ vssd1 vssd1 vccd1 vccd1 _4227_ sky130_fd_sc_hd__and2b_1
XFILLER_69_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6018__A1 _0779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5974_ _0891_ _0920_ _0919_ vssd1 vssd1 vccd1 vccd1 _0970_ sky130_fd_sc_hd__a21bo_1
XFILLER_80_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7713_ _2851_ _2869_ _2871_ vssd1 vssd1 vccd1 vccd1 _2872_ sky130_fd_sc_hd__o21bai_1
XFILLER_100_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4925_ _4077_ _4078_ _4079_ vssd1 vssd1 vccd1 vccd1 _4080_ sky130_fd_sc_hd__o21a_1
XFILLER_40_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4856_ _4009_ _4010_ vssd1 vssd1 vccd1 vccd1 _4011_ sky130_fd_sc_hd__xnor2_1
X_7644_ _2762_ _2795_ vssd1 vssd1 vccd1 vccd1 _2796_ sky130_fd_sc_hd__or2_1
X_7575_ _2704_ _2719_ vssd1 vssd1 vccd1 vccd1 _2720_ sky130_fd_sc_hd__or2_1
X_6526_ _1553_ _1554_ vssd1 vssd1 vccd1 vccd1 _1566_ sky130_fd_sc_hd__xor2_4
X_4787_ _3739_ _3750_ vssd1 vssd1 vccd1 vccd1 _3942_ sky130_fd_sc_hd__or2_1
XFILLER_118_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6457_ _1481_ _1489_ vssd1 vssd1 vccd1 vccd1 _1490_ sky130_fd_sc_hd__xor2_1
X_6388_ _1413_ vssd1 vssd1 vccd1 vccd1 _1414_ sky130_fd_sc_hd__clkbuf_4
X_5408_ _1605_ _3635_ _3651_ _3830_ vssd1 vssd1 vccd1 vccd1 _0381_ sky130_fd_sc_hd__a211o_1
XFILLER_88_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5339_ _0302_ _0310_ vssd1 vssd1 vccd1 vccd1 _0312_ sky130_fd_sc_hd__and2_1
X_8127_ _3200_ _3201_ _3208_ _3254_ _3290_ vssd1 vssd1 vccd1 vccd1 _3323_ sky130_fd_sc_hd__a2111oi_2
X_8058_ _2521_ _3198_ _3207_ vssd1 vssd1 vccd1 vccd1 _3249_ sky130_fd_sc_hd__nand3_2
X_7009_ _2094_ _2096_ vssd1 vssd1 vccd1 vccd1 _2097_ sky130_fd_sc_hd__and2_1
XFILLER_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7757__A1 _1308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7748__A1 _1297_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5690_ _0665_ _0648_ vssd1 vssd1 vccd1 vccd1 _0666_ sky130_fd_sc_hd__or2_1
X_4710_ _3864_ vssd1 vssd1 vccd1 vccd1 _3865_ sky130_fd_sc_hd__buf_2
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4641_ _3793_ _3795_ _3782_ vssd1 vssd1 vccd1 vccd1 _3796_ sky130_fd_sc_hd__or3_1
XFILLER_116_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4572_ _3719_ _3726_ vssd1 vssd1 vccd1 vccd1 _3727_ sky130_fd_sc_hd__nor2_1
X_7360_ _2482_ _2406_ vssd1 vssd1 vccd1 vccd1 _2483_ sky130_fd_sc_hd__xnor2_1
XFILLER_116_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6311_ _1327_ _1328_ vssd1 vssd1 vccd1 vccd1 _1329_ sky130_fd_sc_hd__or2_1
X_7291_ _2399_ _2401_ _2402_ _2405_ _2406_ vssd1 vssd1 vccd1 vccd1 _2407_ sky130_fd_sc_hd__a2111oi_2
XFILLER_115_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6242_ _1251_ _1252_ vssd1 vssd1 vccd1 vccd1 _1254_ sky130_fd_sc_hd__xor2_1
XFILLER_89_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6173_ _1162_ _1174_ _1178_ vssd1 vssd1 vccd1 vccd1 _1179_ sky130_fd_sc_hd__and3_1
XFILLER_69_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5124_ _0094_ _0096_ _0091_ vssd1 vssd1 vccd1 vccd1 _0097_ sky130_fd_sc_hd__o21a_1
X_5055_ _4017_ vssd1 vssd1 vccd1 vccd1 _4210_ sky130_fd_sc_hd__buf_4
XFILLER_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_674 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6411__A1 _0795_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5957_ _0945_ _0947_ vssd1 vssd1 vccd1 vccd1 _0952_ sky130_fd_sc_hd__nand2_1
XFILLER_80_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4908_ _4056_ _4061_ _4062_ vssd1 vssd1 vccd1 vccd1 _4063_ sky130_fd_sc_hd__a21o_1
X_5888_ _0876_ _0877_ _0878_ vssd1 vssd1 vccd1 vccd1 _0879_ sky130_fd_sc_hd__nor3_2
X_7627_ _2731_ _2755_ _2776_ vssd1 vssd1 vccd1 vccd1 _2777_ sky130_fd_sc_hd__o21ai_1
X_4839_ _3992_ _3993_ vssd1 vssd1 vccd1 vccd1 _3994_ sky130_fd_sc_hd__nand2_1
XFILLER_119_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7558_ _2698_ _2699_ _2700_ vssd1 vssd1 vccd1 vccd1 _2701_ sky130_fd_sc_hd__a21o_1
X_6509_ _1545_ _1546_ vssd1 vssd1 vccd1 vccd1 _1547_ sky130_fd_sc_hd__xnor2_2
X_7489_ _2624_ _1539_ vssd1 vssd1 vccd1 vccd1 _2625_ sky130_fd_sc_hd__or2_1
XFILLER_107_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4864__A _4018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6782__C _4089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6860_ _1922_ _1923_ vssd1 vssd1 vccd1 vccd1 _1933_ sky130_fd_sc_hd__or2_1
XFILLER_81_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5811_ _3901_ _0795_ _0634_ _3866_ vssd1 vssd1 vccd1 vccd1 _0796_ sky130_fd_sc_hd__a22o_1
X_6791_ _1845_ _1855_ _1856_ vssd1 vssd1 vccd1 vccd1 _1857_ sky130_fd_sc_hd__o21ai_1
XFILLER_62_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5742_ _3901_ _0722_ _0705_ _0113_ vssd1 vssd1 vccd1 vccd1 _0724_ sky130_fd_sc_hd__a22o_1
X_8530_ clknet_3_4__leaf_clk _0016_ vssd1 vssd1 vccd1 vccd1 in_reg\[13\] sky130_fd_sc_hd__dfxtp_1
X_8461_ in_reg\[7\] posit_add.in1\[7\] _3655_ vssd1 vssd1 vccd1 vccd1 _3664_ sky130_fd_sc_hd__mux2_1
X_5673_ _4043_ _0647_ _3811_ _3812_ _3678_ vssd1 vssd1 vccd1 vccd1 _0648_ sky130_fd_sc_hd__a221o_1
XFILLER_30_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4624_ _3764_ _3778_ vssd1 vssd1 vccd1 vccd1 _3779_ sky130_fd_sc_hd__xnor2_1
X_8392_ _3404_ _3603_ _3416_ vssd1 vssd1 vccd1 vccd1 _3605_ sky130_fd_sc_hd__a21o_1
X_7412_ _2535_ _2539_ vssd1 vssd1 vccd1 vccd1 _2541_ sky130_fd_sc_hd__or2_1
XFILLER_116_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4555_ _1737_ _3706_ _3708_ _3709_ vssd1 vssd1 vccd1 vccd1 _3710_ sky130_fd_sc_hd__a31o_1
X_7343_ _0147_ _2431_ _2437_ _2462_ _2464_ vssd1 vssd1 vccd1 vccd1 _2465_ sky130_fd_sc_hd__o221a_1
XANTENNA__7325__A _3804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7044__B _1531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4486_ _3046_ _3123_ vssd1 vssd1 vccd1 vccd1 _3134_ sky130_fd_sc_hd__or2_2
X_7274_ _2347_ _2359_ _2371_ vssd1 vssd1 vccd1 vccd1 _2389_ sky130_fd_sc_hd__a21oi_2
X_6225_ _0795_ _1164_ _1234_ vssd1 vssd1 vccd1 vccd1 _1235_ sky130_fd_sc_hd__and3_1
X_6156_ _1097_ _1128_ vssd1 vssd1 vccd1 vccd1 _1161_ sky130_fd_sc_hd__and2_1
XFILLER_103_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4684__A _3832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5107_ _4228_ vssd1 vssd1 vccd1 vccd1 _0080_ sky130_fd_sc_hd__buf_4
XFILLER_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6087_ _0802_ _3739_ _1082_ _1086_ _1087_ vssd1 vssd1 vccd1 vccd1 _1088_ sky130_fd_sc_hd__o221a_1
XFILLER_57_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5038_ _4191_ _4192_ vssd1 vssd1 vccd1 vccd1 _4193_ sky130_fd_sc_hd__nor2_1
XFILLER_72_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8385__A1 _3182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5199__A1 _3816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6989_ _2072_ _2073_ _2074_ _2068_ vssd1 vssd1 vccd1 vccd1 _2075_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_80_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7648__A0 _3771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7351__A2 _2412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4340_ posit_add.in2\[12\] _1352_ _1374_ _1396_ _1264_ vssd1 vssd1 vccd1 vccd1 _1528_
+ sky130_fd_sc_hd__o41a_2
XFILLER_113_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4271_ last_SCLK net2 vssd1 vssd1 vccd1 vccd1 _0786_ sky130_fd_sc_hd__nor2b_1
XFILLER_4_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6010_ _0802_ vssd1 vssd1 vccd1 vccd1 _1007_ sky130_fd_sc_hd__inv_2
XFILLER_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7961_ _3084_ _3108_ _3006_ vssd1 vssd1 vccd1 vccd1 _3144_ sky130_fd_sc_hd__mux2_1
XFILLER_27_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6912_ _1985_ _1986_ vssd1 vssd1 vccd1 vccd1 _1991_ sky130_fd_sc_hd__nand2_1
XFILLER_82_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7892_ _3067_ vssd1 vssd1 vccd1 vccd1 _3069_ sky130_fd_sc_hd__clkinv_2
X_6843_ _1850_ _1914_ vssd1 vssd1 vccd1 vccd1 _1915_ sky130_fd_sc_hd__xnor2_1
XANTENNA__8367__A1 _3577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6774_ _1831_ _1835_ _1837_ vssd1 vssd1 vccd1 vccd1 _1839_ sky130_fd_sc_hd__nand3_1
XFILLER_22_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5725_ _4222_ _0684_ _0692_ vssd1 vssd1 vccd1 vccd1 _0705_ sky130_fd_sc_hd__o21ai_1
X_8513_ _3697_ vssd1 vssd1 vccd1 vccd1 _0074_ sky130_fd_sc_hd__clkbuf_1
XFILLER_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5656_ _0616_ _0607_ _3801_ _3717_ vssd1 vssd1 vccd1 vccd1 _0629_ sky130_fd_sc_hd__a211o_1
X_8444_ net4 cmd\[0\] _3637_ net1 vssd1 vssd1 vccd1 vccd1 _3653_ sky130_fd_sc_hd__or4b_1
XANTENNA__5782__B _0762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6878__B _1538_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4607_ _3761_ vssd1 vssd1 vccd1 vccd1 _3762_ sky130_fd_sc_hd__clkbuf_4
X_8375_ _0521_ _3363_ _3429_ vssd1 vssd1 vccd1 vccd1 _3587_ sky130_fd_sc_hd__a21o_1
X_5587_ _0477_ _0544_ _0480_ vssd1 vssd1 vccd1 vccd1 _0560_ sky130_fd_sc_hd__mux2_1
XFILLER_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4538_ _1682_ _3635_ _3665_ _2408_ vssd1 vssd1 vccd1 vccd1 _3671_ sky130_fd_sc_hd__a211o_1
X_7326_ _2414_ _2444_ _2438_ _2335_ _2445_ vssd1 vssd1 vccd1 vccd1 _2446_ sky130_fd_sc_hd__a221oi_2
XFILLER_117_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4469_ _2661_ _2936_ vssd1 vssd1 vccd1 vccd1 _2947_ sky130_fd_sc_hd__xnor2_1
X_7257_ _2365_ _2369_ vssd1 vssd1 vccd1 vccd1 _2370_ sky130_fd_sc_hd__nor2_1
X_6208_ _1164_ _1215_ vssd1 vssd1 vccd1 vccd1 _1216_ sky130_fd_sc_hd__xor2_1
XFILLER_89_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7188_ _2292_ _2293_ vssd1 vssd1 vccd1 vccd1 _2294_ sky130_fd_sc_hd__and2_1
X_6139_ _0795_ _1102_ _1104_ _1142_ vssd1 vssd1 vccd1 vccd1 _1143_ sky130_fd_sc_hd__a31o_1
XFILLER_100_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5408__A2 _3635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_422 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5895__A2 _0706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4552__C1 _1913_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6979__A _1401_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5510_ _0282_ _0324_ vssd1 vssd1 vccd1 vccd1 _0483_ sky130_fd_sc_hd__xor2_1
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6490_ _1505_ _1525_ vssd1 vssd1 vccd1 vccd1 _1526_ sky130_fd_sc_hd__nor2_1
XFILLER_9_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5441_ _0405_ _0412_ vssd1 vssd1 vccd1 vccd1 _0414_ sky130_fd_sc_hd__and2_1
X_8160_ _3356_ _3357_ vssd1 vssd1 vccd1 vccd1 _3358_ sky130_fd_sc_hd__or2_1
X_5372_ _0343_ _0344_ vssd1 vssd1 vccd1 vccd1 _0345_ sky130_fd_sc_hd__nand2_1
X_7111_ _2189_ _2208_ vssd1 vssd1 vccd1 vccd1 _2209_ sky130_fd_sc_hd__and2_1
X_4323_ posit_add.in2\[0\] posit_add.in2\[1\] posit_add.in2\[3\] posit_add.in2\[2\]
+ vssd1 vssd1 vccd1 vccd1 _1341_ sky130_fd_sc_hd__or4_1
X_8091_ _3252_ _3207_ _3198_ _2521_ vssd1 vssd1 vccd1 vccd1 _3284_ sky130_fd_sc_hd__and4b_2
XFILLER_113_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7042_ _4089_ _1676_ _1537_ _2086_ vssd1 vssd1 vccd1 vccd1 _2134_ sky130_fd_sc_hd__or4_1
XFILLER_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5123__A _0092_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7944_ _2894_ _3034_ vssd1 vssd1 vccd1 vccd1 _3126_ sky130_fd_sc_hd__nor2_1
XFILLER_70_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7875_ _3042_ _3048_ _3041_ _3049_ vssd1 vssd1 vccd1 vccd1 _3050_ sky130_fd_sc_hd__a22o_1
XFILLER_23_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_422 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6826_ _1840_ _1895_ vssd1 vssd1 vccd1 vccd1 _1896_ sky130_fd_sc_hd__xnor2_1
X_6757_ _1818_ _1819_ vssd1 vssd1 vccd1 vccd1 _1820_ sky130_fd_sc_hd__nor2_1
XFILLER_11_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5708_ _3718_ _0612_ _0685_ _0617_ vssd1 vssd1 vccd1 vccd1 _0686_ sky130_fd_sc_hd__a31o_1
XFILLER_10_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8512__A1 in_reg\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6688_ _1739_ _1743_ vssd1 vssd1 vccd1 vccd1 _1744_ sky130_fd_sc_hd__xor2_1
XANTENNA__7315__A2 _2412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5639_ _3900_ _0609_ vssd1 vssd1 vccd1 vccd1 _0612_ sky130_fd_sc_hd__nand2_1
X_8427_ in_reg\[1\] _0679_ mode vssd1 vssd1 vccd1 vccd1 _3640_ sky130_fd_sc_hd__a21oi_1
X_8358_ _3502_ _3528_ _3568_ vssd1 vssd1 vccd1 vccd1 _3569_ sky130_fd_sc_hd__and3_1
XFILLER_88_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7309_ _2399_ _2401_ _2402_ _2405_ _2406_ vssd1 vssd1 vccd1 vccd1 _2427_ sky130_fd_sc_hd__a2111o_4
X_8289_ out_reg\[8\] _3316_ _1231_ out_reg\[9\] vssd1 vssd1 vccd1 vccd1 _3496_ sky130_fd_sc_hd__a22o_1
XANTENNA__6129__A _1128_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6799__A _1401_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7306__A2 _2412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8267__B1 _3471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5990_ _0984_ _0985_ vssd1 vssd1 vccd1 vccd1 _0986_ sky130_fd_sc_hd__and2b_1
XFILLER_52_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4941_ _4090_ _4092_ vssd1 vssd1 vccd1 vccd1 _4096_ sky130_fd_sc_hd__xnor2_1
X_4872_ _4012_ _4026_ vssd1 vssd1 vccd1 vccd1 _4027_ sky130_fd_sc_hd__xnor2_1
X_7660_ _2799_ _2800_ vssd1 vssd1 vccd1 vccd1 _2813_ sky130_fd_sc_hd__nand2_1
X_6611_ _1654_ _1658_ vssd1 vssd1 vccd1 vccd1 _1659_ sky130_fd_sc_hd__xnor2_1
X_7591_ _2704_ _2736_ vssd1 vssd1 vccd1 vccd1 _2737_ sky130_fd_sc_hd__nor2_1
XANTENNA__6502__A _0082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6542_ _1530_ _1582_ vssd1 vssd1 vccd1 vccd1 _1584_ sky130_fd_sc_hd__nor2_1
X_6473_ _1191_ _1226_ _1305_ _1309_ vssd1 vssd1 vccd1 vccd1 _1508_ sky130_fd_sc_hd__o31a_1
X_8212_ _1220_ _3413_ vssd1 vssd1 vccd1 vccd1 _0026_ sky130_fd_sc_hd__nor2_1
X_5424_ _0351_ _0396_ vssd1 vssd1 vccd1 vccd1 _0397_ sky130_fd_sc_hd__xnor2_2
X_8143_ _3265_ _3309_ _3338_ vssd1 vssd1 vccd1 vccd1 _3341_ sky130_fd_sc_hd__a21o_1
XFILLER_99_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5355_ _0209_ _0327_ _0206_ vssd1 vssd1 vccd1 vccd1 _0328_ sky130_fd_sc_hd__a21oi_1
XFILLER_102_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4306_ in_reg\[14\] in_reg\[15\] _0819_ vssd1 vssd1 vccd1 vccd1 _1156_ sky130_fd_sc_hd__mux2_1
X_5286_ _0258_ _0232_ vssd1 vssd1 vccd1 vccd1 _0259_ sky130_fd_sc_hd__xnor2_1
XANTENNA__4676__B _3830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8074_ _3265_ _3266_ vssd1 vssd1 vccd1 vccd1 _3267_ sky130_fd_sc_hd__or2_1
X_7025_ _2113_ _2114_ vssd1 vssd1 vccd1 vccd1 _2115_ sky130_fd_sc_hd__or2b_1
XFILLER_68_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5788__A _3763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6891__B _3930_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7927_ _3092_ _3106_ _2842_ vssd1 vssd1 vccd1 vccd1 _3107_ sky130_fd_sc_hd__mux2_1
XFILLER_90_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7858_ _3006_ _3020_ vssd1 vssd1 vccd1 vccd1 _3031_ sky130_fd_sc_hd__or2_1
XFILLER_23_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6809_ _1863_ _1875_ vssd1 vssd1 vccd1 vccd1 _1877_ sky130_fd_sc_hd__and2_1
XFILLER_51_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7789_ _0370_ _2340_ _2721_ vssd1 vssd1 vccd1 vccd1 _2955_ sky130_fd_sc_hd__mux2_1
XFILLER_109_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7227__B _2335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5028__A _3828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5901__A2_N _3832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5210__B _3817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_440 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5140_ _0112_ vssd1 vssd1 vccd1 vccd1 _0113_ sky130_fd_sc_hd__buf_4
XFILLER_69_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5071_ _4218_ _4225_ vssd1 vssd1 vccd1 vccd1 _4226_ sky130_fd_sc_hd__xor2_1
XFILLER_84_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5973_ _0965_ _0966_ _0963_ vssd1 vssd1 vccd1 vccd1 _0969_ sky130_fd_sc_hd__o21ai_1
XFILLER_92_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4924_ _4074_ _4076_ vssd1 vssd1 vccd1 vccd1 _4079_ sky130_fd_sc_hd__nand2_1
X_7712_ _2811_ _2802_ vssd1 vssd1 vccd1 vccd1 _2871_ sky130_fd_sc_hd__and2_1
XFILLER_40_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4855_ _3860_ _3888_ vssd1 vssd1 vccd1 vccd1 _4010_ sky130_fd_sc_hd__nand2_1
XFILLER_20_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7643_ _2756_ _2794_ _2748_ vssd1 vssd1 vccd1 vccd1 _2795_ sky130_fd_sc_hd__mux2_1
XFILLER_33_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4786_ _3897_ _3902_ vssd1 vssd1 vccd1 vccd1 _3941_ sky130_fd_sc_hd__xnor2_1
X_7574_ _2706_ _2711_ _2712_ _2718_ vssd1 vssd1 vccd1 vccd1 _2719_ sky130_fd_sc_hd__o22a_1
XFILLER_118_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6525_ _1543_ _1563_ _1564_ vssd1 vssd1 vccd1 vccd1 _1565_ sky130_fd_sc_hd__a21bo_1
XFILLER_20_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5790__B _0773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6456_ _1487_ _1488_ vssd1 vssd1 vccd1 vccd1 _1489_ sky130_fd_sc_hd__xor2_1
X_6387_ _1405_ _1412_ vssd1 vssd1 vccd1 vccd1 _1413_ sky130_fd_sc_hd__nor2_1
XFILLER_88_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5407_ _3594_ _3156_ _3746_ _3748_ vssd1 vssd1 vccd1 vccd1 _0380_ sky130_fd_sc_hd__nand4_2
XFILLER_102_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7063__A _1531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5338_ _0302_ _0310_ vssd1 vssd1 vccd1 vccd1 _0311_ sky130_fd_sc_hd__nor2_1
X_8126_ _3319_ _3321_ vssd1 vssd1 vccd1 vccd1 _3322_ sky130_fd_sc_hd__xor2_4
XFILLER_102_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8057_ _1319_ _3247_ vssd1 vssd1 vccd1 vccd1 _3248_ sky130_fd_sc_hd__and2_1
XANTENNA__7998__A _1253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7008_ _2051_ _2095_ vssd1 vssd1 vccd1 vccd1 _2096_ sky130_fd_sc_hd__nor2_1
XFILLER_87_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5269_ _0240_ _0225_ _0238_ vssd1 vssd1 vccd1 vccd1 _0242_ sky130_fd_sc_hd__and3_1
XFILLER_28_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7937__S _2937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7238__A _2980_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4640_ _3794_ vssd1 vssd1 vccd1 vccd1 _3795_ sky130_fd_sc_hd__clkbuf_4
XFILLER_30_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6310_ _1324_ _1326_ vssd1 vssd1 vccd1 vccd1 _1328_ sky130_fd_sc_hd__and2_1
X_4571_ _3725_ vssd1 vssd1 vccd1 vccd1 _3726_ sky130_fd_sc_hd__buf_2
XFILLER_116_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7290_ _2400_ _2388_ vssd1 vssd1 vccd1 vccd1 _2406_ sky130_fd_sc_hd__xnor2_2
XFILLER_116_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6241_ _1211_ _1216_ vssd1 vssd1 vccd1 vccd1 _1252_ sky130_fd_sc_hd__xnor2_1
XFILLER_115_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6172_ _1175_ _1029_ _1176_ vssd1 vssd1 vccd1 vccd1 _1178_ sky130_fd_sc_hd__a21o_1
XFILLER_103_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5123_ _0092_ _0075_ _0093_ vssd1 vssd1 vccd1 vccd1 _0096_ sky130_fd_sc_hd__nor3_1
XFILLER_111_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5054_ _4207_ _4208_ vssd1 vssd1 vccd1 vccd1 _4209_ sky130_fd_sc_hd__xor2_1
XFILLER_38_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5956_ _0933_ _0950_ vssd1 vssd1 vccd1 vccd1 _0951_ sky130_fd_sc_hd__nor2_1
XFILLER_80_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5887_ _3738_ _0860_ vssd1 vssd1 vccd1 vccd1 _0878_ sky130_fd_sc_hd__xnor2_1
XFILLER_52_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4907_ _4057_ _4060_ vssd1 vssd1 vccd1 vccd1 _4062_ sky130_fd_sc_hd__nor2_1
XFILLER_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4838_ _3818_ _3842_ vssd1 vssd1 vccd1 vccd1 _3993_ sky130_fd_sc_hd__and2_1
X_7626_ _2712_ _2775_ vssd1 vssd1 vccd1 vccd1 _2776_ sky130_fd_sc_hd__or2_1
X_4769_ _3923_ vssd1 vssd1 vccd1 vccd1 _3924_ sky130_fd_sc_hd__clkbuf_4
X_7557_ _0425_ _2693_ vssd1 vssd1 vccd1 vccd1 _2700_ sky130_fd_sc_hd__xnor2_1
X_6508_ _1353_ _1354_ _3986_ vssd1 vssd1 vccd1 vccd1 _1546_ sky130_fd_sc_hd__and3_1
X_7488_ _3035_ vssd1 vssd1 vccd1 vccd1 _2624_ sky130_fd_sc_hd__inv_2
X_6439_ _0080_ _1423_ vssd1 vssd1 vccd1 vccd1 _1470_ sky130_fd_sc_hd__nor2_1
XFILLER_106_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7224__C _2333_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8109_ _3295_ _3301_ _3302_ _3303_ vssd1 vssd1 vccd1 vccd1 _3304_ sky130_fd_sc_hd__a211o_1
XFILLER_102_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5438__B1 _2980_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7418__A1 _1531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7577__S _2721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5810_ _0633_ vssd1 vssd1 vccd1 vccd1 _0795_ sky130_fd_sc_hd__clkbuf_4
X_6790_ _1852_ _1854_ vssd1 vssd1 vccd1 vccd1 _1856_ sky130_fd_sc_hd__nand2_1
XFILLER_62_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5741_ _0700_ vssd1 vssd1 vccd1 vccd1 _0722_ sky130_fd_sc_hd__inv_2
XFILLER_34_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8460_ _3663_ vssd1 vssd1 vccd1 vccd1 _0049_ sky130_fd_sc_hd__clkbuf_1
X_5672_ _1990_ _3713_ _3715_ _3774_ vssd1 vssd1 vccd1 vccd1 _0647_ sky130_fd_sc_hd__a31o_1
X_7411_ _2538_ _2525_ _2454_ vssd1 vssd1 vccd1 vccd1 _2539_ sky130_fd_sc_hd__mux2_1
X_4623_ _3773_ _3777_ vssd1 vssd1 vccd1 vccd1 _3778_ sky130_fd_sc_hd__xor2_1
X_8391_ _2604_ _3580_ vssd1 vssd1 vccd1 vccd1 _3603_ sky130_fd_sc_hd__nor2_1
XFILLER_116_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6510__A _1400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4554_ posit_add.in2\[0\] _2408_ _2221_ vssd1 vssd1 vccd1 vccd1 _3709_ sky130_fd_sc_hd__and3_1
X_7342_ _2442_ _2458_ vssd1 vssd1 vccd1 vccd1 _2464_ sky130_fd_sc_hd__or2_1
XFILLER_116_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7273_ _2358_ _2387_ vssd1 vssd1 vccd1 vccd1 _2388_ sky130_fd_sc_hd__xnor2_4
XFILLER_116_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6224_ _1193_ _1228_ _1232_ _1233_ vssd1 vssd1 vccd1 vccd1 _1234_ sky130_fd_sc_hd__o22ai_1
X_4485_ _3079_ _3112_ vssd1 vssd1 vccd1 vccd1 _3123_ sky130_fd_sc_hd__nand2_1
XFILLER_106_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7044__C _1537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6155_ _0702_ _1095_ _1102_ _0762_ vssd1 vssd1 vccd1 vccd1 _1160_ sky130_fd_sc_hd__a2bb2o_1
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6086_ _3770_ _3739_ _0787_ vssd1 vssd1 vccd1 vccd1 _1087_ sky130_fd_sc_hd__a21o_1
XFILLER_85_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4684__B _3838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5106_ _4246_ _0078_ vssd1 vssd1 vccd1 vccd1 _0079_ sky130_fd_sc_hd__nand2_1
X_5037_ _4190_ _3994_ _4171_ vssd1 vssd1 vccd1 vccd1 _4192_ sky130_fd_sc_hd__and3_1
XFILLER_73_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5199__A2 _3988_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7593__A0 _0113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6988_ _2072_ _2073_ vssd1 vssd1 vccd1 vccd1 _2074_ sky130_fd_sc_hd__xor2_1
XFILLER_53_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5939_ _0931_ _0932_ vssd1 vssd1 vccd1 vccd1 _0933_ sky130_fd_sc_hd__nor2_1
XFILLER_15_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7609_ _2676_ _2753_ _2756_ _2748_ vssd1 vssd1 vccd1 vccd1 _2757_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__6420__A _1446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7648__A1 _3703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6320__B2 _0722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6320__A1 _0762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6139__A1 _0795_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4270_ _0765_ vssd1 vssd1 vccd1 vccd1 _0002_ sky130_fd_sc_hd__clkbuf_1
XFILLER_97_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7960_ _3132_ _3142_ _3021_ vssd1 vssd1 vccd1 vccd1 _3143_ sky130_fd_sc_hd__mux2_1
XFILLER_39_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6911_ _1988_ _1963_ vssd1 vssd1 vccd1 vccd1 _1989_ sky130_fd_sc_hd__xnor2_1
X_7891_ _3066_ _2921_ _2971_ vssd1 vssd1 vccd1 vccd1 _3067_ sky130_fd_sc_hd__mux2_1
X_6842_ _1408_ _1409_ _1782_ vssd1 vssd1 vccd1 vccd1 _1914_ sky130_fd_sc_hd__and3_1
XFILLER_35_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6773_ _1831_ _1835_ _1837_ vssd1 vssd1 vccd1 vccd1 _1838_ sky130_fd_sc_hd__a21o_1
X_5724_ _3762_ _0693_ _0703_ vssd1 vssd1 vccd1 vccd1 _0704_ sky130_fd_sc_hd__or3b_1
X_8512_ _1275_ in_reg\[15\] _3676_ vssd1 vssd1 vccd1 vccd1 _3697_ sky130_fd_sc_hd__mux2_1
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5655_ _3864_ _0619_ _3699_ _0111_ vssd1 vssd1 vccd1 vccd1 _0628_ sky130_fd_sc_hd__a211o_1
X_8443_ counter\[4\] _3648_ _3652_ vssd1 vssd1 vccd1 vccd1 _0042_ sky130_fd_sc_hd__o21ba_1
X_4606_ _3759_ _3760_ vssd1 vssd1 vccd1 vccd1 _3761_ sky130_fd_sc_hd__nand2_2
X_8374_ _3582_ _3585_ vssd1 vssd1 vccd1 vccd1 _3586_ sky130_fd_sc_hd__xnor2_1
X_7325_ _3804_ _2431_ vssd1 vssd1 vccd1 vccd1 _2445_ sky130_fd_sc_hd__nor2_1
X_5586_ _0491_ _0471_ _0480_ vssd1 vssd1 vccd1 vccd1 _0559_ sky130_fd_sc_hd__mux2_1
XFILLER_89_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4537_ _1726_ _2353_ _2364_ _1946_ vssd1 vssd1 vccd1 vccd1 _3665_ sky130_fd_sc_hd__o211a_1
XFILLER_117_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4468_ posit_add.in1\[3\] _2925_ vssd1 vssd1 vccd1 vccd1 _2936_ sky130_fd_sc_hd__xor2_4
X_7256_ _2367_ _2368_ vssd1 vssd1 vccd1 vccd1 _2369_ sky130_fd_sc_hd__nand2_2
X_6207_ _1213_ _1214_ vssd1 vssd1 vccd1 vccd1 _1215_ sky130_fd_sc_hd__xor2_1
XFILLER_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7187_ _2289_ _2291_ vssd1 vssd1 vccd1 vccd1 _2293_ sky130_fd_sc_hd__nand2_1
X_6138_ _1095_ _1106_ vssd1 vssd1 vccd1 vccd1 _1142_ sky130_fd_sc_hd__and2b_1
X_4399_ _1781_ _1451_ vssd1 vssd1 vccd1 vccd1 _2177_ sky130_fd_sc_hd__nor2_1
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6069_ _3892_ _1019_ _1064_ vssd1 vssd1 vccd1 vccd1 _1069_ sky130_fd_sc_hd__a21oi_1
XFILLER_93_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6979__B _1537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5440_ _0405_ _0412_ vssd1 vssd1 vccd1 vccd1 _0413_ sky130_fd_sc_hd__nor2_1
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5371_ _3328_ _3318_ vssd1 vssd1 vccd1 vccd1 _0344_ sky130_fd_sc_hd__nand2_1
XFILLER_113_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7110_ _2186_ _2187_ _2185_ vssd1 vssd1 vccd1 vccd1 _2208_ sky130_fd_sc_hd__o21ai_1
X_8090_ _1220_ _3283_ vssd1 vssd1 vccd1 vccd1 _0022_ sky130_fd_sc_hd__nor2_1
X_4322_ _1319_ vssd1 vssd1 vccd1 vccd1 _1330_ sky130_fd_sc_hd__clkbuf_4
X_7041_ _2098_ _2124_ _2130_ vssd1 vssd1 vccd1 vccd1 _2132_ sky130_fd_sc_hd__a21o_1
XANTENNA__7493__C1 _2969_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4946__C _3930_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7943_ _3107_ _3114_ _2998_ vssd1 vssd1 vccd1 vccd1 _3125_ sky130_fd_sc_hd__mux2_1
XFILLER_27_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7874_ _3042_ _2937_ vssd1 vssd1 vccd1 vccd1 _3049_ sky130_fd_sc_hd__nor2_1
X_6825_ _1886_ _1892_ _1894_ vssd1 vssd1 vccd1 vccd1 _1895_ sky130_fd_sc_hd__a21oi_2
XFILLER_50_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6756_ _1808_ _1817_ vssd1 vssd1 vccd1 vccd1 _1819_ sky130_fd_sc_hd__and2_1
XFILLER_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5707_ _3762_ _3900_ vssd1 vssd1 vccd1 vccd1 _0685_ sky130_fd_sc_hd__nand2_1
XFILLER_50_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7066__A _4126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6687_ _1741_ _1742_ vssd1 vssd1 vccd1 vccd1 _1743_ sky130_fd_sc_hd__xor2_1
X_5638_ _3762_ _0605_ _0606_ _0608_ _0610_ vssd1 vssd1 vccd1 vccd1 _0611_ sky130_fd_sc_hd__a32o_1
X_8426_ _0635_ _3638_ _0701_ vssd1 vssd1 vccd1 vccd1 _3639_ sky130_fd_sc_hd__or3b_1
XFILLER_117_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8357_ _2611_ _3567_ _3416_ vssd1 vssd1 vccd1 vccd1 _3568_ sky130_fd_sc_hd__a21oi_2
X_5569_ _4139_ _4143_ vssd1 vssd1 vccd1 vccd1 _0542_ sky130_fd_sc_hd__xnor2_1
XFILLER_104_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7308_ _2393_ _2395_ vssd1 vssd1 vccd1 vccd1 _2426_ sky130_fd_sc_hd__xor2_4
XFILLER_104_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8288_ _3479_ _3480_ _3494_ vssd1 vssd1 vccd1 vccd1 _3495_ sky130_fd_sc_hd__a21oi_2
XFILLER_104_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7239_ _2349_ vssd1 vssd1 vccd1 vccd1 _2350_ sky130_fd_sc_hd__inv_2
XFILLER_92_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5014__A1 _3800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6799__B _1510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4525__B1 _3189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4940_ _4070_ _4094_ vssd1 vssd1 vccd1 vccd1 _4095_ sky130_fd_sc_hd__nand2_1
XFILLER_33_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4871_ _4014_ _4025_ vssd1 vssd1 vccd1 vccd1 _4026_ sky130_fd_sc_hd__xor2_1
XANTENNA__5894__A _3792_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6610_ _1656_ _1657_ vssd1 vssd1 vccd1 vccd1 _1658_ sky130_fd_sc_hd__xor2_2
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7590_ _2731_ _2732_ _2735_ vssd1 vssd1 vccd1 vccd1 _2736_ sky130_fd_sc_hd__o21ai_1
X_6541_ _1565_ _1580_ _1581_ vssd1 vssd1 vccd1 vccd1 _1582_ sky130_fd_sc_hd__a21oi_1
XFILLER_20_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6502__B _1538_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6472_ _1490_ _1491_ vssd1 vssd1 vccd1 vccd1 _1507_ sky130_fd_sc_hd__xnor2_1
X_8211_ _3195_ _3411_ _3412_ vssd1 vssd1 vccd1 vccd1 _3413_ sky130_fd_sc_hd__o21ba_1
X_5423_ _0364_ _0394_ _0395_ vssd1 vssd1 vccd1 vccd1 _0396_ sky130_fd_sc_hd__a21o_1
X_5354_ _0250_ _0325_ _0326_ vssd1 vssd1 vccd1 vccd1 _0327_ sky130_fd_sc_hd__o21bai_1
X_8142_ _3265_ _3309_ _3338_ vssd1 vssd1 vccd1 vccd1 _3340_ sky130_fd_sc_hd__nand3_1
XFILLER_114_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4305_ _1135_ vssd1 vssd1 vccd1 vccd1 _0017_ sky130_fd_sc_hd__clkbuf_1
XFILLER_101_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5285_ _3800_ _3615_ vssd1 vssd1 vccd1 vccd1 _0258_ sky130_fd_sc_hd__nor2_1
XANTENNA__4676__C _1748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8073_ _3258_ _3263_ vssd1 vssd1 vccd1 vccd1 _3266_ sky130_fd_sc_hd__and2_1
XFILLER_114_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7024_ _2109_ _2110_ vssd1 vssd1 vccd1 vccd1 _2114_ sky130_fd_sc_hd__xor2_1
XFILLER_68_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5788__B _0702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7926_ _3044_ _3076_ _3105_ vssd1 vssd1 vccd1 vccd1 _3106_ sky130_fd_sc_hd__a21oi_1
XFILLER_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7857_ _3023_ _3029_ vssd1 vssd1 vccd1 vccd1 _3030_ sky130_fd_sc_hd__xnor2_2
XFILLER_23_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6808_ _1863_ _1875_ vssd1 vssd1 vccd1 vccd1 _1876_ sky130_fd_sc_hd__nor2_1
XANTENNA__8194__B1 _3182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7788_ _2918_ _2926_ _2951_ _2953_ _2895_ vssd1 vssd1 vccd1 vccd1 _2954_ sky130_fd_sc_hd__o32ai_4
XFILLER_109_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6739_ _1798_ _1799_ vssd1 vssd1 vccd1 vccd1 _1800_ sky130_fd_sc_hd__xnor2_1
XFILLER_99_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5028__B _3750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8409_ _3621_ _3622_ _0635_ vssd1 vssd1 vccd1 vccd1 _0034_ sky130_fd_sc_hd__a21oi_1
XFILLER_117_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4883__A _2540_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8421__A1 io_out[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8488__A1 in_reg\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4269__S _0712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5070_ _4219_ _4212_ _4224_ vssd1 vssd1 vccd1 vccd1 _4225_ sky130_fd_sc_hd__o21ai_1
XFILLER_84_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5972_ _0963_ _0965_ _0966_ vssd1 vssd1 vccd1 vccd1 _0968_ sky130_fd_sc_hd__or3_1
XFILLER_80_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4923_ _3793_ _3725_ _3959_ vssd1 vssd1 vccd1 vccd1 _4078_ sky130_fd_sc_hd__or3_1
X_7711_ _2856_ _2868_ vssd1 vssd1 vccd1 vccd1 _2869_ sky130_fd_sc_hd__nor2_1
X_4854_ _3996_ _4008_ vssd1 vssd1 vccd1 vccd1 _4009_ sky130_fd_sc_hd__xnor2_1
X_7642_ _2775_ _2792_ _2731_ vssd1 vssd1 vccd1 vccd1 _2794_ sky130_fd_sc_hd__mux2_1
XFILLER_119_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4785_ _3910_ _3911_ vssd1 vssd1 vccd1 vccd1 _3940_ sky130_fd_sc_hd__xnor2_1
X_7573_ _2708_ _2714_ _2717_ vssd1 vssd1 vccd1 vccd1 _2718_ sky130_fd_sc_hd__o21ai_1
XFILLER_119_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6524_ _1559_ _1562_ vssd1 vssd1 vccd1 vccd1 _1564_ sky130_fd_sc_hd__or2b_1
XFILLER_20_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6455_ _1474_ _1477_ vssd1 vssd1 vccd1 vccd1 _1488_ sky130_fd_sc_hd__xor2_1
X_6386_ _1329_ _1306_ _1310_ vssd1 vssd1 vccd1 vccd1 _1412_ sky130_fd_sc_hd__and3_1
X_5406_ _3520_ _0377_ _0378_ _3721_ vssd1 vssd1 vccd1 vccd1 _0379_ sky130_fd_sc_hd__o31ai_4
XFILLER_114_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5337_ _2540_ _0303_ _0308_ _0309_ vssd1 vssd1 vccd1 vccd1 _0310_ sky130_fd_sc_hd__o31a_1
XFILLER_0_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8125_ _2611_ _2576_ _3320_ vssd1 vssd1 vccd1 vccd1 _3321_ sky130_fd_sc_hd__a21oi_4
XFILLER_114_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5268_ _0225_ _0238_ _0240_ vssd1 vssd1 vccd1 vccd1 _0241_ sky130_fd_sc_hd__a21oi_1
X_8056_ _3200_ _3201_ _3208_ vssd1 vssd1 vccd1 vccd1 _3247_ sky130_fd_sc_hd__a21o_1
XFILLER_102_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5799__A _3792_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7007_ _1454_ _1664_ vssd1 vssd1 vccd1 vccd1 _2095_ sky130_fd_sc_hd__or2_1
XFILLER_87_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5199_ _3816_ _3988_ _0167_ vssd1 vssd1 vccd1 vccd1 _0172_ sky130_fd_sc_hd__o21a_1
XANTENNA__8175__A _3182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6965__A1 _1510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4425__C1 posit_add.in2\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7909_ _2908_ _2911_ _2971_ vssd1 vssd1 vccd1 vccd1 _3087_ sky130_fd_sc_hd__mux2_1
XFILLER_12_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7238__B _0082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7381__A1 _4217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4570_ _3722_ _3724_ vssd1 vssd1 vccd1 vccd1 _3725_ sky130_fd_sc_hd__nand2_2
XFILLER_30_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6240_ _1237_ _1249_ _1250_ vssd1 vssd1 vccd1 vccd1 _1251_ sky130_fd_sc_hd__a21boi_1
XFILLER_115_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6171_ _0706_ _1017_ _1028_ _1101_ vssd1 vssd1 vccd1 vccd1 _1176_ sky130_fd_sc_hd__and4_1
XFILLER_97_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5122_ _0091_ _0094_ vssd1 vssd1 vccd1 vccd1 _0095_ sky130_fd_sc_hd__nor2_1
XFILLER_111_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6508__A _1353_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5053_ _4042_ _4151_ _4040_ vssd1 vssd1 vccd1 vccd1 _4208_ sky130_fd_sc_hd__o21ai_1
XFILLER_38_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_635 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5955_ _0931_ _0932_ vssd1 vssd1 vccd1 vccd1 _0950_ sky130_fd_sc_hd__and2_1
XFILLER_80_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5886_ _0866_ _0875_ _0874_ vssd1 vssd1 vccd1 vccd1 _0877_ sky130_fd_sc_hd__a21oi_1
X_4906_ _4057_ _4060_ vssd1 vssd1 vccd1 vccd1 _4061_ sky130_fd_sc_hd__xor2_1
XFILLER_40_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4837_ _3987_ _3991_ vssd1 vssd1 vccd1 vccd1 _3992_ sky130_fd_sc_hd__xor2_1
X_7625_ _2763_ _2774_ _2707_ vssd1 vssd1 vccd1 vccd1 _2775_ sky130_fd_sc_hd__mux2_1
X_4768_ _3917_ _3922_ _3876_ _3729_ vssd1 vssd1 vccd1 vccd1 _3923_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_5_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7556_ _0433_ _2690_ vssd1 vssd1 vccd1 vccd1 _2699_ sky130_fd_sc_hd__or2_1
XFILLER_107_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6507_ _1383_ _1401_ vssd1 vssd1 vccd1 vccd1 _1545_ sky130_fd_sc_hd__or2_1
X_4699_ _3845_ _3853_ vssd1 vssd1 vccd1 vccd1 _3854_ sky130_fd_sc_hd__nor2_1
X_7487_ _3328_ _0347_ vssd1 vssd1 vccd1 vccd1 _2623_ sky130_fd_sc_hd__nand2_1
XFILLER_106_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6438_ _4232_ _1410_ vssd1 vssd1 vccd1 vccd1 _1469_ sky130_fd_sc_hd__or2_1
XFILLER_20_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6369_ _0995_ _1391_ _1392_ vssd1 vssd1 vccd1 vccd1 _1393_ sky130_fd_sc_hd__a21o_1
X_8108_ cmd\[7\] cmd\[6\] _3188_ vssd1 vssd1 vccd1 vccd1 _3303_ sky130_fd_sc_hd__or3_2
XFILLER_102_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6418__A _1446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8039_ _3180_ _3033_ _3165_ vssd1 vssd1 vccd1 vccd1 _3229_ sky130_fd_sc_hd__and3b_1
XFILLER_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7418__A2 _3804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5740_ _3719_ _3815_ _0702_ _0693_ vssd1 vssd1 vccd1 vccd1 _0721_ sky130_fd_sc_hd__or4_2
XFILLER_96_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4282__S _0830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5671_ _0619_ _0614_ _3761_ vssd1 vssd1 vccd1 vccd1 _0645_ sky130_fd_sc_hd__a21oi_1
XFILLER_30_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7410_ _2442_ _2536_ _2537_ _2416_ vssd1 vssd1 vccd1 vccd1 _2538_ sky130_fd_sc_hd__o22ai_1
XANTENNA__7572__C_N _2702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7354__A1 _3986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7593__S _2721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4622_ _3722_ _3754_ _3776_ vssd1 vssd1 vccd1 vccd1 _3777_ sky130_fd_sc_hd__and3_1
X_8390_ _3166_ _3582_ vssd1 vssd1 vccd1 vccd1 _3602_ sky130_fd_sc_hd__or2_1
XFILLER_116_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4553_ _1946_ _2221_ _3707_ _2408_ vssd1 vssd1 vccd1 vccd1 _3708_ sky130_fd_sc_hd__a211o_1
XANTENNA__6510__B _1454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7341_ _1771_ _2461_ vssd1 vssd1 vccd1 vccd1 _2462_ sky130_fd_sc_hd__xnor2_1
XFILLER_116_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4484_ _2661_ _3101_ vssd1 vssd1 vccd1 vccd1 _3112_ sky130_fd_sc_hd__xor2_2
X_7272_ _2347_ _2354_ _2352_ vssd1 vssd1 vccd1 vccd1 _2387_ sky130_fd_sc_hd__a21boi_2
XFILLER_116_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6223_ _1097_ _1164_ vssd1 vssd1 vccd1 vccd1 _1233_ sky130_fd_sc_hd__nand2_1
XFILLER_106_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6154_ _0892_ _1095_ _1119_ vssd1 vssd1 vccd1 vccd1 _1159_ sky130_fd_sc_hd__or3_1
XFILLER_97_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6085_ _1073_ _1083_ _1084_ _1066_ _1085_ vssd1 vssd1 vccd1 vccd1 _1086_ sky130_fd_sc_hd__o221a_1
XFILLER_97_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5105_ _4247_ _0077_ vssd1 vssd1 vccd1 vccd1 _0078_ sky130_fd_sc_hd__xnor2_1
X_5036_ _3994_ _4171_ _4190_ vssd1 vssd1 vccd1 vccd1 _4191_ sky130_fd_sc_hd__a21oi_1
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6987_ _2030_ _2038_ vssd1 vssd1 vccd1 vccd1 _2073_ sky130_fd_sc_hd__xnor2_1
XFILLER_25_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7593__A1 _4153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5938_ _0923_ _0924_ vssd1 vssd1 vccd1 vccd1 _0932_ sky130_fd_sc_hd__xnor2_1
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5869_ _3719_ _0755_ vssd1 vssd1 vccd1 vccd1 _0859_ sky130_fd_sc_hd__nor2_1
X_8588_ clknet_3_3__leaf_clk _0074_ vssd1 vssd1 vccd1 vccd1 posit_add.in2\[15\] sky130_fd_sc_hd__dfxtp_1
X_7608_ _2734_ _2755_ _2731_ vssd1 vssd1 vccd1 vccd1 _2756_ sky130_fd_sc_hd__mux2_1
XFILLER_119_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6420__B _1401_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7539_ _2679_ vssd1 vssd1 vccd1 vccd1 _2680_ sky130_fd_sc_hd__inv_2
XFILLER_107_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6155__A1_N _0702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4891__A _4045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_616 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6910_ _1953_ _1954_ vssd1 vssd1 vccd1 vccd1 _1988_ sky130_fd_sc_hd__nand2_1
XFILLER_47_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7890_ _2915_ vssd1 vssd1 vccd1 vccd1 _3066_ sky130_fd_sc_hd__inv_2
X_6841_ _1422_ _3703_ vssd1 vssd1 vccd1 vccd1 _1912_ sky130_fd_sc_hd__or2_1
XFILLER_62_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8511_ _3695_ vssd1 vssd1 vccd1 vccd1 _0073_ sky130_fd_sc_hd__clkbuf_1
X_6772_ _1750_ _1751_ vssd1 vssd1 vccd1 vccd1 _1837_ sky130_fd_sc_hd__xnor2_1
XFILLER_22_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5723_ _2529_ _0702_ vssd1 vssd1 vccd1 vccd1 _0703_ sky130_fd_sc_hd__nor2_1
XFILLER_31_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5654_ _3699_ _0626_ _3923_ vssd1 vssd1 vccd1 vccd1 _0627_ sky130_fd_sc_hd__o21ai_4
XANTENNA__6521__A _0105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8442_ counter\[4\] _3648_ _3639_ _0679_ vssd1 vssd1 vccd1 vccd1 _3652_ sky130_fd_sc_hd__a211o_1
XFILLER_117_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4605_ _1990_ _3730_ _3732_ _1737_ vssd1 vssd1 vccd1 vccd1 _3760_ sky130_fd_sc_hd__o31a_1
X_8373_ _3481_ _3532_ _3572_ _3584_ vssd1 vssd1 vccd1 vccd1 _3585_ sky130_fd_sc_hd__and4bb_1
X_5585_ _0545_ _0556_ _0557_ vssd1 vssd1 vccd1 vccd1 _0558_ sky130_fd_sc_hd__o21ai_1
X_7324_ _2437_ vssd1 vssd1 vccd1 vccd1 _2444_ sky130_fd_sc_hd__clkinv_2
XFILLER_117_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4536_ _1605_ _3635_ _3651_ _2309_ vssd1 vssd1 vccd1 vccd1 _3659_ sky130_fd_sc_hd__a211o_1
XFILLER_89_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4467_ posit_add.in1\[0\] posit_add.in1\[2\] posit_add.in1\[1\] posit_add.in1\[15\]
+ vssd1 vssd1 vccd1 vccd1 _2925_ sky130_fd_sc_hd__o31a_1
XANTENNA__4976__A _2529_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7255_ _2366_ _0462_ vssd1 vssd1 vccd1 vccd1 _2368_ sky130_fd_sc_hd__nand2_1
X_6206_ _0627_ _1168_ vssd1 vssd1 vccd1 vccd1 _1214_ sky130_fd_sc_hd__or2_1
X_4398_ _1616_ _1627_ _2133_ _2144_ _2155_ vssd1 vssd1 vccd1 vccd1 _2166_ sky130_fd_sc_hd__o32a_1
X_7186_ _2289_ _2291_ vssd1 vssd1 vccd1 vccd1 _2292_ sky130_fd_sc_hd__or2_1
X_6137_ _1138_ _1140_ vssd1 vssd1 vccd1 vccd1 _1141_ sky130_fd_sc_hd__or2b_1
XFILLER_100_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6068_ _0787_ _3739_ _0947_ vssd1 vssd1 vccd1 vccd1 _1068_ sky130_fd_sc_hd__or3b_1
XFILLER_85_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5019_ posit_add.in1\[14\] _3013_ _2584_ vssd1 vssd1 vccd1 vccd1 _4174_ sky130_fd_sc_hd__or3_2
XFILLER_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7527__A _0385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5804__A1 _3735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6606__A _0303_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4543__A1 _3690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5370_ _3068_ _3296_ _3328_ _3035_ vssd1 vssd1 vccd1 vccd1 _0343_ sky130_fd_sc_hd__a211o_1
X_4321_ _1308_ vssd1 vssd1 vccd1 vccd1 _1319_ sky130_fd_sc_hd__clkbuf_2
X_7040_ _2098_ _2124_ _2130_ vssd1 vssd1 vccd1 vccd1 _2131_ sky130_fd_sc_hd__nand3_1
XFILLER_99_468 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7172__A _0080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7942_ _3103_ _3064_ _3085_ _3025_ _3122_ vssd1 vssd1 vccd1 vccd1 _3124_ sky130_fd_sc_hd__a221o_1
XFILLER_82_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5420__A _0369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7873_ _3038_ _3047_ vssd1 vssd1 vccd1 vccd1 _3048_ sky130_fd_sc_hd__nor2_1
XANTENNA__7548__B2 _0351_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6824_ _1835_ _1893_ vssd1 vssd1 vccd1 vccd1 _1894_ sky130_fd_sc_hd__nand2_1
X_6755_ _1808_ _1817_ vssd1 vssd1 vccd1 vccd1 _1818_ sky130_fd_sc_hd__nor2_1
X_5706_ _3700_ _0680_ _0683_ _0654_ vssd1 vssd1 vccd1 vccd1 _0684_ sky130_fd_sc_hd__o22a_1
XFILLER_50_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7066__B _1718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6686_ _1541_ _1542_ vssd1 vssd1 vccd1 vccd1 _1742_ sky130_fd_sc_hd__xnor2_1
X_8425_ _3637_ vssd1 vssd1 vccd1 vccd1 _3638_ sky130_fd_sc_hd__inv_2
X_5637_ _3865_ _3900_ _0609_ _3801_ vssd1 vssd1 vccd1 vccd1 _0610_ sky130_fd_sc_hd__a31o_1
XFILLER_12_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8356_ _2569_ _2495_ _3286_ vssd1 vssd1 vccd1 vccd1 _3567_ sky130_fd_sc_hd__o21ai_1
X_5568_ _0540_ _0475_ _0470_ vssd1 vssd1 vccd1 vccd1 _0541_ sky130_fd_sc_hd__mux2_1
XFILLER_117_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4519_ _3477_ vssd1 vssd1 vccd1 vccd1 _3488_ sky130_fd_sc_hd__clkbuf_4
X_8287_ _3212_ _3486_ _3487_ _3493_ vssd1 vssd1 vccd1 vccd1 _3494_ sky130_fd_sc_hd__a31o_1
X_7307_ _2377_ _2378_ vssd1 vssd1 vccd1 vccd1 _2425_ sky130_fd_sc_hd__nand2_2
X_5499_ _4148_ _4095_ vssd1 vssd1 vccd1 vccd1 _0472_ sky130_fd_sc_hd__or2b_1
X_7238_ _2980_ _0082_ _0400_ vssd1 vssd1 vccd1 vccd1 _2349_ sky130_fd_sc_hd__or3_4
XANTENNA__6039__A1 _0706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7169_ _0080_ _1446_ vssd1 vssd1 vccd1 vccd1 _2273_ sky130_fd_sc_hd__or2_1
XFILLER_85_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6426__A _3930_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5330__A _3988_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5014__A2 _3795_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7475__B1 _1308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4870_ _4023_ _4024_ vssd1 vssd1 vccd1 vccd1 _4025_ sky130_fd_sc_hd__xnor2_1
XFILLER_60_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4290__S _0830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6540_ _1579_ _1578_ vssd1 vssd1 vccd1 vccd1 _1581_ sky130_fd_sc_hd__and2b_1
XFILLER_13_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6471_ _1493_ _1504_ vssd1 vssd1 vccd1 vccd1 _1505_ sky130_fd_sc_hd__xnor2_1
XFILLER_9_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8210_ out_reg\[5\] _3316_ _1231_ out_reg\[6\] vssd1 vssd1 vccd1 vccd1 _3412_ sky130_fd_sc_hd__a22o_1
X_5422_ _0363_ _0356_ vssd1 vssd1 vccd1 vccd1 _0395_ sky130_fd_sc_hd__and2b_1
X_5353_ _0247_ _0249_ vssd1 vssd1 vccd1 vccd1 _0326_ sky130_fd_sc_hd__and2b_1
X_8141_ _0584_ _3337_ _3259_ vssd1 vssd1 vccd1 vccd1 _3338_ sky130_fd_sc_hd__mux2_1
XFILLER_99_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4304_ in_reg\[13\] in_reg\[14\] _0819_ vssd1 vssd1 vccd1 vccd1 _1135_ sky130_fd_sc_hd__mux2_1
XFILLER_114_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5284_ _4179_ _4180_ _0256_ vssd1 vssd1 vccd1 vccd1 _0257_ sky130_fd_sc_hd__a21o_1
X_8072_ _3258_ _3263_ vssd1 vssd1 vccd1 vccd1 _3265_ sky130_fd_sc_hd__nor2_2
XFILLER_99_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7023_ _4153_ _2079_ vssd1 vssd1 vccd1 vccd1 _2113_ sky130_fd_sc_hd__nand2_1
XFILLER_87_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7925_ _3044_ _3104_ _3061_ _3038_ vssd1 vssd1 vccd1 vccd1 _3105_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_63_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7856_ _3025_ _3027_ _3028_ vssd1 vssd1 vccd1 vccd1 _3029_ sky130_fd_sc_hd__a21o_1
X_6807_ _1872_ _1874_ _1870_ vssd1 vssd1 vccd1 vccd1 _1875_ sky130_fd_sc_hd__a21oi_1
XFILLER_11_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4999_ _3929_ _3931_ _4026_ _4025_ _4014_ vssd1 vssd1 vccd1 vccd1 _4154_ sky130_fd_sc_hd__a32o_1
XFILLER_11_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7787_ _2952_ _2916_ _2902_ vssd1 vssd1 vccd1 vccd1 _2953_ sky130_fd_sc_hd__a21oi_1
X_6738_ _1710_ _1719_ vssd1 vssd1 vccd1 vccd1 _1799_ sky130_fd_sc_hd__xor2_1
XFILLER_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6669_ _1683_ _1687_ vssd1 vssd1 vccd1 vccd1 _1723_ sky130_fd_sc_hd__nand2_1
XFILLER_99_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8408_ out_reg\[14\] _3197_ vssd1 vssd1 vccd1 vccd1 _3622_ sky130_fd_sc_hd__nand2_1
XFILLER_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8339_ _3190_ _3540_ _3548_ _1177_ vssd1 vssd1 vccd1 vccd1 _3549_ sky130_fd_sc_hd__a211o_1
XFILLER_105_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4883__B _4037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6156__A _1097_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5060__A _3802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5995__A _0991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7932__A1 _2937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5171__A1 _3701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7620__A0 _4045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5971_ _0879_ _0964_ _0917_ _0915_ vssd1 vssd1 vccd1 vccd1 _0966_ sky130_fd_sc_hd__o211a_1
XFILLER_65_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4922_ _4074_ _4076_ vssd1 vssd1 vccd1 vccd1 _4077_ sky130_fd_sc_hd__xnor2_1
X_7710_ _2861_ _2864_ _2867_ vssd1 vssd1 vccd1 vccd1 _2868_ sky130_fd_sc_hd__nand3b_1
X_7641_ _2784_ _2791_ _2708_ vssd1 vssd1 vccd1 vccd1 _2792_ sky130_fd_sc_hd__mux2_1
XFILLER_100_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4853_ _3998_ _4007_ vssd1 vssd1 vccd1 vccd1 _4008_ sky130_fd_sc_hd__xnor2_1
XFILLER_60_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4784_ _3799_ _3938_ vssd1 vssd1 vccd1 vccd1 _3939_ sky130_fd_sc_hd__xnor2_1
XFILLER_20_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7572_ _0391_ _2715_ _2702_ vssd1 vssd1 vccd1 vccd1 _2717_ sky130_fd_sc_hd__or3b_1
X_6523_ _1559_ _1562_ vssd1 vssd1 vccd1 vccd1 _1563_ sky130_fd_sc_hd__xnor2_1
XFILLER_20_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6454_ _4217_ _1482_ _1485_ _1486_ vssd1 vssd1 vccd1 vccd1 _1487_ sky130_fd_sc_hd__a31o_1
XFILLER_118_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5405_ _3819_ _3530_ _3848_ _3446_ vssd1 vssd1 vccd1 vccd1 _0378_ sky130_fd_sc_hd__o211a_1
X_6385_ _4228_ _1410_ vssd1 vssd1 vccd1 vccd1 _1411_ sky130_fd_sc_hd__or2_1
XFILLER_114_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5336_ _0307_ _0304_ vssd1 vssd1 vccd1 vccd1 _0309_ sky130_fd_sc_hd__or2b_1
XFILLER_0_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8124_ _2569_ _2495_ _3286_ _2520_ vssd1 vssd1 vccd1 vccd1 _3320_ sky130_fd_sc_hd__o211a_1
X_5267_ _0195_ _0239_ vssd1 vssd1 vccd1 vccd1 _0240_ sky130_fd_sc_hd__or2b_1
X_8055_ _1220_ _3246_ vssd1 vssd1 vccd1 vccd1 _0021_ sky130_fd_sc_hd__nor2_1
X_7006_ _2092_ _2093_ vssd1 vssd1 vccd1 vccd1 _2094_ sky130_fd_sc_hd__xnor2_1
XFILLER_87_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5198_ _0169_ _0170_ vssd1 vssd1 vccd1 vccd1 _0171_ sky130_fd_sc_hd__nand2_1
XFILLER_95_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7611__A0 _3816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6965__A2 _3703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7908_ _3063_ _3073_ _2999_ vssd1 vssd1 vccd1 vccd1 _3086_ sky130_fd_sc_hd__mux2_1
XFILLER_71_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7839_ _2842_ _2973_ vssd1 vssd1 vccd1 vccd1 _3010_ sky130_fd_sc_hd__or2_1
XFILLER_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5055__A _4017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8158__A1 _1330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_73 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5392__A1 _3690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6170_ _1016_ _1008_ _1017_ vssd1 vssd1 vccd1 vccd1 _1175_ sky130_fd_sc_hd__or3b_1
XFILLER_97_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5121_ _0092_ _0093_ _0075_ vssd1 vssd1 vccd1 vccd1 _0094_ sky130_fd_sc_hd__o21a_1
XFILLER_57_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6508__B _1354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5052_ _4205_ _4206_ vssd1 vssd1 vccd1 vccd1 _4207_ sky130_fd_sc_hd__xnor2_1
XFILLER_65_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5954_ _0945_ _0947_ _0948_ vssd1 vssd1 vccd1 vccd1 _0949_ sky130_fd_sc_hd__and3_1
XFILLER_80_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5885_ _0866_ _0874_ _0875_ vssd1 vssd1 vccd1 vccd1 _0876_ sky130_fd_sc_hd__and3_1
XFILLER_61_691 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4905_ _4058_ _4059_ vssd1 vssd1 vccd1 vccd1 _4060_ sky130_fd_sc_hd__or2_1
X_4836_ _3893_ _3854_ _3990_ vssd1 vssd1 vccd1 vccd1 _3991_ sky130_fd_sc_hd__a21o_1
X_7624_ _3883_ _3776_ _2652_ vssd1 vssd1 vccd1 vccd1 _2774_ sky130_fd_sc_hd__mux2_1
XFILLER_21_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7555_ _0433_ _2690_ vssd1 vssd1 vccd1 vccd1 _2698_ sky130_fd_sc_hd__nand2_1
X_6506_ _1353_ _1354_ _0147_ vssd1 vssd1 vccd1 vccd1 _1544_ sky130_fd_sc_hd__and3_1
X_4767_ _3736_ _3921_ _1748_ vssd1 vssd1 vccd1 vccd1 _3922_ sky130_fd_sc_hd__o21ai_1
X_4698_ _3772_ _3846_ _3851_ _3852_ vssd1 vssd1 vccd1 vccd1 _3853_ sky130_fd_sc_hd__o31a_1
X_7486_ _2610_ _2618_ _2521_ vssd1 vssd1 vccd1 vccd1 _2622_ sky130_fd_sc_hd__a21oi_1
X_6437_ _1464_ _1467_ vssd1 vssd1 vccd1 vccd1 _1468_ sky130_fd_sc_hd__xnor2_1
XFILLER_115_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6368_ _1338_ vssd1 vssd1 vccd1 vccd1 _1392_ sky130_fd_sc_hd__inv_2
XFILLER_96_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5319_ _4168_ _4169_ _4166_ vssd1 vssd1 vccd1 vccd1 _0292_ sky130_fd_sc_hd__o21ba_1
X_8107_ _3295_ _3301_ vssd1 vssd1 vccd1 vccd1 _3302_ sky130_fd_sc_hd__nor2_1
X_6299_ _1002_ _1102_ _1001_ vssd1 vssd1 vccd1 vccd1 _1316_ sky130_fd_sc_hd__a21o_1
XFILLER_88_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6418__B _1384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8038_ _3181_ _3183_ vssd1 vssd1 vccd1 vccd1 _3228_ sky130_fd_sc_hd__and2_1
XFILLER_75_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8388__A1 _3195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6434__A _0218_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4889__A _3729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7712__B _2802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6609__A _1384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5670_ _0642_ _0638_ vssd1 vssd1 vccd1 vccd1 _0644_ sky130_fd_sc_hd__xnor2_1
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4621_ _3775_ vssd1 vssd1 vccd1 vccd1 _3776_ sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_0_clk_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4552_ _1726_ _2353_ _2364_ _1913_ vssd1 vssd1 vccd1 vccd1 _3707_ sky130_fd_sc_hd__o211a_1
X_7340_ _2263_ _2456_ vssd1 vssd1 vccd1 vccd1 _2461_ sky130_fd_sc_hd__nor2_1
X_4483_ posit_add.in1\[11\] _3090_ vssd1 vssd1 vccd1 vccd1 _3101_ sky130_fd_sc_hd__xnor2_4
X_7271_ _2384_ _2354_ vssd1 vssd1 vccd1 vccd1 _2385_ sky130_fd_sc_hd__nand2_1
XFILLER_116_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6222_ _1229_ _1230_ vssd1 vssd1 vccd1 vccd1 _1232_ sky130_fd_sc_hd__xor2_1
X_6153_ _1140_ _1138_ vssd1 vssd1 vccd1 vccd1 _1158_ sky130_fd_sc_hd__xor2_1
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6084_ _1068_ _1070_ vssd1 vssd1 vccd1 vccd1 _1085_ sky130_fd_sc_hd__and2_1
XFILLER_85_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5104_ _0075_ _0076_ vssd1 vssd1 vccd1 vccd1 _0077_ sky130_fd_sc_hd__nand2_1
XFILLER_111_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5035_ _4181_ _4189_ vssd1 vssd1 vccd1 vccd1 _4190_ sky130_fd_sc_hd__xnor2_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6986_ _2062_ _2070_ _2071_ vssd1 vssd1 vccd1 vccd1 _2072_ sky130_fd_sc_hd__o21a_1
XFILLER_53_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5937_ _0762_ _3832_ vssd1 vssd1 vccd1 vccd1 _0931_ sky130_fd_sc_hd__nand2_1
XFILLER_13_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5868_ _0854_ _0856_ _0857_ vssd1 vssd1 vccd1 vccd1 _0858_ sky130_fd_sc_hd__a21bo_1
X_7607_ _2744_ _2754_ _2708_ vssd1 vssd1 vccd1 vccd1 _2755_ sky130_fd_sc_hd__mux2_1
X_5799_ _3792_ _0782_ vssd1 vssd1 vccd1 vccd1 _0783_ sky130_fd_sc_hd__xnor2_1
X_8587_ clknet_3_5__leaf_clk _0073_ vssd1 vssd1 vccd1 vccd1 posit_add.in2\[14\] sky130_fd_sc_hd__dfxtp_4
X_4819_ _3971_ _3973_ vssd1 vssd1 vccd1 vccd1 _3974_ sky130_fd_sc_hd__and2_1
XFILLER_21_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7538_ _0427_ _2656_ _2651_ vssd1 vssd1 vccd1 vccd1 _2679_ sky130_fd_sc_hd__mux2_1
X_7469_ _2600_ _2601_ _2602_ vssd1 vssd1 vccd1 vccd1 _2603_ sky130_fd_sc_hd__a21bo_1
XANTENNA__5108__A1 _0080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6752__A2_N _0121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4891__B _3986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6164__A _0795_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_1__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_113_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6339__A _0627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6840_ _1904_ _1910_ vssd1 vssd1 vccd1 vccd1 _1911_ sky130_fd_sc_hd__xnor2_1
XANTENNA__8221__B1 _2621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6771_ _1833_ _1834_ vssd1 vssd1 vccd1 vccd1 _1835_ sky130_fd_sc_hd__nand2_1
XFILLER_23_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5722_ _0700_ vssd1 vssd1 vccd1 vccd1 _0702_ sky130_fd_sc_hd__clkbuf_4
X_8510_ posit_add.in2\[14\] in_reg\[14\] _3676_ vssd1 vssd1 vccd1 vccd1 _3695_ sky130_fd_sc_hd__mux2_1
X_5653_ _3864_ _0619_ _0112_ vssd1 vssd1 vccd1 vccd1 _0626_ sky130_fd_sc_hd__a21oi_2
X_8441_ _3650_ vssd1 vssd1 vccd1 vccd1 _0041_ sky130_fd_sc_hd__clkbuf_1
XFILLER_30_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4604_ _3757_ _3758_ _2485_ vssd1 vssd1 vccd1 vccd1 _3759_ sky130_fd_sc_hd__a21o_1
X_8372_ _3166_ _3569_ _3570_ vssd1 vssd1 vccd1 vccd1 _3584_ sky130_fd_sc_hd__or3_1
X_5584_ _0494_ vssd1 vssd1 vccd1 vccd1 _0557_ sky130_fd_sc_hd__buf_2
X_4535_ _1726_ _2353_ _2364_ _3643_ vssd1 vssd1 vccd1 vccd1 _3651_ sky130_fd_sc_hd__o211a_1
X_7323_ _2437_ _2438_ _2440_ _2442_ vssd1 vssd1 vccd1 vccd1 _2443_ sky130_fd_sc_hd__o22ai_2
XFILLER_117_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4976__B _4126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4466_ _2661_ _2903_ vssd1 vssd1 vccd1 vccd1 _2914_ sky130_fd_sc_hd__xnor2_1
X_7254_ _2366_ _0462_ vssd1 vssd1 vccd1 vccd1 _2367_ sky130_fd_sc_hd__or2_1
X_6205_ _1194_ _1195_ _1212_ vssd1 vssd1 vccd1 vccd1 _1213_ sky130_fd_sc_hd__o21a_1
XFILLER_89_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4397_ _1781_ _1583_ vssd1 vssd1 vccd1 vccd1 _2155_ sky130_fd_sc_hd__nor2_1
X_7185_ _1622_ _1647_ _2290_ vssd1 vssd1 vccd1 vccd1 _2291_ sky130_fd_sc_hd__a21oi_1
X_6136_ _0627_ _1095_ _1129_ _1139_ vssd1 vssd1 vccd1 vccd1 _1140_ sky130_fd_sc_hd__o31ai_2
XFILLER_58_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6067_ _1057_ _1060_ _1066_ vssd1 vssd1 vccd1 vccd1 _1067_ sky130_fd_sc_hd__a21o_1
XFILLER_100_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5018_ _3881_ _3894_ vssd1 vssd1 vccd1 vccd1 _4173_ sky130_fd_sc_hd__nand2_1
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6969_ _1510_ _4126_ _2050_ _2052_ vssd1 vssd1 vccd1 vccd1 _2053_ sky130_fd_sc_hd__o31ai_1
XFILLER_13_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4537__C1 _1946_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5063__A _3802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5998__A _0795_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8451__A0 in_reg\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6606__B _1510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6622__A _1423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5238__A _3828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4320_ _1297_ vssd1 vssd1 vccd1 vccd1 _1308_ sky130_fd_sc_hd__clkbuf_4
XFILLER_113_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4288__S _0830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7493__A1 posit_add.in1\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_392 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7941_ _3020_ _3121_ vssd1 vssd1 vccd1 vccd1 _3122_ sky130_fd_sc_hd__and2_1
XFILLER_82_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7872_ _3044_ _3045_ vssd1 vssd1 vccd1 vccd1 _3047_ sky130_fd_sc_hd__or2_1
XFILLER_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6823_ _1833_ _1834_ vssd1 vssd1 vccd1 vccd1 _1893_ sky130_fd_sc_hd__or2_1
XFILLER_63_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6754_ _1806_ _1810_ _1811_ _1816_ vssd1 vssd1 vccd1 vccd1 _1817_ sky130_fd_sc_hd__a22oi_2
XFILLER_11_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5705_ _0681_ _0613_ _0663_ _0666_ _0682_ vssd1 vssd1 vccd1 vccd1 _0683_ sky130_fd_sc_hd__a32o_1
X_6685_ _1696_ _1699_ _1740_ vssd1 vssd1 vccd1 vccd1 _1741_ sky130_fd_sc_hd__a21bo_1
XFILLER_31_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5636_ _1748_ _2507_ _3775_ vssd1 vssd1 vccd1 vccd1 _0609_ sky130_fd_sc_hd__a21o_2
XANTENNA__5148__A _4174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8424_ counter\[3\] _3636_ _0668_ counter\[4\] vssd1 vssd1 vccd1 vccd1 _3637_ sky130_fd_sc_hd__or4b_1
XFILLER_12_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8355_ _3563_ _3564_ _3303_ vssd1 vssd1 vccd1 vccd1 _3566_ sky130_fd_sc_hd__a21oi_1
X_5567_ _0539_ _0473_ _0338_ vssd1 vssd1 vccd1 vccd1 _0540_ sky130_fd_sc_hd__mux2_1
XFILLER_117_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8286_ _3489_ _3491_ _3492_ vssd1 vssd1 vccd1 vccd1 _3493_ sky130_fd_sc_hd__a21oi_1
XFILLER_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5498_ _0339_ _0341_ _0470_ vssd1 vssd1 vccd1 vccd1 _0471_ sky130_fd_sc_hd__mux2_1
X_7306_ _1676_ _2412_ _2335_ _2414_ _2423_ vssd1 vssd1 vccd1 vccd1 _2424_ sky130_fd_sc_hd__a221oi_4
X_4518_ _3046_ _3424_ vssd1 vssd1 vccd1 vccd1 _3477_ sky130_fd_sc_hd__or2_2
X_4449_ posit_add.in1\[10\] _2716_ vssd1 vssd1 vccd1 vccd1 _2727_ sky130_fd_sc_hd__xnor2_4
X_7237_ _0351_ _2345_ _2347_ vssd1 vssd1 vccd1 vccd1 _2348_ sky130_fd_sc_hd__o21a_1
XFILLER_104_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7168_ _1588_ _4251_ _1498_ vssd1 vssd1 vccd1 vccd1 _2272_ sky130_fd_sc_hd__and3_1
XFILLER_112_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6119_ _1120_ _1121_ vssd1 vssd1 vccd1 vccd1 _1122_ sky130_fd_sc_hd__xnor2_1
XFILLER_100_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7099_ _2184_ _2195_ vssd1 vssd1 vccd1 vccd1 _2196_ sky130_fd_sc_hd__nor2_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6442__A _1399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5058__A _4210_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4897__A _3892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6617__A _1665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5410__B1 _3690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6470_ _1503_ _1450_ vssd1 vssd1 vccd1 vccd1 _1504_ sky130_fd_sc_hd__xor2_1
XFILLER_9_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5421_ _0375_ _0392_ _0393_ vssd1 vssd1 vccd1 vccd1 _0394_ sky130_fd_sc_hd__a21o_1
X_5352_ _0282_ _0324_ _0280_ vssd1 vssd1 vccd1 vccd1 _0325_ sky130_fd_sc_hd__a21oi_1
X_8140_ _0557_ _0527_ _3306_ vssd1 vssd1 vccd1 vccd1 _3337_ sky130_fd_sc_hd__o21a_1
XFILLER_114_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6269__A2 _1128_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4303_ _1114_ vssd1 vssd1 vccd1 vccd1 _0016_ sky130_fd_sc_hd__clkbuf_1
X_8071_ _3259_ _0585_ _3262_ vssd1 vssd1 vccd1 vccd1 _3263_ sky130_fd_sc_hd__o21ai_1
X_7022_ _2109_ _2110_ vssd1 vssd1 vccd1 vccd1 _2112_ sky130_fd_sc_hd__or2_1
XFILLER_87_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5283_ _3893_ _3854_ _4178_ vssd1 vssd1 vccd1 vccd1 _0256_ sky130_fd_sc_hd__and3_1
XFILLER_59_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6527__A _0080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8415__B1 _2319_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7924_ _2906_ _2908_ _3034_ vssd1 vssd1 vccd1 vccd1 _3104_ sky130_fd_sc_hd__mux2_1
XFILLER_24_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7855_ _2993_ _3020_ vssd1 vssd1 vccd1 vccd1 _3028_ sky130_fd_sc_hd__and2_1
XFILLER_36_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6806_ _1873_ _1849_ vssd1 vssd1 vccd1 vccd1 _1874_ sky130_fd_sc_hd__xnor2_1
XFILLER_23_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4998_ _3838_ vssd1 vssd1 vccd1 vccd1 _4153_ sky130_fd_sc_hd__buf_4
XFILLER_51_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7786_ _2906_ _2908_ vssd1 vssd1 vccd1 vccd1 _2952_ sky130_fd_sc_hd__nor2_1
X_6737_ _1786_ _1796_ _1797_ vssd1 vssd1 vccd1 vccd1 _1798_ sky130_fd_sc_hd__o21ai_2
XFILLER_23_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6668_ _1683_ _1687_ vssd1 vssd1 vccd1 vccd1 _1722_ sky130_fd_sc_hd__nor2_1
X_6599_ _1606_ _1607_ _1645_ vssd1 vssd1 vccd1 vccd1 _1646_ sky130_fd_sc_hd__o21a_1
X_5619_ _0441_ _0455_ _0518_ _0519_ _0557_ vssd1 vssd1 vccd1 vccd1 _0592_ sky130_fd_sc_hd__a32o_1
X_8407_ _3608_ _3613_ _3619_ _3620_ _3195_ vssd1 vssd1 vccd1 vccd1 _3621_ sky130_fd_sc_hd__a32o_1
X_8338_ _3546_ _3547_ vssd1 vssd1 vccd1 vccd1 _3548_ sky130_fd_sc_hd__and2b_1
XFILLER_117_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7457__A1 _2381_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8269_ _3234_ _3233_ _3438_ vssd1 vssd1 vccd1 vccd1 _3474_ sky130_fd_sc_hd__o21ba_1
XANTENNA__7821__A _2980_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7540__B _1781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6156__B _1128_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5060__B _3838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6196__B2 _0706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5171__A2 _4037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5970_ _0915_ _0917_ _0964_ _0879_ vssd1 vssd1 vccd1 vccd1 _0965_ sky130_fd_sc_hd__a211oi_1
XFILLER_52_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7620__A1 _0147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4921_ _3878_ _3907_ _3789_ _4075_ vssd1 vssd1 vccd1 vccd1 _4076_ sky130_fd_sc_hd__a31oi_2
X_4852_ _4005_ _4006_ vssd1 vssd1 vccd1 vccd1 _4007_ sky130_fd_sc_hd__and2_1
X_7640_ _1531_ _3878_ _2713_ vssd1 vssd1 vccd1 vccd1 _2791_ sky130_fd_sc_hd__mux2_1
X_4783_ _3728_ _3806_ vssd1 vssd1 vccd1 vccd1 _3938_ sky130_fd_sc_hd__nand2_1
X_7571_ _3855_ _3802_ _2652_ vssd1 vssd1 vccd1 vccd1 _2715_ sky130_fd_sc_hd__mux2_1
X_6522_ _1449_ _0148_ _1457_ _1560_ vssd1 vssd1 vccd1 vccd1 _1562_ sky130_fd_sc_hd__o211a_1
XFILLER_119_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6453_ _1469_ _1416_ vssd1 vssd1 vccd1 vccd1 _1486_ sky130_fd_sc_hd__nor2_1
XFILLER_9_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7687__A1 _4250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5404_ _2727_ _3530_ _0352_ _3488_ vssd1 vssd1 vccd1 vccd1 _0377_ sky130_fd_sc_hd__o211a_1
X_6384_ _1408_ _1409_ vssd1 vssd1 vccd1 vccd1 _1410_ sky130_fd_sc_hd__nand2_2
X_8123_ _3249_ _3252_ _3289_ vssd1 vssd1 vccd1 vccd1 _3319_ sky130_fd_sc_hd__or3_2
X_5335_ _0304_ _0307_ vssd1 vssd1 vccd1 vccd1 _0308_ sky130_fd_sc_hd__xor2_1
XFILLER_87_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5266_ _0192_ _0194_ vssd1 vssd1 vccd1 vccd1 _0239_ sky130_fd_sc_hd__nand2_1
X_8054_ out_reg\[1\] _3197_ _3245_ vssd1 vssd1 vccd1 vccd1 _3246_ sky130_fd_sc_hd__a21oi_1
X_7005_ _2015_ _2051_ _2050_ vssd1 vssd1 vccd1 vccd1 _2093_ sky130_fd_sc_hd__o21ba_1
X_5197_ _0137_ _0168_ _3875_ _0124_ vssd1 vssd1 vccd1 vccd1 _0170_ sky130_fd_sc_hd__o22ai_1
XFILLER_28_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7611__A1 _1384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7907_ _3065_ _3084_ vssd1 vssd1 vccd1 vccd1 _3085_ sky130_fd_sc_hd__and2_1
XFILLER_24_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7838_ _2974_ _2975_ vssd1 vssd1 vccd1 vccd1 _3009_ sky130_fd_sc_hd__xor2_1
XFILLER_11_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7769_ _2932_ vssd1 vssd1 vccd1 vccd1 _2933_ sky130_fd_sc_hd__inv_2
XFILLER_109_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_704 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5120_ _4254_ _0084_ _4252_ vssd1 vssd1 vccd1 vccd1 _0093_ sky130_fd_sc_hd__o21bai_1
XFILLER_111_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4296__S _0819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5051_ _4036_ _4038_ _4033_ _4035_ vssd1 vssd1 vccd1 vccd1 _4206_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__4655__A1 _1858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6508__C _3986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5953_ _3792_ _0787_ vssd1 vssd1 vccd1 vccd1 _0948_ sky130_fd_sc_hd__nor2_1
XFILLER_80_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5884_ _0838_ _0839_ _0837_ vssd1 vssd1 vccd1 vccd1 _0875_ sky130_fd_sc_hd__a21o_1
XFILLER_61_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4904_ _4053_ _4054_ vssd1 vssd1 vccd1 vccd1 _4059_ sky130_fd_sc_hd__xnor2_1
XFILLER_21_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4835_ _3828_ _3988_ _3989_ _3845_ vssd1 vssd1 vccd1 vccd1 _3990_ sky130_fd_sc_hd__o22a_1
X_7623_ _2770_ _2772_ vssd1 vssd1 vccd1 vccd1 _2773_ sky130_fd_sc_hd__nand2_1
XFILLER_33_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4766_ _3918_ _3920_ _3830_ vssd1 vssd1 vccd1 vccd1 _3921_ sky130_fd_sc_hd__mux2_1
X_7554_ _0416_ _2695_ vssd1 vssd1 vccd1 vccd1 _2697_ sky130_fd_sc_hd__xnor2_1
XFILLER_119_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6505_ _1541_ _1542_ vssd1 vssd1 vccd1 vccd1 _1543_ sky130_fd_sc_hd__nor2_1
XFILLER_119_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4697_ _3772_ _3724_ vssd1 vssd1 vccd1 vccd1 _3852_ sky130_fd_sc_hd__nand2_1
XFILLER_20_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7485_ _2620_ vssd1 vssd1 vccd1 vccd1 _2621_ sky130_fd_sc_hd__buf_2
X_6436_ _1465_ _1466_ vssd1 vssd1 vccd1 vccd1 _1467_ sky130_fd_sc_hd__xnor2_1
XFILLER_88_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6367_ _1387_ _1390_ vssd1 vssd1 vccd1 vccd1 _1391_ sky130_fd_sc_hd__xnor2_1
X_5318_ _0288_ _0290_ vssd1 vssd1 vccd1 vccd1 _0291_ sky130_fd_sc_hd__or2b_1
X_8106_ _3297_ _3300_ vssd1 vssd1 vccd1 vccd1 _3301_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6298_ _1145_ _1148_ _1314_ vssd1 vssd1 vccd1 vccd1 _1315_ sky130_fd_sc_hd__a21oi_1
XFILLER_88_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5843__B1 _3832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5249_ _0217_ _0221_ vssd1 vssd1 vccd1 vccd1 _0222_ sky130_fd_sc_hd__nand2_1
X_8037_ _3226_ vssd1 vssd1 vccd1 vccd1 _3227_ sky130_fd_sc_hd__buf_2
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8388__A2 _3599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6434__B _1353_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6450__A _1423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6609__B _1423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7587__A0 _4153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7305__A_N _2416_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4620_ _1990_ _3713_ _3715_ _3774_ _3678_ vssd1 vssd1 vccd1 vccd1 _3775_ sky130_fd_sc_hd__a311oi_4
X_4551_ _3643_ _2221_ _3705_ _2309_ vssd1 vssd1 vccd1 vccd1 _3706_ sky130_fd_sc_hd__a211o_1
X_4482_ posit_add.in1\[10\] _2573_ _1253_ vssd1 vssd1 vccd1 vccd1 _3090_ sky130_fd_sc_hd__o21ai_2
X_7270_ _0351_ _2345_ _2380_ _2383_ _2347_ vssd1 vssd1 vccd1 vccd1 _2384_ sky130_fd_sc_hd__o2111a_1
XFILLER_116_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6221_ _0702_ _1168_ vssd1 vssd1 vccd1 vccd1 _1230_ sky130_fd_sc_hd__nor2_1
X_6152_ _1154_ _1155_ vssd1 vssd1 vccd1 vccd1 _1157_ sky130_fd_sc_hd__or2_1
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5103_ _4234_ _4248_ _4256_ vssd1 vssd1 vccd1 vccd1 _0076_ sky130_fd_sc_hd__or3_1
X_6083_ _1062_ _1065_ vssd1 vssd1 vccd1 vccd1 _1084_ sky130_fd_sc_hd__nor2_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5034_ _4187_ _4188_ vssd1 vssd1 vccd1 vccd1 _4189_ sky130_fd_sc_hd__nand2_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6985_ _2060_ _2061_ vssd1 vssd1 vccd1 vccd1 _2071_ sky130_fd_sc_hd__or2b_1
XFILLER_53_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5936_ _0888_ _0903_ _0902_ vssd1 vssd1 vccd1 vccd1 _0930_ sky130_fd_sc_hd__a21oi_1
XFILLER_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5867_ _2529_ _0693_ _0855_ vssd1 vssd1 vccd1 vccd1 _0857_ sky130_fd_sc_hd__or3_1
X_7606_ _3986_ _3901_ _2652_ vssd1 vssd1 vccd1 vccd1 _2754_ sky130_fd_sc_hd__mux2_1
X_5798_ _0780_ _0781_ vssd1 vssd1 vccd1 vccd1 _0782_ sky130_fd_sc_hd__nand2_1
X_8586_ clknet_3_5__leaf_clk _0072_ vssd1 vssd1 vccd1 vccd1 posit_add.in2\[13\] sky130_fd_sc_hd__dfxtp_2
X_4818_ _3972_ _3956_ vssd1 vssd1 vccd1 vccd1 _3973_ sky130_fd_sc_hd__and2b_1
X_4749_ _3871_ _3782_ _3870_ vssd1 vssd1 vccd1 vccd1 _3904_ sky130_fd_sc_hd__o21ba_1
X_7537_ _0345_ _0342_ _2651_ vssd1 vssd1 vccd1 vccd1 _2678_ sky130_fd_sc_hd__mux2_1
XFILLER_110_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7468_ _2594_ _2567_ _2514_ vssd1 vssd1 vccd1 vccd1 _2602_ sky130_fd_sc_hd__mux2_1
XFILLER_31_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5108__A2 _3925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6419_ _1447_ _0105_ vssd1 vssd1 vccd1 vccd1 _1448_ sky130_fd_sc_hd__nand2_1
X_7399_ _2425_ _2426_ _2427_ _2443_ vssd1 vssd1 vccd1 vccd1 _2526_ sky130_fd_sc_hd__a31o_1
XFILLER_103_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6164__B _1128_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5752__C1 _3866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7272__A2 _2354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6770_ _1830_ _1774_ vssd1 vssd1 vccd1 vccd1 _1834_ sky130_fd_sc_hd__xnor2_1
XFILLER_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5721_ _3923_ _0694_ _0696_ _0699_ vssd1 vssd1 vccd1 vccd1 _0700_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_50_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5652_ _3901_ _0624_ vssd1 vssd1 vccd1 vccd1 _0625_ sky130_fd_sc_hd__nand2_1
X_8440_ _3648_ _3641_ _3649_ vssd1 vssd1 vccd1 vccd1 _3650_ sky130_fd_sc_hd__and3b_1
XFILLER_31_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4603_ _1913_ _2221_ _2232_ _2408_ vssd1 vssd1 vccd1 vccd1 _3758_ sky130_fd_sc_hd__a211o_1
X_8371_ _3416_ _3580_ _3581_ vssd1 vssd1 vccd1 vccd1 _3582_ sky130_fd_sc_hd__or3b_1
X_5583_ _0510_ _0543_ _0555_ vssd1 vssd1 vccd1 vccd1 _0556_ sky130_fd_sc_hd__a21o_1
XFILLER_30_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4534_ _1660_ vssd1 vssd1 vccd1 vccd1 _3643_ sky130_fd_sc_hd__inv_2
XFILLER_7_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7322_ _2416_ _2431_ vssd1 vssd1 vccd1 vccd1 _2442_ sky130_fd_sc_hd__nand2_1
XFILLER_117_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4465_ posit_add.in1\[4\] _2892_ vssd1 vssd1 vccd1 vccd1 _2903_ sky130_fd_sc_hd__xnor2_4
X_7253_ _0405_ _0412_ vssd1 vssd1 vccd1 vccd1 _2366_ sky130_fd_sc_hd__and2b_1
X_6204_ _1192_ _1193_ vssd1 vssd1 vccd1 vccd1 _1212_ sky130_fd_sc_hd__or2_1
X_4396_ _1506_ _1583_ vssd1 vssd1 vccd1 vccd1 _2144_ sky130_fd_sc_hd__and2_1
X_7184_ _1644_ _1646_ vssd1 vssd1 vccd1 vccd1 _2290_ sky130_fd_sc_hd__nor2_1
X_6135_ _1128_ _1131_ vssd1 vssd1 vccd1 vccd1 _1139_ sky130_fd_sc_hd__nand2_1
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6066_ _1062_ _1065_ vssd1 vssd1 vccd1 vccd1 _1066_ sky130_fd_sc_hd__and2_1
XFILLER_100_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5017_ _3893_ _3854_ vssd1 vssd1 vccd1 vccd1 _4172_ sky130_fd_sc_hd__nand2_1
XFILLER_100_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6968_ _2015_ _2051_ vssd1 vssd1 vccd1 vccd1 _2052_ sky130_fd_sc_hd__or2_1
XFILLER_13_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5919_ _0910_ _0911_ vssd1 vssd1 vccd1 vccd1 _0912_ sky130_fd_sc_hd__xor2_1
X_6899_ _1422_ _4126_ vssd1 vssd1 vccd1 vccd1 _1976_ sky130_fd_sc_hd__nor2_1
XFILLER_108_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8569_ clknet_3_4__leaf_clk _0055_ vssd1 vssd1 vccd1 vccd1 posit_add.in1\[12\] sky130_fd_sc_hd__dfxtp_2
XFILLER_107_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5063__B _4217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6622__B _1401_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7718__B _2780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7714__B1 _2800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5238__B _4037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7940_ _3108_ _3120_ _3006_ vssd1 vssd1 vccd1 vccd1 _3121_ sky130_fd_sc_hd__mux2_1
XFILLER_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7871_ _2933_ _2928_ _3034_ vssd1 vssd1 vccd1 vccd1 _3045_ sky130_fd_sc_hd__mux2_1
XANTENNA__8504__S _3676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5008__A1 _4017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6822_ _1888_ _1890_ vssd1 vssd1 vccd1 vccd1 _1892_ sky130_fd_sc_hd__or2b_1
XFILLER_50_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6753_ _1806_ _1810_ _1815_ vssd1 vssd1 vccd1 vccd1 _1816_ sky130_fd_sc_hd__a21oi_1
XANTENNA__4767__B1 _1748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5704_ _3717_ _3864_ _0614_ vssd1 vssd1 vccd1 vccd1 _0682_ sky130_fd_sc_hd__and3_1
X_6684_ _1697_ _1698_ vssd1 vssd1 vccd1 vccd1 _1740_ sky130_fd_sc_hd__or2b_1
XANTENNA__5429__A _1946_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5635_ _0112_ _0607_ vssd1 vssd1 vccd1 vccd1 _0608_ sky130_fd_sc_hd__nor2_1
X_8423_ mode vssd1 vssd1 vccd1 vccd1 _3636_ sky130_fd_sc_hd__clkinv_2
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5566_ _4115_ _4145_ vssd1 vssd1 vccd1 vccd1 _0539_ sky130_fd_sc_hd__xor2_1
X_8354_ _3563_ _3564_ vssd1 vssd1 vccd1 vccd1 _3565_ sky130_fd_sc_hd__or2_1
XFILLER_117_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4517_ _3339_ _3349_ _2903_ _3360_ vssd1 vssd1 vccd1 vccd1 _3467_ sky130_fd_sc_hd__o211a_1
X_7305_ _2416_ _2422_ vssd1 vssd1 vccd1 vccd1 _2423_ sky130_fd_sc_hd__and2b_1
X_8285_ _3489_ _3491_ _0599_ vssd1 vssd1 vccd1 vccd1 _3492_ sky130_fd_sc_hd__o21bai_1
X_5497_ _0469_ vssd1 vssd1 vccd1 vccd1 _0470_ sky130_fd_sc_hd__clkbuf_4
XFILLER_104_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5164__A _3881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4448_ _1242_ _2573_ vssd1 vssd1 vccd1 vccd1 _2716_ sky130_fd_sc_hd__nand2_2
X_7236_ _0603_ _2343_ _2346_ _2344_ vssd1 vssd1 vccd1 vccd1 _2347_ sky130_fd_sc_hd__a211o_4
XFILLER_98_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4379_ _1429_ _1946_ vssd1 vssd1 vccd1 vccd1 _1957_ sky130_fd_sc_hd__xnor2_1
X_7167_ _2270_ _1628_ _1623_ _1629_ vssd1 vssd1 vccd1 vccd1 _2271_ sky130_fd_sc_hd__a22o_1
X_6118_ _1095_ _1097_ vssd1 vssd1 vccd1 vccd1 _1121_ sky130_fd_sc_hd__or2b_1
X_7098_ _2192_ _2193_ _2194_ vssd1 vssd1 vccd1 vccd1 _2195_ sky130_fd_sc_hd__a21oi_1
XFILLER_86_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6049_ _1000_ _1046_ vssd1 vssd1 vccd1 vccd1 _1048_ sky130_fd_sc_hd__and2_1
XFILLER_86_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6723__A _1353_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6442__B _1428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5058__B _3615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4897__B _3832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5074__A _4228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6633__A _1383_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5420_ _0369_ _0374_ vssd1 vssd1 vccd1 vccd1 _0393_ sky130_fd_sc_hd__nor2_1
XFILLER_114_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5351_ _0301_ _0323_ _0299_ vssd1 vssd1 vccd1 vccd1 _0324_ sky130_fd_sc_hd__o21ai_1
XFILLER_114_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4302_ in_reg\[12\] in_reg\[13\] _0819_ vssd1 vssd1 vccd1 vccd1 _1114_ sky130_fd_sc_hd__mux2_1
X_5282_ _4187_ _0253_ _0254_ vssd1 vssd1 vccd1 vccd1 _0255_ sky130_fd_sc_hd__a21o_1
X_8070_ _0521_ _3261_ vssd1 vssd1 vccd1 vccd1 _3262_ sky130_fd_sc_hd__or2_1
X_7021_ _2068_ _2074_ vssd1 vssd1 vccd1 vccd1 _2110_ sky130_fd_sc_hd__xnor2_1
XFILLER_99_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6527__B _1510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8415__B2 _1330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8415__A1 _1253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7923_ _3031_ vssd1 vssd1 vccd1 vccd1 _3103_ sky130_fd_sc_hd__inv_2
XFILLER_24_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7854_ _2996_ _3015_ _3026_ vssd1 vssd1 vccd1 vccd1 _3027_ sky130_fd_sc_hd__a21o_1
X_6805_ _1422_ _1456_ vssd1 vssd1 vccd1 vccd1 _1873_ sky130_fd_sc_hd__or2_1
X_7785_ _2861_ _2948_ _2950_ _2934_ vssd1 vssd1 vccd1 vccd1 _2951_ sky130_fd_sc_hd__a31oi_2
X_6736_ _1793_ _1795_ vssd1 vssd1 vccd1 vccd1 _1797_ sky130_fd_sc_hd__nand2_1
XFILLER_51_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4997_ _4042_ _4151_ vssd1 vssd1 vccd1 vccd1 _4152_ sky130_fd_sc_hd__xor2_1
XFILLER_23_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4998__A _3838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6667_ _1710_ _1719_ _1720_ vssd1 vssd1 vccd1 vccd1 _1721_ sky130_fd_sc_hd__a21o_1
XANTENNA__7374__A _2412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6598_ _1592_ _1608_ vssd1 vssd1 vccd1 vccd1 _1645_ sky130_fd_sc_hd__nand2_1
X_5618_ _0566_ _0581_ _0590_ vssd1 vssd1 vccd1 vccd1 _0591_ sky130_fd_sc_hd__a21oi_1
X_8406_ out_reg\[13\] _3242_ vssd1 vssd1 vccd1 vccd1 _3620_ sky130_fd_sc_hd__nand2_1
XFILLER_117_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8337_ _1308_ _3545_ _3544_ vssd1 vssd1 vccd1 vccd1 _3547_ sky130_fd_sc_hd__a21o_1
XFILLER_3_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5549_ _0502_ _0445_ _0510_ vssd1 vssd1 vccd1 vccd1 _0522_ sky130_fd_sc_hd__mux2_1
XFILLER_117_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_534 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8268_ _1220_ _3473_ vssd1 vssd1 vccd1 vccd1 _0028_ sky130_fd_sc_hd__nor2_1
XFILLER_48_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8199_ _0601_ _3399_ vssd1 vssd1 vccd1 vccd1 _3400_ sky130_fd_sc_hd__nand2_1
X_7219_ _2302_ vssd1 vssd1 vccd1 vccd1 _2328_ sky130_fd_sc_hd__inv_2
XFILLER_59_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4701__A _3832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6628__A _1353_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_562 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4920_ _3772_ _3771_ _3882_ _3702_ _3792_ vssd1 vssd1 vccd1 vccd1 _4075_ sky130_fd_sc_hd__o32a_1
XFILLER_18_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4851_ _3829_ _3839_ _4004_ vssd1 vssd1 vccd1 vccd1 _4006_ sky130_fd_sc_hd__o21ai_1
XANTENNA__7893__S _2954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4782_ _3914_ _3936_ vssd1 vssd1 vccd1 vccd1 _3937_ sky130_fd_sc_hd__xnor2_2
X_7570_ _0218_ _4222_ _2713_ vssd1 vssd1 vccd1 vccd1 _2714_ sky130_fd_sc_hd__mux2_1
XFILLER_20_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6521_ _0105_ _1455_ _0184_ vssd1 vssd1 vccd1 vccd1 _1560_ sky130_fd_sc_hd__or3_1
XANTENNA__5707__A _3762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6452_ _1469_ _1416_ _1483_ vssd1 vssd1 vccd1 vccd1 _1485_ sky130_fd_sc_hd__o21a_1
XFILLER_9_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7687__A2 _0082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5403_ _3741_ _3743_ _3156_ vssd1 vssd1 vccd1 vccd1 _0376_ sky130_fd_sc_hd__a21oi_2
XANTENNA__5426__B _1781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6383_ _1406_ _1327_ _1405_ vssd1 vssd1 vccd1 vccd1 _1409_ sky130_fd_sc_hd__or3_4
X_8122_ _3314_ _3317_ _0635_ vssd1 vssd1 vccd1 vccd1 _0023_ sky130_fd_sc_hd__a21oi_1
XFILLER_102_504 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5334_ _0287_ _0305_ _4197_ _0306_ vssd1 vssd1 vccd1 vccd1 _0307_ sky130_fd_sc_hd__o31a_1
XFILLER_102_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5265_ _0235_ _0237_ vssd1 vssd1 vccd1 vccd1 _0238_ sky130_fd_sc_hd__nand2_1
X_8053_ _3213_ _3224_ _3241_ _3244_ vssd1 vssd1 vccd1 vccd1 _3245_ sky130_fd_sc_hd__o31a_1
X_7004_ _1509_ _4126_ vssd1 vssd1 vccd1 vccd1 _2092_ sky130_fd_sc_hd__or2_1
XFILLER_87_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5196_ _0124_ _0137_ _0168_ _3875_ vssd1 vssd1 vccd1 vccd1 _0169_ sky130_fd_sc_hd__or4_2
XFILLER_68_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6273__A _0762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7906_ _3083_ vssd1 vssd1 vccd1 vccd1 _3084_ sky130_fd_sc_hd__inv_2
X_7837_ _2979_ _3007_ vssd1 vssd1 vccd1 vccd1 _3008_ sky130_fd_sc_hd__nor2_1
XFILLER_51_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7768_ _2930_ _2931_ vssd1 vssd1 vccd1 vccd1 _2932_ sky130_fd_sc_hd__nand2_1
XFILLER_24_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6720__B _1676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6719_ _1775_ _1777_ vssd1 vssd1 vccd1 vccd1 _1778_ sky130_fd_sc_hd__or2b_1
XFILLER_50_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7699_ _2675_ _2737_ _2855_ _2743_ vssd1 vssd1 vccd1 vccd1 _2856_ sky130_fd_sc_hd__a22o_1
XFILLER_109_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_20 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7366__A1 _2382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8315__B1 _3523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5050_ _4203_ _4204_ vssd1 vssd1 vccd1 vccd1 _4205_ sky130_fd_sc_hd__nor2_1
XANTENNA__7180__C _0121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4655__A2 _2452_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7888__S _2999_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6805__B _1456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5952_ _3770_ _0802_ vssd1 vssd1 vccd1 vccd1 _0947_ sky130_fd_sc_hd__nor2_1
XFILLER_92_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4903_ _3971_ _3973_ vssd1 vssd1 vccd1 vccd1 _4058_ sky130_fd_sc_hd__xnor2_1
XFILLER_52_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_392 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5883_ _0870_ _0871_ _0872_ _0873_ vssd1 vssd1 vccd1 vccd1 _0874_ sky130_fd_sc_hd__a31o_1
XFILLER_21_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8512__S _3676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4834_ posit_add.in1\[14\] _3013_ _2584_ vssd1 vssd1 vccd1 vccd1 _3989_ sky130_fd_sc_hd__nor3_4
X_7622_ _2768_ _2769_ vssd1 vssd1 vccd1 vccd1 _2772_ sky130_fd_sc_hd__nand2_1
X_4765_ _1583_ _3919_ _2452_ vssd1 vssd1 vccd1 vccd1 _3920_ sky130_fd_sc_hd__mux2_1
XFILLER_21_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7553_ _2677_ _2687_ _2688_ _2695_ _0415_ vssd1 vssd1 vccd1 vccd1 _2696_ sky130_fd_sc_hd__a32o_1
XFILLER_119_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4341__A posit_add.in2\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6504_ _1455_ _0184_ vssd1 vssd1 vccd1 vccd1 _1542_ sky130_fd_sc_hd__xor2_2
XANTENNA__4591__A1 _3189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4696_ _3520_ _3850_ vssd1 vssd1 vccd1 vccd1 _3851_ sky130_fd_sc_hd__nor2_1
X_7484_ cmd\[6\] _0092_ cmd\[7\] vssd1 vssd1 vccd1 vccd1 _2620_ sky130_fd_sc_hd__or3b_1
XFILLER_106_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6435_ _1383_ _0303_ vssd1 vssd1 vccd1 vccd1 _1466_ sky130_fd_sc_hd__nor2_1
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6366_ _1389_ vssd1 vssd1 vccd1 vccd1 _1390_ sky130_fd_sc_hd__inv_2
XFILLER_115_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5317_ _0268_ _0289_ vssd1 vssd1 vccd1 vccd1 _0290_ sky130_fd_sc_hd__and2_1
X_8105_ _3148_ _3299_ _3234_ vssd1 vssd1 vccd1 vccd1 _3300_ sky130_fd_sc_hd__mux2_1
XFILLER_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6297_ _1004_ _1313_ vssd1 vssd1 vccd1 vccd1 _1314_ sky130_fd_sc_hd__xnor2_1
XFILLER_102_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8036_ _3225_ _3185_ _2721_ vssd1 vssd1 vccd1 vccd1 _3226_ sky130_fd_sc_hd__mux2_1
X_5248_ _0220_ vssd1 vssd1 vccd1 vccd1 _0221_ sky130_fd_sc_hd__inv_2
XFILLER_29_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5900__A _0762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5179_ _0145_ _0151_ vssd1 vssd1 vccd1 vccd1 _0152_ sky130_fd_sc_hd__xnor2_1
XFILLER_56_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6434__C _1354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_671 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7827__A _2993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7587__A1 _0113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7339__A1 _4089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8000__A2 _0121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4550_ _1726_ _2353_ _2364_ _1682_ vssd1 vssd1 vccd1 vccd1 _3705_ sky130_fd_sc_hd__o211a_1
X_4481_ _2980_ _3068_ vssd1 vssd1 vccd1 vccd1 _3079_ sky130_fd_sc_hd__xnor2_4
XFILLER_7_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6220_ _0762_ _1128_ vssd1 vssd1 vccd1 vccd1 _1229_ sky130_fd_sc_hd__nand2_1
X_6151_ _1137_ _1141_ _1153_ vssd1 vssd1 vccd1 vccd1 _1155_ sky130_fd_sc_hd__and3_1
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5102_ _4234_ _4248_ _4256_ vssd1 vssd1 vccd1 vccd1 _0075_ sky130_fd_sc_hd__o21ai_2
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6082_ _1057_ _1060_ _1066_ vssd1 vssd1 vccd1 vccd1 _1083_ sky130_fd_sc_hd__a21oi_1
XFILLER_85_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5033_ _4185_ _4186_ vssd1 vssd1 vccd1 vccd1 _4188_ sky130_fd_sc_hd__or2_1
XFILLER_57_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8405__B1_N _1177_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6984_ _2069_ vssd1 vssd1 vccd1 vccd1 _2070_ sky130_fd_sc_hd__inv_2
XFILLER_80_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5935_ _0908_ _0906_ _0907_ vssd1 vssd1 vccd1 vccd1 _0929_ sky130_fd_sc_hd__a21o_1
XFILLER_15_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5866_ _2529_ _0773_ _0855_ vssd1 vssd1 vccd1 vccd1 _0856_ sky130_fd_sc_hd__o21ai_1
XANTENNA__6551__A _4228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4817_ _3739_ _3604_ _3794_ _3735_ vssd1 vssd1 vccd1 vccd1 _3972_ sky130_fd_sc_hd__o22a_1
XFILLER_21_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7605_ _2731_ _2732_ vssd1 vssd1 vccd1 vccd1 _2753_ sky130_fd_sc_hd__nand2_1
XANTENNA__6270__B _1128_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5797_ _0721_ _0725_ _0779_ vssd1 vssd1 vccd1 vccd1 _0781_ sky130_fd_sc_hd__nand3_1
X_8585_ clknet_3_4__leaf_clk _0071_ vssd1 vssd1 vccd1 vccd1 posit_add.in2\[12\] sky130_fd_sc_hd__dfxtp_2
XFILLER_21_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4748_ _3897_ _3902_ vssd1 vssd1 vccd1 vccd1 _3903_ sky130_fd_sc_hd__or2_1
X_7536_ _2658_ _2659_ vssd1 vssd1 vccd1 vccd1 _2677_ sky130_fd_sc_hd__xor2_2
X_4679_ _2859_ _3307_ _3371_ _3477_ vssd1 vssd1 vccd1 vccd1 _3834_ sky130_fd_sc_hd__a211o_1
X_7467_ _2522_ _2523_ _2527_ _2486_ vssd1 vssd1 vccd1 vccd1 _2601_ sky130_fd_sc_hd__a211o_1
X_6418_ _1446_ _1384_ vssd1 vssd1 vccd1 vccd1 _1447_ sky130_fd_sc_hd__or2_1
XFILLER_115_470 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7398_ _2437_ _2440_ _2524_ _2335_ vssd1 vssd1 vccd1 vccd1 _2525_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__6069__A1 _3892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6349_ _1357_ _1346_ _1370_ vssd1 vssd1 vccd1 vccd1 _1371_ sky130_fd_sc_hd__o21ai_1
XFILLER_88_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8019_ _2611_ _2588_ _3206_ vssd1 vssd1 vccd1 vccd1 _3207_ sky130_fd_sc_hd__a21boi_2
XFILLER_56_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5077__A _3989_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_674 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5752__B1 _2529_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5720_ _0629_ _0697_ _0688_ _0698_ vssd1 vssd1 vccd1 vccd1 _0699_ sky130_fd_sc_hd__o22a_1
XFILLER_62_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5651_ _4221_ _0611_ _0618_ _0623_ vssd1 vssd1 vccd1 vccd1 _0624_ sky130_fd_sc_hd__a22o_2
XFILLER_31_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4602_ _1682_ _2221_ _3665_ _2298_ vssd1 vssd1 vccd1 vccd1 _3757_ sky130_fd_sc_hd__a211o_1
X_8370_ _3287_ _3502_ _3568_ _3579_ _2604_ vssd1 vssd1 vccd1 vccd1 _3581_ sky130_fd_sc_hd__a311o_1
X_5582_ _0338_ _0542_ _0547_ _0554_ vssd1 vssd1 vccd1 vccd1 _0555_ sky130_fd_sc_hd__a211o_1
X_4533_ _2221_ vssd1 vssd1 vccd1 vccd1 _3635_ sky130_fd_sc_hd__clkbuf_4
X_7321_ _2253_ _2439_ vssd1 vssd1 vccd1 vccd1 _2440_ sky130_fd_sc_hd__xor2_2
XFILLER_7_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_83 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7252_ _2363_ vssd1 vssd1 vccd1 vccd1 _2365_ sky130_fd_sc_hd__clkbuf_2
XFILLER_116_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6203_ _1208_ _1210_ vssd1 vssd1 vccd1 vccd1 _1211_ sky130_fd_sc_hd__xnor2_1
XFILLER_89_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4464_ _1242_ _2551_ vssd1 vssd1 vccd1 vccd1 _2892_ sky130_fd_sc_hd__nand2_1
XFILLER_89_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4395_ _1506_ _1660_ vssd1 vssd1 vccd1 vccd1 _2133_ sky130_fd_sc_hd__xnor2_1
X_7183_ _2271_ _2288_ vssd1 vssd1 vccd1 vccd1 _2289_ sky130_fd_sc_hd__xnor2_1
XFILLER_112_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6134_ _1136_ _1116_ vssd1 vssd1 vccd1 vccd1 _1138_ sky130_fd_sc_hd__xor2_1
XFILLER_112_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6065_ _3892_ _1019_ _1064_ vssd1 vssd1 vccd1 vccd1 _1065_ sky130_fd_sc_hd__and3_1
XFILLER_100_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4765__S _2452_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6546__A _1420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5016_ _3996_ _4008_ vssd1 vssd1 vccd1 vccd1 _4171_ sky130_fd_sc_hd__or2_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4482__B1 _1253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6967_ _0147_ _1813_ vssd1 vssd1 vccd1 vccd1 _2051_ sky130_fd_sc_hd__nand2_1
X_5918_ _3763_ _0787_ vssd1 vssd1 vccd1 vccd1 _0911_ sky130_fd_sc_hd__nor2_1
XFILLER_41_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6898_ _1973_ _1974_ vssd1 vssd1 vccd1 vccd1 _1975_ sky130_fd_sc_hd__nor2_1
X_5849_ _0822_ _0825_ _0824_ vssd1 vssd1 vccd1 vccd1 _0838_ sky130_fd_sc_hd__nand3_1
XFILLER_21_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8568_ clknet_3_7__leaf_clk _0054_ vssd1 vssd1 vccd1 vccd1 posit_add.in1\[11\] sky130_fd_sc_hd__dfxtp_2
XFILLER_108_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7519_ _2653_ _2654_ _2657_ _0399_ vssd1 vssd1 vccd1 vccd1 _2658_ sky130_fd_sc_hd__a31o_2
X_8499_ _3688_ vssd1 vssd1 vccd1 vccd1 _0067_ sky130_fd_sc_hd__clkbuf_1
XFILLER_107_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_390 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6214__B2 _1164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6191__A _0779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7478__A0 _2488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7870_ _2954_ vssd1 vssd1 vccd1 vccd1 _3044_ sky130_fd_sc_hd__buf_2
X_6821_ _1857_ _1859_ _1889_ vssd1 vssd1 vccd1 vccd1 _1890_ sky130_fd_sc_hd__a21bo_1
XFILLER_63_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5413__C1 _0385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4614__A _3736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6752_ _1813_ _0121_ _4228_ _1664_ vssd1 vssd1 vccd1 vccd1 _1815_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__4767__A1 _3736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5703_ _3814_ _3791_ vssd1 vssd1 vccd1 vccd1 _0681_ sky130_fd_sc_hd__nand2_1
X_6683_ _1727_ _1729_ vssd1 vssd1 vccd1 vccd1 _1739_ sky130_fd_sc_hd__nand2_1
XFILLER_50_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5634_ _3759_ _3760_ _3898_ _3899_ vssd1 vssd1 vccd1 vccd1 _0607_ sky130_fd_sc_hd__o2bb2a_2
X_8422_ _3634_ vssd1 vssd1 vccd1 vccd1 _0036_ sky130_fd_sc_hd__clkbuf_1
X_8353_ _3227_ _3538_ _3539_ vssd1 vssd1 vccd1 vccd1 _3564_ sky130_fd_sc_hd__o21ai_1
X_7304_ _2420_ _2421_ _2412_ vssd1 vssd1 vccd1 vccd1 _2422_ sky130_fd_sc_hd__a21oi_1
X_5565_ _0521_ _0528_ _0537_ vssd1 vssd1 vccd1 vccd1 _0538_ sky130_fd_sc_hd__o21ai_1
XANTENNA__5445__A _3830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4516_ _2859_ _3318_ _3371_ _3446_ vssd1 vssd1 vccd1 vccd1 _3456_ sky130_fd_sc_hd__a211o_1
X_8284_ _3465_ _3490_ vssd1 vssd1 vccd1 vccd1 _3491_ sky130_fd_sc_hd__xnor2_2
XFILLER_2_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5496_ _0441_ _0468_ vssd1 vssd1 vccd1 vccd1 _0469_ sky130_fd_sc_hd__or2_2
XANTENNA__5164__B _3776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4447_ _2650_ _2672_ _2694_ vssd1 vssd1 vccd1 vccd1 _2705_ sky130_fd_sc_hd__mux2_1
X_7235_ _0346_ _0350_ vssd1 vssd1 vccd1 vccd1 _2346_ sky130_fd_sc_hd__nor2_2
X_7166_ _1595_ _1597_ _1602_ vssd1 vssd1 vccd1 vccd1 _2270_ sky130_fd_sc_hd__o21a_1
X_6117_ _1118_ _1119_ vssd1 vssd1 vccd1 vccd1 _1120_ sky130_fd_sc_hd__xnor2_1
XFILLER_86_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4378_ posit_add.in2\[6\] _1935_ vssd1 vssd1 vccd1 vccd1 _1946_ sky130_fd_sc_hd__xor2_4
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6276__A _0706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7097_ _2189_ _2191_ vssd1 vssd1 vccd1 vccd1 _2194_ sky130_fd_sc_hd__nor2_1
XFILLER_85_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6048_ _1000_ _1046_ vssd1 vssd1 vccd1 vccd1 _1047_ sky130_fd_sc_hd__nor2_1
XFILLER_46_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6723__B _1354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7999_ _1275_ _4250_ vssd1 vssd1 vccd1 vccd1 _3186_ sky130_fd_sc_hd__nand2_1
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4524__A _2969_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5074__B _3800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6186__A _0722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6633__B _1454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5350_ _0313_ _0322_ _0311_ vssd1 vssd1 vccd1 vccd1 _0323_ sky130_fd_sc_hd__a21oi_1
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4921__A1 _3878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4301_ _1093_ vssd1 vssd1 vccd1 vccd1 _0015_ sky130_fd_sc_hd__clkbuf_1
X_5281_ _0217_ _0221_ vssd1 vssd1 vccd1 vccd1 _0254_ sky130_fd_sc_hd__xnor2_1
XFILLER_114_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7020_ _2088_ _2107_ _2108_ vssd1 vssd1 vccd1 vccd1 _2109_ sky130_fd_sc_hd__a21boi_1
XFILLER_4_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4609__A _3763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8415__A2 _0082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7922_ _3051_ _3099_ _3100_ _3031_ vssd1 vssd1 vccd1 vccd1 _3102_ sky130_fd_sc_hd__o31a_1
XFILLER_70_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7853_ _2993_ _2995_ vssd1 vssd1 vccd1 vccd1 _3026_ sky130_fd_sc_hd__and2_1
X_6804_ _1870_ _1871_ vssd1 vssd1 vccd1 vccd1 _1872_ sky130_fd_sc_hd__nor2_1
XFILLER_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4996_ _4068_ _4149_ _4150_ vssd1 vssd1 vccd1 vccd1 _4151_ sky130_fd_sc_hd__a21oi_1
X_7784_ _2864_ _2949_ vssd1 vssd1 vccd1 vccd1 _2950_ sky130_fd_sc_hd__xnor2_1
X_6735_ _1793_ _1795_ vssd1 vssd1 vccd1 vccd1 _1796_ sky130_fd_sc_hd__nor2_1
XFILLER_23_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6666_ _1706_ _1709_ vssd1 vssd1 vccd1 vccd1 _1720_ sky130_fd_sc_hd__nor2_1
XANTENNA__5175__A _4017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6597_ _1642_ _1643_ vssd1 vssd1 vccd1 vccd1 _1644_ sky130_fd_sc_hd__nand2_1
X_8405_ _0600_ _3618_ _1177_ vssd1 vssd1 vccd1 vccd1 _3619_ sky130_fd_sc_hd__o21ba_1
X_5617_ _0519_ _0580_ _0582_ _0589_ vssd1 vssd1 vccd1 vccd1 _0590_ sky130_fd_sc_hd__o31a_1
XFILLER_105_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8336_ _1319_ _3544_ _3545_ _0599_ vssd1 vssd1 vccd1 vccd1 _3546_ sky130_fd_sc_hd__a31o_1
X_5548_ _0518_ _0467_ vssd1 vssd1 vccd1 vccd1 _0521_ sky130_fd_sc_hd__nor2_4
XFILLER_105_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8267_ out_reg\[8\] _3197_ _3471_ _3472_ vssd1 vssd1 vccd1 vccd1 _3473_ sky130_fd_sc_hd__a22oi_1
XFILLER_3_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5903__A _2529_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5479_ _0446_ _0450_ _0451_ vssd1 vssd1 vccd1 vccd1 _0452_ sky130_fd_sc_hd__o21a_1
X_7218_ _2316_ _2317_ _2326_ vssd1 vssd1 vccd1 vccd1 _2327_ sky130_fd_sc_hd__a21o_1
X_8198_ _3322_ _3355_ _3323_ vssd1 vssd1 vccd1 vccd1 _3399_ sky130_fd_sc_hd__or3b_1
XFILLER_86_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7149_ _2248_ _2249_ _2250_ vssd1 vssd1 vccd1 vccd1 _2251_ sky130_fd_sc_hd__o21a_1
XFILLER_100_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7614__A0 _0147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7090__A1 _4089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7565__A _2319_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4701__B _3855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_496 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6628__B _1354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_3_7__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_7__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_80_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5631__A2 _2507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4850_ _3829_ _3839_ _4004_ vssd1 vssd1 vccd1 vccd1 _4005_ sky130_fd_sc_hd__or3_1
XFILLER_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4781_ _3935_ _3728_ vssd1 vssd1 vccd1 vccd1 _3936_ sky130_fd_sc_hd__xnor2_2
X_6520_ _1549_ _1557_ _1558_ vssd1 vssd1 vccd1 vccd1 _1559_ sky130_fd_sc_hd__o21a_1
XFILLER_9_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6451_ _0218_ _1408_ _1409_ _1414_ _0121_ vssd1 vssd1 vccd1 vccd1 _1483_ sky130_fd_sc_hd__a32o_1
X_6382_ _1327_ _1405_ _1406_ vssd1 vssd1 vccd1 vccd1 _1408_ sky130_fd_sc_hd__o21ai_4
X_5402_ _0370_ _0374_ vssd1 vssd1 vccd1 vccd1 _0375_ sky130_fd_sc_hd__xnor2_4
X_5333_ _4154_ _4198_ vssd1 vssd1 vccd1 vccd1 _0306_ sky130_fd_sc_hd__nand2_1
X_8121_ out_reg\[2\] _3316_ _3197_ out_reg\[3\] vssd1 vssd1 vccd1 vccd1 _3317_ sky130_fd_sc_hd__a22oi_1
XANTENNA__5723__A _2529_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5264_ _0225_ _0236_ vssd1 vssd1 vccd1 vccd1 _0237_ sky130_fd_sc_hd__and2_1
XANTENNA__7844__B1 _2993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8052_ out_reg\[0\] _3242_ _0701_ vssd1 vssd1 vccd1 vccd1 _3244_ sky130_fd_sc_hd__a21bo_1
X_7003_ _2054_ _2057_ _2055_ vssd1 vssd1 vccd1 vccd1 _2091_ sky130_fd_sc_hd__a21o_1
XFILLER_102_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5195_ _3763_ _3840_ _3989_ _3793_ vssd1 vssd1 vccd1 vccd1 _0168_ sky130_fd_sc_hd__o22a_1
XFILLER_68_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_614 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6554__A _4153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6273__B _1164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7905_ _3074_ _3082_ _2998_ vssd1 vssd1 vccd1 vccd1 _3083_ sky130_fd_sc_hd__mux2_1
XFILLER_70_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7836_ _2976_ _2978_ vssd1 vssd1 vccd1 vccd1 _3007_ sky130_fd_sc_hd__and2_1
XFILLER_34_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4979_ _4117_ _4128_ vssd1 vssd1 vccd1 vccd1 _4134_ sky130_fd_sc_hd__nand2_1
X_7767_ _2851_ _2871_ _2869_ _2929_ vssd1 vssd1 vccd1 vccd1 _2931_ sky130_fd_sc_hd__o22ai_1
X_6718_ _1776_ _1725_ vssd1 vssd1 vccd1 vccd1 _1777_ sky130_fd_sc_hd__xnor2_1
X_7698_ _2704_ _2777_ _2854_ vssd1 vssd1 vccd1 vccd1 _2855_ sky130_fd_sc_hd__a21oi_1
XFILLER_109_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5138__B2 _3690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6649_ _1695_ _1700_ vssd1 vssd1 vccd1 vccd1 _1701_ sky130_fd_sc_hd__xnor2_1
XFILLER_118_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8319_ out_reg\[11\] _3197_ vssd1 vssd1 vccd1 vccd1 _3527_ sky130_fd_sc_hd__nand2_1
XFILLER_105_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5310__A1 _4045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6464__A _4250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7295__A _2411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8052__B1_N _0701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5951_ _0773_ _3738_ vssd1 vssd1 vccd1 vccd1 _0945_ sky130_fd_sc_hd__nor2_1
XFILLER_92_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4902_ _3968_ _3975_ vssd1 vssd1 vccd1 vccd1 _4057_ sky130_fd_sc_hd__xnor2_1
XFILLER_33_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5882_ _0867_ _0869_ vssd1 vssd1 vccd1 vccd1 _0873_ sky130_fd_sc_hd__and2_1
X_4833_ _3853_ vssd1 vssd1 vccd1 vccd1 _3988_ sky130_fd_sc_hd__clkbuf_4
X_7621_ _2768_ _2769_ vssd1 vssd1 vccd1 vccd1 _2770_ sky130_fd_sc_hd__or2_1
XANTENNA__5718__A _3762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4764_ posit_add.in2\[9\] _1594_ vssd1 vssd1 vccd1 vccd1 _3919_ sky130_fd_sc_hd__xnor2_1
X_7552_ _2662_ _2689_ _2693_ _0448_ vssd1 vssd1 vccd1 vccd1 _2695_ sky130_fd_sc_hd__a2bb2o_1
X_6503_ _1532_ _0184_ _1534_ _1540_ vssd1 vssd1 vccd1 vccd1 _1541_ sky130_fd_sc_hd__o2bb2a_1
X_7483_ _2521_ _2610_ _2618_ vssd1 vssd1 vccd1 vccd1 _2619_ sky130_fd_sc_hd__and3_1
X_6434_ _0218_ _1353_ _1354_ vssd1 vssd1 vccd1 vccd1 _1465_ sky130_fd_sc_hd__nand3_1
X_4695_ _3446_ _3847_ _3849_ vssd1 vssd1 vccd1 vccd1 _3850_ sky130_fd_sc_hd__a21o_1
XFILLER_115_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6365_ _1097_ _0993_ _1388_ vssd1 vssd1 vccd1 vccd1 _1389_ sky130_fd_sc_hd__a21o_1
XANTENNA__5453__A _3830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6296_ _1033_ _1032_ _1027_ vssd1 vssd1 vccd1 vccd1 _1313_ sky130_fd_sc_hd__a21o_1
X_5316_ _0265_ _0267_ vssd1 vssd1 vccd1 vccd1 _0289_ sky130_fd_sc_hd__nand2_1
X_8104_ _3298_ vssd1 vssd1 vccd1 vccd1 _3299_ sky130_fd_sc_hd__clkinv_2
X_5247_ _0211_ _0219_ vssd1 vssd1 vccd1 vccd1 _0220_ sky130_fd_sc_hd__nand2_1
X_8035_ _1275_ vssd1 vssd1 vccd1 vccd1 _3225_ sky130_fd_sc_hd__inv_2
XFILLER_29_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5178_ _0146_ _0149_ _0150_ vssd1 vssd1 vccd1 vccd1 _0151_ sky130_fd_sc_hd__o21a_1
XFILLER_28_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7819_ _2662_ _2677_ vssd1 vssd1 vccd1 vccd1 _2988_ sky130_fd_sc_hd__xnor2_1
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6087__A2 _3739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5538__A _0440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4480_ posit_add.in1\[12\] _3057_ vssd1 vssd1 vccd1 vccd1 _3068_ sky130_fd_sc_hd__xnor2_4
XFILLER_7_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6150_ _1137_ _1141_ _1153_ vssd1 vssd1 vccd1 vccd1 _1154_ sky130_fd_sc_hd__a21oi_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5101_ _4254_ _4255_ vssd1 vssd1 vccd1 vccd1 _4256_ sky130_fd_sc_hd__and2_1
X_6081_ _1073_ _1067_ _1071_ vssd1 vssd1 vccd1 vccd1 _1082_ sky130_fd_sc_hd__and3b_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5032_ _4185_ _4186_ vssd1 vssd1 vccd1 vccd1 _4187_ sky130_fd_sc_hd__nand2_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6983_ _2064_ _2066_ _2068_ vssd1 vssd1 vccd1 vccd1 _2069_ sky130_fd_sc_hd__a21oi_1
X_5934_ _0908_ _0906_ _0907_ vssd1 vssd1 vccd1 vccd1 _0928_ sky130_fd_sc_hd__nand3_1
XFILLER_15_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5865_ _3735_ _0700_ vssd1 vssd1 vccd1 vccd1 _0855_ sky130_fd_sc_hd__or2_1
XFILLER_80_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6551__B _1383_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4816_ _3816_ _3726_ vssd1 vssd1 vccd1 vccd1 _3971_ sky130_fd_sc_hd__nor2_1
X_7604_ _3881_ _1355_ _2721_ vssd1 vssd1 vccd1 vccd1 _2752_ sky130_fd_sc_hd__mux2_1
XANTENNA__5448__A _1781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5796_ _0721_ _0725_ _0779_ vssd1 vssd1 vccd1 vccd1 _0780_ sky130_fd_sc_hd__a21o_1
X_8584_ clknet_3_7__leaf_clk _0070_ vssd1 vssd1 vccd1 vccd1 posit_add.in2\[11\] sky130_fd_sc_hd__dfxtp_2
XFILLER_119_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4747_ _3901_ _3868_ vssd1 vssd1 vccd1 vccd1 _3902_ sky130_fd_sc_hd__nand2_1
XFILLER_31_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7535_ _0442_ _2670_ vssd1 vssd1 vccd1 vccd1 _2676_ sky130_fd_sc_hd__xnor2_2
XFILLER_119_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4678_ _2694_ _3307_ _3820_ _3435_ vssd1 vssd1 vccd1 vccd1 _3833_ sky130_fd_sc_hd__a211o_1
XANTENNA__7502__A2 _1682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7466_ _2522_ _2581_ _2582_ _2514_ vssd1 vssd1 vccd1 vccd1 _2600_ sky130_fd_sc_hd__a211o_1
XFILLER_107_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6417_ _1445_ vssd1 vssd1 vccd1 vccd1 _1446_ sky130_fd_sc_hd__buf_2
X_7397_ _2085_ _2247_ vssd1 vssd1 vccd1 vccd1 _2524_ sky130_fd_sc_hd__xor2_2
X_6348_ _1368_ _1369_ vssd1 vssd1 vccd1 vccd1 _1370_ sky130_fd_sc_hd__and2_1
XFILLER_1_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6279_ _1271_ _1270_ vssd1 vssd1 vccd1 vccd1 _1294_ sky130_fd_sc_hd__and2b_1
XFILLER_76_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4619__A3 _2452_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8018_ _2514_ _3203_ _3205_ _2611_ vssd1 vssd1 vccd1 vccd1 _3206_ sky130_fd_sc_hd__a211o_1
XFILLER_29_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5650_ _0620_ _0621_ _0622_ _3923_ vssd1 vssd1 vccd1 vccd1 _0623_ sky130_fd_sc_hd__o31a_1
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_31_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4601_ _3735_ _3739_ _3750_ _3755_ vssd1 vssd1 vccd1 vccd1 _3756_ sky130_fd_sc_hd__nor4_2
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5581_ _4131_ _0549_ _0553_ vssd1 vssd1 vccd1 vccd1 _0554_ sky130_fd_sc_hd__a21o_1
XFILLER_30_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4532_ _2485_ _2320_ _2419_ vssd1 vssd1 vccd1 vccd1 _3625_ sky130_fd_sc_hd__and3_1
X_7320_ _2085_ _2247_ _2083_ vssd1 vssd1 vccd1 vccd1 _2439_ sky130_fd_sc_hd__a21oi_1
XFILLER_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4463_ _2837_ _2870_ vssd1 vssd1 vccd1 vccd1 _2881_ sky130_fd_sc_hd__nand2_1
X_7251_ _2361_ _2362_ vssd1 vssd1 vccd1 vccd1 _2363_ sky130_fd_sc_hd__or2_1
X_6202_ _1179_ _1209_ vssd1 vssd1 vccd1 vccd1 _1210_ sky130_fd_sc_hd__nor2_1
XFILLER_89_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4394_ _1495_ _1517_ _1550_ vssd1 vssd1 vccd1 vccd1 _2122_ sky130_fd_sc_hd__a21o_1
X_7182_ _1642_ _2286_ vssd1 vssd1 vccd1 vccd1 _2288_ sky130_fd_sc_hd__xnor2_1
XFILLER_112_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6133_ _1116_ _1136_ vssd1 vssd1 vccd1 vccd1 _1137_ sky130_fd_sc_hd__or2b_1
XFILLER_98_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6064_ _0952_ _1063_ vssd1 vssd1 vccd1 vccd1 _1064_ sky130_fd_sc_hd__and2_1
XFILLER_97_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5015_ _4168_ _4169_ vssd1 vssd1 vccd1 vccd1 _4170_ sky130_fd_sc_hd__xnor2_1
XFILLER_73_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6546__B _1446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4482__A1 posit_add.in1\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6966_ _3817_ _1663_ _2014_ vssd1 vssd1 vccd1 vccd1 _2050_ sky130_fd_sc_hd__o21ba_1
XFILLER_53_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5917_ _0896_ _0898_ vssd1 vssd1 vccd1 vccd1 _0910_ sky130_fd_sc_hd__nand2_1
X_6897_ _1972_ _1966_ vssd1 vssd1 vccd1 vccd1 _1974_ sky130_fd_sc_hd__and2b_1
XFILLER_42_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5848_ _0834_ _0836_ vssd1 vssd1 vccd1 vccd1 _0837_ sky130_fd_sc_hd__xnor2_1
X_5779_ _0624_ vssd1 vssd1 vccd1 vccd1 _0762_ sky130_fd_sc_hd__clkbuf_4
X_8567_ clknet_3_4__leaf_clk _0053_ vssd1 vssd1 vccd1 vccd1 posit_add.in1\[10\] sky130_fd_sc_hd__dfxtp_2
XFILLER_21_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7518_ _2656_ _0427_ _2651_ vssd1 vssd1 vccd1 vccd1 _2657_ sky130_fd_sc_hd__mux2_1
XFILLER_107_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8498_ posit_add.in2\[8\] in_reg\[8\] _3677_ vssd1 vssd1 vccd1 vccd1 _3688_ sky130_fd_sc_hd__mux2_1
X_7449_ _2454_ _2465_ _2580_ vssd1 vssd1 vccd1 vccd1 _2581_ sky130_fd_sc_hd__o21a_1
XFILLER_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8022__A_N cmd\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4257__A net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7568__A _2702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5088__A _3800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5725__A1 _4222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7650__A1 _4126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6820_ _1843_ _1860_ vssd1 vssd1 vccd1 vccd1 _1889_ sky130_fd_sc_hd__or2b_1
XFILLER_35_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6751_ _1812_ vssd1 vssd1 vccd1 vccd1 _1813_ sky130_fd_sc_hd__clkbuf_2
XFILLER_90_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5702_ _0613_ _0648_ _0678_ vssd1 vssd1 vccd1 vccd1 _0680_ sky130_fd_sc_hd__a21oi_1
X_6682_ _1735_ _1736_ vssd1 vssd1 vccd1 vccd1 _1738_ sky130_fd_sc_hd__xor2_1
X_5633_ _3699_ _3814_ _0112_ vssd1 vssd1 vccd1 vccd1 _0606_ sky130_fd_sc_hd__a21o_1
X_8421_ out_reg\[15\] io_out[3] _0819_ vssd1 vssd1 vccd1 vccd1 _3634_ sky130_fd_sc_hd__mux2_1
X_8352_ _3560_ _3561_ vssd1 vssd1 vccd1 vccd1 _3563_ sky130_fd_sc_hd__nor2_1
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5564_ _0519_ _0536_ vssd1 vssd1 vccd1 vccd1 _0537_ sky130_fd_sc_hd__or2_1
X_7303_ _1896_ _2418_ vssd1 vssd1 vccd1 vccd1 _2421_ sky130_fd_sc_hd__nand2_1
X_4515_ _3435_ vssd1 vssd1 vccd1 vccd1 _3446_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__5445__B _3635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8283_ _0521_ _3217_ _3429_ vssd1 vssd1 vccd1 vccd1 _3490_ sky130_fd_sc_hd__a21oi_1
X_5495_ _0456_ _0460_ _0467_ vssd1 vssd1 vccd1 vccd1 _0468_ sky130_fd_sc_hd__o21bai_2
XFILLER_104_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5164__C _3838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4446_ posit_add.in1\[7\] _2683_ vssd1 vssd1 vccd1 vccd1 _2694_ sky130_fd_sc_hd__xor2_2
X_7234_ _0603_ _2343_ _2344_ vssd1 vssd1 vccd1 vccd1 _2345_ sky130_fd_sc_hd__a21oi_1
X_4377_ posit_add.in2\[5\] posit_add.in2\[4\] _1352_ _1264_ vssd1 vssd1 vccd1 vccd1
+ _1935_ sky130_fd_sc_hd__o31a_1
X_7165_ _1648_ _1650_ vssd1 vssd1 vccd1 vccd1 _2269_ sky130_fd_sc_hd__nor2_1
XANTENNA__7660__B _2800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6116_ _1098_ _1100_ _4017_ _0702_ vssd1 vssd1 vccd1 vccd1 _1119_ sky130_fd_sc_hd__a211o_1
XFILLER_98_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6276__B _1128_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7096_ _1703_ _2171_ vssd1 vssd1 vccd1 vccd1 _2193_ sky130_fd_sc_hd__xnor2_1
XFILLER_86_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5180__B _3838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6047_ _1042_ _1045_ vssd1 vssd1 vccd1 vccd1 _1046_ sky130_fd_sc_hd__xor2_1
XFILLER_85_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4805__A _3793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6723__C _1782_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7998_ _1253_ vssd1 vssd1 vccd1 vccd1 _3185_ sky130_fd_sc_hd__inv_2
XFILLER_26_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6949_ _1384_ _1538_ vssd1 vssd1 vccd1 vccd1 _2031_ sky130_fd_sc_hd__nor2_1
XFILLER_26_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4897__D _3868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4300_ in_reg\[11\] in_reg\[12\] _0819_ vssd1 vssd1 vccd1 vccd1 _1093_ sky130_fd_sc_hd__mux2_1
X_5280_ _4181_ _4189_ vssd1 vssd1 vccd1 vccd1 _0253_ sky130_fd_sc_hd__or2_1
XFILLER_5_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6377__A _1400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4609__B _3702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4437__A1 posit_add.in1\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7921_ _3050_ _3058_ _2999_ vssd1 vssd1 vccd1 vccd1 _3100_ sky130_fd_sc_hd__mux2_1
XFILLER_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7852_ _3020_ vssd1 vssd1 vccd1 vccd1 _3025_ sky130_fd_sc_hd__clkinv_2
XFILLER_23_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6803_ _1868_ _1864_ vssd1 vssd1 vccd1 vccd1 _1871_ sky130_fd_sc_hd__and2b_1
XFILLER_51_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4995_ _4047_ _4067_ vssd1 vssd1 vccd1 vccd1 _4150_ sky130_fd_sc_hd__and2b_1
X_7783_ _1308_ _2861_ vssd1 vssd1 vccd1 vccd1 _2949_ sky130_fd_sc_hd__nand2_1
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6734_ _1794_ _1679_ vssd1 vssd1 vccd1 vccd1 _1795_ sky130_fd_sc_hd__xnor2_1
XFILLER_11_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6665_ _0082_ _1718_ vssd1 vssd1 vccd1 vccd1 _1719_ sky130_fd_sc_hd__nor2_1
X_8404_ _3616_ _3617_ vssd1 vssd1 vccd1 vccd1 _3618_ sky130_fd_sc_hd__xnor2_1
X_6596_ _1630_ _1641_ vssd1 vssd1 vccd1 vccd1 _1643_ sky130_fd_sc_hd__or2_1
X_5616_ _0583_ _0584_ _0585_ _0588_ vssd1 vssd1 vccd1 vccd1 _0589_ sky130_fd_sc_hd__or4_1
XANTENNA__5175__B _3795_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8335_ _3462_ _3468_ _3491_ _3519_ vssd1 vssd1 vccd1 vccd1 _3545_ sky130_fd_sc_hd__or4_1
X_5547_ _0496_ _0517_ _0519_ vssd1 vssd1 vccd1 vccd1 _0520_ sky130_fd_sc_hd__mux2_1
XFILLER_117_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8266_ out_reg\[7\] _3242_ _1177_ vssd1 vssd1 vccd1 vccd1 _3472_ sky130_fd_sc_hd__a21bo_1
X_5478_ _0440_ vssd1 vssd1 vccd1 vccd1 _0451_ sky130_fd_sc_hd__clkinv_2
XFILLER_2_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4429_ _1990_ _2320_ _2419_ _2496_ vssd1 vssd1 vccd1 vccd1 _2507_ sky130_fd_sc_hd__a31o_4
X_7217_ _2312_ _2325_ vssd1 vssd1 vccd1 vccd1 _2326_ sky130_fd_sc_hd__xnor2_1
X_8197_ _3396_ _3397_ vssd1 vssd1 vccd1 vccd1 _3398_ sky130_fd_sc_hd__nand2_1
XFILLER_101_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7148_ _1951_ _1997_ vssd1 vssd1 vccd1 vccd1 _2250_ sky130_fd_sc_hd__xor2_1
XFILLER_100_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7079_ _2172_ _2170_ _2173_ vssd1 vssd1 vccd1 vccd1 _2174_ sky130_fd_sc_hd__nand3_1
XFILLER_59_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7614__A1 _4045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8007__A _1177_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6628__C _4089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7520__S _2652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4780_ _3933_ _3934_ vssd1 vssd1 vccd1 vccd1 _3935_ sky130_fd_sc_hd__or2_1
XFILLER_60_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7756__A _1308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4611__C _2452_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6450_ _1423_ vssd1 vssd1 vccd1 vccd1 _1482_ sky130_fd_sc_hd__inv_2
XFILLER_9_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6381_ _1323_ vssd1 vssd1 vccd1 vccd1 _1406_ sky130_fd_sc_hd__inv_2
XANTENNA__4355__B1 _1682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5401_ _3882_ _0373_ _3721_ vssd1 vssd1 vccd1 vccd1 _0374_ sky130_fd_sc_hd__mux2_4
X_5332_ _4191_ _4192_ _4170_ vssd1 vssd1 vccd1 vccd1 _0305_ sky130_fd_sc_hd__o21a_1
X_8120_ _3315_ vssd1 vssd1 vccd1 vccd1 _3316_ sky130_fd_sc_hd__clkbuf_2
XANTENNA__5723__B _0702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5263_ _0224_ _0211_ _0222_ vssd1 vssd1 vccd1 vccd1 _0236_ sky130_fd_sc_hd__nand3_1
X_8051_ _0786_ vssd1 vssd1 vccd1 vccd1 _3242_ sky130_fd_sc_hd__buf_2
X_7002_ _2059_ _2048_ vssd1 vssd1 vccd1 vccd1 _2090_ sky130_fd_sc_hd__xor2_1
X_5194_ _0165_ _0166_ vssd1 vssd1 vccd1 vccd1 _0167_ sky130_fd_sc_hd__or2_1
XFILLER_68_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6835__A _1454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4830__A1 _2540_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7904_ _3075_ _3081_ _2842_ vssd1 vssd1 vccd1 vccd1 _3082_ sky130_fd_sc_hd__mux2_1
XFILLER_51_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7835_ _3003_ _3005_ vssd1 vssd1 vccd1 vccd1 _3006_ sky130_fd_sc_hd__nand2_2
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5386__A2 _3635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4978_ _4100_ _4110_ vssd1 vssd1 vccd1 vccd1 _4133_ sky130_fd_sc_hd__xnor2_1
X_7766_ _2929_ _2851_ _2871_ _2869_ vssd1 vssd1 vccd1 vccd1 _2930_ sky130_fd_sc_hd__or4_1
XFILLER_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6717_ _0303_ _1537_ vssd1 vssd1 vccd1 vccd1 _1776_ sky130_fd_sc_hd__or2_1
XFILLER_50_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7697_ _2704_ _2853_ vssd1 vssd1 vccd1 vccd1 _2854_ sky130_fd_sc_hd__nor2_1
X_6648_ _1696_ _1699_ vssd1 vssd1 vccd1 vccd1 _1700_ sky130_fd_sc_hd__xor2_2
XFILLER_105_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8318_ _1220_ _3526_ vssd1 vssd1 vccd1 vccd1 _0030_ sky130_fd_sc_hd__nor2_1
X_6579_ _1420_ _1446_ vssd1 vssd1 vccd1 vccd1 _1624_ sky130_fd_sc_hd__or2_1
XFILLER_3_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8088__A1 _3256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6099__B1 _4016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8249_ _3448_ _3452_ vssd1 vssd1 vccd1 vccd1 _3453_ sky130_fd_sc_hd__xor2_1
XFILLER_105_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5310__A2 _0121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6464__B _1428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5096__A _4250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6655__A _0080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5950_ _0940_ _0939_ _0927_ vssd1 vssd1 vccd1 vccd1 _0944_ sky130_fd_sc_hd__a21o_1
XFILLER_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4901_ _4053_ _4054_ _4055_ vssd1 vssd1 vccd1 vccd1 _4056_ sky130_fd_sc_hd__a21bo_1
XFILLER_46_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5881_ _0856_ _0857_ _0854_ vssd1 vssd1 vccd1 vccd1 _0872_ sky130_fd_sc_hd__a21o_1
XFILLER_61_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7620_ _4045_ _0147_ _2721_ vssd1 vssd1 vccd1 vccd1 _2769_ sky130_fd_sc_hd__mux2_1
X_4832_ _3901_ _3986_ vssd1 vssd1 vccd1 vccd1 _3987_ sky130_fd_sc_hd__nand2_1
XANTENNA__6390__A _0218_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_526 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4763_ _3643_ _3635_ _3705_ vssd1 vssd1 vccd1 vccd1 _3918_ sky130_fd_sc_hd__a21oi_1
XFILLER_60_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7551_ _0433_ _2690_ _2692_ _2665_ vssd1 vssd1 vccd1 vccd1 _2693_ sky130_fd_sc_hd__a22o_1
X_6502_ _0082_ _1538_ vssd1 vssd1 vccd1 vccd1 _1540_ sky130_fd_sc_hd__or2_1
X_4694_ _3819_ _3530_ _3848_ _3477_ vssd1 vssd1 vccd1 vccd1 _3849_ sky130_fd_sc_hd__o211a_1
X_7482_ _2611_ _2615_ _2616_ vssd1 vssd1 vccd1 vccd1 _2618_ sky130_fd_sc_hd__o21a_1
XFILLER_107_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6433_ _1420_ _1399_ vssd1 vssd1 vccd1 vccd1 _1464_ sky130_fd_sc_hd__or2_1
XANTENNA__5734__A _4045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6364_ _0627_ _0994_ vssd1 vssd1 vccd1 vccd1 _1388_ sky130_fd_sc_hd__and2_1
XFILLER_114_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6295_ _1037_ _1311_ vssd1 vssd1 vccd1 vccd1 _1312_ sky130_fd_sc_hd__nor2_1
XFILLER_88_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5315_ _4191_ _0287_ vssd1 vssd1 vccd1 vccd1 _0288_ sky130_fd_sc_hd__nor2_1
X_8103_ _3025_ _3177_ _3028_ vssd1 vssd1 vccd1 vccd1 _3298_ sky130_fd_sc_hd__a21o_1
XFILLER_115_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5246_ _0218_ _3901_ _3844_ _0210_ vssd1 vssd1 vccd1 vccd1 _0219_ sky130_fd_sc_hd__a31o_1
X_8034_ _0600_ _3222_ _3223_ vssd1 vssd1 vccd1 vccd1 _3224_ sky130_fd_sc_hd__nor3_2
XFILLER_29_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5177_ _3925_ _0105_ _3795_ vssd1 vssd1 vccd1 vccd1 _0150_ sky130_fd_sc_hd__or3_1
XFILLER_68_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7818_ _2939_ _2985_ _2986_ vssd1 vssd1 vccd1 vccd1 _2987_ sky130_fd_sc_hd__o21ai_1
XFILLER_61_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7749_ _2773_ _2910_ vssd1 vssd1 vccd1 vccd1 _2911_ sky130_fd_sc_hd__xor2_2
XFILLER_117_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_695 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5755__C1 _4222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6080_ _0942_ _1080_ _1056_ _1074_ vssd1 vssd1 vccd1 vccd1 _1081_ sky130_fd_sc_hd__a211o_1
XFILLER_111_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5100_ _4249_ _4253_ vssd1 vssd1 vccd1 vccd1 _4255_ sky130_fd_sc_hd__or2_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5031_ _3987_ _3991_ vssd1 vssd1 vccd1 vccd1 _4186_ sky130_fd_sc_hd__nor2_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6385__A _4228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6982_ _2064_ _2036_ vssd1 vssd1 vccd1 vccd1 _2068_ sky130_fd_sc_hd__and2b_1
XFILLER_65_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5933_ _0923_ _0924_ _0926_ vssd1 vssd1 vccd1 vccd1 _0927_ sky130_fd_sc_hd__and3_1
XFILLER_53_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5864_ _3815_ _0676_ vssd1 vssd1 vccd1 vccd1 _0854_ sky130_fd_sc_hd__nor2_1
XFILLER_80_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8583_ clknet_3_5__leaf_clk _0069_ vssd1 vssd1 vccd1 vccd1 posit_add.in2\[10\] sky130_fd_sc_hd__dfxtp_2
X_4815_ _3945_ _3969_ vssd1 vssd1 vccd1 vccd1 _3970_ sky130_fd_sc_hd__xnor2_1
XFILLER_21_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7603_ _2743_ _2750_ vssd1 vssd1 vccd1 vccd1 _2751_ sky130_fd_sc_hd__and2_1
X_5795_ _4016_ _0755_ vssd1 vssd1 vccd1 vccd1 _0779_ sky130_fd_sc_hd__or2_2
X_7534_ _2346_ _2674_ vssd1 vssd1 vccd1 vccd1 _2675_ sky130_fd_sc_hd__xnor2_2
X_4746_ _3900_ vssd1 vssd1 vccd1 vccd1 _3901_ sky130_fd_sc_hd__buf_4
XFILLER_31_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4677_ _3831_ vssd1 vssd1 vccd1 vccd1 _3832_ sky130_fd_sc_hd__clkbuf_4
X_7465_ _2585_ _2588_ _2592_ _2598_ vssd1 vssd1 vccd1 vccd1 _2599_ sky130_fd_sc_hd__nand4_1
XFILLER_119_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6416_ _1443_ _1444_ vssd1 vssd1 vccd1 vccd1 _1445_ sky130_fd_sc_hd__nor2_1
X_7396_ _2446_ _2424_ _2410_ vssd1 vssd1 vccd1 vccd1 _2523_ sky130_fd_sc_hd__mux2_1
X_6347_ _1000_ _1367_ vssd1 vssd1 vccd1 vccd1 _1369_ sky130_fd_sc_hd__nand2_1
XFILLER_115_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8463__A1 posit_add.in1\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6278_ _1288_ _1289_ _1292_ vssd1 vssd1 vccd1 vccd1 _1293_ sky130_fd_sc_hd__o21ai_1
XFILLER_88_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4808__A _3800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5229_ _0199_ _0201_ vssd1 vssd1 vccd1 vccd1 _0202_ sky130_fd_sc_hd__and2b_1
X_8017_ _2494_ _2613_ _3204_ _2486_ vssd1 vssd1 vccd1 vccd1 _3205_ sky130_fd_sc_hd__o211a_1
XFILLER_56_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_423 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5029__A1 _3816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5752__A2 _3901_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5374__A _1781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4600_ _3722_ _3754_ vssd1 vssd1 vccd1 vccd1 _3755_ sky130_fd_sc_hd__nand2_2
XFILLER_31_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7193__A1 _0082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5580_ _4129_ _0550_ _0552_ vssd1 vssd1 vccd1 vccd1 _0553_ sky130_fd_sc_hd__o21ai_1
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4531_ _3604_ vssd1 vssd1 vccd1 vccd1 _3615_ sky130_fd_sc_hd__clkbuf_4
X_4462_ _2661_ _2859_ vssd1 vssd1 vccd1 vccd1 _2870_ sky130_fd_sc_hd__xor2_1
XFILLER_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7250_ _2360_ _0415_ vssd1 vssd1 vccd1 vccd1 _2362_ sky130_fd_sc_hd__and2_1
X_6201_ _1162_ _1174_ _1178_ vssd1 vssd1 vccd1 vccd1 _1209_ sky130_fd_sc_hd__a21oi_1
XFILLER_98_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4393_ _2067_ _2100_ _1968_ vssd1 vssd1 vccd1 vccd1 _2111_ sky130_fd_sc_hd__mux2_2
X_7181_ _2284_ _2285_ vssd1 vssd1 vccd1 vccd1 _2286_ sky130_fd_sc_hd__xnor2_1
X_6132_ _1125_ _1134_ vssd1 vssd1 vccd1 vccd1 _1136_ sky130_fd_sc_hd__nand2_1
XFILLER_98_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6063_ _0945_ _0947_ vssd1 vssd1 vccd1 vccd1 _1063_ sky130_fd_sc_hd__or2_1
XFILLER_85_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5014_ _3800_ _3795_ _4023_ _3928_ _4022_ vssd1 vssd1 vccd1 vccd1 _4169_ sky130_fd_sc_hd__o32a_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6965_ _1510_ _3703_ _2016_ vssd1 vssd1 vccd1 vccd1 _2049_ sky130_fd_sc_hd__o21bai_1
XFILLER_81_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5431__A1 _3690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5916_ _0906_ _0907_ _0908_ vssd1 vssd1 vccd1 vccd1 _0909_ sky130_fd_sc_hd__a21bo_1
X_6896_ _1966_ _1972_ vssd1 vssd1 vccd1 vccd1 _1973_ sky130_fd_sc_hd__and2b_1
XFILLER_21_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5847_ _0641_ _0835_ vssd1 vssd1 vccd1 vccd1 _0836_ sky130_fd_sc_hd__nand2_1
XFILLER_21_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5778_ _0711_ _0718_ _0727_ vssd1 vssd1 vccd1 vccd1 _0761_ sky130_fd_sc_hd__a21o_1
X_8566_ clknet_3_6__leaf_clk _0052_ vssd1 vssd1 vccd1 vccd1 posit_add.in1\[9\] sky130_fd_sc_hd__dfxtp_2
XANTENNA__5195__B1 _3989_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8497_ _3687_ vssd1 vssd1 vccd1 vccd1 _0066_ sky130_fd_sc_hd__clkbuf_1
X_4729_ _3881_ _3883_ vssd1 vssd1 vccd1 vccd1 _3884_ sky130_fd_sc_hd__nand2_1
X_7517_ _0419_ _2655_ vssd1 vssd1 vccd1 vccd1 _2656_ sky130_fd_sc_hd__and2_1
XFILLER_107_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4302__S _0819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7448_ _2425_ _2426_ _2427_ _2477_ vssd1 vssd1 vccd1 vccd1 _2580_ sky130_fd_sc_hd__a31o_1
XFILLER_107_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7379_ _2316_ _2317_ _2326_ vssd1 vssd1 vccd1 vccd1 _2504_ sky130_fd_sc_hd__a21oi_1
XFILLER_115_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4273__A net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5369__A _1781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5088__B _4232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7584__A _2702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8427__A1 in_reg\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6750_ _1300_ _1809_ vssd1 vssd1 vccd1 vccd1 _1812_ sky130_fd_sc_hd__and2_1
XFILLER_90_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5701_ _0112_ _3865_ _3791_ _0614_ _0619_ vssd1 vssd1 vccd1 vccd1 _0678_ sky130_fd_sc_hd__o221a_1
X_6681_ _1570_ _1571_ vssd1 vssd1 vccd1 vccd1 _1736_ sky130_fd_sc_hd__xnor2_1
X_5632_ _3814_ _0604_ _3699_ vssd1 vssd1 vccd1 vccd1 _0605_ sky130_fd_sc_hd__a21o_1
X_8420_ _3633_ vssd1 vssd1 vccd1 vccd1 _0035_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4911__A _2540_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8351_ _3536_ _3559_ _3438_ vssd1 vssd1 vccd1 vccd1 _3561_ sky130_fd_sc_hd__o21bai_1
X_5563_ _0531_ _0534_ _0535_ vssd1 vssd1 vccd1 vccd1 _0536_ sky130_fd_sc_hd__mux2_1
X_7302_ _1896_ _2418_ vssd1 vssd1 vccd1 vccd1 _2420_ sky130_fd_sc_hd__or2_1
X_4514_ _3046_ _3424_ vssd1 vssd1 vccd1 vccd1 _3435_ sky130_fd_sc_hd__nor2_1
X_8282_ _3462_ _3468_ _1319_ vssd1 vssd1 vccd1 vccd1 _3489_ sky130_fd_sc_hd__o21a_1
X_5494_ _0464_ _0466_ vssd1 vssd1 vccd1 vccd1 _0467_ sky130_fd_sc_hd__nand2_2
XFILLER_105_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5164__D _0121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4445_ _1242_ _2562_ vssd1 vssd1 vccd1 vccd1 _2683_ sky130_fd_sc_hd__and2_1
X_7233_ _0356_ _0363_ vssd1 vssd1 vccd1 vccd1 _2344_ sky130_fd_sc_hd__and2_1
X_4376_ _1429_ _1913_ vssd1 vssd1 vccd1 vccd1 _1924_ sky130_fd_sc_hd__xnor2_1
X_7164_ _1653_ _2264_ _2267_ vssd1 vssd1 vccd1 vccd1 _2268_ sky130_fd_sc_hd__o21a_1
XFILLER_112_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6115_ _4017_ _0892_ _0992_ vssd1 vssd1 vccd1 vccd1 _1118_ sky130_fd_sc_hd__or3_1
XANTENNA__6557__B _4232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7095_ _2189_ _2191_ vssd1 vssd1 vccd1 vccd1 _2192_ sky130_fd_sc_hd__xor2_1
XANTENNA__5180__C _0113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6046_ _1004_ _1043_ _1044_ vssd1 vssd1 vccd1 vccd1 _1045_ sky130_fd_sc_hd__o21a_1
XFILLER_86_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4805__B _3817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7997_ _3181_ _3182_ _3183_ vssd1 vssd1 vccd1 vccd1 _3184_ sky130_fd_sc_hd__o21ai_1
X_6948_ _2028_ _2029_ vssd1 vssd1 vccd1 vccd1 _2030_ sky130_fd_sc_hd__xor2_1
XFILLER_53_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6879_ _1384_ _1718_ vssd1 vssd1 vccd1 vccd1 _1954_ sky130_fd_sc_hd__nor2_1
XFILLER_41_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8549_ clknet_3_1__leaf_clk _0035_ vssd1 vssd1 vccd1 vccd1 out_reg\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_10_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6748__A _0218_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5652__A _3901_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8409__A1 _3621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5546__B _0467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6377__B _1401_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4437__A2 posit_add.in1\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4328__D posit_add.in2\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6393__A _3840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7920_ _3064_ _3085_ _3086_ _3098_ _3021_ vssd1 vssd1 vccd1 vccd1 _3099_ sky130_fd_sc_hd__o41a_1
XFILLER_82_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7851_ _2989_ _3022_ vssd1 vssd1 vccd1 vccd1 _3023_ sky130_fd_sc_hd__or2_2
XFILLER_91_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6802_ _1864_ _1868_ vssd1 vssd1 vccd1 vccd1 _1870_ sky130_fd_sc_hd__and2b_1
XFILLER_36_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4994_ _4095_ _4147_ _4148_ vssd1 vssd1 vccd1 vccd1 _4149_ sky130_fd_sc_hd__a21o_1
X_7782_ _2867_ _2946_ vssd1 vssd1 vccd1 vccd1 _2948_ sky130_fd_sc_hd__xnor2_1
X_6733_ _1399_ _1676_ vssd1 vssd1 vccd1 vccd1 _1794_ sky130_fd_sc_hd__nor2_1
X_6664_ _1717_ vssd1 vssd1 vccd1 vccd1 _1718_ sky130_fd_sc_hd__buf_2
XANTENNA__4641__A _3793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8403_ _0601_ _3591_ vssd1 vssd1 vccd1 vccd1 _3617_ sky130_fd_sc_hd__nand2_1
X_5615_ _0521_ _0563_ _0565_ _0587_ vssd1 vssd1 vccd1 vccd1 _0588_ sky130_fd_sc_hd__or4_1
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6595_ _1630_ _1641_ vssd1 vssd1 vccd1 vccd1 _1642_ sky130_fd_sc_hd__nand2_1
X_8334_ _3543_ vssd1 vssd1 vccd1 vccd1 _3544_ sky130_fd_sc_hd__inv_2
XFILLER_3_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5546_ _0518_ _0467_ vssd1 vssd1 vccd1 vccd1 _0519_ sky130_fd_sc_hd__or2_2
X_8265_ _3212_ _3453_ _3470_ _1177_ vssd1 vssd1 vccd1 vccd1 _3471_ sky130_fd_sc_hd__a211o_2
XFILLER_2_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5477_ _0433_ _0435_ vssd1 vssd1 vccd1 vccd1 _0450_ sky130_fd_sc_hd__xor2_4
X_4428_ _2430_ _2452_ _2463_ _2408_ _2485_ vssd1 vssd1 vccd1 vccd1 _2496_ sky130_fd_sc_hd__o2111a_1
X_7216_ _2323_ _2324_ vssd1 vssd1 vccd1 vccd1 _2325_ sky130_fd_sc_hd__nand2_1
X_8196_ _3394_ _3395_ _3303_ vssd1 vssd1 vccd1 vccd1 _3397_ sky130_fd_sc_hd__a21oi_1
XFILLER_98_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7147_ _2009_ _2046_ vssd1 vssd1 vccd1 vccd1 _2249_ sky130_fd_sc_hd__and2_1
X_4359_ _1385_ _1726_ vssd1 vssd1 vccd1 vccd1 _1737_ sky130_fd_sc_hd__or2_2
XFILLER_48_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7078_ _2138_ _2154_ _2169_ vssd1 vssd1 vccd1 vccd1 _2173_ sky130_fd_sc_hd__o21ai_1
XFILLER_86_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6029_ _1015_ _1022_ vssd1 vssd1 vccd1 vccd1 _1027_ sky130_fd_sc_hd__nor2_1
XFILLER_100_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4428__A2 _2452_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4816__A _3816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5625__A1 _1330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4726__A _3866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7102__A _0147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6380_ _1306_ _1310_ _1329_ vssd1 vssd1 vccd1 vccd1 _1405_ sky130_fd_sc_hd__a21oi_2
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5400_ _3520_ _3833_ _3834_ _0371_ _0372_ vssd1 vssd1 vccd1 vccd1 _0373_ sky130_fd_sc_hd__a32oi_4
X_5331_ _0292_ _0293_ vssd1 vssd1 vccd1 vccd1 _0304_ sky130_fd_sc_hd__xnor2_1
XFILLER_88_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8050_ _3190_ _3239_ _3240_ _0701_ vssd1 vssd1 vccd1 vccd1 _3241_ sky130_fd_sc_hd__a31o_1
X_7001_ _2086_ _2064_ _2087_ vssd1 vssd1 vccd1 vccd1 _2088_ sky130_fd_sc_hd__and3b_1
X_5262_ _0229_ _0234_ vssd1 vssd1 vccd1 vccd1 _0235_ sky130_fd_sc_hd__xor2_1
XFILLER_102_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5193_ _3893_ _0121_ vssd1 vssd1 vccd1 vccd1 _0166_ sky130_fd_sc_hd__nand2_1
XFILLER_95_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6835__B _1510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8108__A cmd\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7903_ _3080_ _3047_ _3038_ vssd1 vssd1 vccd1 vccd1 _3081_ sky130_fd_sc_hd__mux2_1
XFILLER_36_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4830__A2 _3615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7834_ _3004_ vssd1 vssd1 vccd1 vccd1 _3005_ sky130_fd_sc_hd__inv_2
X_7765_ _1253_ _1275_ vssd1 vssd1 vccd1 vccd1 _2929_ sky130_fd_sc_hd__xnor2_2
XFILLER_24_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6716_ _0080_ _1718_ vssd1 vssd1 vccd1 vccd1 _1775_ sky130_fd_sc_hd__or2_1
X_4977_ _2529_ _3703_ vssd1 vssd1 vccd1 vccd1 _4132_ sky130_fd_sc_hd__or2_1
XFILLER_51_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7696_ _2792_ _2852_ _2731_ vssd1 vssd1 vccd1 vccd1 _2853_ sky130_fd_sc_hd__mux2_1
X_6647_ _1697_ _1698_ vssd1 vssd1 vccd1 vccd1 _1699_ sky130_fd_sc_hd__xnor2_1
X_6578_ _1497_ _4213_ _4219_ vssd1 vssd1 vccd1 vccd1 _1623_ sky130_fd_sc_hd__and3b_1
XFILLER_117_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8317_ out_reg\[10\] _3197_ _3524_ _3525_ vssd1 vssd1 vccd1 vccd1 _3526_ sky130_fd_sc_hd__a22oi_1
XFILLER_3_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8088__A2 _3270_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5529_ _0499_ _0501_ _0336_ vssd1 vssd1 vccd1 vccd1 _0502_ sky130_fd_sc_hd__mux2_1
XFILLER_105_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5846__A1 _4045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8248_ _3419_ _3450_ _3451_ vssd1 vssd1 vccd1 vccd1 _3452_ sky130_fd_sc_hd__a21oi_2
X_8179_ out_reg\[4\] _3316_ _3197_ out_reg\[5\] vssd1 vssd1 vccd1 vccd1 _3379_ sky130_fd_sc_hd__a22oi_1
XANTENNA__5930__A _3770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6271__A1 _0706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4282__A0 in_reg\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5096__B _3988_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5840__A _0754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6655__B _1538_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5880_ _0854_ _0856_ _0857_ vssd1 vssd1 vccd1 vccd1 _0871_ sky130_fd_sc_hd__nand3_1
XANTENNA__6671__A _1446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4900_ _4051_ _4052_ vssd1 vssd1 vccd1 vccd1 _4055_ sky130_fd_sc_hd__nand2_1
XFILLER_18_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4831_ _3894_ vssd1 vssd1 vccd1 vccd1 _3986_ sky130_fd_sc_hd__buf_6
XANTENNA__6390__B _1414_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4762_ _3736_ _3808_ _3810_ vssd1 vssd1 vccd1 vccd1 _3917_ sky130_fd_sc_hd__and3_1
XANTENNA__4622__C _3776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7550_ _2691_ _2679_ vssd1 vssd1 vccd1 vccd1 _2692_ sky130_fd_sc_hd__xnor2_1
X_6501_ _1537_ vssd1 vssd1 vccd1 vccd1 _1538_ sky130_fd_sc_hd__clkbuf_4
X_4693_ _3079_ _3296_ _2760_ _3046_ vssd1 vssd1 vccd1 vccd1 _3848_ sky130_fd_sc_hd__a211o_1
X_7481_ _2600_ _2601_ _2520_ vssd1 vssd1 vccd1 vccd1 _2616_ sky130_fd_sc_hd__a21o_1
X_6432_ _0082_ _1423_ vssd1 vssd1 vccd1 vccd1 _1463_ sky130_fd_sc_hd__nor2_1
XFILLER_106_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7007__A _1454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6363_ _1362_ _1359_ vssd1 vssd1 vccd1 vccd1 _1387_ sky130_fd_sc_hd__or2b_1
X_8102_ _3229_ _3235_ _3276_ vssd1 vssd1 vccd1 vccd1 _3297_ sky130_fd_sc_hd__and3_1
XFILLER_115_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6294_ _1000_ _1036_ vssd1 vssd1 vccd1 vccd1 _1311_ sky130_fd_sc_hd__and2_1
XFILLER_88_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5314_ _4170_ _4193_ vssd1 vssd1 vccd1 vccd1 _0287_ sky130_fd_sc_hd__and2b_1
XANTENNA__5828__A1 _3792_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5245_ _4228_ vssd1 vssd1 vccd1 vccd1 _0218_ sky130_fd_sc_hd__inv_4
X_8033_ _1330_ _3214_ _3220_ vssd1 vssd1 vccd1 vccd1 _3223_ sky130_fd_sc_hd__a21oi_1
XFILLER_114_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5176_ _4222_ _0147_ _0148_ vssd1 vssd1 vccd1 vccd1 _0149_ sky130_fd_sc_hd__a21oi_1
XFILLER_96_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4366__A _1781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7817_ _2662_ _2664_ vssd1 vssd1 vccd1 vccd1 _2986_ sky130_fd_sc_hd__xnor2_1
X_7748_ _1297_ _2878_ _2909_ vssd1 vssd1 vccd1 vccd1 _2910_ sky130_fd_sc_hd__a21oi_1
X_7679_ _2675_ _2720_ _2722_ vssd1 vssd1 vccd1 vccd1 _2834_ sky130_fd_sc_hd__or3b_1
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5819__A1 _4222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8447__S _3655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4558__A1 _1803_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5835__A _3792_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5030_ _4183_ _4184_ vssd1 vssd1 vccd1 vccd1 _4185_ sky130_fd_sc_hd__and2_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6981_ _1954_ _2065_ _2036_ vssd1 vssd1 vccd1 vccd1 _2066_ sky130_fd_sc_hd__o21ai_1
XFILLER_26_619 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5932_ _2529_ _0787_ vssd1 vssd1 vccd1 vccd1 _0926_ sky130_fd_sc_hd__nor2_1
XFILLER_93_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6786__A2 _1782_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5863_ _0851_ _0852_ vssd1 vssd1 vccd1 vccd1 _0853_ sky130_fd_sc_hd__nor2_1
XFILLER_80_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5794_ _0761_ _0777_ vssd1 vssd1 vccd1 vccd1 _0778_ sky130_fd_sc_hd__xnor2_1
X_8582_ clknet_3_7__leaf_clk _0068_ vssd1 vssd1 vccd1 vccd1 posit_add.in2\[9\] sky130_fd_sc_hd__dfxtp_2
X_4814_ _3815_ _3702_ vssd1 vssd1 vccd1 vccd1 _3969_ sky130_fd_sc_hd__nor2_1
XFILLER_61_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7602_ _2709_ _2747_ _2748_ vssd1 vssd1 vccd1 vccd1 _2750_ sky130_fd_sc_hd__mux2_1
X_4745_ _3898_ _3899_ vssd1 vssd1 vccd1 vccd1 _3900_ sky130_fd_sc_hd__nor2_4
X_7533_ _0442_ _2670_ _2673_ _0395_ vssd1 vssd1 vccd1 vccd1 _2674_ sky130_fd_sc_hd__o2bb2ai_2
X_4676_ _3690_ _3830_ _1748_ _3696_ vssd1 vssd1 vccd1 vccd1 _3831_ sky130_fd_sc_hd__and4_1
X_7464_ _2594_ _2597_ _2486_ vssd1 vssd1 vccd1 vccd1 _2598_ sky130_fd_sc_hd__mux2_1
X_6415_ _1437_ _1438_ _1442_ vssd1 vssd1 vccd1 vccd1 _1444_ sky130_fd_sc_hd__a21oi_1
X_7395_ _2494_ vssd1 vssd1 vccd1 vccd1 _2522_ sky130_fd_sc_hd__buf_2
X_6346_ _1000_ _1367_ vssd1 vssd1 vccd1 vccd1 _1368_ sky130_fd_sc_hd__or2_1
XFILLER_115_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6277_ _1239_ _1291_ _1282_ _1019_ _1164_ vssd1 vssd1 vccd1 vccd1 _1292_ sky130_fd_sc_hd__o2111a_1
XANTENNA__7484__C_N cmd\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8016_ _2392_ _2494_ vssd1 vssd1 vccd1 vccd1 _3204_ sky130_fd_sc_hd__nand2_1
XFILLER_69_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5228_ _0178_ _0191_ _0200_ vssd1 vssd1 vccd1 vccd1 _0201_ sky130_fd_sc_hd__a21bo_1
XFILLER_84_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5159_ _0101_ _0131_ vssd1 vssd1 vccd1 vccd1 _0132_ sky130_fd_sc_hd__nand2_1
XANTENNA__6226__A1 _0795_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5029__A2 _4037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7870__A _2954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4476__B1 _1253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6933__B _3986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7193__A2 _1446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4530_ _3167_ _3509_ _3573_ _3594_ vssd1 vssd1 vccd1 vccd1 _3604_ sky130_fd_sc_hd__a211o_1
XFILLER_116_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4461_ posit_add.in1\[5\] _2848_ vssd1 vssd1 vccd1 vccd1 _2859_ sky130_fd_sc_hd__xnor2_4
XFILLER_116_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6200_ _1196_ _1206_ _1207_ vssd1 vssd1 vccd1 vccd1 _1208_ sky130_fd_sc_hd__a21oi_1
X_7180_ _1593_ _1596_ _0121_ vssd1 vssd1 vccd1 vccd1 _2285_ sky130_fd_sc_hd__and3_1
X_6131_ _1132_ _1133_ vssd1 vssd1 vccd1 vccd1 _1134_ sky130_fd_sc_hd__nand2_1
X_4392_ _2078_ _2089_ _1869_ _1957_ vssd1 vssd1 vccd1 vccd1 _2100_ sky130_fd_sc_hd__a31o_1
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6062_ _0955_ _1061_ vssd1 vssd1 vccd1 vccd1 _1062_ sky130_fd_sc_hd__nor2_1
XFILLER_100_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_498 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7004__B _4126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5013_ _4166_ _4167_ vssd1 vssd1 vccd1 vccd1 _4168_ sky130_fd_sc_hd__or2_1
XFILLER_66_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7405__B1 _2412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6964_ _2019_ _2021_ vssd1 vssd1 vccd1 vccd1 _2048_ sky130_fd_sc_hd__xnor2_1
XFILLER_93_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5915_ _0905_ _0900_ _0901_ vssd1 vssd1 vccd1 vccd1 _0908_ sky130_fd_sc_hd__nand3_1
X_6895_ _1665_ _1905_ _1967_ _1971_ vssd1 vssd1 vccd1 vccd1 _1972_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_81_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5431__A2 _3830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5846_ _4045_ _0624_ _0640_ _0639_ vssd1 vssd1 vccd1 vccd1 _0835_ sky130_fd_sc_hd__a22o_1
X_5777_ _0729_ _0759_ vssd1 vssd1 vccd1 vccd1 _0760_ sky130_fd_sc_hd__and2b_1
X_8565_ clknet_3_7__leaf_clk _0051_ vssd1 vssd1 vccd1 vccd1 posit_add.in1\[8\] sky130_fd_sc_hd__dfxtp_2
XANTENNA__5195__A1 _3763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5195__B2 _3793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8496_ posit_add.in2\[7\] in_reg\[7\] _3677_ vssd1 vssd1 vccd1 vccd1 _3687_ sky130_fd_sc_hd__mux2_1
X_4728_ _3772_ _3882_ vssd1 vssd1 vccd1 vccd1 _3883_ sky130_fd_sc_hd__nor2_4
X_7516_ _0347_ _3635_ _3830_ vssd1 vssd1 vccd1 vccd1 _2655_ sky130_fd_sc_hd__a21o_1
XFILLER_5_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4659_ _3813_ vssd1 vssd1 vccd1 vccd1 _3814_ sky130_fd_sc_hd__buf_2
X_7447_ _2577_ _2578_ _2494_ vssd1 vssd1 vccd1 vccd1 _2579_ sky130_fd_sc_hd__mux2_1
XFILLER_107_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7378_ _2315_ _2502_ vssd1 vssd1 vccd1 vccd1 _2503_ sky130_fd_sc_hd__xor2_1
XFILLER_115_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6329_ _1337_ _1047_ _1348_ vssd1 vssd1 vccd1 vccd1 _1349_ sky130_fd_sc_hd__o21a_1
XFILLER_89_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7947__A1 _2937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4554__A posit_add.in2\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5369__B _2452_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4729__A _3881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5700_ _3719_ _0676_ vssd1 vssd1 vccd1 vccd1 _0677_ sky130_fd_sc_hd__nor2_1
XFILLER_90_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6680_ _1654_ _1658_ _1694_ _1695_ _1700_ vssd1 vssd1 vccd1 vccd1 _1735_ sky130_fd_sc_hd__a32oi_4
X_5631_ _1737_ _2507_ _3775_ vssd1 vssd1 vccd1 vccd1 _0604_ sky130_fd_sc_hd__a21oi_4
XANTENNA__4911__B _3817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8350_ _3508_ _3535_ _3559_ vssd1 vssd1 vccd1 vccd1 _3560_ sky130_fd_sc_hd__and3_1
XANTENNA__8115__A1 _1330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5562_ _0494_ vssd1 vssd1 vccd1 vccd1 _0535_ sky130_fd_sc_hd__inv_2
X_4513_ _2782_ _3414_ _3123_ vssd1 vssd1 vccd1 vccd1 _3424_ sky130_fd_sc_hd__a21oi_2
X_7301_ _2417_ _2260_ _2004_ vssd1 vssd1 vccd1 vccd1 _2418_ sky130_fd_sc_hd__a21oi_1
X_8281_ _3481_ _3485_ vssd1 vssd1 vccd1 vccd1 _3487_ sky130_fd_sc_hd__or2_1
XFILLER_8_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5493_ _0457_ _0458_ _0465_ _0439_ _0440_ vssd1 vssd1 vccd1 vccd1 _0466_ sky130_fd_sc_hd__a2111o_1
X_7232_ _0370_ _2338_ _2340_ _2341_ vssd1 vssd1 vccd1 vccd1 _2343_ sky130_fd_sc_hd__a2bb2o_2
X_4444_ _2661_ _2639_ vssd1 vssd1 vccd1 vccd1 _2672_ sky130_fd_sc_hd__nor2_1
XFILLER_98_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4375_ posit_add.in2\[5\] _1902_ vssd1 vssd1 vccd1 vccd1 _1913_ sky130_fd_sc_hd__xnor2_4
X_7163_ _1620_ _2266_ _1651_ vssd1 vssd1 vccd1 vccd1 _2267_ sky130_fd_sc_hd__a21o_1
X_6114_ _1008_ _1016_ _1031_ vssd1 vssd1 vccd1 vccd1 _1117_ sky130_fd_sc_hd__a21o_1
XFILLER_100_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7094_ _2165_ _2190_ vssd1 vssd1 vccd1 vccd1 _2191_ sky130_fd_sc_hd__or2_1
XFILLER_86_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6045_ _1013_ _1024_ vssd1 vssd1 vccd1 vccd1 _1044_ sky130_fd_sc_hd__or2b_1
XFILLER_85_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7996_ _3165_ _3180_ vssd1 vssd1 vccd1 vccd1 _3183_ sky130_fd_sc_hd__xor2_1
XANTENNA__7659__A_N _2802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6947_ _1981_ _1983_ vssd1 vssd1 vccd1 vccd1 _2029_ sky130_fd_sc_hd__xnor2_1
X_6878_ _1428_ _1538_ vssd1 vssd1 vccd1 vccd1 _1953_ sky130_fd_sc_hd__nor2_1
XFILLER_22_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5829_ _0761_ _0777_ vssd1 vssd1 vccd1 vccd1 _0816_ sky130_fd_sc_hd__nand2_1
XFILLER_10_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8548_ clknet_3_0__leaf_clk _0034_ vssd1 vssd1 vccd1 vccd1 out_reg\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_10_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8479_ net4 cmd\[0\] _3638_ net1 vssd1 vssd1 vccd1 vccd1 _3675_ sky130_fd_sc_hd__and4b_1
XFILLER_5_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7624__S _2652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4549__A _3701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8455__S _3655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6930__C _3804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6939__A _1414_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7850_ _2988_ _2666_ _2987_ vssd1 vssd1 vccd1 vccd1 _3022_ sky130_fd_sc_hd__and3_1
XFILLER_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6801_ _1810_ _1865_ _1866_ _1867_ vssd1 vssd1 vccd1 vccd1 _1868_ sky130_fd_sc_hd__a22o_1
XFILLER_63_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4993_ _4070_ _4094_ vssd1 vssd1 vccd1 vccd1 _4148_ sky130_fd_sc_hd__nor2_1
X_7781_ _2858_ _2860_ _2864_ _2929_ vssd1 vssd1 vccd1 vccd1 _2946_ sky130_fd_sc_hd__a31o_1
X_6732_ _1668_ _1787_ _1791_ vssd1 vssd1 vccd1 vccd1 _1793_ sky130_fd_sc_hd__o21ai_1
XFILLER_51_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6663_ _1714_ _1716_ vssd1 vssd1 vccd1 vccd1 _1717_ sky130_fd_sc_hd__or2_1
XANTENNA__4641__B _3795_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8402_ _0521_ _3384_ _3614_ _3429_ vssd1 vssd1 vccd1 vccd1 _3616_ sky130_fd_sc_hd__a31o_1
X_5614_ _0495_ _0586_ _0561_ _0536_ vssd1 vssd1 vccd1 vccd1 _0587_ sky130_fd_sc_hd__or4_1
X_6594_ _1637_ _1640_ vssd1 vssd1 vccd1 vccd1 _1641_ sky130_fd_sc_hd__and2_1
XANTENNA__4373__A2 _1858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6849__A _1414_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8333_ _3518_ _3542_ vssd1 vssd1 vccd1 vccd1 _3543_ sky130_fd_sc_hd__xnor2_1
X_5545_ _0456_ _0460_ vssd1 vssd1 vccd1 vccd1 _0518_ sky130_fd_sc_hd__nand2_1
XFILLER_105_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8264_ _3460_ _3461_ _3469_ _0600_ vssd1 vssd1 vccd1 vccd1 _3470_ sky130_fd_sc_hd__o22ai_1
X_5476_ _0448_ _0437_ vssd1 vssd1 vccd1 vccd1 _0449_ sky130_fd_sc_hd__xnor2_2
XANTENNA__4369__A _1275_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4427_ _2474_ vssd1 vssd1 vccd1 vccd1 _2485_ sky130_fd_sc_hd__buf_2
X_8195_ _3394_ _3395_ vssd1 vssd1 vccd1 vccd1 _3396_ sky130_fd_sc_hd__or2_1
X_7215_ _2318_ _2306_ _2322_ vssd1 vssd1 vccd1 vccd1 _2324_ sky130_fd_sc_hd__nand3_1
X_7146_ _2044_ _2043_ vssd1 vssd1 vccd1 vccd1 _2248_ sky130_fd_sc_hd__and2b_1
XFILLER_48_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input4_A rst vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4358_ _1561_ _1638_ _1715_ vssd1 vssd1 vccd1 vccd1 _1726_ sky130_fd_sc_hd__nand3_4
XFILLER_59_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7077_ _1456_ _1538_ _1705_ _2171_ vssd1 vssd1 vccd1 vccd1 _2172_ sky130_fd_sc_hd__o211a_1
X_4289_ _0967_ vssd1 vssd1 vccd1 vccd1 _0009_ sky130_fd_sc_hd__clkbuf_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6028_ _1004_ _1025_ vssd1 vssd1 vccd1 vccd1 _1026_ sky130_fd_sc_hd__xnor2_1
XFILLER_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7979_ _3157_ _3163_ _3021_ vssd1 vssd1 vccd1 vccd1 _3164_ sky130_fd_sc_hd__mux2_1
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4832__A _3901_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5330_ _3988_ vssd1 vssd1 vccd1 vccd1 _0303_ sky130_fd_sc_hd__clkbuf_4
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5261_ _3800_ _3615_ _0232_ _0233_ vssd1 vssd1 vccd1 vccd1 _0234_ sky130_fd_sc_hd__o31ai_2
XFILLER_114_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7000_ _1454_ _1537_ vssd1 vssd1 vccd1 vccd1 _2087_ sky130_fd_sc_hd__nor2_1
X_5192_ _3901_ _3838_ vssd1 vssd1 vccd1 vccd1 _0165_ sky130_fd_sc_hd__nand2_1
XFILLER_68_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8254__B1 _3182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7902_ _3078_ vssd1 vssd1 vccd1 vccd1 _3080_ sky130_fd_sc_hd__clkinv_2
XANTENNA__8108__B cmd\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7833_ _2995_ _3001_ vssd1 vssd1 vccd1 vccd1 _3004_ sky130_fd_sc_hd__nor2_1
XFILLER_36_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7764_ _2856_ _2927_ vssd1 vssd1 vccd1 vccd1 _2928_ sky130_fd_sc_hd__xnor2_1
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6715_ _1702_ _1732_ vssd1 vssd1 vccd1 vccd1 _1774_ sky130_fd_sc_hd__xnor2_1
XANTENNA__5240__B1 _3750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4976_ _2529_ _4126_ _4130_ vssd1 vssd1 vccd1 vccd1 _4131_ sky130_fd_sc_hd__or3_1
XANTENNA__4371__B _1858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7695_ _2708_ _2803_ vssd1 vssd1 vccd1 vccd1 _2852_ sky130_fd_sc_hd__nor2_1
X_6646_ _1548_ _1547_ vssd1 vssd1 vccd1 vccd1 _1698_ sky130_fd_sc_hd__xor2_1
X_6577_ _1587_ _1590_ _1621_ vssd1 vssd1 vccd1 vccd1 _1622_ sky130_fd_sc_hd__a21o_1
XANTENNA__6579__A _1420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8316_ out_reg\[9\] _3242_ _1177_ vssd1 vssd1 vccd1 vccd1 _3525_ sky130_fd_sc_hd__a21bo_1
X_5528_ _0099_ _0334_ vssd1 vssd1 vccd1 vccd1 _0501_ sky130_fd_sc_hd__or2_1
XFILLER_3_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8247_ _3419_ _3450_ _3416_ vssd1 vssd1 vccd1 vccd1 _3451_ sky130_fd_sc_hd__o21bai_1
X_5459_ _0430_ _0431_ vssd1 vssd1 vccd1 vccd1 _0432_ sky130_fd_sc_hd__and2_1
XFILLER_105_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8178_ _3358_ _3369_ _3377_ _3195_ vssd1 vssd1 vccd1 vccd1 _3378_ sky130_fd_sc_hd__a31o_2
XANTENNA__5930__B _0773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7129_ _1531_ _2079_ vssd1 vssd1 vccd1 vccd1 _2229_ sky130_fd_sc_hd__nand2_1
XFILLER_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6271__A2 _1164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4282__A1 in_reg\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8034__A _0600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5393__A _1748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7287__A1 _2349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6936__B _3703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4737__A _3729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6671__B _0548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8003__A3 _3182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4830_ _2540_ _3615_ _3984_ _3983_ _3955_ vssd1 vssd1 vccd1 vccd1 _3985_ sky130_fd_sc_hd__o32a_1
XFILLER_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4761_ _3906_ _3909_ vssd1 vssd1 vccd1 vccd1 _3916_ sky130_fd_sc_hd__or2b_1
XANTENNA__7783__A _1308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6500_ _1535_ _1536_ vssd1 vssd1 vccd1 vccd1 _1537_ sky130_fd_sc_hd__nand2_4
X_4692_ _2826_ _3307_ _3740_ vssd1 vssd1 vccd1 vccd1 _3847_ sky130_fd_sc_hd__a21o_1
X_7480_ _2579_ _2614_ _2486_ vssd1 vssd1 vccd1 vccd1 _2615_ sky130_fd_sc_hd__mux2_1
XFILLER_119_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6431_ _1435_ _1448_ _1453_ _1460_ vssd1 vssd1 vccd1 vccd1 _1461_ sky130_fd_sc_hd__a31o_1
XANTENNA__6399__A _1400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6362_ _1383_ _1384_ vssd1 vssd1 vccd1 vccd1 _1386_ sky130_fd_sc_hd__nor2_2
X_5313_ _0271_ _0270_ vssd1 vssd1 vccd1 vccd1 _0286_ sky130_fd_sc_hd__xor2_1
X_8101_ _3227_ _3294_ vssd1 vssd1 vccd1 vccd1 _3295_ sky130_fd_sc_hd__or2_1
XFILLER_114_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6293_ _1307_ _1309_ _1155_ vssd1 vssd1 vccd1 vccd1 _1310_ sky130_fd_sc_hd__a21o_1
XFILLER_114_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5244_ _0215_ _0216_ vssd1 vssd1 vccd1 vccd1 _0217_ sky130_fd_sc_hd__and2_1
X_8032_ _0601_ _3214_ _3220_ vssd1 vssd1 vccd1 vccd1 _3222_ sky130_fd_sc_hd__and3_1
X_5175_ _4017_ _3795_ vssd1 vssd1 vccd1 vccd1 _0148_ sky130_fd_sc_hd__nor2_1
XANTENNA__7023__A _4153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8119__A _0701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4366__B _1803_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5478__A _0440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7816_ _2945_ _2982_ _2984_ vssd1 vssd1 vccd1 vccd1 _2985_ sky130_fd_sc_hd__o21a_1
XFILLER_51_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4959_ _4097_ _4112_ _4113_ vssd1 vssd1 vccd1 vccd1 _4114_ sky130_fd_sc_hd__a21oi_1
X_7747_ _1297_ _2819_ vssd1 vssd1 vccd1 vccd1 _2909_ sky130_fd_sc_hd__nor2_1
XFILLER_20_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7678_ _2741_ _2831_ _2832_ vssd1 vssd1 vccd1 vccd1 _2833_ sky130_fd_sc_hd__a21oi_1
X_6629_ _1677_ _1678_ vssd1 vssd1 vccd1 vccd1 _1679_ sky130_fd_sc_hd__xnor2_1
XFILLER_20_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8463__S _3655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5755__A1 _0113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7542__S _2652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6980_ _1401_ _1538_ vssd1 vssd1 vccd1 vccd1 _2065_ sky130_fd_sc_hd__nor2_1
XFILLER_81_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5931_ _3735_ _0676_ vssd1 vssd1 vccd1 vccd1 _0924_ sky130_fd_sc_hd__nor2_1
XFILLER_81_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5862_ _0849_ _0850_ _0827_ _0829_ vssd1 vssd1 vccd1 vccd1 _0852_ sky130_fd_sc_hd__a211oi_1
X_5793_ _0770_ _0776_ vssd1 vssd1 vccd1 vccd1 _0777_ sky130_fd_sc_hd__xor2_1
X_8581_ clknet_3_7__leaf_clk _0067_ vssd1 vssd1 vccd1 vccd1 posit_add.in2\[8\] sky130_fd_sc_hd__dfxtp_2
X_4813_ _3958_ _3960_ vssd1 vssd1 vccd1 vccd1 _3968_ sky130_fd_sc_hd__xnor2_1
XFILLER_21_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7601_ _2676_ _2702_ vssd1 vssd1 vccd1 vccd1 _2748_ sky130_fd_sc_hd__and2_2
XFILLER_33_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4744_ _2485_ _3766_ _3767_ _3678_ vssd1 vssd1 vccd1 vccd1 _3899_ sky130_fd_sc_hd__a31o_1
X_7532_ _0356_ _2651_ _2671_ vssd1 vssd1 vccd1 vccd1 _2673_ sky130_fd_sc_hd__a21oi_2
XFILLER_119_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4675_ _2408_ vssd1 vssd1 vccd1 vccd1 _3830_ sky130_fd_sc_hd__clkbuf_4
X_7463_ _2451_ _2512_ _2596_ vssd1 vssd1 vccd1 vccd1 _2597_ sky130_fd_sc_hd__a21oi_1
X_6414_ _1437_ _1438_ _1442_ vssd1 vssd1 vccd1 vccd1 _1443_ sky130_fd_sc_hd__and3_1
X_7394_ _2487_ _2515_ _2520_ vssd1 vssd1 vccd1 vccd1 _2521_ sky130_fd_sc_hd__mux2_2
X_6345_ _1365_ _1366_ vssd1 vssd1 vccd1 vccd1 _1367_ sky130_fd_sc_hd__nand2_1
XANTENNA__6857__A _1420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6276_ _0706_ _1128_ vssd1 vssd1 vccd1 vccd1 _1291_ sky130_fd_sc_hd__nor2_1
XANTENNA__5761__A _0113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5227_ _0153_ _0169_ _0176_ vssd1 vssd1 vccd1 vccd1 _0200_ sky130_fd_sc_hd__or3_1
X_8015_ _2451_ _2578_ _2590_ vssd1 vssd1 vccd1 vccd1 _3203_ sky130_fd_sc_hd__a21o_1
XFILLER_88_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5158_ _0118_ _0130_ _0128_ vssd1 vssd1 vccd1 vccd1 _0131_ sky130_fd_sc_hd__a21o_1
XANTENNA__6226__A2 _1164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5089_ _3800_ _4232_ _4242_ vssd1 vssd1 vccd1 vccd1 _4244_ sky130_fd_sc_hd__o21ai_1
XFILLER_71_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5434__B1 _2980_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5001__A _3719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_450 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6188__B_N _1097_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4460_ posit_add.in1\[4\] _2551_ _1242_ vssd1 vssd1 vccd1 vccd1 _2848_ sky130_fd_sc_hd__o21ai_2
XFILLER_116_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4391_ _1506_ _1858_ vssd1 vssd1 vccd1 vccd1 _2089_ sky130_fd_sc_hd__or2_1
X_6130_ _1123_ _1124_ vssd1 vssd1 vccd1 vccd1 _1133_ sky130_fd_sc_hd__xnor2_1
XFILLER_98_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6061_ _0951_ _0954_ vssd1 vssd1 vccd1 vccd1 _1061_ sky130_fd_sc_hd__nor2_1
XFILLER_100_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5012_ _4005_ _4155_ _4165_ vssd1 vssd1 vccd1 vccd1 _4167_ sky130_fd_sc_hd__and3_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6963_ _2009_ _2046_ vssd1 vssd1 vccd1 vccd1 _2047_ sky130_fd_sc_hd__xnor2_1
XFILLER_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5914_ _0889_ _0890_ vssd1 vssd1 vccd1 vccd1 _0907_ sky130_fd_sc_hd__xor2_1
X_6894_ _1907_ _1969_ _1970_ vssd1 vssd1 vccd1 vccd1 _1971_ sky130_fd_sc_hd__a21o_1
XANTENNA__5431__A3 _3635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5845_ _0831_ _0833_ vssd1 vssd1 vccd1 vccd1 _0834_ sky130_fd_sc_hd__nand2_1
XFILLER_22_612 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5776_ _0729_ _0730_ _0758_ vssd1 vssd1 vccd1 vccd1 _0759_ sky130_fd_sc_hd__or3_1
X_8564_ clknet_3_7__leaf_clk _0050_ vssd1 vssd1 vccd1 vccd1 posit_add.in1\[7\] sky130_fd_sc_hd__dfxtp_2
XANTENNA__5195__A2 _3840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8495_ _3686_ vssd1 vssd1 vccd1 vccd1 _0065_ sky130_fd_sc_hd__clkbuf_1
X_4727_ _3145_ _3783_ _3785_ _3787_ vssd1 vssd1 vccd1 vccd1 _3882_ sky130_fd_sc_hd__a31oi_4
X_7515_ _0348_ _0349_ _2651_ vssd1 vssd1 vccd1 vccd1 _2654_ sky130_fd_sc_hd__mux2_2
X_4658_ _3811_ _3812_ vssd1 vssd1 vccd1 vccd1 _3813_ sky130_fd_sc_hd__nand2_2
X_7446_ _2506_ _2511_ _2410_ vssd1 vssd1 vccd1 vccd1 _2578_ sky130_fd_sc_hd__mux2_1
X_4589_ _3741_ _3743_ vssd1 vssd1 vccd1 vccd1 _3744_ sky130_fd_sc_hd__nand2_1
XFILLER_1_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7377_ _2297_ _2497_ _2295_ vssd1 vssd1 vccd1 vccd1 _2502_ sky130_fd_sc_hd__o21a_1
XFILLER_107_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6328_ _1346_ _1347_ vssd1 vssd1 vccd1 vccd1 _1348_ sky130_fd_sc_hd__nor2_1
XFILLER_89_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6259_ _1262_ _1270_ _1271_ vssd1 vssd1 vccd1 vccd1 _1272_ sky130_fd_sc_hd__a21oi_1
XFILLER_88_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7211__A _4250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4630__A1 _3232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5385__B _2452_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6497__A _4157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4729__B _3883_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8348__C1 _0600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7571__A0 _3855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5630_ _0356_ _0363_ vssd1 vssd1 vccd1 vccd1 _0603_ sky130_fd_sc_hd__or2_1
X_5561_ _0532_ _0533_ _0480_ vssd1 vssd1 vccd1 vccd1 _0534_ sky130_fd_sc_hd__mux2_1
XFILLER_117_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7300_ _2085_ _2247_ _2253_ _2255_ vssd1 vssd1 vccd1 vccd1 _2417_ sky130_fd_sc_hd__a31o_1
X_4512_ _2881_ _3403_ _2705_ vssd1 vssd1 vccd1 vccd1 _3414_ sky130_fd_sc_hd__o21ai_1
X_8280_ _3481_ _3485_ vssd1 vssd1 vccd1 vccd1 _3486_ sky130_fd_sc_hd__nand2_1
X_5492_ _0461_ _0401_ vssd1 vssd1 vccd1 vccd1 _0465_ sky130_fd_sc_hd__nor2_1
XFILLER_105_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7323__B1 _2440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7231_ _0369_ _2338_ vssd1 vssd1 vccd1 vccd1 _2341_ sky130_fd_sc_hd__xnor2_1
XFILLER_104_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4443_ _2606_ vssd1 vssd1 vccd1 vccd1 _2661_ sky130_fd_sc_hd__buf_4
XFILLER_98_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4374_ posit_add.in2\[4\] _1352_ _1264_ vssd1 vssd1 vccd1 vccd1 _1902_ sky130_fd_sc_hd__o21ai_2
X_7162_ _1584_ _1618_ vssd1 vssd1 vccd1 vccd1 _2266_ sky130_fd_sc_hd__nand2_1
XFILLER_112_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6113_ _1107_ _1115_ vssd1 vssd1 vccd1 vccd1 _1116_ sky130_fd_sc_hd__xor2_1
X_7093_ _2128_ _2164_ vssd1 vssd1 vccd1 vccd1 _2190_ sky130_fd_sc_hd__and2_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6044_ _1013_ _1023_ _1033_ vssd1 vssd1 vccd1 vccd1 _1043_ sky130_fd_sc_hd__and3_1
XFILLER_58_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7995_ _1275_ _1253_ _2721_ vssd1 vssd1 vccd1 vccd1 _3182_ sky130_fd_sc_hd__mux2_4
XFILLER_26_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6946_ _2011_ _2026_ _2027_ vssd1 vssd1 vccd1 vccd1 _2028_ sky130_fd_sc_hd__a21oi_1
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4612__A1 _1803_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8339__C1 _1177_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6877_ _1944_ _1941_ vssd1 vssd1 vccd1 vccd1 _1952_ sky130_fd_sc_hd__xor2_1
XANTENNA__5486__A _0440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5828_ _3792_ _0782_ _0780_ vssd1 vssd1 vccd1 vccd1 _0815_ sky130_fd_sc_hd__o21ai_1
XANTENNA__6365__A1 _1097_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5759_ _0666_ _0667_ _3865_ vssd1 vssd1 vccd1 vccd1 _0741_ sky130_fd_sc_hd__a21o_1
X_8547_ clknet_3_2__leaf_clk _0033_ vssd1 vssd1 vccd1 vccd1 out_reg\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_10_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8478_ _3674_ vssd1 vssd1 vccd1 vccd1 _0058_ sky130_fd_sc_hd__clkbuf_1
XFILLER_118_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7429_ _2522_ _2447_ _2558_ vssd1 vssd1 vccd1 vccd1 _2559_ sky130_fd_sc_hd__or3_1
XANTENNA__4549__B _3703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8290__A1 _3195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8471__S _3654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4603__A1 _1913_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7595__B _2702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4367__B1 _1275_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6939__B _1531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4475__A posit_add.in1\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8033__A1 _1330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6800_ _1810_ _1865_ vssd1 vssd1 vccd1 vccd1 _1867_ sky130_fd_sc_hd__xor2_1
XFILLER_63_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4992_ _4115_ _4145_ _4146_ vssd1 vssd1 vccd1 vccd1 _4147_ sky130_fd_sc_hd__a21o_1
X_7780_ _2942_ _2944_ vssd1 vssd1 vccd1 vccd1 _2945_ sky130_fd_sc_hd__and2b_1
XFILLER_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6731_ _1789_ _1790_ vssd1 vssd1 vccd1 vccd1 _1791_ sky130_fd_sc_hd__nand2_1
X_6662_ _1304_ _1711_ _1713_ vssd1 vssd1 vccd1 vccd1 _1716_ sky130_fd_sc_hd__and3_1
Xclkbuf_3_2__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_8401_ _3553_ _3554_ _3587_ vssd1 vssd1 vccd1 vccd1 _3614_ sky130_fd_sc_hd__or3_1
X_5613_ _0492_ _0508_ _0494_ vssd1 vssd1 vccd1 vccd1 _0586_ sky130_fd_sc_hd__mux2_1
X_6593_ _1639_ _1636_ vssd1 vssd1 vccd1 vccd1 _1640_ sky130_fd_sc_hd__or2_1
X_8332_ _3259_ _3308_ _3429_ vssd1 vssd1 vccd1 vccd1 _3542_ sky130_fd_sc_hd__o21bai_1
XFILLER_117_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6849__B _1782_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5544_ _0509_ _0516_ _0494_ vssd1 vssd1 vccd1 vccd1 _0517_ sky130_fd_sc_hd__mux2_1
X_8263_ _3463_ _3468_ vssd1 vssd1 vccd1 vccd1 _3469_ sky130_fd_sc_hd__xor2_1
X_5475_ _0425_ vssd1 vssd1 vccd1 vccd1 _0448_ sky130_fd_sc_hd__inv_2
XANTENNA__7026__A _4217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4426_ _1759_ _1979_ _1561_ vssd1 vssd1 vccd1 vccd1 _2474_ sky130_fd_sc_hd__o21a_1
X_8194_ _3334_ _3374_ _3182_ vssd1 vssd1 vccd1 vccd1 _3395_ sky130_fd_sc_hd__o21a_1
X_7214_ _2318_ _2306_ _2322_ vssd1 vssd1 vccd1 vccd1 _2323_ sky130_fd_sc_hd__a21o_1
X_7145_ _2118_ _2120_ _2151_ _2244_ _2246_ vssd1 vssd1 vccd1 vccd1 _2247_ sky130_fd_sc_hd__a41o_2
XFILLER_113_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4357_ _1693_ _1704_ vssd1 vssd1 vccd1 vccd1 _1715_ sky130_fd_sc_hd__nor2_1
XFILLER_59_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7076_ _1676_ _1718_ vssd1 vssd1 vccd1 vccd1 _2171_ sky130_fd_sc_hd__nor2_1
X_4288_ in_reg\[5\] in_reg\[6\] _0830_ vssd1 vssd1 vccd1 vccd1 _0967_ sky130_fd_sc_hd__mux2_1
XFILLER_59_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6027_ _1013_ _1024_ vssd1 vssd1 vccd1 vccd1 _1025_ sky130_fd_sc_hd__xnor2_1
XANTENNA__4385__A posit_add.in2\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7978_ _3003_ _3141_ _3004_ vssd1 vssd1 vccd1 vccd1 _3163_ sky130_fd_sc_hd__a21o_1
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4832__B _3986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6929_ _0218_ _1711_ _1950_ vssd1 vssd1 vccd1 vccd1 _2009_ sky130_fd_sc_hd__and3_1
XFILLER_42_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6338__B2 _1097_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6338__A1 _0722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_448 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5552__A2 _0440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5260_ _0230_ _0231_ vssd1 vssd1 vccd1 vccd1 _0233_ sky130_fd_sc_hd__or2b_1
XFILLER_114_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5191_ _0134_ _0162_ vssd1 vssd1 vccd1 vccd1 _0164_ sky130_fd_sc_hd__xor2_1
XFILLER_95_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7901_ _3044_ _3060_ _3077_ vssd1 vssd1 vccd1 vccd1 _3078_ sky130_fd_sc_hd__a21oi_1
XFILLER_36_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7832_ _2995_ _3001_ vssd1 vssd1 vccd1 vccd1 _3003_ sky130_fd_sc_hd__nand2_1
XFILLER_24_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4975_ _4117_ _4129_ vssd1 vssd1 vccd1 vccd1 _4130_ sky130_fd_sc_hd__xnor2_1
XFILLER_51_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7763_ _1308_ _2868_ vssd1 vssd1 vccd1 vccd1 _2927_ sky130_fd_sc_hd__and2_1
XANTENNA__5240__A1 _3827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5240__B2 _3763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6714_ _1653_ _1772_ vssd1 vssd1 vccd1 vccd1 _1773_ sky130_fd_sc_hd__or2_1
X_7694_ _2811_ _2802_ vssd1 vssd1 vccd1 vccd1 _2851_ sky130_fd_sc_hd__nor2_1
X_6645_ _1655_ _1551_ _1656_ _1657_ vssd1 vssd1 vccd1 vccd1 _1697_ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6576_ _1499_ _1591_ vssd1 vssd1 vccd1 vccd1 _1621_ sky130_fd_sc_hd__and2b_1
XANTENNA__6579__B _1446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8315_ _3212_ _3506_ _3507_ _3523_ vssd1 vssd1 vccd1 vccd1 _3524_ sky130_fd_sc_hd__a31o_1
X_5527_ _0498_ _0499_ _0338_ vssd1 vssd1 vccd1 vccd1 _0500_ sky130_fd_sc_hd__mux2_1
XFILLER_105_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8246_ _3449_ vssd1 vssd1 vccd1 vccd1 _3450_ sky130_fd_sc_hd__buf_2
X_5458_ _0426_ _0429_ vssd1 vssd1 vccd1 vccd1 _0431_ sky130_fd_sc_hd__nand2_1
X_4409_ _1495_ _1517_ _1638_ vssd1 vssd1 vccd1 vccd1 _2287_ sky130_fd_sc_hd__a21oi_1
X_5389_ _1748_ _2507_ vssd1 vssd1 vccd1 vccd1 _0362_ sky130_fd_sc_hd__nor2_1
X_8177_ _3374_ _3375_ _3376_ vssd1 vssd1 vccd1 vccd1 _3377_ sky130_fd_sc_hd__a21o_1
XFILLER_115_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7128_ _2211_ _2227_ vssd1 vssd1 vccd1 vccd1 _2228_ sky130_fd_sc_hd__or2_1
XFILLER_59_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7059_ _2123_ _2147_ vssd1 vssd1 vccd1 vccd1 _2152_ sky130_fd_sc_hd__xnor2_1
XFILLER_86_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5004__A _4157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7220__A2 _0092_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8484__A1 in_reg\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6495__B1 _1531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7995__A0 _1275_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4760_ _3896_ _3905_ vssd1 vssd1 vccd1 vccd1 _3915_ sky130_fd_sc_hd__nand2_1
XFILLER_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4691_ _3751_ _3752_ _3167_ vssd1 vssd1 vccd1 vccd1 _3846_ sky130_fd_sc_hd__a21oi_2
X_6430_ _1457_ _1459_ vssd1 vssd1 vccd1 vccd1 _1460_ sky130_fd_sc_hd__and2b_1
X_6361_ _3615_ vssd1 vssd1 vccd1 vccd1 _1384_ sky130_fd_sc_hd__buf_4
XANTENNA__6399__B _1384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5312_ _4228_ _2540_ vssd1 vssd1 vccd1 vccd1 _0285_ sky130_fd_sc_hd__or2_1
X_8100_ _3228_ _3238_ _3277_ vssd1 vssd1 vccd1 vccd1 _3294_ sky130_fd_sc_hd__and3_1
XFILLER_114_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6292_ _1158_ _1190_ vssd1 vssd1 vccd1 vccd1 _1309_ sky130_fd_sc_hd__or2_1
XANTENNA__8475__A1 posit_add.in1\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5243_ _0214_ _4175_ _0212_ vssd1 vssd1 vccd1 vccd1 _0216_ sky130_fd_sc_hd__or3_1
X_8031_ _0595_ _3219_ vssd1 vssd1 vccd1 vccd1 _3220_ sky130_fd_sc_hd__xnor2_1
X_5174_ _3943_ vssd1 vssd1 vccd1 vccd1 _0147_ sky130_fd_sc_hd__buf_4
XFILLER_96_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4663__A _3816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7815_ _2939_ _2983_ vssd1 vssd1 vccd1 vccd1 _2984_ sky130_fd_sc_hd__nor2_1
XFILLER_101_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5213__A1 _4222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4958_ _4099_ _4111_ vssd1 vssd1 vccd1 vccd1 _4113_ sky130_fd_sc_hd__and2b_1
X_7746_ _2845_ _2907_ vssd1 vssd1 vccd1 vccd1 _2908_ sky130_fd_sc_hd__xor2_2
X_4889_ _3729_ _4043_ vssd1 vssd1 vccd1 vccd1 _4044_ sky130_fd_sc_hd__nor2_1
X_7677_ _2729_ _2737_ _2740_ vssd1 vssd1 vccd1 vccd1 _2832_ sky130_fd_sc_hd__and3_1
X_6628_ _1353_ _1354_ _4089_ vssd1 vssd1 vccd1 vccd1 _1678_ sky130_fd_sc_hd__nand3_1
XFILLER_20_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6559_ _1598_ _1601_ vssd1 vssd1 vccd1 vccd1 _1602_ sky130_fd_sc_hd__xor2_1
XFILLER_3_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5819__A3 _0113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8229_ _3428_ _3430_ vssd1 vssd1 vccd1 vccd1 _3432_ sky130_fd_sc_hd__nand2_1
XFILLER_105_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6952__A1 _1384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4715__B1 _3615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8209__A1 _0600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7778__B _2937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5930_ _3770_ _0773_ vssd1 vssd1 vccd1 vccd1 _0923_ sky130_fd_sc_hd__nor2_1
XFILLER_53_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4483__A posit_add.in1\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5861_ _0827_ _0829_ _0849_ _0850_ vssd1 vssd1 vccd1 vccd1 _0851_ sky130_fd_sc_hd__o211a_1
XFILLER_61_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7794__A _2954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7600_ _2712_ _2718_ _2746_ vssd1 vssd1 vccd1 vccd1 _2747_ sky130_fd_sc_hd__a21oi_1
X_5792_ _0771_ _0775_ vssd1 vssd1 vccd1 vccd1 _0776_ sky130_fd_sc_hd__xnor2_1
X_8580_ clknet_3_7__leaf_clk _0066_ vssd1 vssd1 vccd1 vccd1 posit_add.in2\[7\] sky130_fd_sc_hd__dfxtp_1
X_4812_ _3949_ _3966_ vssd1 vssd1 vccd1 vccd1 _3967_ sky130_fd_sc_hd__or2_1
XFILLER_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4743_ _3808_ _3810_ _2485_ vssd1 vssd1 vccd1 vccd1 _3898_ sky130_fd_sc_hd__a21oi_2
XFILLER_21_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7531_ _0363_ _2651_ vssd1 vssd1 vccd1 vccd1 _2671_ sky130_fd_sc_hd__nor2_1
XFILLER_119_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7462_ _2382_ _2454_ _2489_ _2494_ vssd1 vssd1 vccd1 vccd1 _2596_ sky130_fd_sc_hd__o211a_1
XFILLER_107_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6413_ _0795_ _1392_ _1441_ vssd1 vssd1 vccd1 vccd1 _1442_ sky130_fd_sc_hd__a21o_1
X_4674_ _3827_ _3828_ vssd1 vssd1 vccd1 vccd1 _3829_ sky130_fd_sc_hd__or2_1
X_7393_ _2519_ vssd1 vssd1 vccd1 vccd1 _2520_ sky130_fd_sc_hd__buf_2
X_6344_ _1358_ _1364_ vssd1 vssd1 vccd1 vccd1 _1366_ sky130_fd_sc_hd__nand2_1
XANTENNA__6857__B _1538_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6275_ _1288_ _1289_ vssd1 vssd1 vccd1 vccd1 _1290_ sky130_fd_sc_hd__nand2_1
XFILLER_103_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7034__A _1782_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5226_ _0197_ _0198_ vssd1 vssd1 vccd1 vccd1 _0199_ sky130_fd_sc_hd__or2_1
X_8014_ _1319_ _3200_ _3201_ vssd1 vssd1 vccd1 vccd1 _3202_ sky130_fd_sc_hd__and3_1
XFILLER_84_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5157_ _0128_ _0129_ vssd1 vssd1 vccd1 vccd1 _0130_ sky130_fd_sc_hd__nor2_1
X_5088_ _3800_ _4232_ _4242_ vssd1 vssd1 vccd1 vccd1 _4243_ sky130_fd_sc_hd__or3_1
XFILLER_84_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5001__B _3817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7908__S _2999_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7729_ _1297_ _2841_ _2888_ vssd1 vssd1 vccd1 vccd1 _2889_ sky130_fd_sc_hd__o21bai_1
XFILLER_40_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5952__A _3770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4390_ _1506_ _1913_ vssd1 vssd1 vccd1 vccd1 _2078_ sky130_fd_sc_hd__xor2_1
XFILLER_7_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4478__A _2980_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6060_ _1058_ _1059_ _0949_ vssd1 vssd1 vccd1 vccd1 _1060_ sky130_fd_sc_hd__o21bai_1
XFILLER_98_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5011_ _4005_ _4155_ _4165_ vssd1 vssd1 vccd1 vccd1 _4166_ sky130_fd_sc_hd__a21oi_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6962_ _2043_ _2044_ vssd1 vssd1 vccd1 vccd1 _2046_ sky130_fd_sc_hd__xnor2_1
XFILLER_81_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5913_ _0900_ _0901_ _0905_ vssd1 vssd1 vccd1 vccd1 _0906_ sky130_fd_sc_hd__a21o_1
X_6893_ _1665_ _1905_ vssd1 vssd1 vccd1 vccd1 _1970_ sky130_fd_sc_hd__nor2_1
X_5844_ _3776_ _0624_ _0831_ _0832_ vssd1 vssd1 vccd1 vccd1 _0833_ sky130_fd_sc_hd__nand4_1
XFILLER_22_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8563_ clknet_3_2__leaf_clk _0049_ vssd1 vssd1 vccd1 vccd1 posit_add.in1\[6\] sky130_fd_sc_hd__dfxtp_2
XFILLER_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4927__B1 _3930_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5775_ _3735_ _0757_ vssd1 vssd1 vccd1 vccd1 _0758_ sky130_fd_sc_hd__xnor2_1
XANTENNA__8118__B1 _3195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7514_ _0420_ _0410_ _2652_ vssd1 vssd1 vccd1 vccd1 _2653_ sky130_fd_sc_hd__mux2_2
X_8494_ posit_add.in2\[6\] in_reg\[6\] _3677_ vssd1 vssd1 vccd1 vccd1 _3686_ sky130_fd_sc_hd__mux2_1
X_4726_ _3866_ vssd1 vssd1 vccd1 vccd1 _3881_ sky130_fd_sc_hd__clkbuf_4
XFILLER_21_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4657_ _2485_ _3766_ _3767_ _3678_ vssd1 vssd1 vccd1 vccd1 _3812_ sky130_fd_sc_hd__a31oi_2
X_7445_ _2473_ _2501_ _2410_ vssd1 vssd1 vccd1 vccd1 _2577_ sky130_fd_sc_hd__mux2_1
XFILLER_107_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7376_ _4153_ _2431_ _2499_ _2416_ _2500_ vssd1 vssd1 vccd1 vccd1 _2501_ sky130_fd_sc_hd__o221a_1
X_6327_ _1345_ _1000_ vssd1 vssd1 vccd1 vccd1 _1347_ sky130_fd_sc_hd__and2b_1
XFILLER_89_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4588_ _2903_ _3307_ _3742_ _3477_ vssd1 vssd1 vccd1 vccd1 _3743_ sky130_fd_sc_hd__a211o_1
XFILLER_1_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4388__A posit_add.in2\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6258_ _1263_ _1265_ _1269_ vssd1 vssd1 vccd1 vccd1 _1271_ sky130_fd_sc_hd__and3_1
XFILLER_88_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6189_ _1194_ _1195_ vssd1 vssd1 vccd1 vccd1 _1196_ sky130_fd_sc_hd__xor2_1
XFILLER_88_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5209_ _0146_ _0181_ vssd1 vssd1 vccd1 vccd1 _0182_ sky130_fd_sc_hd__xnor2_1
XFILLER_57_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7211__B _3989_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8469__S _3654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5646__B2 _2507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7571__A1 _3802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5560_ _0476_ _0339_ _0470_ vssd1 vssd1 vccd1 vccd1 _0533_ sky130_fd_sc_hd__mux2_1
X_4511_ _2958_ _3392_ vssd1 vssd1 vccd1 vccd1 _3403_ sky130_fd_sc_hd__nor2_1
X_5491_ _0462_ _0439_ _0463_ vssd1 vssd1 vccd1 vccd1 _0464_ sky130_fd_sc_hd__nand3_1
XANTENNA__7791__B _2941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4442_ _2606_ _2639_ vssd1 vssd1 vccd1 vccd1 _2650_ sky130_fd_sc_hd__and2_1
X_7230_ _3722_ _3788_ _2339_ vssd1 vssd1 vccd1 vccd1 _2340_ sky130_fd_sc_hd__o21a_1
XFILLER_113_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4373_ _1429_ _1858_ _1880_ vssd1 vssd1 vccd1 vccd1 _1891_ sky130_fd_sc_hd__o21a_1
X_7161_ _2262_ _2263_ _1769_ vssd1 vssd1 vccd1 vccd1 _2264_ sky130_fd_sc_hd__o21ai_1
X_6112_ _1112_ _1113_ vssd1 vssd1 vccd1 vccd1 _1115_ sky130_fd_sc_hd__or2b_1
XFILLER_98_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7092_ _2185_ _2186_ _2187_ vssd1 vssd1 vccd1 vccd1 _2189_ sky130_fd_sc_hd__or3_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6043_ _1004_ _1041_ vssd1 vssd1 vccd1 vccd1 _1042_ sky130_fd_sc_hd__xnor2_1
XFILLER_86_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7312__A _2333_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7994_ _3033_ _3172_ _3180_ vssd1 vssd1 vccd1 vccd1 _3181_ sky130_fd_sc_hd__a21o_1
X_6945_ _2024_ _2025_ vssd1 vssd1 vccd1 vccd1 _2027_ sky130_fd_sc_hd__and2_1
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4612__A2 _3635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6876_ _1711_ _0121_ _1950_ vssd1 vssd1 vccd1 vccd1 _1951_ sky130_fd_sc_hd__and3_1
XFILLER_50_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5827_ _0810_ _0813_ vssd1 vssd1 vccd1 vccd1 _0814_ sky130_fd_sc_hd__xnor2_1
XANTENNA__4390__B _1913_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5758_ _3866_ _0667_ _0738_ _0739_ vssd1 vssd1 vccd1 vccd1 _0740_ sky130_fd_sc_hd__a31o_1
X_8546_ clknet_3_2__leaf_clk _0032_ vssd1 vssd1 vccd1 vccd1 out_reg\[12\] sky130_fd_sc_hd__dfxtp_1
X_4709_ _3863_ vssd1 vssd1 vccd1 vccd1 _3864_ sky130_fd_sc_hd__buf_2
X_8477_ in_reg\[15\] _1253_ _3654_ vssd1 vssd1 vccd1 vccd1 _3674_ sky130_fd_sc_hd__mux2_1
X_5689_ _4043_ _3791_ vssd1 vssd1 vccd1 vccd1 _0665_ sky130_fd_sc_hd__nor2_1
X_7428_ _2454_ _2538_ _2557_ _2431_ vssd1 vssd1 vccd1 vccd1 _2558_ sky130_fd_sc_hd__a22o_1
XFILLER_118_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7921__S _2999_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7359_ _2402_ _2405_ vssd1 vssd1 vccd1 vccd1 _2482_ sky130_fd_sc_hd__nor2_1
XANTENNA__4846__A _3763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7222__A _3925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8290__A2 _3495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8502__A0 posit_add.in2\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6277__D1 _1164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7132__A _3804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4475__B posit_add.in1\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6971__A _1414_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6730_ _1423_ _1454_ vssd1 vssd1 vccd1 vccd1 _1790_ sky130_fd_sc_hd__nor2_1
XFILLER_51_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4991_ _4114_ _4096_ vssd1 vssd1 vccd1 vccd1 _4146_ sky130_fd_sc_hd__and2b_1
XFILLER_23_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6661_ _1304_ _1711_ _1713_ vssd1 vssd1 vccd1 vccd1 _1714_ sky130_fd_sc_hd__a21oi_1
X_6592_ _1632_ _1633_ vssd1 vssd1 vccd1 vccd1 _1639_ sky130_fd_sc_hd__nand2_1
X_5612_ _0571_ _0564_ _0535_ vssd1 vssd1 vccd1 vccd1 _0585_ sky130_fd_sc_hd__mux2_1
X_8400_ _2993_ _3610_ _3611_ _3612_ _3303_ vssd1 vssd1 vccd1 vccd1 _3613_ sky130_fd_sc_hd__a311o_1
X_8331_ _3538_ _3539_ vssd1 vssd1 vccd1 vccd1 _3540_ sky130_fd_sc_hd__xor2_1
X_5543_ _0512_ _0514_ _0515_ vssd1 vssd1 vccd1 vccd1 _0516_ sky130_fd_sc_hd__mux2_1
X_8262_ _3465_ _3466_ vssd1 vssd1 vccd1 vccd1 _3468_ sky130_fd_sc_hd__and2_1
X_5474_ _0446_ vssd1 vssd1 vccd1 vccd1 _0447_ sky130_fd_sc_hd__inv_2
X_4425_ _2012_ _2111_ _2210_ posit_add.in2\[0\] vssd1 vssd1 vccd1 vccd1 _2463_ sky130_fd_sc_hd__a211o_1
X_8193_ _3391_ _3393_ vssd1 vssd1 vccd1 vccd1 _3394_ sky130_fd_sc_hd__nor2_1
X_7213_ _2302_ _2321_ vssd1 vssd1 vccd1 vccd1 _2322_ sky130_fd_sc_hd__xor2_1
X_7144_ _2118_ _2245_ _2119_ vssd1 vssd1 vccd1 vccd1 _2246_ sky130_fd_sc_hd__a21oi_1
X_4356_ _1429_ _1660_ _1682_ vssd1 vssd1 vccd1 vccd1 _1704_ sky130_fd_sc_hd__o21a_1
XFILLER_113_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7042__A _4089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7075_ _2138_ _2154_ _2169_ vssd1 vssd1 vccd1 vccd1 _2170_ sky130_fd_sc_hd__or3_1
XFILLER_86_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4287_ _0946_ vssd1 vssd1 vccd1 vccd1 _0008_ sky130_fd_sc_hd__clkbuf_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6026_ _1015_ _1022_ _1023_ vssd1 vssd1 vccd1 vccd1 _1024_ sky130_fd_sc_hd__a21bo_1
XFILLER_86_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4385__B _1275_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7977_ _3149_ _3161_ _3030_ vssd1 vssd1 vccd1 vccd1 _3162_ sky130_fd_sc_hd__o21a_1
XFILLER_14_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6928_ _1773_ _2007_ vssd1 vssd1 vccd1 vccd1 _2008_ sky130_fd_sc_hd__or2b_1
XANTENNA__4597__A1 _3189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6859_ _1930_ _1931_ vssd1 vssd1 vccd1 vccd1 _1932_ sky130_fd_sc_hd__or2_1
XFILLER_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8529_ clknet_3_5__leaf_clk _0015_ vssd1 vssd1 vccd1 vccd1 in_reg\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_6_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4588__A1 _2903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5190_ _0134_ _0162_ vssd1 vssd1 vccd1 vccd1 _0163_ sky130_fd_sc_hd__or2b_1
XFILLER_95_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7900_ _2954_ _3076_ vssd1 vssd1 vccd1 vccd1 _3077_ sky130_fd_sc_hd__and2b_1
XANTENNA__8006__A2 _0600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7831_ _2985_ _3000_ vssd1 vssd1 vccd1 vccd1 _3001_ sky130_fd_sc_hd__or2_1
XFILLER_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6206__A _0627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4974_ _4128_ _4124_ vssd1 vssd1 vccd1 vccd1 _4129_ sky130_fd_sc_hd__or2_1
XFILLER_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7762_ _2921_ _2924_ vssd1 vssd1 vccd1 vccd1 _2926_ sky130_fd_sc_hd__nand2_1
XFILLER_24_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5110__A _4228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5240__A2 _3793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6713_ _1768_ _1771_ vssd1 vssd1 vccd1 vccd1 _1772_ sky130_fd_sc_hd__or2b_1
X_7693_ _2801_ _2813_ vssd1 vssd1 vccd1 vccd1 _2850_ sky130_fd_sc_hd__and2b_1
X_6644_ _1678_ _1545_ _1685_ _1686_ vssd1 vssd1 vccd1 vccd1 _1696_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_32_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6575_ _1615_ _1617_ vssd1 vssd1 vccd1 vccd1 _1620_ sky130_fd_sc_hd__or2_1
X_8314_ _3513_ _3514_ _3522_ _0701_ vssd1 vssd1 vccd1 vccd1 _3523_ sky130_fd_sc_hd__a211o_1
X_5526_ _0331_ _0333_ vssd1 vssd1 vccd1 vccd1 _0499_ sky130_fd_sc_hd__xor2_1
XFILLER_105_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6876__A _1711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8245_ _2604_ _2515_ vssd1 vssd1 vccd1 vccd1 _3449_ sky130_fd_sc_hd__or2_1
X_5457_ _0426_ _0429_ vssd1 vssd1 vccd1 vccd1 _0430_ sky130_fd_sc_hd__or2_1
XFILLER_105_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4408_ _1968_ _2243_ _2254_ _2265_ vssd1 vssd1 vccd1 vccd1 _2276_ sky130_fd_sc_hd__o31ai_1
X_5388_ _1451_ _3830_ _0360_ _3736_ vssd1 vssd1 vccd1 vccd1 _0361_ sky130_fd_sc_hd__a211o_1
XFILLER_59_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8176_ _3374_ _3375_ _3190_ vssd1 vssd1 vccd1 vccd1 _3376_ sky130_fd_sc_hd__o21ai_1
XFILLER_101_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7127_ _2160_ _2209_ vssd1 vssd1 vccd1 vccd1 _2227_ sky130_fd_sc_hd__nor2_1
X_4339_ _1506_ _1451_ _1484_ vssd1 vssd1 vccd1 vccd1 _1517_ sky130_fd_sc_hd__nand3_2
XFILLER_101_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7058_ _2150_ vssd1 vssd1 vccd1 vccd1 _2151_ sky130_fd_sc_hd__inv_2
XFILLER_86_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4267__A0 in_reg\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6009_ _4017_ _0802_ _0773_ _0992_ vssd1 vssd1 vccd1 vccd1 _1006_ sky130_fd_sc_hd__or4_2
XFILLER_91_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5767__B1 _3792_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5020__A _3776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6192__B1 _4016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8477__S _3654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7995__A1 _1253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5865__A _3735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4690_ _3739_ vssd1 vssd1 vccd1 vccd1 _3845_ sky130_fd_sc_hd__buf_2
X_6360_ _1382_ vssd1 vssd1 vccd1 vccd1 _1383_ sky130_fd_sc_hd__buf_2
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5311_ _0277_ _0283_ vssd1 vssd1 vccd1 vccd1 _0284_ sky130_fd_sc_hd__nand2_1
X_6291_ _1154_ vssd1 vssd1 vccd1 vccd1 _1307_ sky130_fd_sc_hd__inv_2
X_8030_ _0583_ _3218_ _0519_ vssd1 vssd1 vccd1 vccd1 _3219_ sky130_fd_sc_hd__mux2_1
XFILLER_88_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5242_ _4175_ _0212_ _0214_ vssd1 vssd1 vccd1 vccd1 _0215_ sky130_fd_sc_hd__o21ai_1
X_5173_ _3802_ _3986_ vssd1 vssd1 vccd1 vccd1 _0146_ sky130_fd_sc_hd__nand2_1
XFILLER_96_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput1 io_in[0] vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__clkbuf_2
XANTENNA__4663__B _3817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7814_ _2665_ _2938_ vssd1 vssd1 vccd1 vccd1 _2983_ sky130_fd_sc_hd__and2_1
XANTENNA__5213__A2 _3883_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5775__A _3735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4957_ _4099_ _4111_ vssd1 vssd1 vccd1 vccd1 _4112_ sky130_fd_sc_hd__xnor2_1
XANTENNA__8148__D1 _1177_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7745_ _2821_ _2880_ _1297_ vssd1 vssd1 vccd1 vccd1 _2907_ sky130_fd_sc_hd__mux2_1
X_4888_ _1990_ _2320_ _2419_ _2496_ vssd1 vssd1 vccd1 vccd1 _4043_ sky130_fd_sc_hd__a31oi_2
X_7676_ _2751_ _2752_ _2830_ vssd1 vssd1 vccd1 vccd1 _2831_ sky130_fd_sc_hd__a21bo_1
X_6627_ _1382_ _1456_ vssd1 vssd1 vccd1 vccd1 _1677_ sky130_fd_sc_hd__or2_1
X_6558_ _1593_ _1600_ vssd1 vssd1 vccd1 vccd1 _1601_ sky130_fd_sc_hd__xnor2_1
XFILLER_106_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6489_ _1522_ _1523_ _1524_ vssd1 vssd1 vccd1 vccd1 _1525_ sky130_fd_sc_hd__a21oi_1
X_5509_ _0301_ _0323_ vssd1 vssd1 vccd1 vccd1 _0482_ sky130_fd_sc_hd__xor2_1
XFILLER_105_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5819__A4 _0706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8228_ _3428_ _3430_ vssd1 vssd1 vccd1 vccd1 _3431_ sky130_fd_sc_hd__or2_1
XFILLER_99_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8159_ _0601_ _3350_ _3355_ _2621_ vssd1 vssd1 vccd1 vccd1 _3357_ sky130_fd_sc_hd__a31o_1
XFILLER_87_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7729__A1 _1297_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6952__A2 _1538_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4715__A1 _3771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4715__B2 _3793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7272__B1_N _2352_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5860_ _0759_ _0848_ _0847_ _0844_ vssd1 vssd1 vccd1 vccd1 _0850_ sky130_fd_sc_hd__a211o_1
XFILLER_80_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4811_ _3947_ _3948_ vssd1 vssd1 vccd1 vccd1 _3966_ sky130_fd_sc_hd__and2_1
X_5791_ _0772_ _0774_ vssd1 vssd1 vccd1 vccd1 _0775_ sky130_fd_sc_hd__xnor2_1
XFILLER_21_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4742_ _3839_ _3895_ _3896_ vssd1 vssd1 vccd1 vccd1 _3897_ sky130_fd_sc_hd__a21o_1
XFILLER_21_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7530_ _2668_ _2669_ _0375_ vssd1 vssd1 vccd1 vccd1 _2670_ sky130_fd_sc_hd__mux2_1
X_4673_ _3735_ vssd1 vssd1 vccd1 vccd1 _3828_ sky130_fd_sc_hd__clkbuf_4
X_7461_ _2522_ _2508_ _2593_ vssd1 vssd1 vccd1 vccd1 _2594_ sky130_fd_sc_hd__a21oi_1
XFILLER_119_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6412_ _1387_ _1390_ _1439_ _1338_ vssd1 vssd1 vccd1 vccd1 _1441_ sky130_fd_sc_hd__o211a_1
X_7392_ _2516_ _2396_ _2517_ vssd1 vssd1 vccd1 vccd1 _2519_ sky130_fd_sc_hd__or3b_1
X_6343_ _1358_ _1364_ vssd1 vssd1 vccd1 vccd1 _1365_ sky130_fd_sc_hd__or2_1
X_6274_ _1281_ _1285_ vssd1 vssd1 vccd1 vccd1 _1289_ sky130_fd_sc_hd__xor2_1
XFILLER_0_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5225_ _0196_ _0175_ _0195_ vssd1 vssd1 vccd1 vccd1 _0198_ sky130_fd_sc_hd__nor3_1
X_8013_ _2521_ _2618_ vssd1 vssd1 vccd1 vccd1 _3201_ sky130_fd_sc_hd__or2_1
XFILLER_102_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5156_ _0127_ _0123_ _0125_ vssd1 vssd1 vccd1 vccd1 _0129_ sky130_fd_sc_hd__and3_1
XFILLER_29_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4674__A _3827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5087_ _4240_ _4241_ vssd1 vssd1 vccd1 vccd1 _4242_ sky130_fd_sc_hd__nand2_1
XFILLER_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6631__A1 _1400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5989_ _0983_ _0982_ _0851_ vssd1 vssd1 vccd1 vccd1 _0985_ sky130_fd_sc_hd__or3_1
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7728_ _2844_ _2886_ _2887_ _1286_ vssd1 vssd1 vccd1 vccd1 _2888_ sky130_fd_sc_hd__o211a_1
X_7659_ _2802_ _2811_ vssd1 vssd1 vccd1 vccd1 _2812_ sky130_fd_sc_hd__and2b_1
XFILLER_108_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7398__A2_N _2440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7135__A _1782_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7638__A0 _3893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5010_ _4156_ _4164_ vssd1 vssd1 vccd1 vccd1 _4165_ sky130_fd_sc_hd__xnor2_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6861__A1 _0303_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4467__A3 posit_add.in1\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6961_ _1965_ _1994_ vssd1 vssd1 vccd1 vccd1 _2044_ sky130_fd_sc_hd__xnor2_1
XFILLER_81_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5912_ _0888_ _0902_ _0903_ vssd1 vssd1 vccd1 vccd1 _0905_ sky130_fd_sc_hd__and3_1
X_6892_ _1300_ _1355_ _1809_ vssd1 vssd1 vccd1 vccd1 _1969_ sky130_fd_sc_hd__and3_1
XFILLER_81_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5843_ _3877_ _0631_ _3832_ _0633_ vssd1 vssd1 vccd1 vccd1 _0832_ sky130_fd_sc_hd__a22o_1
XFILLER_61_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8413__B _4250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8562_ clknet_3_2__leaf_clk _0048_ vssd1 vssd1 vccd1 vccd1 posit_add.in1\[5\] sky130_fd_sc_hd__dfxtp_2
XANTENNA__4927__B2 _3828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5774_ _0731_ _0756_ vssd1 vssd1 vccd1 vccd1 _0757_ sky130_fd_sc_hd__xor2_1
X_7513_ _2651_ vssd1 vssd1 vccd1 vccd1 _2652_ sky130_fd_sc_hd__clkbuf_4
X_8493_ _3685_ vssd1 vssd1 vccd1 vccd1 _0064_ sky130_fd_sc_hd__clkbuf_1
X_4725_ _3875_ _3879_ vssd1 vssd1 vccd1 vccd1 _3880_ sky130_fd_sc_hd__xor2_1
X_4656_ _3808_ _3810_ _2485_ vssd1 vssd1 vccd1 vccd1 _3811_ sky130_fd_sc_hd__a21o_1
X_7444_ _2480_ _2513_ _2569_ vssd1 vssd1 vccd1 vccd1 _2576_ sky130_fd_sc_hd__mux2_1
X_4587_ _3339_ _3349_ _2859_ _3360_ vssd1 vssd1 vccd1 vccd1 _3742_ sky130_fd_sc_hd__o211a_1
X_7375_ _2335_ _2470_ vssd1 vssd1 vccd1 vccd1 _2500_ sky130_fd_sc_hd__nand2_1
X_6326_ _1000_ _1345_ vssd1 vssd1 vccd1 vccd1 _1346_ sky130_fd_sc_hd__and2b_1
XFILLER_89_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6257_ _1263_ _1265_ _1269_ vssd1 vssd1 vccd1 vccd1 _1270_ sky130_fd_sc_hd__a21o_1
XFILLER_88_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6188_ _1168_ _1097_ vssd1 vssd1 vccd1 vccd1 _1195_ sky130_fd_sc_hd__or2b_1
X_5208_ _0180_ _0149_ vssd1 vssd1 vccd1 vccd1 _0181_ sky130_fd_sc_hd__nor2_1
X_5139_ _0111_ vssd1 vssd1 vccd1 vccd1 _0112_ sky130_fd_sc_hd__clkbuf_4
XFILLER_69_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4579__A _3729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8348__A1 _1330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4510_ _2969_ _2980_ _3199_ _3381_ vssd1 vssd1 vccd1 vccd1 _3392_ sky130_fd_sc_hd__o211a_1
XFILLER_7_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5490_ _0457_ _0458_ _0461_ vssd1 vssd1 vccd1 vccd1 _0463_ sky130_fd_sc_hd__a21bo_1
X_4441_ posit_add.in1\[8\] _2628_ vssd1 vssd1 vccd1 vccd1 _2639_ sky130_fd_sc_hd__xor2_2
XFILLER_7_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7160_ _1761_ _1767_ vssd1 vssd1 vccd1 vccd1 _2263_ sky130_fd_sc_hd__and2b_1
X_6111_ _1108_ _1111_ vssd1 vssd1 vccd1 vccd1 _1113_ sky130_fd_sc_hd__nand2_1
X_4372_ posit_add.in2\[3\] _1825_ vssd1 vssd1 vccd1 vccd1 _1880_ sky130_fd_sc_hd__xor2_1
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7091_ _4089_ _2158_ _2164_ vssd1 vssd1 vccd1 vccd1 _2187_ sky130_fd_sc_hd__a21oi_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6042_ _1039_ _1040_ vssd1 vssd1 vccd1 vccd1 _1041_ sky130_fd_sc_hd__nor2_1
XFILLER_86_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7993_ _3173_ _3179_ _3030_ vssd1 vssd1 vccd1 vccd1 _3180_ sky130_fd_sc_hd__mux2_1
XANTENNA__7739__S _1297_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6944_ _2024_ _2025_ vssd1 vssd1 vccd1 vccd1 _2026_ sky130_fd_sc_hd__xor2_1
XFILLER_81_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6875_ _1257_ _1302_ vssd1 vssd1 vccd1 vccd1 _1950_ sky130_fd_sc_hd__nand2_2
X_5826_ _2529_ _0812_ vssd1 vssd1 vccd1 vccd1 _0813_ sky130_fd_sc_hd__xnor2_1
XFILLER_22_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6879__A _1384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5757_ _2507_ _3815_ _0670_ _3866_ vssd1 vssd1 vccd1 vccd1 _0739_ sky130_fd_sc_hd__a211oi_1
X_8545_ clknet_3_2__leaf_clk _0031_ vssd1 vssd1 vccd1 vccd1 out_reg\[11\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__5783__A _3901_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8476_ _3673_ vssd1 vssd1 vccd1 vccd1 _0057_ sky130_fd_sc_hd__clkbuf_1
X_4708_ _3759_ _3760_ vssd1 vssd1 vccd1 vccd1 _3863_ sky130_fd_sc_hd__and2_1
X_5688_ _0613_ _0663_ vssd1 vssd1 vccd1 vccd1 _0664_ sky130_fd_sc_hd__nor2_1
X_7427_ _2203_ _2542_ _2550_ _2556_ vssd1 vssd1 vccd1 vccd1 _2557_ sky130_fd_sc_hd__a211o_1
XANTENNA__4399__A _1781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4639_ _3721_ _3788_ vssd1 vssd1 vccd1 vccd1 _3794_ sky130_fd_sc_hd__nand2_1
XFILLER_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7358_ _2426_ _2427_ vssd1 vssd1 vccd1 vccd1 _2481_ sky130_fd_sc_hd__nand2_1
XFILLER_103_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6309_ _1324_ _1326_ vssd1 vssd1 vccd1 vccd1 _1327_ sky130_fd_sc_hd__nor2_2
XFILLER_89_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8275__B1 _1308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7289_ _2403_ _2404_ vssd1 vssd1 vccd1 vccd1 _2405_ sky130_fd_sc_hd__xnor2_2
XFILLER_77_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4846__B _3817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7222__B _3828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4862__A _4016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6971__B _3804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4772__A _3924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4990_ _4140_ _4143_ _4144_ vssd1 vssd1 vccd1 vccd1 _4145_ sky130_fd_sc_hd__a21o_1
XFILLER_51_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6660_ _1712_ _1226_ vssd1 vssd1 vccd1 vccd1 _1713_ sky130_fd_sc_hd__or2_1
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6752__B1 _4228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6591_ _1632_ _1633_ _1636_ vssd1 vssd1 vccd1 vccd1 _1637_ sky130_fd_sc_hd__a21bo_1
X_5611_ _0531_ _0524_ _0494_ vssd1 vssd1 vccd1 vccd1 _0584_ sky130_fd_sc_hd__mux2_1
X_8330_ _3460_ _3478_ _3511_ _3226_ vssd1 vssd1 vccd1 vccd1 _3539_ sky130_fd_sc_hd__a31o_1
X_5542_ _0480_ vssd1 vssd1 vccd1 vccd1 _0515_ sky130_fd_sc_hd__clkbuf_4
XFILLER_117_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8261_ _3429_ _3464_ _3431_ vssd1 vssd1 vccd1 vccd1 _3466_ sky130_fd_sc_hd__o21ai_1
X_5473_ _0397_ _0443_ _0444_ _0445_ vssd1 vssd1 vccd1 vccd1 _0446_ sky130_fd_sc_hd__or4_2
X_4424_ _2441_ vssd1 vssd1 vccd1 vccd1 _2452_ sky130_fd_sc_hd__buf_4
X_8192_ _3388_ _3390_ vssd1 vssd1 vccd1 vccd1 _3393_ sky130_fd_sc_hd__nor2_1
X_7212_ _2273_ _2319_ vssd1 vssd1 vccd1 vccd1 _2321_ sky130_fd_sc_hd__nand2_1
X_7143_ _2121_ _2149_ vssd1 vssd1 vccd1 vccd1 _2245_ sky130_fd_sc_hd__or2_1
X_4355_ _1506_ _1660_ _1682_ vssd1 vssd1 vccd1 vccd1 _1693_ sky130_fd_sc_hd__a21oi_1
X_7074_ _2128_ _2129_ _2159_ _2168_ vssd1 vssd1 vccd1 vccd1 _2169_ sky130_fd_sc_hd__o31a_1
XFILLER_59_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7042__B _1676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4286_ in_reg\[4\] in_reg\[5\] _0830_ vssd1 vssd1 vccd1 vccd1 _0946_ sky130_fd_sc_hd__mux2_1
XFILLER_58_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6025_ _1006_ _1018_ vssd1 vssd1 vccd1 vccd1 _1023_ sky130_fd_sc_hd__nand2_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7976_ _3152_ _3154_ _3158_ _3160_ vssd1 vssd1 vccd1 vccd1 _3161_ sky130_fd_sc_hd__or4_1
XFILLER_14_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6927_ _1900_ _2004_ _2006_ vssd1 vssd1 vccd1 vccd1 _2007_ sky130_fd_sc_hd__a21o_1
X_6858_ _1428_ _1718_ vssd1 vssd1 vccd1 vccd1 _1931_ sky130_fd_sc_hd__or2_1
X_5809_ _3802_ _0762_ vssd1 vssd1 vccd1 vccd1 _0794_ sky130_fd_sc_hd__nand2_1
XFILLER_10_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8528_ clknet_3_5__leaf_clk _0014_ vssd1 vssd1 vccd1 vccd1 in_reg\[11\] sky130_fd_sc_hd__dfxtp_1
X_6789_ _1852_ _1854_ vssd1 vssd1 vccd1 vccd1 _1855_ sky130_fd_sc_hd__nor2_1
XANTENNA__6402__A _1383_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5018__A _3881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8459_ in_reg\[6\] posit_add.in1\[6\] _3655_ vssd1 vssd1 vccd1 vccd1 _3663_ sky130_fd_sc_hd__mux2_1
XFILLER_2_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7462__A1 _2382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7830_ _2984_ _2945_ _2982_ vssd1 vssd1 vccd1 vccd1 _3000_ sky130_fd_sc_hd__nor3_1
XFILLER_64_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4973_ _4127_ vssd1 vssd1 vccd1 vccd1 _4128_ sky130_fd_sc_hd__inv_2
XFILLER_51_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7761_ _2923_ vssd1 vssd1 vccd1 vccd1 _2924_ sky130_fd_sc_hd__inv_2
XFILLER_51_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6712_ _1765_ _1769_ vssd1 vssd1 vccd1 vccd1 _1771_ sky130_fd_sc_hd__xnor2_1
X_7692_ _2790_ _2816_ vssd1 vssd1 vccd1 vccd1 _2849_ sky130_fd_sc_hd__or2_1
XANTENNA__5110__B _4250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6643_ _1692_ _1694_ vssd1 vssd1 vccd1 vccd1 _1695_ sky130_fd_sc_hd__xnor2_2
XFILLER_20_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7318__A _2416_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6574_ _1584_ _1618_ vssd1 vssd1 vccd1 vccd1 _1619_ sky130_fd_sc_hd__xnor2_1
X_8313_ _3515_ _3519_ _3521_ vssd1 vssd1 vccd1 vccd1 _3522_ sky130_fd_sc_hd__o21a_1
X_5525_ _0330_ _0497_ vssd1 vssd1 vccd1 vccd1 _0498_ sky130_fd_sc_hd__nor2_1
XFILLER_118_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8244_ _3421_ _3415_ _0601_ vssd1 vssd1 vccd1 vccd1 _3448_ sky130_fd_sc_hd__o21a_1
X_5456_ _3488_ _0428_ _0344_ vssd1 vssd1 vccd1 vccd1 _0429_ sky130_fd_sc_hd__mux2_1
XANTENNA__6876__B _0121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4407_ _1957_ _1924_ vssd1 vssd1 vccd1 vccd1 _2265_ sky130_fd_sc_hd__nor2_1
XFILLER_99_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5387_ _3830_ _0359_ vssd1 vssd1 vccd1 vccd1 _0360_ sky130_fd_sc_hd__nor2_1
X_8175_ _3182_ _3334_ vssd1 vssd1 vccd1 vccd1 _3375_ sky130_fd_sc_hd__and2_1
XFILLER_113_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7126_ _1782_ _2079_ _2225_ vssd1 vssd1 vccd1 vccd1 _2226_ sky130_fd_sc_hd__a21oi_1
X_4338_ _1429_ vssd1 vssd1 vccd1 vccd1 _1506_ sky130_fd_sc_hd__buf_2
XFILLER_115_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7057_ _2121_ _2149_ vssd1 vssd1 vccd1 vccd1 _2150_ sky130_fd_sc_hd__xnor2_1
X_4269_ in_reg\[7\] cmd\[7\] _0712_ vssd1 vssd1 vccd1 vccd1 _0765_ sky130_fd_sc_hd__mux2_1
XANTENNA__4267__A1 cmd\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input2_A io_in[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6008_ _0634_ _0994_ _0996_ _0997_ vssd1 vssd1 vccd1 vccd1 _1005_ sky130_fd_sc_hd__a22o_1
XFILLER_27_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5767__A1 _2507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7959_ _3140_ _3141_ _3065_ vssd1 vssd1 vccd1 vccd1 _3142_ sky130_fd_sc_hd__mux2_1
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5020__B _3878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5211__A _4017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5758__A1 _3866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6290_ _1157_ _1191_ _1226_ _1305_ vssd1 vssd1 vccd1 vccd1 _1306_ sky130_fd_sc_hd__or4_2
X_5310_ _4045_ _0121_ _0276_ vssd1 vssd1 vccd1 vccd1 _0283_ sky130_fd_sc_hd__a21o_1
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5241_ _0124_ _3875_ _0213_ vssd1 vssd1 vccd1 vccd1 _0214_ sky130_fd_sc_hd__o21ba_1
X_5172_ _0109_ _0144_ vssd1 vssd1 vccd1 vccd1 _0145_ sky130_fd_sc_hd__nand2_1
XFILLER_28_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput2 io_in[1] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_1
XFILLER_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7813_ _2960_ _2979_ _2981_ vssd1 vssd1 vccd1 vccd1 _2982_ sky130_fd_sc_hd__o21a_1
XFILLER_36_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7744_ _2829_ _2905_ vssd1 vssd1 vccd1 vccd1 _2906_ sky130_fd_sc_hd__xnor2_2
XFILLER_51_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4956_ _4100_ _4110_ vssd1 vssd1 vccd1 vccd1 _4111_ sky130_fd_sc_hd__and2b_1
X_4887_ _4040_ _4041_ vssd1 vssd1 vccd1 vccd1 _4042_ sky130_fd_sc_hd__nand2_1
XFILLER_20_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7675_ _2823_ _2829_ vssd1 vssd1 vccd1 vccd1 _2830_ sky130_fd_sc_hd__or2b_1
X_6626_ _3703_ vssd1 vssd1 vccd1 vccd1 _1676_ sky130_fd_sc_hd__buf_4
X_6557_ _1599_ _4232_ vssd1 vssd1 vccd1 vccd1 _1600_ sky130_fd_sc_hd__or2_1
X_5508_ _0471_ _0477_ _0480_ vssd1 vssd1 vccd1 vccd1 _0481_ sky130_fd_sc_hd__mux2_1
XFILLER_105_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6488_ _1507_ _1521_ vssd1 vssd1 vccd1 vccd1 _1524_ sky130_fd_sc_hd__and2b_1
XFILLER_106_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8227_ _0521_ _0517_ _3429_ vssd1 vssd1 vccd1 vccd1 _3430_ sky130_fd_sc_hd__a21o_1
X_5439_ _3772_ _0406_ _0411_ vssd1 vssd1 vccd1 vccd1 _0412_ sky130_fd_sc_hd__mux2_1
XFILLER_105_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8158_ _1330_ _3350_ _3355_ vssd1 vssd1 vccd1 vccd1 _3356_ sky130_fd_sc_hd__a21oi_1
X_7109_ _2192_ _2193_ vssd1 vssd1 vccd1 vccd1 _2207_ sky130_fd_sc_hd__xor2_1
XFILLER_59_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8089_ out_reg\[2\] _3197_ _3282_ vssd1 vssd1 vccd1 vccd1 _3283_ sky130_fd_sc_hd__a21oi_1
XFILLER_47_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6127__A _0627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_718 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4412__A1 _1913_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4715__A2 _3840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5206__A _3800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4651__A1 _3800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5876__A _3892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4810_ _3727_ _3962_ vssd1 vssd1 vccd1 vccd1 _3965_ sky130_fd_sc_hd__xnor2_1
XFILLER_33_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5790_ _3700_ _0773_ vssd1 vssd1 vccd1 vccd1 _0774_ sky130_fd_sc_hd__nor2_1
XFILLER_61_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4741_ _3893_ _3832_ _3838_ _3894_ vssd1 vssd1 vccd1 vccd1 _3896_ sky130_fd_sc_hd__and4_1
XFILLER_14_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4672_ _3825_ _3826_ _3594_ vssd1 vssd1 vccd1 vccd1 _3827_ sky130_fd_sc_hd__mux2_4
X_7460_ _2450_ _2475_ _2478_ vssd1 vssd1 vccd1 vccd1 _2593_ sky130_fd_sc_hd__and3_1
X_6411_ _0795_ _0993_ _1388_ vssd1 vssd1 vccd1 vccd1 _1439_ sky130_fd_sc_hd__a21o_1
X_7391_ _2402_ _2405_ _2406_ vssd1 vssd1 vccd1 vccd1 _2517_ sky130_fd_sc_hd__or3_1
X_6342_ _1359_ _1362_ vssd1 vssd1 vccd1 vccd1 _1364_ sky130_fd_sc_hd__xor2_1
XFILLER_103_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6273_ _0762_ _1164_ vssd1 vssd1 vccd1 vccd1 _1288_ sky130_fd_sc_hd__and2_1
XFILLER_88_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5224_ _0175_ _0195_ _0196_ vssd1 vssd1 vccd1 vccd1 _0197_ sky130_fd_sc_hd__o21a_1
X_8012_ _2521_ _3198_ vssd1 vssd1 vccd1 vccd1 _3200_ sky130_fd_sc_hd__nand2_2
XFILLER_69_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5155_ _0123_ _0125_ _0127_ vssd1 vssd1 vccd1 vccd1 _0128_ sky130_fd_sc_hd__a21oi_1
XFILLER_110_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4674__B _3828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5086_ _4238_ _4239_ vssd1 vssd1 vccd1 vccd1 _4241_ sky130_fd_sc_hd__nand2_1
XFILLER_84_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6631__A2 _1676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5988_ _0982_ _0851_ _0983_ vssd1 vssd1 vccd1 vccd1 _0984_ sky130_fd_sc_hd__o21a_1
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4690__A _3739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4939_ _4071_ _4072_ _4088_ _4093_ vssd1 vssd1 vccd1 vccd1 _4094_ sky130_fd_sc_hd__o31a_1
X_7727_ _2743_ _2797_ _2838_ vssd1 vssd1 vccd1 vccd1 _2887_ sky130_fd_sc_hd__a21o_1
X_7658_ _2729_ _2720_ _2810_ vssd1 vssd1 vccd1 vccd1 _2811_ sky130_fd_sc_hd__o21bai_1
X_6609_ _1384_ _1423_ vssd1 vssd1 vccd1 vccd1 _1657_ sky130_fd_sc_hd__nor2_1
XFILLER_106_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7589_ _2712_ _2734_ vssd1 vssd1 vccd1 vccd1 _2735_ sky130_fd_sc_hd__or2_1
XFILLER_118_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4865__A _3701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7638__A1 _3868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6861__A2 _1718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6960_ _2040_ _2041_ _2042_ _2033_ vssd1 vssd1 vccd1 vccd1 _2043_ sky130_fd_sc_hd__a22o_1
XFILLER_66_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5911_ _0885_ _0887_ _0886_ vssd1 vssd1 vccd1 vccd1 _0903_ sky130_fd_sc_hd__a21o_1
X_6891_ _1509_ _3930_ vssd1 vssd1 vccd1 vccd1 _1967_ sky130_fd_sc_hd__or2_1
X_5842_ _0627_ _3770_ _3738_ _0631_ vssd1 vssd1 vccd1 vccd1 _0831_ sky130_fd_sc_hd__or4b_1
XFILLER_61_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5773_ _3924_ _0755_ vssd1 vssd1 vccd1 vccd1 _0756_ sky130_fd_sc_hd__nor2_1
X_8561_ clknet_3_3__leaf_clk _0047_ vssd1 vssd1 vccd1 vccd1 posit_add.in1\[4\] sky130_fd_sc_hd__dfxtp_2
XFILLER_61_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4927__A2 _3817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4724_ _3878_ _3855_ vssd1 vssd1 vccd1 vccd1 _3879_ sky130_fd_sc_hd__nand2_1
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7512_ _2649_ vssd1 vssd1 vccd1 vccd1 _2651_ sky130_fd_sc_hd__clkbuf_4
X_8492_ posit_add.in2\[5\] in_reg\[5\] _3677_ vssd1 vssd1 vccd1 vccd1 _3685_ sky130_fd_sc_hd__mux2_1
XFILLER_30_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4655_ _1858_ _2452_ _3809_ _2309_ vssd1 vssd1 vccd1 vccd1 _3810_ sky130_fd_sc_hd__o211ai_2
X_7443_ _2541_ _2574_ _2522_ vssd1 vssd1 vccd1 vccd1 _2575_ sky130_fd_sc_hd__mux2_1
X_4586_ _2826_ _3318_ _3740_ _3446_ vssd1 vssd1 vccd1 vccd1 _3741_ sky130_fd_sc_hd__a211o_1
X_7374_ _2412_ _2498_ vssd1 vssd1 vccd1 vccd1 _2499_ sky130_fd_sc_hd__or2_1
X_6325_ _1343_ _1344_ vssd1 vssd1 vccd1 vccd1 _1345_ sky130_fd_sc_hd__xnor2_1
XFILLER_115_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6256_ _1266_ _1267_ _1268_ vssd1 vssd1 vccd1 vccd1 _1269_ sky130_fd_sc_hd__a21bo_1
X_6187_ _1192_ _1193_ vssd1 vssd1 vccd1 vccd1 _1194_ sky130_fd_sc_hd__xnor2_1
XFILLER_97_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5207_ _0150_ vssd1 vssd1 vccd1 vccd1 _0180_ sky130_fd_sc_hd__inv_2
X_5138_ _3716_ _3711_ _3710_ _3690_ vssd1 vssd1 vccd1 vccd1 _0111_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_57_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xposit_unit_5 vssd1 vssd1 vccd1 vccd1 posit_unit_5/HI io_out[0] sky130_fd_sc_hd__conb_1
X_5069_ _4220_ _4223_ vssd1 vssd1 vccd1 vccd1 _4224_ sky130_fd_sc_hd__nand2_1
XFILLER_45_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7859__A1 _2999_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4440_ _1242_ _2617_ vssd1 vssd1 vccd1 vccd1 _2628_ sky130_fd_sc_hd__nand2_1
X_6110_ _1108_ _1111_ vssd1 vssd1 vccd1 vccd1 _1112_ sky130_fd_sc_hd__nor2_1
X_4371_ _1506_ _1858_ vssd1 vssd1 vccd1 vccd1 _1869_ sky130_fd_sc_hd__nand2_1
X_7090_ _4089_ _1813_ _2156_ vssd1 vssd1 vccd1 vccd1 _2186_ sky130_fd_sc_hd__a21boi_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6041_ _1006_ _1038_ vssd1 vssd1 vccd1 vccd1 _1040_ sky130_fd_sc_hd__and2_1
XFILLER_86_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4845__A1 _3827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7992_ _3174_ _3177_ _3021_ vssd1 vssd1 vccd1 vccd1 _3179_ sky130_fd_sc_hd__mux2_1
XFILLER_27_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6943_ _1975_ _1977_ vssd1 vssd1 vccd1 vccd1 _2025_ sky130_fd_sc_hd__xor2_1
XFILLER_93_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6225__A _0795_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6874_ _1947_ _1901_ vssd1 vssd1 vccd1 vccd1 _1949_ sky130_fd_sc_hd__xor2_1
XFILLER_34_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5825_ _0764_ _0769_ _0811_ vssd1 vssd1 vccd1 vccd1 _0812_ sky130_fd_sc_hd__a21oi_1
XFILLER_34_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6879__B _1718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5756_ _0365_ _3900_ _2518_ vssd1 vssd1 vccd1 vccd1 _0738_ sky130_fd_sc_hd__or3_1
X_8544_ clknet_3_3__leaf_clk _0030_ vssd1 vssd1 vccd1 vccd1 out_reg\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_22_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5687_ _0616_ _0609_ vssd1 vssd1 vccd1 vccd1 _0663_ sky130_fd_sc_hd__nand2_1
X_4707_ _3860_ _3861_ vssd1 vssd1 vccd1 vccd1 _3862_ sky130_fd_sc_hd__and2_1
X_8475_ in_reg\[14\] posit_add.in1\[14\] _3654_ vssd1 vssd1 vccd1 vccd1 _3673_ sky130_fd_sc_hd__mux2_1
X_7426_ _2554_ _2555_ _2416_ vssd1 vssd1 vccd1 vccd1 _2556_ sky130_fd_sc_hd__mux2_1
X_4638_ _3792_ vssd1 vssd1 vccd1 vccd1 _3793_ sky130_fd_sc_hd__buf_2
XFILLER_104_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4569_ _2969_ _3530_ _3723_ _3167_ _3488_ vssd1 vssd1 vccd1 vccd1 _3724_ sky130_fd_sc_hd__o2111a_1
XFILLER_1_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7357_ _2451_ _2467_ _2479_ vssd1 vssd1 vccd1 vccd1 _2480_ sky130_fd_sc_hd__a21oi_1
X_6308_ _1143_ _1152_ _1325_ vssd1 vssd1 vccd1 vccd1 _1326_ sky130_fd_sc_hd__a21boi_1
XFILLER_103_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5089__A1 _3800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7288_ _2347_ _2354_ vssd1 vssd1 vccd1 vccd1 _2404_ sky130_fd_sc_hd__xor2_2
X_6239_ _1247_ _1248_ vssd1 vssd1 vccd1 vccd1 _1250_ sky130_fd_sc_hd__nand2_1
XFILLER_103_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4836__A1 _3893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7222__C _3771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5304__A _2540_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6589__A1 _0080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6135__A _1128_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5261__A1 _3800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6513__A1 _1420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4772__B _3702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6590_ _1634_ _1635_ vssd1 vssd1 vccd1 vccd1 _1636_ sky130_fd_sc_hd__and2_1
X_5610_ _0567_ _0559_ _0535_ vssd1 vssd1 vccd1 vccd1 _0583_ sky130_fd_sc_hd__mux2_1
X_5541_ _0445_ _0510_ _0513_ vssd1 vssd1 vccd1 vccd1 _0514_ sky130_fd_sc_hd__o21ai_1
XFILLER_117_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8260_ _3431_ _3464_ vssd1 vssd1 vccd1 vccd1 _3465_ sky130_fd_sc_hd__or2_1
XFILLER_117_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5472_ _0390_ _0337_ vssd1 vssd1 vccd1 vccd1 _0445_ sky130_fd_sc_hd__xnor2_2
X_7211_ _4250_ _3989_ vssd1 vssd1 vccd1 vccd1 _2319_ sky130_fd_sc_hd__nor2_4
X_4423_ _2012_ _2111_ _2210_ vssd1 vssd1 vccd1 vccd1 _2441_ sky130_fd_sc_hd__a21oi_1
X_8191_ _3388_ _3390_ vssd1 vssd1 vccd1 vccd1 _3391_ sky130_fd_sc_hd__and2_1
X_7142_ _2181_ _2241_ _2242_ vssd1 vssd1 vccd1 vccd1 _2244_ sky130_fd_sc_hd__a21o_1
X_4354_ posit_add.in2\[7\] _1671_ vssd1 vssd1 vccd1 vccd1 _1682_ sky130_fd_sc_hd__xor2_4
XFILLER_98_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7073_ _2163_ _2167_ vssd1 vssd1 vccd1 vccd1 _2168_ sky130_fd_sc_hd__or2b_1
XANTENNA__8419__B _3630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6024_ _1006_ _1018_ _1021_ vssd1 vssd1 vccd1 vccd1 _1022_ sky130_fd_sc_hd__a21oi_1
XFILLER_86_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4285_ _0925_ vssd1 vssd1 vccd1 vccd1 _0007_ sky130_fd_sc_hd__clkbuf_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7042__C _1537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6881__C _1531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7975_ _3155_ _3159_ _3025_ vssd1 vssd1 vccd1 vccd1 _3160_ sky130_fd_sc_hd__mux2_1
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6926_ _1838_ _2005_ _1898_ vssd1 vssd1 vccd1 vccd1 _2006_ sky130_fd_sc_hd__a21oi_1
XFILLER_82_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6857_ _1420_ _1538_ vssd1 vssd1 vccd1 vccd1 _1930_ sky130_fd_sc_hd__or2_1
X_5808_ _0715_ _0767_ _0792_ vssd1 vssd1 vccd1 vccd1 _0793_ sky130_fd_sc_hd__o21a_1
X_6788_ _1853_ _1785_ vssd1 vssd1 vccd1 vccd1 _1854_ sky130_fd_sc_hd__xnor2_2
XFILLER_50_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5739_ _3700_ _0676_ vssd1 vssd1 vccd1 vccd1 _0720_ sky130_fd_sc_hd__nor2_1
X_8527_ clknet_3_5__leaf_clk _0013_ vssd1 vssd1 vccd1 vccd1 in_reg\[10\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__6402__B _1428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8496__A1 in_reg\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8458_ _3662_ vssd1 vssd1 vccd1 vccd1 _0048_ sky130_fd_sc_hd__clkbuf_1
X_8389_ _1220_ _3601_ vssd1 vssd1 vccd1 vccd1 _0033_ sky130_fd_sc_hd__nor2_1
X_7409_ _2534_ vssd1 vssd1 vccd1 vccd1 _2537_ sky130_fd_sc_hd__inv_2
XFILLER_89_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7424__A _2536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8239__A1 _3182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4972_ _4119_ _4118_ _4121_ vssd1 vssd1 vccd1 vccd1 _4127_ sky130_fd_sc_hd__or3_1
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7760_ _2850_ _2922_ vssd1 vssd1 vccd1 vccd1 _2923_ sky130_fd_sc_hd__xor2_2
X_6711_ _1530_ _1582_ vssd1 vssd1 vccd1 vccd1 _1769_ sky130_fd_sc_hd__xor2_1
X_7691_ _2846_ vssd1 vssd1 vccd1 vccd1 _2847_ sky130_fd_sc_hd__inv_2
X_6642_ _1566_ _1567_ vssd1 vssd1 vccd1 vccd1 _1694_ sky130_fd_sc_hd__xor2_2
XFILLER_20_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7318__B _2412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6573_ _1615_ _1617_ vssd1 vssd1 vccd1 vccd1 _1618_ sky130_fd_sc_hd__xor2_1
X_8312_ _3515_ _3519_ _0599_ vssd1 vssd1 vccd1 vccd1 _3521_ sky130_fd_sc_hd__a21oi_1
XANTENNA__5119__A _4210_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5524_ _0329_ _0328_ vssd1 vssd1 vccd1 vccd1 _0497_ sky130_fd_sc_hd__and2b_1
X_8243_ _3445_ _3447_ _0635_ vssd1 vssd1 vccd1 vccd1 _0027_ sky130_fd_sc_hd__a21oi_1
X_5455_ _0427_ vssd1 vssd1 vccd1 vccd1 _0428_ sky130_fd_sc_hd__clkinv_2
XANTENNA__6876__C _1950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4406_ posit_add.in2\[0\] _1781_ _1803_ _2034_ vssd1 vssd1 vccd1 vccd1 _2254_ sky130_fd_sc_hd__and4_1
XFILLER_59_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8174_ _3329_ _3373_ vssd1 vssd1 vccd1 vccd1 _3374_ sky130_fd_sc_hd__xnor2_1
XFILLER_113_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7125_ _2214_ _2224_ vssd1 vssd1 vccd1 vccd1 _2225_ sky130_fd_sc_hd__nor2_1
X_5386_ _1583_ _3635_ _0358_ vssd1 vssd1 vccd1 vccd1 _0359_ sky130_fd_sc_hd__o21ai_1
XFILLER_99_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4337_ _1429_ _1451_ _1484_ vssd1 vssd1 vccd1 vccd1 _1495_ sky130_fd_sc_hd__or3_2
XFILLER_115_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6892__B _1355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7056_ _2123_ _2147_ _2148_ vssd1 vssd1 vccd1 vccd1 _2149_ sky130_fd_sc_hd__a21oi_1
X_4268_ _0744_ vssd1 vssd1 vccd1 vccd1 _0001_ sky130_fd_sc_hd__clkbuf_1
X_6007_ _1003_ vssd1 vssd1 vccd1 vccd1 _1004_ sky130_fd_sc_hd__buf_2
XFILLER_74_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_451 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5767__A2 _3815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7958_ _3009_ _3008_ _2999_ vssd1 vssd1 vccd1 vccd1 _3141_ sky130_fd_sc_hd__mux2_1
X_6909_ _1985_ _1986_ vssd1 vssd1 vccd1 vccd1 _1987_ sky130_fd_sc_hd__xor2_1
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5020__C _3855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7889_ _3006_ vssd1 vssd1 vccd1 vccd1 _3065_ sky130_fd_sc_hd__clkbuf_4
XFILLER_10_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8469__A1 posit_add.in1\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5211__B _3930_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5240_ _3827_ _3793_ _3750_ _3763_ vssd1 vssd1 vccd1 vccd1 _0213_ sky130_fd_sc_hd__o22a_1
XFILLER_102_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5171_ _3701_ _4037_ _0108_ vssd1 vssd1 vccd1 vccd1 _0144_ sky130_fd_sc_hd__o21ai_1
XFILLER_83_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7601__B _2702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput3 io_in[2] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__clkbuf_1
XFILLER_49_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7812_ _2942_ _2944_ vssd1 vssd1 vccd1 vccd1 _2981_ sky130_fd_sc_hd__xnor2_1
XFILLER_101_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4955_ _4104_ _4108_ _4109_ vssd1 vssd1 vccd1 vccd1 _4110_ sky130_fd_sc_hd__a21boi_1
X_7743_ _2823_ _2883_ _1297_ vssd1 vssd1 vccd1 vccd1 _2905_ sky130_fd_sc_hd__mux2_1
XFILLER_24_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4886_ _4039_ _3985_ vssd1 vssd1 vccd1 vccd1 _4041_ sky130_fd_sc_hd__or2b_1
X_7674_ _2825_ _2828_ vssd1 vssd1 vccd1 vccd1 _2829_ sky130_fd_sc_hd__nand2_1
XFILLER_32_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6625_ _1659_ _1674_ vssd1 vssd1 vccd1 vccd1 _1675_ sky130_fd_sc_hd__xor2_1
X_6556_ _1353_ _1354_ vssd1 vssd1 vccd1 vccd1 _1599_ sky130_fd_sc_hd__nand2_1
XFILLER_20_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5507_ _0468_ _0479_ vssd1 vssd1 vccd1 vccd1 _0480_ sky130_fd_sc_hd__nor2_4
XFILLER_105_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6487_ _1457_ _1459_ vssd1 vssd1 vccd1 vccd1 _1523_ sky130_fd_sc_hd__xnor2_1
XANTENNA__5134__B1 _0105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8226_ _0440_ _0521_ vssd1 vssd1 vccd1 vccd1 _3429_ sky130_fd_sc_hd__nor2_2
XFILLER_105_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5438_ _0407_ _0410_ _2980_ vssd1 vssd1 vccd1 vccd1 _0411_ sky130_fd_sc_hd__a21o_1
XFILLER_114_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8157_ _3351_ _3354_ vssd1 vssd1 vccd1 vccd1 _3355_ sky130_fd_sc_hd__xnor2_2
XANTENNA__7999__A _1275_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5369_ _1781_ _2452_ vssd1 vssd1 vccd1 vccd1 _0342_ sky130_fd_sc_hd__xnor2_1
X_7108_ _2196_ _2205_ vssd1 vssd1 vccd1 vccd1 _2206_ sky130_fd_sc_hd__or2_1
X_8088_ _3256_ _3270_ _3280_ _3281_ vssd1 vssd1 vccd1 vccd1 _3282_ sky130_fd_sc_hd__o31a_1
X_7039_ _2126_ _2128_ _2129_ vssd1 vssd1 vccd1 vccd1 _2130_ sky130_fd_sc_hd__nor3_1
XFILLER_87_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5312__A _4228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6937__A1 _1665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7239__A _2349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5206__B _4037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4651__A2 _3703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4740_ _3893_ _3894_ vssd1 vssd1 vccd1 vccd1 _3895_ sky130_fd_sc_hd__nand2_1
XFILLER_14_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4671_ _3541_ _3562_ _3520_ vssd1 vssd1 vccd1 vccd1 _3826_ sky130_fd_sc_hd__a21o_1
X_6410_ _1378_ _1380_ _1397_ _1373_ vssd1 vssd1 vccd1 vccd1 _1438_ sky130_fd_sc_hd__a211o_1
X_7390_ _2399_ _2401_ vssd1 vssd1 vccd1 vccd1 _2516_ sky130_fd_sc_hd__nand2_1
X_6341_ _0994_ _1361_ vssd1 vssd1 vccd1 vccd1 _1362_ sky130_fd_sc_hd__nand2_1
XFILLER_115_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6272_ _1281_ _1285_ vssd1 vssd1 vccd1 vccd1 _1287_ sky130_fd_sc_hd__nand2_1
XFILLER_103_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5223_ _0155_ _0141_ vssd1 vssd1 vccd1 vccd1 _0196_ sky130_fd_sc_hd__xnor2_1
X_8011_ _2611_ _2615_ _2616_ _2609_ vssd1 vssd1 vccd1 vccd1 _3198_ sky130_fd_sc_hd__o211a_1
XFILLER_102_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5154_ _4246_ _0126_ vssd1 vssd1 vccd1 vccd1 _0127_ sky130_fd_sc_hd__or2_1
XFILLER_111_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5132__A _4017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5085_ _4238_ _4239_ vssd1 vssd1 vccd1 vccd1 _4240_ sky130_fd_sc_hd__or2_1
XFILLER_112_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5987_ _0789_ _0785_ vssd1 vssd1 vccd1 vccd1 _0983_ sky130_fd_sc_hd__xnor2_1
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7726_ _2723_ _2885_ _2724_ vssd1 vssd1 vccd1 vccd1 _2886_ sky130_fd_sc_hd__a21oi_1
X_4938_ _4090_ _4092_ vssd1 vssd1 vccd1 vccd1 _4093_ sky130_fd_sc_hd__or2b_1
X_4869_ _3719_ _3795_ vssd1 vssd1 vccd1 vccd1 _4024_ sky130_fd_sc_hd__nor2_1
X_7657_ _2704_ _2808_ _2809_ _2742_ vssd1 vssd1 vccd1 vccd1 _2810_ sky130_fd_sc_hd__o211a_1
X_6608_ _1655_ _1551_ vssd1 vssd1 vccd1 vccd1 _1656_ sky130_fd_sc_hd__xor2_2
XFILLER_20_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7588_ _2715_ _2733_ _2707_ vssd1 vssd1 vccd1 vccd1 _2734_ sky130_fd_sc_hd__mux2_1
X_6539_ _1578_ _1579_ vssd1 vssd1 vccd1 vccd1 _1580_ sky130_fd_sc_hd__xnor2_1
XFILLER_106_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8209_ _0600_ _3387_ _3398_ _3410_ vssd1 vssd1 vccd1 vccd1 _3411_ sky130_fd_sc_hd__o211a_1
XFILLER_0_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4865__B _3930_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4618__C1 _3771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4881__A _4033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4267__S _0712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5910_ _3770_ _0892_ vssd1 vssd1 vccd1 vccd1 _0902_ sky130_fd_sc_hd__nor2_1
XFILLER_81_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4791__A _3816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6890_ _1906_ _1909_ vssd1 vssd1 vccd1 vccd1 _1966_ sky130_fd_sc_hd__xnor2_1
XFILLER_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5841_ _3770_ _0828_ vssd1 vssd1 vccd1 vccd1 _0829_ sky130_fd_sc_hd__nor2_1
X_5772_ _3700_ _0737_ _0745_ _0754_ vssd1 vssd1 vccd1 vccd1 _0755_ sky130_fd_sc_hd__a31oi_4
X_8560_ clknet_3_2__leaf_clk _0046_ vssd1 vssd1 vccd1 vccd1 posit_add.in1\[3\] sky130_fd_sc_hd__dfxtp_2
X_4723_ _3877_ vssd1 vssd1 vccd1 vccd1 _3878_ sky130_fd_sc_hd__clkbuf_4
X_8491_ _3683_ vssd1 vssd1 vccd1 vccd1 _0063_ sky130_fd_sc_hd__clkbuf_1
X_7511_ _2623_ _2625_ _2647_ _2648_ vssd1 vssd1 vccd1 vccd1 _2649_ sky130_fd_sc_hd__a31o_1
X_7442_ _2569_ _2558_ _2572_ _2447_ vssd1 vssd1 vccd1 vccd1 _2574_ sky130_fd_sc_hd__a211o_1
XANTENNA__7326__B2 _2335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4654_ _2012_ _2111_ _2210_ _1836_ vssd1 vssd1 vccd1 vccd1 _3809_ sky130_fd_sc_hd__a211o_1
XFILLER_30_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4585_ _3339_ _3349_ _2694_ _3360_ vssd1 vssd1 vccd1 vccd1 _3740_ sky130_fd_sc_hd__o211a_1
X_7373_ _2297_ _2497_ vssd1 vssd1 vccd1 vccd1 _2498_ sky130_fd_sc_hd__xor2_1
XFILLER_115_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6324_ _1004_ _1040_ _1039_ vssd1 vssd1 vccd1 vccd1 _1344_ sky130_fd_sc_hd__o21ba_1
XANTENNA__4560__A1 _1858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8341__A2_N _3549_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6255_ _0802_ _0787_ _1094_ _1127_ vssd1 vssd1 vccd1 vccd1 _1268_ sky130_fd_sc_hd__or4b_1
X_5206_ _3800_ _4037_ vssd1 vssd1 vccd1 vccd1 _0179_ sky130_fd_sc_hd__nor2_1
X_6186_ _0722_ _1127_ vssd1 vssd1 vccd1 vccd1 _1193_ sky130_fd_sc_hd__nand2_1
XFILLER_57_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5137_ _0106_ _0109_ vssd1 vssd1 vccd1 vccd1 _0110_ sky130_fd_sc_hd__nand2_1
X_5068_ _4222_ _3838_ vssd1 vssd1 vccd1 vccd1 _4223_ sky130_fd_sc_hd__nand2_1
Xposit_unit_6 vssd1 vssd1 vccd1 vccd1 posit_unit_6/HI io_out[1] sky130_fd_sc_hd__conb_1
XFILLER_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7709_ _2743_ _2750_ _2866_ vssd1 vssd1 vccd1 vccd1 _2867_ sky130_fd_sc_hd__o21ai_2
XFILLER_21_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4370_ posit_add.in2\[4\] _1847_ vssd1 vssd1 vccd1 vccd1 _1858_ sky130_fd_sc_hd__xor2_4
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6040_ _1006_ _1011_ _1038_ vssd1 vssd1 vccd1 vccd1 _1039_ sky130_fd_sc_hd__a21oi_1
XFILLER_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4845__A2 _3771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7991_ _3175_ _3176_ _3065_ vssd1 vssd1 vccd1 vccd1 _3177_ sky130_fd_sc_hd__mux2_1
X_6942_ _2019_ _2021_ _2022_ vssd1 vssd1 vccd1 vccd1 _2024_ sky130_fd_sc_hd__a21o_1
XFILLER_81_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6506__A _1353_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6225__B _1164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6873_ _1901_ _1947_ vssd1 vssd1 vccd1 vccd1 _1948_ sky130_fd_sc_hd__and2b_1
X_5824_ _0770_ _0776_ vssd1 vssd1 vccd1 vccd1 _0811_ sky130_fd_sc_hd__nor2_1
X_5755_ _0113_ _0733_ _0734_ _0736_ _4222_ vssd1 vssd1 vccd1 vccd1 _0737_ sky130_fd_sc_hd__a311o_1
X_8543_ clknet_3_2__leaf_clk _0029_ vssd1 vssd1 vccd1 vccd1 out_reg\[9\] sky130_fd_sc_hd__dfxtp_1
X_5686_ _0651_ _0661_ _0613_ vssd1 vssd1 vccd1 vccd1 _0662_ sky130_fd_sc_hd__o21a_1
X_4706_ _3843_ _3859_ vssd1 vssd1 vccd1 vccd1 _3861_ sky130_fd_sc_hd__nand2_1
X_8474_ _3672_ vssd1 vssd1 vccd1 vccd1 _0056_ sky130_fd_sc_hd__clkbuf_1
X_7425_ _2552_ _2241_ vssd1 vssd1 vccd1 vccd1 _2555_ sky130_fd_sc_hd__xnor2_1
X_4637_ _3791_ vssd1 vssd1 vccd1 vccd1 _3792_ sky130_fd_sc_hd__buf_4
XFILLER_104_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4568_ _3079_ _3296_ _3232_ _3046_ vssd1 vssd1 vccd1 vccd1 _3723_ sky130_fd_sc_hd__a211o_1
X_7356_ _2475_ _2478_ _2451_ vssd1 vssd1 vccd1 vccd1 _2479_ sky130_fd_sc_hd__a21oi_1
X_6307_ _1150_ _1151_ vssd1 vssd1 vccd1 vccd1 _1325_ sky130_fd_sc_hd__nand2_1
XFILLER_89_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4499_ _2837_ _3264_ _2793_ vssd1 vssd1 vccd1 vccd1 _3275_ sky130_fd_sc_hd__a21oi_2
XANTENNA__5089__A2 _4232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7287_ _2349_ _2391_ _2384_ vssd1 vssd1 vccd1 vccd1 _2403_ sky130_fd_sc_hd__a21oi_2
XFILLER_103_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6238_ _1247_ _1248_ vssd1 vssd1 vccd1 vccd1 _1249_ sky130_fd_sc_hd__xor2_1
XFILLER_89_468 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6169_ _1160_ _1159_ _1161_ vssd1 vssd1 vccd1 vccd1 _1174_ sky130_fd_sc_hd__a21o_1
XFILLER_103_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5304__B _4232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6589__A2 _1400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5261__A2 _3615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7247__A _2354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4280__S _0830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5540_ _0444_ _0510_ vssd1 vssd1 vccd1 vccd1 _0513_ sky130_fd_sc_hd__or2b_1
X_5471_ _0375_ _0392_ vssd1 vssd1 vccd1 vccd1 _0444_ sky130_fd_sc_hd__xor2_2
XFILLER_117_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4422_ posit_add.in2\[1\] _2023_ vssd1 vssd1 vccd1 vccd1 _2430_ sky130_fd_sc_hd__xnor2_1
X_7210_ _2299_ _2302_ _2303_ vssd1 vssd1 vccd1 vccd1 _2318_ sky130_fd_sc_hd__or3_1
X_8190_ _3234_ _3143_ _3389_ vssd1 vssd1 vccd1 vccd1 _3390_ sky130_fd_sc_hd__o21a_1
X_7141_ _2152_ _2180_ vssd1 vssd1 vccd1 vccd1 _2242_ sky130_fd_sc_hd__nor2_1
X_4353_ posit_add.in2\[5\] posit_add.in2\[4\] posit_add.in2\[6\] _1352_ _1264_ vssd1
+ vssd1 vccd1 vccd1 _1671_ sky130_fd_sc_hd__o41a_2
X_7072_ _2129_ _2165_ vssd1 vssd1 vccd1 vccd1 _2167_ sky130_fd_sc_hd__xnor2_1
X_4284_ in_reg\[3\] in_reg\[4\] _0830_ vssd1 vssd1 vccd1 vccd1 _0925_ sky130_fd_sc_hd__mux2_1
X_6023_ _0803_ _0993_ _1008_ _1020_ vssd1 vssd1 vccd1 vccd1 _1021_ sky130_fd_sc_hd__o211a_1
XFILLER_100_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7974_ _3100_ _3086_ _3065_ vssd1 vssd1 vccd1 vccd1 _3159_ sky130_fd_sc_hd__mux2_1
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6925_ _1840_ _1895_ vssd1 vssd1 vccd1 vccd1 _2005_ sky130_fd_sc_hd__nand2_1
XFILLER_42_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6856_ _1927_ _1928_ vssd1 vssd1 vccd1 vccd1 _1929_ sky130_fd_sc_hd__xnor2_1
XFILLER_50_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5807_ _0766_ _0768_ vssd1 vssd1 vccd1 vccd1 _0792_ sky130_fd_sc_hd__or2b_1
X_6787_ _1399_ _4126_ vssd1 vssd1 vccd1 vccd1 _1853_ sky130_fd_sc_hd__or2_1
XFILLER_10_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7067__A _1676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5738_ _0711_ _0718_ vssd1 vssd1 vccd1 vccd1 _0719_ sky130_fd_sc_hd__xor2_1
X_8526_ clknet_3_7__leaf_clk _0012_ vssd1 vssd1 vccd1 vccd1 in_reg\[9\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__4754__A1 _3881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5669_ _0638_ _0642_ vssd1 vssd1 vccd1 vccd1 _0643_ sky130_fd_sc_hd__or2b_1
X_8457_ in_reg\[5\] posit_add.in1\[5\] _3655_ vssd1 vssd1 vccd1 vccd1 _3662_ sky130_fd_sc_hd__mux2_1
X_7408_ _2151_ _2244_ vssd1 vssd1 vccd1 vccd1 _2536_ sky130_fd_sc_hd__xnor2_2
X_8388_ _3195_ _3599_ _3600_ vssd1 vssd1 vccd1 vccd1 _3601_ sky130_fd_sc_hd__o21ba_1
X_7339_ _4089_ _2431_ _2437_ _2458_ _2459_ vssd1 vssd1 vccd1 vccd1 _2460_ sky130_fd_sc_hd__o221a_1
XFILLER_1_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7456__B1 _2382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4971_ _3726_ vssd1 vssd1 vccd1 vccd1 _4126_ sky130_fd_sc_hd__buf_4
X_6710_ _1761_ _1767_ vssd1 vssd1 vccd1 vccd1 _1768_ sky130_fd_sc_hd__xor2_1
X_7690_ _2783_ _2818_ vssd1 vssd1 vccd1 vccd1 _2846_ sky130_fd_sc_hd__nand2_1
XFILLER_32_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6641_ _1654_ _1658_ vssd1 vssd1 vccd1 vccd1 _1692_ sky130_fd_sc_hd__nand2_1
XFILLER_20_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6572_ _1461_ _1527_ _1526_ vssd1 vssd1 vccd1 vccd1 _1617_ sky130_fd_sc_hd__a21oi_1
X_8311_ _0440_ _0521_ _3516_ _3517_ _3518_ vssd1 vssd1 vccd1 vccd1 _3519_ sky130_fd_sc_hd__o221a_1
XANTENNA__5119__B _3989_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5523_ _0495_ vssd1 vssd1 vccd1 vccd1 _0496_ sky130_fd_sc_hd__clkinv_2
XFILLER_117_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8242_ out_reg\[6\] _3316_ _3197_ out_reg\[7\] vssd1 vssd1 vccd1 vccd1 _3447_ sky130_fd_sc_hd__a22oi_1
XANTENNA__7686__B1 _1297_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5454_ _3488_ _0408_ _0409_ vssd1 vssd1 vccd1 vccd1 _0427_ sky130_fd_sc_hd__o21a_1
X_4405_ _2034_ _2045_ vssd1 vssd1 vccd1 vccd1 _2243_ sky130_fd_sc_hd__nor2_1
X_5385_ _1484_ _2452_ vssd1 vssd1 vccd1 vccd1 _0358_ sky130_fd_sc_hd__or2_1
X_8173_ _3152_ _3372_ _3234_ vssd1 vssd1 vccd1 vccd1 _3373_ sky130_fd_sc_hd__mux2_1
X_7124_ _2207_ _2211_ vssd1 vssd1 vccd1 vccd1 _2224_ sky130_fd_sc_hd__nor2_1
X_4336_ posit_add.in2\[11\] _1473_ vssd1 vssd1 vccd1 vccd1 _1484_ sky130_fd_sc_hd__xnor2_4
XFILLER_5_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7055_ _2146_ _2145_ vssd1 vssd1 vccd1 vccd1 _2148_ sky130_fd_sc_hd__and2b_1
X_4267_ in_reg\[6\] cmd\[6\] _0712_ vssd1 vssd1 vccd1 vccd1 _0744_ sky130_fd_sc_hd__mux2_1
XFILLER_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8446__A _3654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7350__A _2335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6006_ _4210_ _0993_ _1002_ vssd1 vssd1 vccd1 vccd1 _1003_ sky130_fd_sc_hd__or3_1
XFILLER_74_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6413__A1 _0795_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7957_ _3139_ _3011_ _2999_ vssd1 vssd1 vccd1 vccd1 _3140_ sky130_fd_sc_hd__mux2_1
X_6908_ _1920_ _1925_ vssd1 vssd1 vccd1 vccd1 _1986_ sky130_fd_sc_hd__xor2_1
XFILLER_70_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5020__D _4174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7888_ _3058_ _3063_ _2999_ vssd1 vssd1 vccd1 vccd1 _3064_ sky130_fd_sc_hd__mux2_1
X_6839_ _1865_ _1905_ _1906_ _1909_ vssd1 vssd1 vccd1 vccd1 _1910_ sky130_fd_sc_hd__a22o_1
XFILLER_7_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8509_ _3694_ vssd1 vssd1 vccd1 vccd1 _0072_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5170_ _0138_ _0142_ vssd1 vssd1 vccd1 vccd1 _0143_ sky130_fd_sc_hd__xnor2_1
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7170__A _4250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput4 rst vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__clkbuf_2
XFILLER_96_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7811_ _2976_ _2978_ vssd1 vssd1 vccd1 vccd1 _2979_ sky130_fd_sc_hd__nor2_1
XFILLER_101_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4954_ _4083_ _4084_ vssd1 vssd1 vccd1 vccd1 _4109_ sky130_fd_sc_hd__xnor2_1
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7742_ _2895_ _2902_ vssd1 vssd1 vccd1 vccd1 _2904_ sky130_fd_sc_hd__or2_1
XFILLER_24_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4885_ _3985_ _4039_ vssd1 vssd1 vccd1 vccd1 _4040_ sky130_fd_sc_hd__or2b_1
X_7673_ _2827_ vssd1 vssd1 vccd1 vccd1 _2828_ sky130_fd_sc_hd__inv_2
XFILLER_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6624_ _1667_ _1673_ _1420_ _1666_ vssd1 vssd1 vccd1 vccd1 _1674_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_118_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6555_ _0303_ _1400_ vssd1 vssd1 vccd1 vccd1 _1598_ sky130_fd_sc_hd__or2_1
X_5506_ _0478_ _0455_ vssd1 vssd1 vccd1 vccd1 _0479_ sky130_fd_sc_hd__xor2_2
X_6486_ _1507_ _1521_ vssd1 vssd1 vccd1 vccd1 _1522_ sky130_fd_sc_hd__xnor2_1
XANTENNA__5134__A1 _3925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8225_ _3340_ _3364_ _3385_ vssd1 vssd1 vccd1 vccd1 _3428_ sky130_fd_sc_hd__or3_1
X_5437_ _3167_ _0409_ vssd1 vssd1 vccd1 vccd1 _0410_ sky130_fd_sc_hd__xnor2_2
XFILLER_99_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8156_ _2604_ _2592_ _3353_ vssd1 vssd1 vccd1 vccd1 _3354_ sky130_fd_sc_hd__o21ai_2
XANTENNA__7999__B _4250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5368_ _4209_ _0340_ _0338_ vssd1 vssd1 vccd1 vccd1 _0341_ sky130_fd_sc_hd__mux2_1
XFILLER_114_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7107_ _2184_ _2195_ vssd1 vssd1 vccd1 vccd1 _2205_ sky130_fd_sc_hd__and2_1
XFILLER_87_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5299_ _0270_ _0271_ vssd1 vssd1 vccd1 vccd1 _0272_ sky130_fd_sc_hd__and2b_1
X_4319_ _1286_ vssd1 vssd1 vccd1 vccd1 _1297_ sky130_fd_sc_hd__clkbuf_4
X_8087_ out_reg\[1\] _3242_ _0701_ vssd1 vssd1 vccd1 vccd1 _3281_ sky130_fd_sc_hd__a21bo_1
XFILLER_101_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7038_ _2094_ _2096_ vssd1 vssd1 vccd1 vccd1 _2129_ sky130_fd_sc_hd__xnor2_1
XFILLER_59_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5312__B _2540_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6424__A _3795_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8311__A1 _0440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5428__A2 _0121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6334__A _4037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4670_ _3509_ _3824_ _3156_ vssd1 vssd1 vccd1 vccd1 _3825_ sky130_fd_sc_hd__mux2_1
XANTENNA__4789__A _3893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6340_ _0995_ _1338_ _1360_ vssd1 vssd1 vccd1 vccd1 _1361_ sky130_fd_sc_hd__o21ai_1
XFILLER_115_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6271_ _0706_ _1164_ _1283_ _1284_ vssd1 vssd1 vccd1 vccd1 _1285_ sky130_fd_sc_hd__a31o_1
X_5222_ _0192_ _0194_ vssd1 vssd1 vccd1 vccd1 _0195_ sky130_fd_sc_hd__nor2_1
X_8010_ _1231_ vssd1 vssd1 vccd1 vccd1 _3197_ sky130_fd_sc_hd__buf_2
X_5153_ _4227_ _4231_ _4245_ vssd1 vssd1 vccd1 vccd1 _0126_ sky130_fd_sc_hd__nor3_1
XFILLER_111_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4627__B1 _3771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5084_ _4220_ _4223_ _4225_ _4218_ vssd1 vssd1 vccd1 vccd1 _4239_ sky130_fd_sc_hd__o22a_1
XFILLER_49_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5986_ _0849_ vssd1 vssd1 vccd1 vccd1 _0982_ sky130_fd_sc_hd__inv_2
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4937_ _4071_ _4091_ vssd1 vssd1 vccd1 vccd1 _4092_ sky130_fd_sc_hd__xnor2_1
X_7725_ _2739_ _2740_ _2884_ vssd1 vssd1 vccd1 vccd1 _2885_ sky130_fd_sc_hd__o21a_1
X_4868_ _4022_ _3928_ vssd1 vssd1 vccd1 vccd1 _4023_ sky130_fd_sc_hd__xnor2_1
X_7656_ _2704_ _2766_ vssd1 vssd1 vccd1 vccd1 _2809_ sky130_fd_sc_hd__nand2_1
X_6607_ _1428_ _1410_ vssd1 vssd1 vccd1 vccd1 _1655_ sky130_fd_sc_hd__or2_2
XFILLER_118_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4799_ _3937_ _3953_ vssd1 vssd1 vccd1 vccd1 _3954_ sky130_fd_sc_hd__xnor2_1
X_7587_ _4153_ _0113_ _2652_ vssd1 vssd1 vccd1 vccd1 _2733_ sky130_fd_sc_hd__mux2_1
X_6538_ _1522_ _1523_ vssd1 vssd1 vccd1 vccd1 _1579_ sky130_fd_sc_hd__xnor2_1
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6469_ _1496_ _1502_ vssd1 vssd1 vccd1 vccd1 _1503_ sky130_fd_sc_hd__xor2_1
XFILLER_106_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8208_ _3400_ _3408_ _3409_ vssd1 vssd1 vccd1 vccd1 _3410_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8139_ _3305_ _3310_ vssd1 vssd1 vccd1 vccd1 _3336_ sky130_fd_sc_hd__nor2_1
XFILLER_102_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_503 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4791__B _3702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5840_ _0754_ _0826_ vssd1 vssd1 vccd1 vccd1 _0828_ sky130_fd_sc_hd__xor2_1
XFILLER_34_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6999__A _1456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5771_ _0749_ _0753_ _3802_ vssd1 vssd1 vccd1 vccd1 _0754_ sky130_fd_sc_hd__o21a_2
X_4722_ _3729_ _3876_ vssd1 vssd1 vccd1 vccd1 _3877_ sky130_fd_sc_hd__nor2_1
X_8490_ posit_add.in2\[4\] in_reg\[4\] _3677_ vssd1 vssd1 vccd1 vccd1 _3683_ sky130_fd_sc_hd__mux2_1
X_7510_ _3328_ _0347_ vssd1 vssd1 vccd1 vccd1 _2648_ sky130_fd_sc_hd__nor2_1
XANTENNA__5337__A1 _2540_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7441_ _2454_ _2525_ _2526_ vssd1 vssd1 vccd1 vccd1 _2572_ sky130_fd_sc_hd__o21a_1
X_4653_ _1946_ _3635_ _3707_ _2309_ vssd1 vssd1 vccd1 vccd1 _3808_ sky130_fd_sc_hd__a211o_1
X_4584_ _3738_ vssd1 vssd1 vccd1 vccd1 _3739_ sky130_fd_sc_hd__clkbuf_4
X_7372_ _2008_ _2261_ _2268_ vssd1 vssd1 vccd1 vccd1 _2497_ sky130_fd_sc_hd__and3_1
X_6323_ _1004_ _1342_ vssd1 vssd1 vccd1 vccd1 _1343_ sky130_fd_sc_hd__xor2_1
XFILLER_107_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6254_ _0787_ _1095_ _1128_ _1007_ vssd1 vssd1 vccd1 vccd1 _1267_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6837__A1 _4217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5205_ _0169_ _0177_ vssd1 vssd1 vccd1 vccd1 _0178_ sky130_fd_sc_hd__xnor2_1
X_6185_ _0892_ _1094_ vssd1 vssd1 vccd1 vccd1 _1192_ sky130_fd_sc_hd__or2_1
X_5136_ _3701_ _3750_ _0108_ vssd1 vssd1 vccd1 vccd1 _0109_ sky130_fd_sc_hd__or3_1
X_5067_ _4221_ vssd1 vssd1 vccd1 vccd1 _4222_ sky130_fd_sc_hd__buf_4
XFILLER_84_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xposit_unit_7 vssd1 vssd1 vccd1 vccd1 posit_unit_7/HI io_out[2] sky130_fd_sc_hd__conb_1
XFILLER_65_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5969_ _0876_ _0877_ _0878_ vssd1 vssd1 vccd1 vccd1 _0964_ sky130_fd_sc_hd__o21a_1
XANTENNA__5576__A1 _2540_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7708_ _2704_ _2786_ _2865_ _2762_ vssd1 vssd1 vccd1 vccd1 _2866_ sky130_fd_sc_hd__a211o_1
X_7639_ _2788_ _2789_ vssd1 vssd1 vccd1 vccd1 _2790_ sky130_fd_sc_hd__and2_1
XFILLER_106_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6612__A _1420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4542__A2 _2452_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4278__S _0830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5898__A _3815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7990_ _3026_ _3008_ _2996_ vssd1 vssd1 vccd1 vccd1 _3176_ sky130_fd_sc_hd__o21ai_1
XANTENNA__7795__A2 _2721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6941_ _2013_ _2018_ vssd1 vssd1 vccd1 vccd1 _2022_ sky130_fd_sc_hd__and2b_1
XFILLER_93_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6506__B _1354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6872_ _1903_ _1940_ _1945_ vssd1 vssd1 vccd1 vccd1 _1947_ sky130_fd_sc_hd__o21ai_2
XFILLER_62_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5823_ _0801_ _0809_ vssd1 vssd1 vccd1 vccd1 _0810_ sky130_fd_sc_hd__xnor2_1
X_8542_ clknet_3_2__leaf_clk _0028_ vssd1 vssd1 vccd1 vccd1 out_reg\[8\] sky130_fd_sc_hd__dfxtp_1
X_5754_ _0687_ _0735_ _3718_ vssd1 vssd1 vccd1 vccd1 _0736_ sky130_fd_sc_hd__o21a_1
X_5685_ _3814_ _3791_ _2518_ vssd1 vssd1 vccd1 vccd1 _0661_ sky130_fd_sc_hd__a21oi_1
X_4705_ _3843_ _3859_ vssd1 vssd1 vccd1 vccd1 _3860_ sky130_fd_sc_hd__or2_1
X_8473_ in_reg\[13\] posit_add.in1\[13\] _3654_ vssd1 vssd1 vccd1 vccd1 _3672_ sky130_fd_sc_hd__mux2_1
XFILLER_118_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7424_ _2536_ _2553_ vssd1 vssd1 vccd1 vccd1 _2554_ sky130_fd_sc_hd__nand2_1
X_4636_ _3690_ _3713_ _3715_ _3774_ _3678_ vssd1 vssd1 vccd1 vccd1 _3791_ sky130_fd_sc_hd__a311o_2
XANTENNA__4977__A _2529_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7355_ _2379_ _2396_ _2407_ _2477_ vssd1 vssd1 vccd1 vccd1 _2478_ sky130_fd_sc_hd__or4_1
X_6306_ _1316_ _1318_ vssd1 vssd1 vccd1 vccd1 _1324_ sky130_fd_sc_hd__xnor2_1
XFILLER_89_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4567_ _3721_ vssd1 vssd1 vccd1 vccd1 _3722_ sky130_fd_sc_hd__clkbuf_4
XFILLER_104_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4498_ _2914_ _3253_ _2870_ vssd1 vssd1 vccd1 vccd1 _3264_ sky130_fd_sc_hd__o21ai_1
XFILLER_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7286_ _2377_ _2378_ _2384_ vssd1 vssd1 vccd1 vccd1 _2402_ sky130_fd_sc_hd__a21o_1
X_6237_ _1196_ _1206_ vssd1 vssd1 vccd1 vccd1 _1248_ sky130_fd_sc_hd__xor2_1
XFILLER_103_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6168_ _1168_ _1170_ vssd1 vssd1 vccd1 vccd1 _1173_ sky130_fd_sc_hd__xnor2_1
XFILLER_97_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5119_ _4210_ _3989_ vssd1 vssd1 vccd1 vccd1 _0092_ sky130_fd_sc_hd__or2_4
X_6099_ _1098_ _1100_ _4016_ vssd1 vssd1 vccd1 vccd1 _1101_ sky130_fd_sc_hd__a21oi_1
XFILLER_84_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5549__A1 _0445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6432__A _0082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7962__S _2999_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5048__A _4045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4288__A1 in_reg\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6607__A _1428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4763__A2 _3635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5470_ _0442_ _0394_ vssd1 vssd1 vccd1 vccd1 _0443_ sky130_fd_sc_hd__xnor2_2
XFILLER_117_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4421_ _1880_ _2221_ _2386_ _2408_ vssd1 vssd1 vccd1 vccd1 _2419_ sky130_fd_sc_hd__a211o_1
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7140_ _2203_ _2239_ _2240_ vssd1 vssd1 vccd1 vccd1 _2241_ sky130_fd_sc_hd__a21bo_1
X_4352_ posit_add.in2\[8\] _1649_ vssd1 vssd1 vccd1 vccd1 _1660_ sky130_fd_sc_hd__xnor2_2
X_7071_ _2128_ _2164_ vssd1 vssd1 vccd1 vccd1 _2165_ sky130_fd_sc_hd__nor2_1
X_4283_ _0904_ vssd1 vssd1 vccd1 vccd1 _0006_ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6022_ _1019_ _0993_ vssd1 vssd1 vccd1 vccd1 _1020_ sky130_fd_sc_hd__nand2_1
XFILLER_100_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7973_ _3155_ _3157_ _3021_ vssd1 vssd1 vccd1 vccd1 _3158_ sky130_fd_sc_hd__mux2_1
XFILLER_54_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6924_ _1948_ _2000_ _2003_ vssd1 vssd1 vccd1 vccd1 _2004_ sky130_fd_sc_hd__o21a_1
XFILLER_81_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4451__A1 posit_add.in1\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6855_ _1878_ _1881_ vssd1 vssd1 vccd1 vccd1 _1928_ sky130_fd_sc_hd__xnor2_1
XFILLER_22_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5806_ _0760_ _0784_ _0790_ vssd1 vssd1 vccd1 vccd1 _0791_ sky130_fd_sc_hd__o21a_1
X_6786_ _1482_ _1782_ _1849_ _1851_ vssd1 vssd1 vccd1 vccd1 _1852_ sky130_fd_sc_hd__a31o_1
XANTENNA__7067__B _1537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5737_ _0713_ _0717_ vssd1 vssd1 vccd1 vccd1 _0718_ sky130_fd_sc_hd__xor2_1
X_8525_ clknet_3_7__leaf_clk _0011_ vssd1 vssd1 vccd1 vccd1 in_reg\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_22_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8456_ _3661_ vssd1 vssd1 vccd1 vccd1 _0047_ sky130_fd_sc_hd__clkbuf_1
X_5668_ _0639_ _0641_ vssd1 vssd1 vccd1 vccd1 _0642_ sky130_fd_sc_hd__nand2_1
XFILLER_89_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7407_ _2444_ _2524_ _2534_ _2416_ vssd1 vssd1 vccd1 vccd1 _2535_ sky130_fd_sc_hd__a22o_1
X_4619_ _3765_ _2309_ _2452_ _2474_ vssd1 vssd1 vccd1 vccd1 _3774_ sky130_fd_sc_hd__o31a_2
X_8387_ out_reg\[12\] _3316_ _1231_ out_reg\[13\] vssd1 vssd1 vccd1 vccd1 _3600_ sky130_fd_sc_hd__a22o_1
X_5599_ _0526_ _0522_ _0515_ vssd1 vssd1 vccd1 vccd1 _0572_ sky130_fd_sc_hd__mux2_1
XFILLER_116_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7338_ _2416_ _2432_ vssd1 vssd1 vccd1 vccd1 _2459_ sky130_fd_sc_hd__nand2_1
XFILLER_8_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7269_ _2381_ _2382_ vssd1 vssd1 vccd1 vccd1 _2383_ sky130_fd_sc_hd__nor2_1
XFILLER_104_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6427__A _4250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7957__S _2999_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4970_ _4117_ _4124_ vssd1 vssd1 vccd1 vccd1 _4125_ sky130_fd_sc_hd__nand2_1
XFILLER_17_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6640_ _1675_ _1689_ _1690_ vssd1 vssd1 vccd1 vccd1 _1691_ sky130_fd_sc_hd__a21oi_1
XANTENNA__5394__C1 _3736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6571_ _1585_ _1614_ vssd1 vssd1 vccd1 vccd1 _1615_ sky130_fd_sc_hd__xnor2_1
XFILLER_32_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8310_ _3516_ _3517_ vssd1 vssd1 vccd1 vccd1 _3518_ sky130_fd_sc_hd__nand2_1
X_5522_ _0481_ _0492_ _0494_ vssd1 vssd1 vccd1 vccd1 _0495_ sky130_fd_sc_hd__mux2_1
XFILLER_117_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8241_ _3425_ _3436_ _3444_ _3195_ vssd1 vssd1 vccd1 vccd1 _3445_ sky130_fd_sc_hd__a31o_1
X_5453_ _3830_ _0348_ vssd1 vssd1 vccd1 vccd1 _0426_ sky130_fd_sc_hd__xnor2_1
X_4404_ _2012_ _2111_ _2210_ _1858_ vssd1 vssd1 vccd1 vccd1 _2232_ sky130_fd_sc_hd__a211oi_1
X_5384_ _3736_ _3659_ _3671_ vssd1 vssd1 vccd1 vccd1 _0357_ sky130_fd_sc_hd__nand3_1
X_8172_ _3370_ vssd1 vssd1 vccd1 vccd1 _3372_ sky130_fd_sc_hd__clkinv_2
XANTENNA__4320__A _1297_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7123_ _2216_ _2222_ vssd1 vssd1 vccd1 vccd1 _2223_ sky130_fd_sc_hd__nand2_1
XFILLER_87_704 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4335_ _1341_ _1374_ _1462_ _1264_ vssd1 vssd1 vccd1 vccd1 _1473_ sky130_fd_sc_hd__o31a_1
XFILLER_115_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7631__A _2780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5449__A0 _3736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7054_ _2145_ _2146_ vssd1 vssd1 vccd1 vccd1 _2147_ sky130_fd_sc_hd__xnor2_1
X_4266_ _0723_ vssd1 vssd1 vccd1 vccd1 _0000_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6661__A2 _1711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6005_ _1000_ _1001_ vssd1 vssd1 vccd1 vccd1 _1002_ sky130_fd_sc_hd__nor2_1
XANTENNA__6247__A _0722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5151__A _3827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7956_ _3129_ _3138_ _3042_ vssd1 vssd1 vccd1 vccd1 _3139_ sky130_fd_sc_hd__mux2_1
X_6907_ _1981_ _1983_ _1984_ vssd1 vssd1 vccd1 vccd1 _1985_ sky130_fd_sc_hd__a21o_1
X_7887_ _3042_ _3062_ _3056_ _3049_ vssd1 vssd1 vccd1 vccd1 _3063_ sky130_fd_sc_hd__a22o_1
XFILLER_23_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6838_ _1865_ _1905_ _1908_ vssd1 vssd1 vccd1 vccd1 _1909_ sky130_fd_sc_hd__a21oi_1
XFILLER_10_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8508_ posit_add.in2\[13\] in_reg\[13\] _3676_ vssd1 vssd1 vccd1 vccd1 _3694_ sky130_fd_sc_hd__mux2_1
X_6769_ _1778_ _1800_ _1832_ vssd1 vssd1 vccd1 vccd1 _1833_ sky130_fd_sc_hd__o21ai_1
XFILLER_6_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8439_ counter\[2\] _3644_ counter\[3\] vssd1 vssd1 vccd1 vccd1 _3649_ sky130_fd_sc_hd__a21o_1
XFILLER_2_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7365__B1 _2488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8314__C1 _0701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4286__S _0830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7170__B _0303_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7810_ _2960_ _2977_ vssd1 vssd1 vccd1 vccd1 _2978_ sky130_fd_sc_hd__or2_1
XFILLER_37_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4953_ _4106_ _4107_ vssd1 vssd1 vccd1 vccd1 _4108_ sky130_fd_sc_hd__nand2_1
XFILLER_51_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7741_ _2899_ _2901_ vssd1 vssd1 vccd1 vccd1 _2902_ sky130_fd_sc_hd__or2_1
XFILLER_24_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7672_ _2824_ _2752_ vssd1 vssd1 vccd1 vccd1 _2827_ sky130_fd_sc_hd__and2_1
X_6623_ _1670_ _1672_ vssd1 vssd1 vccd1 vccd1 _1673_ sky130_fd_sc_hd__xnor2_1
X_4884_ _4036_ _4038_ vssd1 vssd1 vccd1 vccd1 _4039_ sky130_fd_sc_hd__xor2_1
XFILLER_20_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6554_ _4153_ _1596_ _1467_ vssd1 vssd1 vccd1 vccd1 _1597_ sky130_fd_sc_hd__and3_1
XFILLER_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6485_ _1519_ _1520_ _1516_ vssd1 vssd1 vccd1 vccd1 _1521_ sky130_fd_sc_hd__a21o_1
X_5505_ _0447_ _0441_ vssd1 vssd1 vccd1 vccd1 _0478_ sky130_fd_sc_hd__nor2_1
XFILLER_118_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5436_ _3424_ _0408_ vssd1 vssd1 vccd1 vccd1 _0409_ sky130_fd_sc_hd__nand2_1
XFILLER_10_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8224_ _3166_ _3426_ vssd1 vssd1 vccd1 vccd1 _3427_ sky130_fd_sc_hd__or2_1
XFILLER_105_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5134__A2 _3615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5367_ _0319_ _0321_ vssd1 vssd1 vccd1 vccd1 _0340_ sky130_fd_sc_hd__xor2_1
X_8155_ _2569_ _3352_ _3286_ _2520_ vssd1 vssd1 vccd1 vccd1 _3353_ sky130_fd_sc_hd__o211ai_1
XFILLER_101_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7106_ _2198_ _2201_ _2200_ vssd1 vssd1 vccd1 vccd1 _2204_ sky130_fd_sc_hd__o21ai_1
X_5298_ _0257_ _0259_ _0263_ vssd1 vssd1 vccd1 vccd1 _0271_ sky130_fd_sc_hd__a21bo_1
XFILLER_59_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8086_ _3190_ _3278_ _3279_ _0701_ vssd1 vssd1 vccd1 vccd1 _3280_ sky130_fd_sc_hd__a31o_1
X_4318_ _1253_ _1275_ vssd1 vssd1 vccd1 vccd1 _1286_ sky130_fd_sc_hd__xor2_2
X_7037_ _2096_ _2127_ vssd1 vssd1 vccd1 vccd1 _2128_ sky130_fd_sc_hd__or2_1
XFILLER_87_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7939_ _3114_ _3119_ _2998_ vssd1 vssd1 vccd1 vccd1 _3120_ sky130_fd_sc_hd__mux2_1
XFILLER_27_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5056__A _4210_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4636__A1 _3690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7586__A0 _2319_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5876__D _3832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6270_ _1019_ _1128_ _1282_ vssd1 vssd1 vccd1 vccd1 _1284_ sky130_fd_sc_hd__and3_1
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5221_ _0175_ _0193_ vssd1 vssd1 vccd1 vccd1 _0194_ sky130_fd_sc_hd__or2_1
X_5152_ _3816_ _3989_ _0124_ vssd1 vssd1 vccd1 vccd1 _0125_ sky130_fd_sc_hd__or3_1
XFILLER_111_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5083_ _4233_ _4237_ vssd1 vssd1 vccd1 vccd1 _4238_ sky130_fd_sc_hd__xnor2_1
XFILLER_84_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7577__A0 _3802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5985_ _0962_ _0973_ _0979_ _0980_ vssd1 vssd1 vccd1 vccd1 _0981_ sky130_fd_sc_hd__o31ai_4
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7724_ _2739_ _2740_ _2825_ _2883_ _2827_ vssd1 vssd1 vccd1 vccd1 _2884_ sky130_fd_sc_hd__a221o_1
X_4936_ _4072_ _4088_ vssd1 vssd1 vccd1 vccd1 _4091_ sky130_fd_sc_hd__nor2_1
XFILLER_40_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4867_ _4020_ _4021_ vssd1 vssd1 vccd1 vccd1 _4022_ sky130_fd_sc_hd__nand2_1
X_7655_ _2712_ _2806_ _2807_ vssd1 vssd1 vccd1 vccd1 _2808_ sky130_fd_sc_hd__o21ai_1
X_6606_ _0303_ _1510_ vssd1 vssd1 vccd1 vccd1 _1654_ sky130_fd_sc_hd__nor2_2
XFILLER_20_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7586_ _2319_ _2714_ _2707_ vssd1 vssd1 vccd1 vccd1 _2732_ sky130_fd_sc_hd__mux2_1
XANTENNA__4699__B _3853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4798_ _3939_ _3951_ _3952_ vssd1 vssd1 vccd1 vccd1 _3953_ sky130_fd_sc_hd__a21bo_1
X_6537_ _1575_ _1576_ _1577_ vssd1 vssd1 vccd1 vccd1 _1578_ sky130_fd_sc_hd__a21o_1
XFILLER_118_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6468_ _1497_ _4211_ _1501_ vssd1 vssd1 vccd1 vccd1 _1502_ sky130_fd_sc_hd__a21o_1
X_6399_ _1400_ _1384_ vssd1 vssd1 vccd1 vccd1 _1426_ sky130_fd_sc_hd__nor2_1
X_8207_ _3400_ _3408_ _2621_ vssd1 vssd1 vccd1 vccd1 _3409_ sky130_fd_sc_hd__a21oi_1
X_5419_ _0391_ _0337_ _0389_ vssd1 vssd1 vccd1 vccd1 _0392_ sky130_fd_sc_hd__a21o_1
XFILLER_102_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4866__A1 _3701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8138_ _3190_ _3333_ _3334_ vssd1 vssd1 vccd1 vccd1 _3335_ sky130_fd_sc_hd__and3_1
XFILLER_0_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6419__B _0105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_718 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_675 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8069_ _0572_ _3260_ _0557_ vssd1 vssd1 vccd1 vccd1 _3261_ sky130_fd_sc_hd__mux2_1
XANTENNA__6435__A _1383_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6620__A1_N _1355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8036__S _2721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8220__A1 _1330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5770_ _0613_ _0750_ _0752_ vssd1 vssd1 vccd1 vccd1 _0753_ sky130_fd_sc_hd__a21oi_1
XFILLER_34_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4721_ _2485_ _3768_ vssd1 vssd1 vccd1 vccd1 _3876_ sky130_fd_sc_hd__or2_1
XANTENNA__5337__A2 _0303_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4652_ _3728_ _3799_ _3806_ vssd1 vssd1 vccd1 vccd1 _3807_ sky130_fd_sc_hd__and3_1
X_7440_ _2528_ _2560_ _2568_ _2570_ vssd1 vssd1 vccd1 vccd1 _2571_ sky130_fd_sc_hd__o31a_1
XFILLER_116_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4583_ _3737_ vssd1 vssd1 vccd1 vccd1 _3738_ sky130_fd_sc_hd__clkbuf_2
X_7371_ _2490_ _2492_ _2494_ vssd1 vssd1 vccd1 vccd1 _2495_ sky130_fd_sc_hd__mux2_1
X_6322_ _1338_ _1340_ vssd1 vssd1 vccd1 vccd1 _1342_ sky130_fd_sc_hd__nand2_1
XFILLER_115_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6253_ _0773_ _1168_ vssd1 vssd1 vccd1 vccd1 _1266_ sky130_fd_sc_hd__nor2_1
XFILLER_115_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5204_ _0153_ _0176_ vssd1 vssd1 vccd1 vccd1 _0177_ sky130_fd_sc_hd__nor2_1
XANTENNA__5424__A _0351_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6184_ _1158_ _1190_ vssd1 vssd1 vccd1 vccd1 _1191_ sky130_fd_sc_hd__xnor2_1
XFILLER_69_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5135_ _0106_ _0107_ vssd1 vssd1 vccd1 vccd1 _0108_ sky130_fd_sc_hd__nand2_1
XFILLER_96_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5066_ _3917_ _3922_ _3769_ _1748_ vssd1 vssd1 vccd1 vccd1 _4221_ sky130_fd_sc_hd__o22a_1
XFILLER_57_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5797__C _0779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8211__A1 _3195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5968_ _0910_ _0911_ vssd1 vssd1 vccd1 vccd1 _0963_ sky130_fd_sc_hd__nand2_1
XFILLER_80_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5576__A2 _0548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4919_ _3892_ _3883_ _4073_ vssd1 vssd1 vccd1 vccd1 _4074_ sky130_fd_sc_hd__and3_1
X_7707_ _2806_ _2862_ vssd1 vssd1 vccd1 vccd1 _2865_ sky130_fd_sc_hd__and2b_1
X_5899_ _0889_ _0890_ vssd1 vssd1 vccd1 vccd1 _0891_ sky130_fd_sc_hd__and2_1
XFILLER_20_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7638_ _3893_ _3868_ _2713_ vssd1 vssd1 vccd1 vccd1 _2789_ sky130_fd_sc_hd__mux2_1
XFILLER_119_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7569_ _2652_ vssd1 vssd1 vccd1 vccd1 _2713_ sky130_fd_sc_hd__clkbuf_4
XFILLER_4_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6612__B _1510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6940_ _2020_ _2010_ vssd1 vssd1 vccd1 vccd1 _2021_ sky130_fd_sc_hd__xnor2_1
XANTENNA__4294__S _0830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6506__C _0147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6871_ _1941_ _1944_ vssd1 vssd1 vccd1 vccd1 _1945_ sky130_fd_sc_hd__or2b_1
XFILLER_62_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5822_ _0806_ _0807_ vssd1 vssd1 vccd1 vccd1 _0809_ sky130_fd_sc_hd__xnor2_1
XFILLER_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5753_ _0616_ _0648_ _3762_ vssd1 vssd1 vccd1 vccd1 _0735_ sky130_fd_sc_hd__a21oi_1
X_8541_ clknet_3_0__leaf_clk _0027_ vssd1 vssd1 vccd1 vccd1 out_reg\[7\] sky130_fd_sc_hd__dfxtp_1
X_4704_ _3857_ _3858_ vssd1 vssd1 vccd1 vccd1 _3859_ sky130_fd_sc_hd__nand2_1
X_5684_ _3700_ _0652_ _0654_ _0659_ vssd1 vssd1 vccd1 vccd1 _0660_ sky130_fd_sc_hd__o22a_1
XANTENNA__4323__A posit_add.in2\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8472_ _3670_ vssd1 vssd1 vccd1 vccd1 _0055_ sky130_fd_sc_hd__clkbuf_1
XFILLER_30_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7423_ _2552_ _2542_ vssd1 vssd1 vccd1 vccd1 _2553_ sky130_fd_sc_hd__xnor2_1
X_4635_ _3782_ _3789_ vssd1 vssd1 vccd1 vccd1 _3790_ sky130_fd_sc_hd__xnor2_1
XFILLER_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4566_ _3720_ vssd1 vssd1 vccd1 vccd1 _3721_ sky130_fd_sc_hd__clkbuf_4
X_7354_ _3986_ _2431_ _2442_ _2462_ _2476_ vssd1 vssd1 vccd1 vccd1 _2477_ sky130_fd_sc_hd__o221a_1
X_6305_ _1321_ _1322_ vssd1 vssd1 vccd1 vccd1 _1323_ sky130_fd_sc_hd__or2b_1
XANTENNA__4977__B _3703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4497_ _3199_ _3243_ _2947_ vssd1 vssd1 vccd1 vccd1 _3253_ sky130_fd_sc_hd__a21oi_1
X_7285_ _2392_ _2388_ _2398_ _2400_ vssd1 vssd1 vccd1 vccd1 _2401_ sky130_fd_sc_hd__a211o_1
XFILLER_103_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6236_ _1238_ _1245_ _1246_ vssd1 vssd1 vccd1 vccd1 _1247_ sky130_fd_sc_hd__o21ai_1
X_6167_ _0795_ _1128_ _1163_ _1171_ vssd1 vssd1 vccd1 vccd1 _1172_ sky130_fd_sc_hd__a31o_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5118_ _0087_ _0086_ vssd1 vssd1 vccd1 vccd1 _0091_ sky130_fd_sc_hd__or2_1
X_6098_ _1099_ _0986_ vssd1 vssd1 vccd1 vccd1 _1100_ sky130_fd_sc_hd__xnor2_2
XANTENNA__5246__A1 _0218_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_698 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5049_ _4045_ _4153_ _4202_ vssd1 vssd1 vccd1 vccd1 _4204_ sky130_fd_sc_hd__a21oi_1
XFILLER_84_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6746__A1 _1665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6432__B _1423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5048__B _4153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5064__A _4210_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5999__A _4016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5239__A _3881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4420_ _2397_ vssd1 vssd1 vccd1 vccd1 _2408_ sky130_fd_sc_hd__buf_2
XFILLER_8_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5712__A2 _0687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4351_ _1352_ _1374_ _1264_ vssd1 vssd1 vccd1 vccd1 _1649_ sky130_fd_sc_hd__o21a_1
XANTENNA__4920__B1 _3702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7070_ _2156_ _2157_ _2126_ vssd1 vssd1 vccd1 vccd1 _2164_ sky130_fd_sc_hd__o21a_1
X_4282_ in_reg\[2\] in_reg\[3\] _0830_ vssd1 vssd1 vccd1 vccd1 _0904_ sky130_fd_sc_hd__mux2_1
XFILLER_101_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6021_ _3701_ _0737_ _0745_ _0754_ vssd1 vssd1 vccd1 vccd1 _1019_ sky130_fd_sc_hd__a31o_2
XFILLER_86_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8414__A1 cmd\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8414__B2 cmd\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7972_ _3131_ _3140_ _3065_ vssd1 vssd1 vccd1 vccd1 _3157_ sky130_fd_sc_hd__mux2_1
XANTENNA__4318__A _1253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6923_ _1895_ _2002_ vssd1 vssd1 vccd1 vccd1 _2003_ sky130_fd_sc_hd__nor2_2
XFILLER_54_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8178__B1 _3195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6854_ _1920_ _1925_ _1926_ vssd1 vssd1 vccd1 vccd1 _1927_ sky130_fd_sc_hd__a21bo_1
X_5805_ _0785_ _0789_ vssd1 vssd1 vccd1 vccd1 _0790_ sky130_fd_sc_hd__or2b_1
X_6785_ _1787_ _1850_ vssd1 vssd1 vccd1 vccd1 _1851_ sky130_fd_sc_hd__nor2_1
XANTENNA__5149__A _3881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5736_ _0714_ _0715_ _0716_ vssd1 vssd1 vccd1 vccd1 _0717_ sky130_fd_sc_hd__o21ai_1
X_8524_ clknet_3_3__leaf_clk _0010_ vssd1 vssd1 vccd1 vccd1 in_reg\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_10_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5667_ _4045_ _0639_ _0624_ _0640_ vssd1 vssd1 vccd1 vccd1 _0641_ sky130_fd_sc_hd__nand4_1
X_8455_ in_reg\[4\] posit_add.in1\[4\] _3655_ vssd1 vssd1 vccd1 vccd1 _3661_ sky130_fd_sc_hd__mux2_1
X_7406_ _2530_ _2532_ _2533_ vssd1 vssd1 vccd1 vccd1 _2534_ sky130_fd_sc_hd__o21a_1
X_4618_ _3167_ _3744_ _3749_ _3771_ _3772_ vssd1 vssd1 vccd1 vccd1 _3773_ sky130_fd_sc_hd__a2111oi_2
X_8386_ _2621_ _3586_ _3592_ _3598_ vssd1 vssd1 vccd1 vccd1 _3599_ sky130_fd_sc_hd__o211a_1
X_5598_ _0523_ _0529_ _0515_ vssd1 vssd1 vccd1 vccd1 _0571_ sky130_fd_sc_hd__mux2_1
XFILLER_104_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4549_ _3701_ _3703_ vssd1 vssd1 vccd1 vccd1 _3704_ sky130_fd_sc_hd__nor2_1
X_7337_ _2456_ _2457_ vssd1 vssd1 vccd1 vccd1 _2458_ sky130_fd_sc_hd__nor2_1
XFILLER_89_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7268_ _0374_ _2341_ vssd1 vssd1 vccd1 vccd1 _2382_ sky130_fd_sc_hd__xnor2_2
XFILLER_104_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6219_ _0892_ _1168_ vssd1 vssd1 vccd1 vccd1 _1228_ sky130_fd_sc_hd__or2_1
XFILLER_89_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5467__A1 _4250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8405__A1 _0600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7199_ _2279_ _2282_ _2305_ vssd1 vssd1 vccd1 vccd1 _2306_ sky130_fd_sc_hd__o21ai_1
XFILLER_58_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6427__B _0147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6443__A _4217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_584 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5394__B1 _3729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6570_ _1612_ _1613_ vssd1 vssd1 vccd1 vccd1 _1614_ sky130_fd_sc_hd__and2b_1
X_5521_ _0456_ _0493_ _0468_ vssd1 vssd1 vccd1 vccd1 _0494_ sky130_fd_sc_hd__a21o_2
XFILLER_118_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8240_ _3182_ _3396_ _3442_ _3443_ _3303_ vssd1 vssd1 vccd1 vccd1 _3444_ sky130_fd_sc_hd__a311o_1
XANTENNA__4601__A _3735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5452_ _0423_ _0424_ vssd1 vssd1 vccd1 vccd1 _0425_ sky130_fd_sc_hd__nor2_2
XFILLER_117_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4403_ _2012_ _2111_ _2210_ vssd1 vssd1 vccd1 vccd1 _2221_ sky130_fd_sc_hd__a21o_2
X_5383_ _3754_ _0355_ _3721_ vssd1 vssd1 vccd1 vccd1 _0356_ sky130_fd_sc_hd__mux2_4
X_8171_ _3025_ _3230_ _3028_ vssd1 vssd1 vccd1 vccd1 _3370_ sky130_fd_sc_hd__a21o_1
XFILLER_99_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7122_ _2213_ _2215_ vssd1 vssd1 vccd1 vccd1 _2222_ sky130_fd_sc_hd__or2_1
X_4334_ posit_add.in2\[9\] posit_add.in2\[8\] posit_add.in2\[10\] vssd1 vssd1 vccd1
+ vccd1 _1462_ sky130_fd_sc_hd__or3_1
X_7053_ _2088_ _2107_ vssd1 vssd1 vccd1 vccd1 _2146_ sky130_fd_sc_hd__xnor2_1
XFILLER_87_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6004_ _0996_ _0998_ _0995_ vssd1 vssd1 vccd1 vccd1 _1001_ sky130_fd_sc_hd__a21oi_1
X_4265_ in_reg\[0\] cmd\[0\] _0712_ vssd1 vssd1 vccd1 vccd1 _0723_ sky130_fd_sc_hd__mux2_1
XANTENNA__6247__B _1164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5151__B _3763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7955_ _3044_ _3115_ _3137_ _3059_ vssd1 vssd1 vccd1 vccd1 _3138_ sky130_fd_sc_hd__a211o_1
X_6906_ _1978_ _1980_ vssd1 vssd1 vccd1 vccd1 _1984_ sky130_fd_sc_hd__nor2_1
XFILLER_70_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7886_ _3059_ _3061_ vssd1 vssd1 vccd1 vccd1 _3062_ sky130_fd_sc_hd__nor2_1
X_6837_ _4217_ _1813_ _1907_ vssd1 vssd1 vccd1 vccd1 _1908_ sky130_fd_sc_hd__a21oi_1
XFILLER_50_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8507_ _3693_ vssd1 vssd1 vccd1 vccd1 _0071_ sky130_fd_sc_hd__clkbuf_1
X_6768_ _1798_ _1799_ vssd1 vssd1 vccd1 vccd1 _1832_ sky130_fd_sc_hd__nand2_1
XFILLER_10_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5719_ _3699_ _3718_ vssd1 vssd1 vccd1 vccd1 _0698_ sky130_fd_sc_hd__nand2_1
XANTENNA__7126__A1 _1782_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6699_ _1738_ _1744_ _1755_ vssd1 vssd1 vccd1 vccd1 _1756_ sky130_fd_sc_hd__a21o_1
XFILLER_6_219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8323__B1 _1308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8438_ counter\[3\] counter\[2\] _3644_ vssd1 vssd1 vccd1 vccd1 _3648_ sky130_fd_sc_hd__and3_1
X_8369_ _2604_ _3579_ _3502_ _3528_ _3568_ vssd1 vssd1 vccd1 vccd1 _3580_ sky130_fd_sc_hd__o2111a_1
XFILLER_104_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6438__A _4232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5342__A _2540_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7269__A _2381_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_252 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4952_ _4101_ _4103_ vssd1 vssd1 vccd1 vccd1 _4107_ sky130_fd_sc_hd__xnor2_1
XFILLER_51_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7740_ _2726_ _2900_ vssd1 vssd1 vccd1 vccd1 _2901_ sky130_fd_sc_hd__xnor2_1
X_4883_ _2540_ _4037_ vssd1 vssd1 vccd1 vccd1 _4038_ sky130_fd_sc_hd__nor2_1
X_7671_ _2824_ _2752_ vssd1 vssd1 vccd1 vccd1 _2825_ sky130_fd_sc_hd__or2_1
XANTENNA__8502__S _3676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6622_ _1423_ _1401_ vssd1 vssd1 vccd1 vccd1 _1672_ sky130_fd_sc_hd__or2_1
XFILLER_32_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6553_ _1400_ vssd1 vssd1 vccd1 vccd1 _1596_ sky130_fd_sc_hd__inv_2
XFILLER_118_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6484_ _1404_ _1433_ vssd1 vssd1 vccd1 vccd1 _1520_ sky130_fd_sc_hd__xor2_1
X_5504_ _0475_ _0476_ _0469_ vssd1 vssd1 vccd1 vccd1 _0477_ sky130_fd_sc_hd__mux2_1
XFILLER_118_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8223_ _3380_ _3386_ vssd1 vssd1 vccd1 vccd1 _3426_ sky130_fd_sc_hd__nor2_1
X_5435_ _0343_ vssd1 vssd1 vccd1 vccd1 _0408_ sky130_fd_sc_hd__inv_2
XFILLER_10_49 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8154_ _2522_ _2613_ _3204_ vssd1 vssd1 vccd1 vccd1 _3352_ sky130_fd_sc_hd__o21a_1
X_5366_ _4152_ _4209_ _0338_ vssd1 vssd1 vccd1 vccd1 _0339_ sky130_fd_sc_hd__mux2_1
XFILLER_113_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7105_ _2182_ _2197_ _2202_ vssd1 vssd1 vccd1 vccd1 _2203_ sky130_fd_sc_hd__nand3_1
X_4317_ _1264_ vssd1 vssd1 vccd1 vccd1 _1275_ sky130_fd_sc_hd__buf_4
X_5297_ _0252_ _0269_ vssd1 vssd1 vccd1 vccd1 _0270_ sky130_fd_sc_hd__xnor2_1
X_8085_ _3227_ _3271_ _3277_ vssd1 vssd1 vccd1 vccd1 _3279_ sky130_fd_sc_hd__or3_1
XFILLER_113_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7036_ _2051_ _2095_ vssd1 vssd1 vccd1 vccd1 _2127_ sky130_fd_sc_hd__and2_1
XFILLER_87_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7938_ _3113_ _3118_ _2842_ vssd1 vssd1 vccd1 vccd1 _3119_ sky130_fd_sc_hd__mux2_1
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7869_ _3037_ _3041_ _3042_ vssd1 vssd1 vccd1 vccd1 _3043_ sky130_fd_sc_hd__mux2_1
XANTENNA__6721__A _1400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_3__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_51_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5056__B _3615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7271__B _2354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6086__A1 _3770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5220_ _0174_ _0173_ vssd1 vssd1 vccd1 vccd1 _0193_ sky130_fd_sc_hd__and2b_1
XFILLER_102_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5151_ _3827_ _3763_ vssd1 vssd1 vccd1 vccd1 _0124_ sky130_fd_sc_hd__or2_1
XFILLER_111_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5082_ _4234_ _4236_ vssd1 vssd1 vccd1 vccd1 _4237_ sky130_fd_sc_hd__nor2_1
XFILLER_96_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7577__A1 _4217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5984_ _0971_ _0977_ _0978_ vssd1 vssd1 vccd1 vccd1 _0980_ sky130_fd_sc_hd__o21bai_1
X_7723_ _2845_ _2880_ _2882_ vssd1 vssd1 vccd1 vccd1 _2883_ sky130_fd_sc_hd__a21o_1
X_4935_ _4045_ _4089_ vssd1 vssd1 vccd1 vccd1 _4090_ sky130_fd_sc_hd__nand2_1
XFILLER_40_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4866_ _3701_ _3930_ _4019_ vssd1 vssd1 vccd1 vccd1 _4021_ sky130_fd_sc_hd__o21ai_1
XFILLER_20_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7654_ _2712_ _2785_ vssd1 vssd1 vccd1 vccd1 _2807_ sky130_fd_sc_hd__nand2_1
X_4797_ _3950_ _3940_ vssd1 vssd1 vccd1 vccd1 _3952_ sky130_fd_sc_hd__or2b_1
X_6605_ _1619_ _1652_ vssd1 vssd1 vccd1 vccd1 _1653_ sky130_fd_sc_hd__or2_1
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7585_ _2730_ vssd1 vssd1 vccd1 vccd1 _2731_ sky130_fd_sc_hd__buf_2
XANTENNA__5760__B1 _3762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6536_ _1573_ _1574_ vssd1 vssd1 vccd1 vccd1 _1577_ sky130_fd_sc_hd__nor2_1
XFILLER_21_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6467_ _1499_ _1500_ vssd1 vssd1 vccd1 vccd1 _1501_ sky130_fd_sc_hd__nand2_1
X_6398_ _1411_ _1415_ _1419_ _1424_ vssd1 vssd1 vccd1 vccd1 _1425_ sky130_fd_sc_hd__o22a_1
X_8206_ _3402_ _3405_ _3407_ vssd1 vssd1 vccd1 vccd1 _3408_ sky130_fd_sc_hd__a21o_1
X_5418_ _0390_ vssd1 vssd1 vccd1 vccd1 _0391_ sky130_fd_sc_hd__inv_2
XFILLER_99_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4866__A2 _3930_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5349_ _0319_ _0321_ _0317_ vssd1 vssd1 vccd1 vccd1 _0322_ sky130_fd_sc_hd__o21ai_1
X_8137_ _3331_ _3332_ vssd1 vssd1 vccd1 vccd1 _3334_ sky130_fd_sc_hd__or2_1
XFILLER_87_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8068_ _0440_ _0398_ _0515_ vssd1 vssd1 vccd1 vccd1 _3260_ sky130_fd_sc_hd__mux2_1
X_7019_ _2106_ _2105_ vssd1 vssd1 vccd1 vccd1 _2108_ sky130_fd_sc_hd__or2b_1
XFILLER_101_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6716__A _0080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6435__B _0303_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5751__B1 _3762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4306__A1 in_reg\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6626__A _3703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8508__A0 posit_add.in2\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6361__A _3615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4720_ _3874_ vssd1 vssd1 vccd1 vccd1 _3875_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4651_ _3800_ _3703_ _3805_ vssd1 vssd1 vccd1 vccd1 _3806_ sky130_fd_sc_hd__o21ai_1
XFILLER_116_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4582_ _3736_ _2309_ _3729_ _3696_ vssd1 vssd1 vccd1 vccd1 _3737_ sky130_fd_sc_hd__or4b_1
X_7370_ _2493_ vssd1 vssd1 vccd1 vccd1 _2494_ sky130_fd_sc_hd__buf_2
XFILLER_115_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6321_ _1097_ _0994_ _1339_ vssd1 vssd1 vccd1 vccd1 _1340_ sky130_fd_sc_hd__a21o_1
XFILLER_115_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6252_ _1241_ _1240_ _1239_ vssd1 vssd1 vccd1 vccd1 _1265_ sky130_fd_sc_hd__a21o_1
XANTENNA__7495__B1 _1803_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6183_ _1172_ _1187_ _1189_ vssd1 vssd1 vccd1 vccd1 _1190_ sky130_fd_sc_hd__a21oi_1
X_5203_ _3800_ _3840_ _0152_ vssd1 vssd1 vccd1 vccd1 _0176_ sky130_fd_sc_hd__o21a_1
X_5134_ _3925_ _3615_ _0105_ vssd1 vssd1 vccd1 vccd1 _0107_ sky130_fd_sc_hd__o21ai_1
XFILLER_69_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5065_ _4210_ _4037_ vssd1 vssd1 vccd1 vccd1 _4220_ sky130_fd_sc_hd__or2_1
XFILLER_53_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8211__A2 _3411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5967_ _0942_ _0960_ _0961_ vssd1 vssd1 vccd1 vccd1 _0962_ sky130_fd_sc_hd__a21oi_2
XFILLER_12_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_468 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4918_ _3739_ _3702_ vssd1 vssd1 vccd1 vccd1 _4073_ sky130_fd_sc_hd__nor2_1
X_7706_ _2743_ _2757_ _2863_ vssd1 vssd1 vccd1 vccd1 _2864_ sky130_fd_sc_hd__o21ai_2
X_5898_ _3815_ _0787_ vssd1 vssd1 vccd1 vccd1 _0890_ sky130_fd_sc_hd__nor2_1
XFILLER_21_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7637_ _2675_ _2748_ _2709_ _2787_ vssd1 vssd1 vccd1 vccd1 _2788_ sky130_fd_sc_hd__a31o_1
X_4849_ _4002_ _4003_ vssd1 vssd1 vccd1 vccd1 _4004_ sky130_fd_sc_hd__or2_1
XFILLER_21_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7568_ _2702_ _2706_ vssd1 vssd1 vccd1 vccd1 _2712_ sky130_fd_sc_hd__nand2_2
XFILLER_106_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6519_ _1555_ _1556_ vssd1 vssd1 vccd1 vccd1 _1558_ sky130_fd_sc_hd__nand2_1
X_7499_ _2859_ _2629_ _2634_ _2635_ vssd1 vssd1 vccd1 vccd1 _2636_ sky130_fd_sc_hd__o22a_1
XFILLER_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7277__A _2349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6870_ _1933_ _1942_ _1943_ vssd1 vssd1 vccd1 vccd1 _1944_ sky130_fd_sc_hd__o21ai_1
X_5821_ _0772_ _0774_ _0775_ _0771_ vssd1 vssd1 vccd1 vccd1 _0807_ sky130_fd_sc_hd__o2bb2ai_1
X_5752_ _0365_ _3901_ _2529_ _3866_ vssd1 vssd1 vccd1 vccd1 _0734_ sky130_fd_sc_hd__a211o_1
X_8540_ clknet_3_1__leaf_clk _0026_ vssd1 vssd1 vccd1 vccd1 out_reg\[6\] sky130_fd_sc_hd__dfxtp_1
X_4703_ _3816_ _3795_ vssd1 vssd1 vccd1 vccd1 _3858_ sky130_fd_sc_hd__nor2_1
X_5683_ _3762_ _0655_ _0656_ _0658_ vssd1 vssd1 vccd1 vccd1 _0659_ sky130_fd_sc_hd__o211a_1
X_8471_ in_reg\[12\] posit_add.in1\[12\] _3654_ vssd1 vssd1 vccd1 vccd1 _3670_ sky130_fd_sc_hd__mux2_1
XANTENNA__8510__S _3676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7422_ _2242_ _2181_ vssd1 vssd1 vccd1 vccd1 _2552_ sky130_fd_sc_hd__or2b_1
X_4634_ _3721_ _3776_ _3788_ vssd1 vssd1 vccd1 vccd1 _3789_ sky130_fd_sc_hd__and3_1
X_4565_ _2793_ _3134_ _2617_ vssd1 vssd1 vccd1 vccd1 _3720_ sky130_fd_sc_hd__or3b_1
X_7353_ _2444_ _2471_ vssd1 vssd1 vccd1 vccd1 _2476_ sky130_fd_sc_hd__nand2_1
X_6304_ _1315_ _1320_ _1312_ vssd1 vssd1 vccd1 vccd1 _1322_ sky130_fd_sc_hd__o21ai_1
XFILLER_116_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4496_ _3210_ _3232_ _2606_ vssd1 vssd1 vccd1 vccd1 _3243_ sky130_fd_sc_hd__mux2_1
X_7284_ _2384_ _2354_ _2376_ _2350_ vssd1 vssd1 vccd1 vccd1 _2400_ sky130_fd_sc_hd__o2bb2a_1
X_6235_ _1244_ _1243_ vssd1 vssd1 vccd1 vccd1 _1246_ sky130_fd_sc_hd__or2b_1
XFILLER_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6166_ _1168_ _1170_ vssd1 vssd1 vccd1 vccd1 _1171_ sky130_fd_sc_hd__and2b_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6097_ _0884_ _0981_ _0987_ vssd1 vssd1 vccd1 vccd1 _1099_ sky130_fd_sc_hd__a21oi_1
XFILLER_57_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5117_ _0079_ _0089_ vssd1 vssd1 vccd1 vccd1 _0090_ sky130_fd_sc_hd__nor2_1
X_5048_ _4045_ _4153_ _4202_ vssd1 vssd1 vccd1 vccd1 _4203_ sky130_fd_sc_hd__and3_1
XANTENNA__5246__A2 _3901_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7640__A0 _1531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8481__A _3676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6999_ _1456_ _1717_ vssd1 vssd1 vccd1 vccd1 _2086_ sky130_fd_sc_hd__or2_1
XFILLER_13_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5064__B _3840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5080__A _4210_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5239__B _3986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4350_ _1616_ _1627_ vssd1 vssd1 vccd1 vccd1 _1638_ sky130_fd_sc_hd__nor2_2
XFILLER_113_524 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4920__B2 _3792_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4281_ _0883_ vssd1 vssd1 vccd1 vccd1 _0005_ sky130_fd_sc_hd__clkbuf_1
XFILLER_4_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6020_ _1008_ _1016_ _1017_ vssd1 vssd1 vccd1 vccd1 _1018_ sky130_fd_sc_hd__o21ai_1
XFILLER_101_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7971_ _3097_ _3125_ _3065_ vssd1 vssd1 vccd1 vccd1 _3155_ sky130_fd_sc_hd__mux2_1
XANTENNA__4318__B _1275_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6922_ _1886_ _1892_ _1894_ vssd1 vssd1 vccd1 vccd1 _2002_ sky130_fd_sc_hd__and3_1
XFILLER_47_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6853_ _1918_ _1919_ vssd1 vssd1 vccd1 vccd1 _1926_ sky130_fd_sc_hd__nand2_1
X_5804_ _3735_ _0757_ _0788_ vssd1 vssd1 vccd1 vccd1 _0789_ sky130_fd_sc_hd__o21ai_1
XFILLER_90_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6784_ _1413_ _4089_ vssd1 vssd1 vccd1 vccd1 _1850_ sky130_fd_sc_hd__nand2_1
XFILLER_22_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5735_ _3775_ _0633_ _0631_ _4044_ vssd1 vssd1 vccd1 vccd1 _0716_ sky130_fd_sc_hd__a22o_1
X_8523_ clknet_3_3__leaf_clk _0009_ vssd1 vssd1 vccd1 vccd1 in_reg\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_50_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5149__B _0121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5666_ _0633_ _3878_ _0631_ _3892_ vssd1 vssd1 vccd1 vccd1 _0640_ sky130_fd_sc_hd__a22o_1
X_8454_ _3660_ vssd1 vssd1 vccd1 vccd1 _0046_ sky130_fd_sc_hd__clkbuf_1
X_7405_ _2530_ _2532_ _2412_ vssd1 vssd1 vccd1 vccd1 _2533_ sky130_fd_sc_hd__a21oi_1
X_4617_ _3594_ vssd1 vssd1 vccd1 vccd1 _3772_ sky130_fd_sc_hd__buf_4
XANTENNA__5165__A _3855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8385_ _3182_ _3565_ _3595_ _3597_ vssd1 vssd1 vccd1 vccd1 _3598_ sky130_fd_sc_hd__a31o_1
X_5597_ _0567_ _0569_ _0494_ vssd1 vssd1 vccd1 vccd1 _0570_ sky130_fd_sc_hd__mux2_1
XFILLER_89_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4548_ _3702_ vssd1 vssd1 vccd1 vccd1 _3703_ sky130_fd_sc_hd__clkbuf_4
X_7336_ _1768_ _2455_ vssd1 vssd1 vccd1 vccd1 _2457_ sky130_fd_sc_hd__and2_1
XFILLER_89_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4479_ _1253_ _3013_ vssd1 vssd1 vccd1 vccd1 _3057_ sky130_fd_sc_hd__nand2_1
X_7267_ _0388_ _2336_ vssd1 vssd1 vccd1 vccd1 _2381_ sky130_fd_sc_hd__xor2_2
X_6218_ _1223_ _1222_ vssd1 vssd1 vccd1 vccd1 _1227_ sky130_fd_sc_hd__xor2_1
XFILLER_77_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5467__A2 _0082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_611 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7198_ _2299_ _2304_ vssd1 vssd1 vccd1 vccd1 _2305_ sky130_fd_sc_hd__xnor2_1
X_6149_ _1143_ _1152_ vssd1 vssd1 vccd1 vccd1 _1153_ sky130_fd_sc_hd__xnor2_1
XFILLER_58_666 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6724__A _1383_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8169__A1 _1330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6443__B _1353_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8341__B2 _3195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5803__A _3924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7604__A0 _3881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6319__D_N _1097_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5520_ _0478_ _0455_ _0453_ vssd1 vssd1 vccd1 vccd1 _0493_ sky130_fd_sc_hd__a21bo_1
XFILLER_117_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4601__B _3739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5451_ _0417_ _0422_ vssd1 vssd1 vccd1 vccd1 _0424_ sky130_fd_sc_hd__and2_1
X_4402_ _2122_ _2166_ _2199_ vssd1 vssd1 vccd1 vccd1 _2210_ sky130_fd_sc_hd__o21ai_2
X_5382_ _3850_ _0354_ _3156_ vssd1 vssd1 vccd1 vccd1 _0355_ sky130_fd_sc_hd__mux2_1
X_8170_ _1330_ _3359_ _3367_ _3368_ _0600_ vssd1 vssd1 vccd1 vccd1 _3369_ sky130_fd_sc_hd__a311o_1
X_7121_ _2218_ _2219_ vssd1 vssd1 vccd1 vccd1 _2220_ sky130_fd_sc_hd__nor2_1
X_4333_ posit_add.in2\[12\] _1440_ vssd1 vssd1 vccd1 vccd1 _1451_ sky130_fd_sc_hd__xnor2_4
XFILLER_113_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7052_ _2104_ _2139_ _2140_ _2142_ _2143_ vssd1 vssd1 vccd1 vccd1 _2145_ sky130_fd_sc_hd__a32o_1
XFILLER_101_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4264_ _0635_ _0690_ _0701_ vssd1 vssd1 vccd1 vccd1 _0712_ sky130_fd_sc_hd__or3b_2
XFILLER_113_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6003_ _0999_ vssd1 vssd1 vccd1 vccd1 _1000_ sky130_fd_sc_hd__clkbuf_2
XFILLER_39_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4329__A posit_add.in2\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8399__A1 _2993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7954_ _3136_ vssd1 vssd1 vccd1 vccd1 _3137_ sky130_fd_sc_hd__inv_2
XFILLER_27_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6905_ _1982_ _1960_ vssd1 vssd1 vccd1 vccd1 _1983_ sky130_fd_sc_hd__xnor2_1
XFILLER_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7885_ _3060_ _3045_ _3044_ vssd1 vssd1 vccd1 vccd1 _3061_ sky130_fd_sc_hd__mux2_1
XFILLER_23_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6836_ _3840_ _1664_ vssd1 vssd1 vccd1 vccd1 _1907_ sky130_fd_sc_hd__nor2_1
XFILLER_50_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6767_ _1774_ _1830_ vssd1 vssd1 vccd1 vccd1 _1831_ sky130_fd_sc_hd__or2b_1
XFILLER_23_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5718_ _3762_ _0614_ vssd1 vssd1 vccd1 vccd1 _0697_ sky130_fd_sc_hd__nor2_1
X_8506_ posit_add.in2\[12\] in_reg\[12\] _3676_ vssd1 vssd1 vccd1 vccd1 _3693_ sky130_fd_sc_hd__mux2_1
XFILLER_10_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7375__A _2335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6698_ _1735_ _1736_ vssd1 vssd1 vccd1 vccd1 _1755_ sky130_fd_sc_hd__nor2_1
X_5649_ _3717_ _0607_ _3699_ vssd1 vssd1 vccd1 vccd1 _0622_ sky130_fd_sc_hd__a21o_1
X_8437_ counter\[2\] _3644_ _3647_ vssd1 vssd1 vccd1 vccd1 _0040_ sky130_fd_sc_hd__a21oi_1
XFILLER_117_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8368_ _2569_ _3352_ _3286_ vssd1 vssd1 vccd1 vccd1 _3579_ sky130_fd_sc_hd__o21a_1
X_7319_ _2256_ _2258_ vssd1 vssd1 vccd1 vccd1 _2438_ sky130_fd_sc_hd__xnor2_2
XFILLER_104_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7314__S _2416_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8299_ _3481_ _3499_ _3505_ vssd1 vssd1 vccd1 vccd1 _3506_ sky130_fd_sc_hd__o21ai_1
XANTENNA__5342__B _3988_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7269__B _2382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6364__A _0627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4951_ _4074_ _4105_ vssd1 vssd1 vccd1 vccd1 _4106_ sky130_fd_sc_hd__nor2_1
XFILLER_45_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4882_ _3750_ vssd1 vssd1 vccd1 vccd1 _4037_ sky130_fd_sc_hd__clkbuf_4
XFILLER_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7670_ _2743_ _2750_ vssd1 vssd1 vccd1 vccd1 _2824_ sky130_fd_sc_hd__nand2_1
X_6621_ _1655_ _1668_ _1669_ vssd1 vssd1 vccd1 vccd1 _1670_ sky130_fd_sc_hd__o21ba_1
XFILLER_32_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6552_ _1593_ _1475_ vssd1 vssd1 vccd1 vccd1 _1595_ sky130_fd_sc_hd__and2b_1
XFILLER_118_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6483_ _1516_ _1518_ vssd1 vssd1 vccd1 vccd1 _1519_ sky130_fd_sc_hd__nor2_1
XANTENNA__5427__B _4210_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5503_ _0474_ _4152_ _0337_ vssd1 vssd1 vccd1 vccd1 _0476_ sky130_fd_sc_hd__mux2_1
XFILLER_106_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5434_ _3424_ _3530_ _2980_ vssd1 vssd1 vccd1 vccd1 _0407_ sky130_fd_sc_hd__a21o_1
X_8222_ _3422_ _3423_ vssd1 vssd1 vccd1 vccd1 _3425_ sky130_fd_sc_hd__or2_1
XFILLER_10_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8153_ _3289_ _3321_ _3284_ vssd1 vssd1 vccd1 vccd1 _3351_ sky130_fd_sc_hd__or3b_1
XFILLER_99_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7104_ _2198_ _2200_ _2201_ vssd1 vssd1 vccd1 vccd1 _2202_ sky130_fd_sc_hd__or3_1
X_5365_ _0337_ vssd1 vssd1 vccd1 vccd1 _0338_ sky130_fd_sc_hd__clkbuf_4
XFILLER_101_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5296_ _0255_ _0268_ vssd1 vssd1 vccd1 vccd1 _0269_ sky130_fd_sc_hd__and2_1
X_4316_ posit_add.in2\[15\] vssd1 vssd1 vccd1 vccd1 _1264_ sky130_fd_sc_hd__buf_2
X_8084_ _3227_ _3271_ _3277_ vssd1 vssd1 vccd1 vccd1 _3278_ sky130_fd_sc_hd__o21ai_1
X_7035_ _2095_ _2125_ vssd1 vssd1 vccd1 vccd1 _2126_ sky130_fd_sc_hd__or2_1
XFILLER_19_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8241__B1 _3195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7089__B _1782_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7937_ _3117_ _3048_ _2937_ vssd1 vssd1 vccd1 vccd1 _3118_ sky130_fd_sc_hd__mux2_1
XFILLER_70_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7868_ _2842_ vssd1 vssd1 vccd1 vccd1 _3042_ sky130_fd_sc_hd__clkbuf_4
XFILLER_35_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6819_ _1886_ _1887_ vssd1 vssd1 vccd1 vccd1 _1888_ sky130_fd_sc_hd__nand2_1
XFILLER_11_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6721__B _0548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7799_ _2965_ _2915_ _2908_ vssd1 vssd1 vccd1 vccd1 _2966_ sky130_fd_sc_hd__a21oi_1
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6086__A2 _3739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_672 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4432__A _2529_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5150_ _0120_ _0122_ vssd1 vssd1 vccd1 vccd1 _0123_ sky130_fd_sc_hd__or2b_1
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5081_ _4222_ _3855_ _4235_ vssd1 vssd1 vccd1 vccd1 _4236_ sky130_fd_sc_hd__a21oi_1
XFILLER_110_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_388 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6094__A _0762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5983_ _0977_ _0978_ vssd1 vssd1 vccd1 vccd1 _0979_ sky130_fd_sc_hd__or2_1
XFILLER_64_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4934_ _3883_ vssd1 vssd1 vccd1 vccd1 _4089_ sky130_fd_sc_hd__buf_4
XFILLER_24_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7722_ _2743_ _2757_ _2759_ vssd1 vssd1 vccd1 vccd1 _2882_ sky130_fd_sc_hd__a21oi_1
X_4865_ _3701_ _3930_ _4019_ vssd1 vssd1 vccd1 vccd1 _4020_ sky130_fd_sc_hd__or3_1
X_7653_ _2708_ _2791_ _2805_ vssd1 vssd1 vccd1 vccd1 _2806_ sky130_fd_sc_hd__o21ai_1
X_4796_ _3940_ _3950_ vssd1 vssd1 vccd1 vccd1 _3951_ sky130_fd_sc_hd__xnor2_1
X_6604_ _1620_ _1651_ vssd1 vssd1 vccd1 vccd1 _1652_ sky130_fd_sc_hd__xnor2_1
X_7584_ _2702_ _2706_ vssd1 vssd1 vccd1 vccd1 _2730_ sky130_fd_sc_hd__and2_1
X_6535_ _1543_ _1563_ vssd1 vssd1 vccd1 vccd1 _1576_ sky130_fd_sc_hd__xor2_1
XFILLER_21_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7501__A2 _1682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6466_ _1497_ _4211_ _1449_ vssd1 vssd1 vccd1 vccd1 _1500_ sky130_fd_sc_hd__or3_1
X_8205_ _3289_ _3406_ _3284_ vssd1 vssd1 vccd1 vccd1 _3407_ sky130_fd_sc_hd__and3b_1
X_6397_ _1420_ _1423_ vssd1 vssd1 vccd1 vccd1 _1424_ sky130_fd_sc_hd__or2_2
XANTENNA__5173__A _3802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5417_ _0386_ _0389_ vssd1 vssd1 vccd1 vccd1 _0390_ sky130_fd_sc_hd__or2_2
XFILLER_114_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5348_ _4207_ _4208_ _0320_ vssd1 vssd1 vccd1 vccd1 _0321_ sky130_fd_sc_hd__a21oi_1
X_8136_ _3331_ _3332_ vssd1 vssd1 vccd1 vccd1 _3333_ sky130_fd_sc_hd__nand2_1
XFILLER_102_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8067_ _0519_ vssd1 vssd1 vccd1 vccd1 _3259_ sky130_fd_sc_hd__clkbuf_4
X_7018_ _2105_ _2106_ vssd1 vssd1 vccd1 vccd1 _2107_ sky130_fd_sc_hd__xnor2_1
XFILLER_87_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5279_ _0238_ _0251_ vssd1 vssd1 vccd1 vccd1 _0252_ sky130_fd_sc_hd__nand2_1
XANTENNA__6716__B _1718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5579__A1 _3878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7563__A _2702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8453__A0 in_reg\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7223__A_N _0698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4650_ _3802_ _3804_ vssd1 vssd1 vccd1 vccd1 _3805_ sky130_fd_sc_hd__nand2_1
XFILLER_14_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5742__A1 _3901_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5742__B2 _0113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6320_ _0762_ _0993_ _0994_ _0722_ vssd1 vssd1 vccd1 vccd1 _1339_ sky130_fd_sc_hd__a22o_1
X_4581_ _2485_ vssd1 vssd1 vccd1 vccd1 _3736_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__8149__B1_N _1177_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6251_ _1241_ _1239_ _1240_ vssd1 vssd1 vccd1 vccd1 _1263_ sky130_fd_sc_hd__nand3_1
XANTENNA__7495__B2 _3189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6182_ _1184_ _1186_ vssd1 vssd1 vccd1 vccd1 _1189_ sky130_fd_sc_hd__nor2_1
XFILLER_88_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5202_ _0173_ _0174_ vssd1 vssd1 vccd1 vccd1 _0175_ sky130_fd_sc_hd__and2b_1
XFILLER_69_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5133_ _3925_ _3615_ _0105_ vssd1 vssd1 vccd1 vccd1 _0106_ sky130_fd_sc_hd__or3_1
XFILLER_111_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8508__S _3676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5064_ _4210_ _3840_ vssd1 vssd1 vccd1 vccd1 _4219_ sky130_fd_sc_hd__or2_1
XFILLER_84_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5966_ _0921_ _0922_ _0941_ vssd1 vssd1 vccd1 vccd1 _0961_ sky130_fd_sc_hd__and3_1
XFILLER_80_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5430__B1 _1748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5897_ _0885_ _0888_ vssd1 vssd1 vccd1 vccd1 _0889_ sky130_fd_sc_hd__nand2_1
X_4917_ _4056_ _4061_ vssd1 vssd1 vccd1 vccd1 _4072_ sky130_fd_sc_hd__xnor2_1
X_7705_ _2704_ _2794_ _2852_ _2862_ _2762_ vssd1 vssd1 vccd1 vccd1 _2863_ sky130_fd_sc_hd__a221o_1
XFILLER_33_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4848_ _3999_ _4000_ _4001_ vssd1 vssd1 vccd1 vccd1 _4003_ sky130_fd_sc_hd__a21oi_1
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7636_ _2676_ _2747_ _2786_ _2704_ _2743_ vssd1 vssd1 vccd1 vccd1 _2787_ sky130_fd_sc_hd__o221a_1
XFILLER_21_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4779_ _3915_ _3916_ _3932_ vssd1 vssd1 vccd1 vccd1 _3934_ sky130_fd_sc_hd__and3_1
XANTENNA__4536__A2 _3635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7567_ _2319_ _2708_ vssd1 vssd1 vccd1 vccd1 _2711_ sky130_fd_sc_hd__nand2_1
XFILLER_119_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6518_ _1555_ _1556_ vssd1 vssd1 vccd1 vccd1 _1557_ sky130_fd_sc_hd__xnor2_1
X_7498_ _2859_ _2629_ _1858_ _2903_ vssd1 vssd1 vccd1 vccd1 _2635_ sky130_fd_sc_hd__a22o_1
X_6449_ _1427_ _1430_ _1426_ _1431_ vssd1 vssd1 vccd1 vccd1 _1481_ sky130_fd_sc_hd__a22o_1
XFILLER_106_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8119_ _0701_ _0786_ vssd1 vssd1 vccd1 vccd1 _3315_ sky130_fd_sc_hd__and2_1
XFILLER_102_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7410__B2 _2416_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5078__A _4228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7477__A1 _2381_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5820_ _0803_ _0805_ vssd1 vssd1 vccd1 vccd1 _0806_ sky130_fd_sc_hd__xnor2_1
XFILLER_62_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5751_ _0666_ _0732_ _3762_ vssd1 vssd1 vccd1 vccd1 _0733_ sky130_fd_sc_hd__a21o_1
XFILLER_62_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8470_ _3669_ vssd1 vssd1 vccd1 vccd1 _0054_ sky130_fd_sc_hd__clkbuf_1
X_4702_ _3844_ _3854_ _3856_ vssd1 vssd1 vccd1 vccd1 _3857_ sky130_fd_sc_hd__o21ba_1
X_7421_ _2545_ _2547_ _2549_ vssd1 vssd1 vccd1 vccd1 _2550_ sky130_fd_sc_hd__or3b_1
X_5682_ _0604_ _0607_ _0112_ vssd1 vssd1 vccd1 vccd1 _0658_ sky130_fd_sc_hd__a21oi_1
X_4633_ _3156_ _3783_ _3785_ _3787_ vssd1 vssd1 vccd1 vccd1 _3788_ sky130_fd_sc_hd__a31o_1
XFILLER_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4564_ _3718_ vssd1 vssd1 vccd1 vccd1 _3719_ sky130_fd_sc_hd__clkbuf_4
X_7352_ _2425_ _2426_ _2427_ _2473_ vssd1 vssd1 vccd1 vccd1 _2475_ sky130_fd_sc_hd__a31o_1
XFILLER_116_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6303_ _1312_ _1315_ _1320_ vssd1 vssd1 vccd1 vccd1 _1321_ sky130_fd_sc_hd__nor3_1
X_7283_ _2385_ _2388_ _2398_ _2392_ vssd1 vssd1 vccd1 vccd1 _2399_ sky130_fd_sc_hd__o211ai_4
X_6234_ _1243_ _1244_ vssd1 vssd1 vccd1 vccd1 _1245_ sky130_fd_sc_hd__xor2_1
XFILLER_89_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4495_ posit_add.in1\[1\] _3221_ vssd1 vssd1 vccd1 vccd1 _3232_ sky130_fd_sc_hd__xnor2_4
XANTENNA__5479__B1 _0451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6165_ _1163_ _1169_ vssd1 vssd1 vccd1 vccd1 _1170_ sky130_fd_sc_hd__xnor2_1
XANTENNA__4766__S _3830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6096_ _1053_ _1078_ _1092_ _1090_ _1089_ vssd1 vssd1 vccd1 vccd1 _1098_ sky130_fd_sc_hd__a2111o_1
XFILLER_97_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5116_ _0086_ _0088_ vssd1 vssd1 vccd1 vccd1 _0089_ sky130_fd_sc_hd__xor2_1
XFILLER_111_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5047_ _4199_ _4201_ vssd1 vssd1 vccd1 vccd1 _4202_ sky130_fd_sc_hd__xor2_1
XANTENNA__7640__A1 _3878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6998_ _2083_ _2084_ vssd1 vssd1 vccd1 vccd1 _2085_ sky130_fd_sc_hd__nor2_2
XFILLER_53_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5949_ _0927_ _0940_ _0939_ vssd1 vssd1 vccd1 vccd1 _0943_ sky130_fd_sc_hd__nand3_1
XFILLER_40_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7619_ _2762_ _2767_ vssd1 vssd1 vccd1 vccd1 _2768_ sky130_fd_sc_hd__or2_1
XFILLER_107_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5626__A _0092_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8002__A cmd\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5999__C _0702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7560__B _2702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5080__B _3840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6904__B _0548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4920__A2 _3771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4280_ in_reg\[1\] in_reg\[2\] _0830_ vssd1 vssd1 vccd1 vccd1 _0883_ sky130_fd_sc_hd__mux2_1
XFILLER_4_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7970_ _3144_ _3153_ _3025_ vssd1 vssd1 vccd1 vccd1 _3154_ sky130_fd_sc_hd__mux2_1
XFILLER_39_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6921_ _1949_ _1999_ vssd1 vssd1 vccd1 vccd1 _2000_ sky130_fd_sc_hd__and2b_1
XFILLER_47_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4615__A _1748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6852_ _1922_ _1923_ vssd1 vssd1 vccd1 vccd1 _1925_ sky130_fd_sc_hd__xor2_1
XFILLER_81_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5803_ _3924_ _0731_ _0787_ vssd1 vssd1 vccd1 vccd1 _0788_ sky130_fd_sc_hd__or3_1
XFILLER_50_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6783_ _1846_ _1848_ vssd1 vssd1 vccd1 vccd1 _1849_ sky130_fd_sc_hd__xnor2_1
X_8522_ clknet_3_3__leaf_clk _0008_ vssd1 vssd1 vccd1 vccd1 in_reg\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_50_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5734_ _4045_ _0633_ vssd1 vssd1 vccd1 vccd1 _0715_ sky130_fd_sc_hd__nand2_1
XFILLER_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5665_ _0627_ _3734_ _3770_ _0631_ vssd1 vssd1 vccd1 vccd1 _0639_ sky130_fd_sc_hd__or4b_1
X_8453_ in_reg\[3\] posit_add.in1\[3\] _3655_ vssd1 vssd1 vccd1 vccd1 _3660_ sky130_fd_sc_hd__mux2_1
X_7404_ _2245_ _2531_ vssd1 vssd1 vccd1 vccd1 _2532_ sky130_fd_sc_hd__and2_1
X_4616_ _3770_ vssd1 vssd1 vccd1 vccd1 _3771_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__5446__A _1781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8384_ _3190_ _3596_ vssd1 vssd1 vccd1 vccd1 _3597_ sky130_fd_sc_hd__nand2_1
X_7335_ _1768_ _2455_ vssd1 vssd1 vccd1 vccd1 _2456_ sky130_fd_sc_hd__nor2_1
X_5596_ _0568_ _0503_ _0515_ vssd1 vssd1 vccd1 vccd1 _0569_ sky130_fd_sc_hd__mux2_1
XFILLER_116_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4547_ _3541_ _3562_ _3594_ _3520_ vssd1 vssd1 vccd1 vccd1 _3702_ sky130_fd_sc_hd__a211o_4
XFILLER_116_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4478_ _2980_ _3035_ vssd1 vssd1 vccd1 vccd1 _3046_ sky130_fd_sc_hd__xnor2_4
X_7266_ _2343_ _0442_ vssd1 vssd1 vccd1 vccd1 _2380_ sky130_fd_sc_hd__xnor2_1
X_6217_ _1221_ _1224_ _1225_ vssd1 vssd1 vccd1 vccd1 _1226_ sky130_fd_sc_hd__and3_1
XFILLER_104_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7197_ _2302_ _2303_ vssd1 vssd1 vccd1 vccd1 _2304_ sky130_fd_sc_hd__nor2_1
X_6148_ _1150_ _1151_ vssd1 vssd1 vccd1 vccd1 _1152_ sky130_fd_sc_hd__xor2_1
XFILLER_58_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6427__D _1456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4509__B _3232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6079_ _0961_ _0960_ vssd1 vssd1 vccd1 vccd1 _1080_ sky130_fd_sc_hd__nor2_1
XFILLER_58_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6724__B _3703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6443__C _1354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5388__C1 _3736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_634 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7604__A1 _1355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4435__A posit_add.in1\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5394__A2 _3830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5450_ _0417_ _0422_ vssd1 vssd1 vccd1 vccd1 _0423_ sky130_fd_sc_hd__nor2_1
XFILLER_117_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4401_ _2177_ _2188_ _1550_ vssd1 vssd1 vccd1 vccd1 _2199_ sky130_fd_sc_hd__or3_1
XANTENNA__4601__C _3750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5381_ _3068_ _0353_ _3446_ vssd1 vssd1 vccd1 vccd1 _0354_ sky130_fd_sc_hd__mux2_1
XFILLER_113_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7120_ _2202_ _2204_ _2217_ vssd1 vssd1 vccd1 vccd1 _2219_ sky130_fd_sc_hd__a21oi_1
X_4332_ _1341_ _1374_ _1396_ _1264_ vssd1 vssd1 vccd1 vccd1 _1440_ sky130_fd_sc_hd__o31a_1
XFILLER_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7051_ _4089_ _1676_ _1538_ _2086_ vssd1 vssd1 vccd1 vccd1 _2143_ sky130_fd_sc_hd__nor4_1
XFILLER_87_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4263_ net1 vssd1 vssd1 vccd1 vccd1 _0701_ sky130_fd_sc_hd__clkbuf_4
X_6002_ _0995_ _0996_ _0998_ vssd1 vssd1 vccd1 vccd1 _0999_ sky130_fd_sc_hd__and3_1
XFILLER_86_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7953_ _2890_ _2894_ _3034_ vssd1 vssd1 vccd1 vccd1 _3136_ sky130_fd_sc_hd__mux2_1
X_6904_ _1599_ _0548_ vssd1 vssd1 vccd1 vccd1 _1982_ sky130_fd_sc_hd__nor2_1
XANTENNA__4345__A posit_add.in2\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7884_ _2921_ _2924_ _3034_ vssd1 vssd1 vccd1 vccd1 _3060_ sky130_fd_sc_hd__mux2_1
X_6835_ _1454_ _1510_ vssd1 vssd1 vccd1 vccd1 _1906_ sky130_fd_sc_hd__nor2_1
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6766_ _1801_ _1828_ _1829_ vssd1 vssd1 vccd1 vccd1 _1830_ sky130_fd_sc_hd__a21o_1
XFILLER_11_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5717_ _3699_ _0626_ _0695_ _3923_ vssd1 vssd1 vccd1 vccd1 _0696_ sky130_fd_sc_hd__o31a_1
X_8505_ _3692_ vssd1 vssd1 vccd1 vccd1 _0070_ sky130_fd_sc_hd__clkbuf_1
XFILLER_109_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6697_ _1739_ _1743_ _1753_ vssd1 vssd1 vccd1 vccd1 _1754_ sky130_fd_sc_hd__o21ai_1
XFILLER_40_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5648_ _3865_ _0619_ vssd1 vssd1 vccd1 vccd1 _0621_ sky130_fd_sc_hd__nor2_1
X_8436_ counter\[2\] _3644_ _3641_ vssd1 vssd1 vccd1 vccd1 _3647_ sky130_fd_sc_hd__o21ai_1
X_5579_ _3878_ _3804_ _4073_ _0551_ _4122_ vssd1 vssd1 vccd1 vccd1 _0552_ sky130_fd_sc_hd__a2111oi_1
XANTENNA__4896__A1 _3792_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8367_ _3577_ _3578_ _1220_ vssd1 vssd1 vccd1 vccd1 _0032_ sky130_fd_sc_hd__o21ba_1
XANTENNA__5904__A _3770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8298_ _3502_ _3504_ vssd1 vssd1 vccd1 vccd1 _3505_ sky130_fd_sc_hd__and2b_1
X_7318_ _2416_ _2412_ vssd1 vssd1 vccd1 vccd1 _2437_ sky130_fd_sc_hd__or2_2
X_7249_ _2360_ _0415_ vssd1 vssd1 vccd1 vccd1 _2361_ sky130_fd_sc_hd__nor2_1
XFILLER_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_442 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4950_ _3845_ _3795_ _3702_ _3828_ vssd1 vssd1 vccd1 vccd1 _4105_ sky130_fd_sc_hd__o22a_1
X_4881_ _4033_ _4035_ vssd1 vssd1 vccd1 vccd1 _4036_ sky130_fd_sc_hd__xor2_1
XFILLER_17_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6620_ _1355_ _1414_ _1410_ _1384_ vssd1 vssd1 vccd1 vccd1 _1669_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_20_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6551_ _4228_ _1383_ vssd1 vssd1 vccd1 vccd1 _1593_ sky130_fd_sc_hd__or2_1
X_5502_ _0473_ _0474_ _0338_ vssd1 vssd1 vccd1 vccd1 _0475_ sky130_fd_sc_hd__mux2_1
X_6482_ _1511_ _1513_ _1515_ vssd1 vssd1 vccd1 vccd1 _1518_ sky130_fd_sc_hd__a21oi_1
XFILLER_118_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5433_ _3328_ _2826_ _3772_ vssd1 vssd1 vccd1 vccd1 _0406_ sky130_fd_sc_hd__o21ai_1
X_8221_ _0601_ _3421_ _3415_ _2621_ vssd1 vssd1 vccd1 vccd1 _3423_ sky130_fd_sc_hd__a31o_1
XANTENNA__5724__A _3762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8152_ _3322_ _3323_ vssd1 vssd1 vccd1 vccd1 _3350_ sky130_fd_sc_hd__or2b_1
X_5364_ _0099_ _0334_ _0336_ vssd1 vssd1 vccd1 vccd1 _0337_ sky130_fd_sc_hd__a21o_2
X_7103_ _2174_ _2183_ _2196_ vssd1 vssd1 vccd1 vccd1 _2201_ sky130_fd_sc_hd__a21oi_1
X_4315_ _1242_ vssd1 vssd1 vccd1 vccd1 _1253_ sky130_fd_sc_hd__buf_4
X_5295_ _0265_ _0267_ vssd1 vssd1 vccd1 vccd1 _0268_ sky130_fd_sc_hd__or2_1
X_8083_ _3236_ _3276_ vssd1 vssd1 vccd1 vccd1 _3277_ sky130_fd_sc_hd__xor2_1
X_7034_ _1782_ _1813_ vssd1 vssd1 vccd1 vccd1 _2125_ sky130_fd_sc_hd__nand2_1
XFILLER_19_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6555__A _0303_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_615 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7089__C _4126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7936_ _3038_ _3078_ _3116_ vssd1 vssd1 vccd1 vccd1 _3117_ sky130_fd_sc_hd__a21o_1
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_26 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7867_ _3038_ _3040_ vssd1 vssd1 vccd1 vccd1 _3041_ sky130_fd_sc_hd__nor2_1
XFILLER_35_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6818_ _1841_ _1885_ vssd1 vssd1 vccd1 vccd1 _1887_ sky130_fd_sc_hd__nand2_1
XFILLER_51_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7798_ _2911_ vssd1 vssd1 vccd1 vccd1 _2965_ sky130_fd_sc_hd__inv_2
X_6749_ _1384_ _1510_ vssd1 vssd1 vccd1 vccd1 _1811_ sky130_fd_sc_hd__nor2_1
XFILLER_51_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8419_ _0635_ _3630_ _3632_ vssd1 vssd1 vccd1 vccd1 _3633_ sky130_fd_sc_hd__and3b_1
XFILLER_105_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7995__S _2721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5809__A _3802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5080_ _4210_ _3840_ vssd1 vssd1 vccd1 vccd1 _4235_ sky130_fd_sc_hd__nor2_1
XFILLER_110_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6375__A _1399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6094__B _0722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5982_ _0976_ _0975_ _0968_ _0974_ vssd1 vssd1 vccd1 vccd1 _0978_ sky130_fd_sc_hd__o211a_1
XFILLER_92_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4933_ _4080_ _4086_ _4087_ vssd1 vssd1 vccd1 vccd1 _4088_ sky130_fd_sc_hd__o21a_1
X_7721_ _2770_ _2878_ _2879_ vssd1 vssd1 vccd1 vccd1 _2880_ sky130_fd_sc_hd__a21o_1
XFILLER_32_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4864_ _4018_ _3927_ vssd1 vssd1 vccd1 vccd1 _4019_ sky130_fd_sc_hd__xor2_1
XFILLER_32_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7652_ _2708_ _2803_ vssd1 vssd1 vccd1 vccd1 _2805_ sky130_fd_sc_hd__nand2_1
XFILLER_119_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4795_ _3941_ _3946_ _3949_ vssd1 vssd1 vccd1 vccd1 _3950_ sky130_fd_sc_hd__o21ba_1
X_6603_ _1648_ _1650_ vssd1 vssd1 vccd1 vccd1 _1651_ sky130_fd_sc_hd__xnor2_1
XFILLER_20_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7583_ _2675_ vssd1 vssd1 vccd1 vccd1 _2729_ sky130_fd_sc_hd__inv_2
XFILLER_32_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6534_ _1573_ _1574_ vssd1 vssd1 vccd1 vccd1 _1575_ sky130_fd_sc_hd__xor2_1
X_6465_ _1498_ _1447_ _0105_ vssd1 vssd1 vccd1 vccd1 _1499_ sky130_fd_sc_hd__or3_1
XFILLER_9_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8204_ _3321_ _3405_ _3354_ vssd1 vssd1 vccd1 vccd1 _3406_ sky130_fd_sc_hd__nor3b_1
X_5416_ _0387_ _0388_ vssd1 vssd1 vccd1 vccd1 _0389_ sky130_fd_sc_hd__and2_1
X_6396_ _1422_ vssd1 vssd1 vccd1 vccd1 _1423_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__5173__B _3986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5347_ _4206_ _4205_ vssd1 vssd1 vccd1 vccd1 _0320_ sky130_fd_sc_hd__and2b_1
X_8135_ _3294_ _3301_ _3226_ vssd1 vssd1 vccd1 vccd1 _3332_ sky130_fd_sc_hd__a21oi_1
XFILLER_102_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5278_ _0235_ _0237_ vssd1 vssd1 vccd1 vccd1 _0251_ sky130_fd_sc_hd__or2_1
X_8066_ _0595_ _3219_ vssd1 vssd1 vccd1 vccd1 _3258_ sky130_fd_sc_hd__or2b_1
X_7017_ _2062_ _2070_ vssd1 vssd1 vccd1 vccd1 _2106_ sky130_fd_sc_hd__xnor2_1
XFILLER_101_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5579__A2 _3804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7919_ _3065_ _3097_ vssd1 vssd1 vccd1 vccd1 _3098_ sky130_fd_sc_hd__and2_1
XANTENNA__6118__B_N _1097_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5200__A1 _3988_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8150__B1 _3346_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4490__A2 posit_add.in1\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4580_ _3734_ vssd1 vssd1 vccd1 vccd1 _3735_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__5742__A2 _0722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4950__B1 _3702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6250_ _1228_ _1259_ vssd1 vssd1 vccd1 vccd1 _1262_ sky130_fd_sc_hd__xor2_1
X_6181_ _1184_ _1186_ vssd1 vssd1 vccd1 vccd1 _1187_ sky130_fd_sc_hd__xor2_1
X_5201_ _4182_ _0140_ vssd1 vssd1 vccd1 vccd1 _0174_ sky130_fd_sc_hd__xor2_1
XFILLER_97_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5132_ _4017_ _3755_ vssd1 vssd1 vccd1 vccd1 _0105_ sky130_fd_sc_hd__or2_2
XFILLER_97_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5258__A1 _4157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5063_ _3802_ _4217_ vssd1 vssd1 vccd1 vccd1 _4218_ sky130_fd_sc_hd__nand2_1
XFILLER_53_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5965_ _0943_ _0944_ _0959_ vssd1 vssd1 vccd1 vccd1 _0960_ sky130_fd_sc_hd__and3_1
XFILLER_80_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5896_ _0885_ _0886_ _0887_ vssd1 vssd1 vccd1 vccd1 _0888_ sky130_fd_sc_hd__nand3_1
X_4916_ _4049_ _4063_ vssd1 vssd1 vccd1 vccd1 _4071_ sky130_fd_sc_hd__xor2_1
X_7704_ _2703_ _2706_ vssd1 vssd1 vccd1 vccd1 _2862_ sky130_fd_sc_hd__nor2_1
XFILLER_40_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4847_ _3999_ _4000_ _4001_ vssd1 vssd1 vccd1 vccd1 _4002_ sky130_fd_sc_hd__and3_1
XFILLER_21_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7635_ _2764_ _2785_ _2731_ vssd1 vssd1 vccd1 vccd1 _2786_ sky130_fd_sc_hd__mux2_1
XFILLER_20_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4778_ _3915_ _3916_ _3932_ vssd1 vssd1 vccd1 vccd1 _3933_ sky130_fd_sc_hd__a21oi_1
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7566_ _2675_ _2704_ _2709_ vssd1 vssd1 vccd1 vccd1 _2710_ sky130_fd_sc_hd__or3b_2
X_6517_ _1402_ _1403_ vssd1 vssd1 vccd1 vccd1 _1556_ sky130_fd_sc_hd__xor2_1
X_7497_ _2903_ _1858_ _2631_ _2632_ _2633_ vssd1 vssd1 vccd1 vccd1 _2634_ sky130_fd_sc_hd__o221a_1
XFILLER_106_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6448_ _1463_ _1479_ vssd1 vssd1 vccd1 vccd1 _1480_ sky130_fd_sc_hd__xnor2_1
X_6379_ _1356_ _1386_ _1402_ _1403_ vssd1 vssd1 vccd1 vccd1 _1404_ sky130_fd_sc_hd__a22o_1
X_8118_ _3293_ _3304_ _3313_ _3195_ vssd1 vssd1 vccd1 vccd1 _3314_ sky130_fd_sc_hd__a31o_1
XFILLER_102_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6727__B _1401_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8049_ _3227_ _3228_ _3238_ vssd1 vssd1 vccd1 vccd1 _3240_ sky130_fd_sc_hd__o21ai_1
XFILLER_29_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7410__A2 _2536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4263__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5078__B _3701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5094__A _3701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4438__A posit_add.in1\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5750_ _0647_ _4044_ _3814_ vssd1 vssd1 vccd1 vccd1 _0732_ sky130_fd_sc_hd__a21o_1
XFILLER_22_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5681_ _2507_ _3864_ _3813_ vssd1 vssd1 vccd1 vccd1 _0656_ sky130_fd_sc_hd__or3_1
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4701_ _3832_ _3855_ _3844_ vssd1 vssd1 vccd1 vccd1 _3856_ sky130_fd_sc_hd__and3_1
XFILLER_15_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7420_ _2548_ _2238_ _2220_ vssd1 vssd1 vccd1 vccd1 _2549_ sky130_fd_sc_hd__mux2_1
X_4632_ _3520_ _3786_ vssd1 vssd1 vccd1 vccd1 _3787_ sky130_fd_sc_hd__and2_1
XANTENNA__7484__A cmd\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4563_ _3717_ vssd1 vssd1 vccd1 vccd1 _3718_ sky130_fd_sc_hd__buf_2
X_7351_ _1428_ _2412_ _2444_ _2470_ _2472_ vssd1 vssd1 vccd1 vccd1 _2473_ sky130_fd_sc_hd__a221oi_4
XFILLER_116_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6302_ _1316_ _1318_ vssd1 vssd1 vccd1 vccd1 _1320_ sky130_fd_sc_hd__and2_1
X_4494_ posit_add.in1\[0\] _1242_ vssd1 vssd1 vccd1 vccd1 _3221_ sky130_fd_sc_hd__nand2_1
X_7282_ _2365_ _2389_ vssd1 vssd1 vccd1 vccd1 _2398_ sky130_fd_sc_hd__xnor2_2
XFILLER_116_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6233_ _1197_ _1201_ vssd1 vssd1 vccd1 vccd1 _1244_ sky130_fd_sc_hd__xnor2_1
XANTENNA__5732__A _3866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6164_ _0795_ _1128_ vssd1 vssd1 vccd1 vccd1 _1169_ sky130_fd_sc_hd__nand2_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6095_ _0634_ vssd1 vssd1 vccd1 vccd1 _1097_ sky130_fd_sc_hd__buf_2
XFILLER_69_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5115_ _0075_ _0087_ vssd1 vssd1 vccd1 vccd1 _0088_ sky130_fd_sc_hd__nand2_1
XFILLER_85_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5046_ _4028_ _4030_ _4200_ vssd1 vssd1 vccd1 vccd1 _4201_ sky130_fd_sc_hd__a21oi_1
XFILLER_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6997_ _2047_ _2082_ vssd1 vssd1 vccd1 vccd1 _2084_ sky130_fd_sc_hd__and2_1
XFILLER_53_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5948_ _0921_ _0922_ _0941_ vssd1 vssd1 vccd1 vccd1 _0942_ sky130_fd_sc_hd__a21o_1
XFILLER_80_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5879_ _0867_ _0869_ vssd1 vssd1 vccd1 vccd1 _0870_ sky130_fd_sc_hd__xor2_1
XFILLER_21_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7618_ _2719_ _2766_ _2748_ vssd1 vssd1 vccd1 vccd1 _2767_ sky130_fd_sc_hd__mux2_1
XFILLER_119_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5626__B cmd\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8002__B cmd\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7549_ _2681_ _2678_ vssd1 vssd1 vccd1 vccd1 _2691_ sky130_fd_sc_hd__or2b_1
XANTENNA__6116__C1 _0702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5999__D _0991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7569__A _2652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7288__B _2354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5817__A _4016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5698__S _3924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6920_ _1951_ _1997_ _1998_ vssd1 vssd1 vccd1 vccd1 _1999_ sky130_fd_sc_hd__a21o_1
XFILLER_35_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6851_ _1779_ _1844_ vssd1 vssd1 vccd1 vccd1 _1923_ sky130_fd_sc_hd__xnor2_1
XANTENNA__7386__A1 _2381_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5802_ _0755_ vssd1 vssd1 vccd1 vccd1 _0787_ sky130_fd_sc_hd__buf_2
XFILLER_90_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6782_ _1408_ _1409_ _4089_ vssd1 vssd1 vccd1 vccd1 _1848_ sky130_fd_sc_hd__and3_1
X_8521_ clknet_3_3__leaf_clk _0007_ vssd1 vssd1 vccd1 vccd1 in_reg\[4\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__4334__C posit_add.in2\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5733_ _3775_ _0634_ vssd1 vssd1 vccd1 vccd1 _0714_ sky130_fd_sc_hd__nand2_1
X_5664_ _0625_ _0637_ vssd1 vssd1 vccd1 vccd1 _0638_ sky130_fd_sc_hd__xnor2_1
X_8452_ _3658_ vssd1 vssd1 vccd1 vccd1 _0045_ sky130_fd_sc_hd__clkbuf_1
XFILLER_30_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7403_ _2151_ _2244_ vssd1 vssd1 vccd1 vccd1 _2531_ sky130_fd_sc_hd__nand2_1
X_4615_ _1748_ _3769_ vssd1 vssd1 vccd1 vccd1 _3770_ sky130_fd_sc_hd__nand2_4
X_8383_ _3182_ _3565_ _3595_ vssd1 vssd1 vccd1 vccd1 _3596_ sky130_fd_sc_hd__a21o_1
X_5595_ _0514_ vssd1 vssd1 vccd1 vccd1 _0568_ sky130_fd_sc_hd__clkinv_2
X_4546_ _3700_ vssd1 vssd1 vccd1 vccd1 _3701_ sky130_fd_sc_hd__clkbuf_4
X_7334_ _1900_ _2417_ _2260_ _2007_ vssd1 vssd1 vccd1 vccd1 _2455_ sky130_fd_sc_hd__a31oi_1
X_4477_ posit_add.in1\[13\] _3024_ vssd1 vssd1 vccd1 vccd1 _3035_ sky130_fd_sc_hd__xnor2_4
XFILLER_1_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7265_ _2377_ _2378_ vssd1 vssd1 vccd1 vccd1 _2379_ sky130_fd_sc_hd__and2_1
X_6216_ _1172_ _1187_ vssd1 vssd1 vccd1 vccd1 _1225_ sky130_fd_sc_hd__xnor2_1
XFILLER_89_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7196_ _1634_ _2301_ vssd1 vssd1 vccd1 vccd1 _2303_ sky130_fd_sc_hd__and2_1
X_6147_ _1107_ _1113_ _1112_ vssd1 vssd1 vccd1 vccd1 _1151_ sky130_fd_sc_hd__a21o_1
XFILLER_85_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6078_ _1056_ _1074_ vssd1 vssd1 vccd1 vccd1 _1079_ sky130_fd_sc_hd__nand2_1
X_5029_ _3816_ _4037_ _3829_ vssd1 vssd1 vccd1 vccd1 _4184_ sky130_fd_sc_hd__o21ai_1
XFILLER_54_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8087__B1_N _0701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4716__A _3776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4435__B posit_add.in1\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6931__A _1414_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8317__B1 _3524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4400_ _1506_ _1451_ vssd1 vssd1 vccd1 vccd1 _2188_ sky130_fd_sc_hd__and2_1
X_5380_ _2727_ _3530_ _0352_ vssd1 vssd1 vccd1 vccd1 _0353_ sky130_fd_sc_hd__o21a_1
X_4331_ posit_add.in2\[14\] _1418_ vssd1 vssd1 vccd1 vccd1 _1429_ sky130_fd_sc_hd__xnor2_4
X_7050_ _2139_ _2141_ vssd1 vssd1 vccd1 vccd1 _2142_ sky130_fd_sc_hd__xnor2_1
X_4262_ _0646_ _0657_ _0679_ vssd1 vssd1 vccd1 vccd1 _0690_ sky130_fd_sc_hd__o21ai_1
X_6001_ _0634_ _0994_ _0996_ _0997_ vssd1 vssd1 vccd1 vccd1 _0998_ sky130_fd_sc_hd__nand4_2
XFILLER_101_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4626__A _3763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7952_ _3103_ _3086_ _3098_ _3025_ _3133_ vssd1 vssd1 vccd1 vccd1 _3135_ sky130_fd_sc_hd__a221o_1
XFILLER_27_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6903_ _1978_ _1980_ vssd1 vssd1 vccd1 vccd1 _1981_ sky130_fd_sc_hd__xor2_1
XANTENNA__4290__A0 in_reg\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7883_ _2937_ _2941_ vssd1 vssd1 vccd1 vccd1 _3059_ sky130_fd_sc_hd__or2_1
XFILLER_35_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6834_ _1300_ _4153_ _1809_ vssd1 vssd1 vccd1 vccd1 _1905_ sky130_fd_sc_hd__and3_1
XFILLER_63_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6765_ _1802_ _1827_ vssd1 vssd1 vccd1 vccd1 _1829_ sky130_fd_sc_hd__nor2_1
XFILLER_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5716_ _0111_ _3864_ _0619_ vssd1 vssd1 vccd1 vccd1 _0695_ sky130_fd_sc_hd__and3_1
X_8504_ posit_add.in2\[11\] in_reg\[11\] _3676_ vssd1 vssd1 vccd1 vccd1 _3692_ sky130_fd_sc_hd__mux2_1
XFILLER_50_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4593__A1 _2969_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6696_ _1742_ _1741_ vssd1 vssd1 vccd1 vccd1 _1753_ sky130_fd_sc_hd__or2b_1
X_8435_ _3646_ vssd1 vssd1 vccd1 vccd1 _0039_ sky130_fd_sc_hd__clkbuf_1
XFILLER_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5647_ _3865_ _0619_ vssd1 vssd1 vccd1 vccd1 _0620_ sky130_fd_sc_hd__and2_1
X_5578_ _3845_ _0548_ vssd1 vssd1 vccd1 vccd1 _0551_ sky130_fd_sc_hd__nor2_1
X_8366_ out_reg\[11\] _3316_ _3197_ out_reg\[12\] vssd1 vssd1 vccd1 vccd1 _3578_ sky130_fd_sc_hd__a22o_1
XFILLER_117_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5904__B _0773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4529_ _3583_ vssd1 vssd1 vccd1 vccd1 _3594_ sky130_fd_sc_hd__clkbuf_4
X_8297_ _3419_ _3450_ _3482_ _3503_ vssd1 vssd1 vccd1 vccd1 _3504_ sky130_fd_sc_hd__a31o_1
X_7317_ _2410_ _2424_ _2435_ vssd1 vssd1 vccd1 vccd1 _2436_ sky130_fd_sc_hd__o21a_1
XFILLER_116_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4300__S _0819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5192__A _3901_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7248_ _0422_ _0417_ vssd1 vssd1 vccd1 vccd1 _2360_ sky130_fd_sc_hd__and2b_1
XFILLER_104_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7611__S _2721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7179_ _2282_ _2283_ vssd1 vssd1 vccd1 vccd1 _2284_ sky130_fd_sc_hd__or2_1
XFILLER_58_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5836__A1 _3815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4446__A posit_add.in1\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4880_ _3807_ _3954_ _4034_ vssd1 vssd1 vccd1 vccd1 _4035_ sky130_fd_sc_hd__a21boi_1
XFILLER_60_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6550_ _1499_ _1591_ vssd1 vssd1 vccd1 vccd1 _1592_ sky130_fd_sc_hd__xnor2_1
XANTENNA__5772__B1 _0754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5501_ _4068_ _4149_ vssd1 vssd1 vccd1 vccd1 _0474_ sky130_fd_sc_hd__xor2_1
XFILLER_9_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7492__A _1913_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6481_ _1511_ _1513_ _1515_ vssd1 vssd1 vccd1 vccd1 _1516_ sky130_fd_sc_hd__and3_1
X_5432_ _3729_ _0403_ _0404_ vssd1 vssd1 vccd1 vccd1 _0405_ sky130_fd_sc_hd__mux2_1
X_8220_ _1330_ _3415_ _3421_ vssd1 vssd1 vccd1 vccd1 _3422_ sky130_fd_sc_hd__a21oi_1
X_8151_ _1220_ _3348_ vssd1 vssd1 vccd1 vccd1 _0024_ sky130_fd_sc_hd__nor2_1
X_5363_ _0090_ _0098_ _0335_ vssd1 vssd1 vccd1 vccd1 _0336_ sky130_fd_sc_hd__a21o_1
XFILLER_114_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7102_ _0147_ _2079_ vssd1 vssd1 vccd1 vccd1 _2200_ sky130_fd_sc_hd__nand2_1
X_4314_ posit_add.in1\[15\] vssd1 vssd1 vccd1 vccd1 _1242_ sky130_fd_sc_hd__clkbuf_4
XFILLER_87_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5294_ _0255_ _0266_ vssd1 vssd1 vccd1 vccd1 _0267_ sky130_fd_sc_hd__nand2_1
XFILLER_59_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8082_ _3135_ _3274_ _3030_ vssd1 vssd1 vccd1 vccd1 _3276_ sky130_fd_sc_hd__mux2_1
X_7033_ _2058_ _2091_ _2097_ vssd1 vssd1 vccd1 vccd1 _2124_ sky130_fd_sc_hd__a21o_1
XFILLER_101_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5740__A _3719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6836__A _3840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6555__B _1400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7935_ _3115_ _3104_ _3044_ vssd1 vssd1 vccd1 vccd1 _3116_ sky130_fd_sc_hd__mux2_1
XFILLER_35_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7866_ _2954_ _3039_ vssd1 vssd1 vccd1 vccd1 _3040_ sky130_fd_sc_hd__or2_1
X_6817_ _1841_ _1885_ vssd1 vssd1 vccd1 vccd1 _1886_ sky130_fd_sc_hd__or2_1
XFILLER_11_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7797_ _2923_ _2963_ _2921_ vssd1 vssd1 vccd1 vccd1 _2964_ sky130_fd_sc_hd__o21a_1
XFILLER_23_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6748_ _0218_ _1300_ _1809_ vssd1 vssd1 vccd1 vccd1 _1810_ sky130_fd_sc_hd__and3_1
XFILLER_51_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6679_ _1702_ _1732_ _1733_ vssd1 vssd1 vccd1 vccd1 _1734_ sky130_fd_sc_hd__a21oi_1
XANTENNA__7606__S _2652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8418_ out_reg\[14\] _0797_ _3631_ out_reg\[15\] vssd1 vssd1 vccd1 vccd1 _3632_ sky130_fd_sc_hd__o22a_1
X_8349_ _3234_ _3326_ vssd1 vssd1 vccd1 vccd1 _3559_ sky130_fd_sc_hd__or2_1
XFILLER_116_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5818__A1 _3719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5809__B _0762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5097__A _4228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7284__A2_N _2354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5981_ _0974_ _0968_ _0975_ _0976_ vssd1 vssd1 vccd1 vccd1 _0977_ sky130_fd_sc_hd__a211oi_1
XANTENNA__6391__A _0303_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4932_ _4081_ _4085_ vssd1 vssd1 vccd1 vccd1 _4087_ sky130_fd_sc_hd__nand2_1
XFILLER_18_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7720_ _2768_ _2769_ vssd1 vssd1 vccd1 vccd1 _2879_ sky130_fd_sc_hd__and2_1
X_7651_ _3726_ _3845_ _2713_ vssd1 vssd1 vccd1 vccd1 _2803_ sky130_fd_sc_hd__mux2_1
XFILLER_33_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4863_ _4017_ _3725_ vssd1 vssd1 vccd1 vccd1 _4018_ sky130_fd_sc_hd__nor2_2
X_6602_ _1585_ _1613_ _1612_ vssd1 vssd1 vccd1 vccd1 _1650_ sky130_fd_sc_hd__a21oi_1
XFILLER_20_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4794_ _3947_ _3948_ vssd1 vssd1 vccd1 vccd1 _3949_ sky130_fd_sc_hd__nor2_1
X_7582_ _2726_ vssd1 vssd1 vccd1 vccd1 _2728_ sky130_fd_sc_hd__inv_2
X_6533_ _1519_ _1520_ vssd1 vssd1 vccd1 vccd1 _1574_ sky130_fd_sc_hd__xnor2_1
XANTENNA__7426__S _2416_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7498__B1 _1858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6464_ _4250_ _1428_ vssd1 vssd1 vccd1 vccd1 _1498_ sky130_fd_sc_hd__nor2_1
XANTENNA__8111__A _0451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5415_ _0376_ _0379_ _0380_ vssd1 vssd1 vccd1 vccd1 _0388_ sky130_fd_sc_hd__o21ai_4
X_8203_ _2598_ _3404_ _2520_ vssd1 vssd1 vccd1 vccd1 _3405_ sky130_fd_sc_hd__mux2_1
X_6395_ _1335_ _1421_ vssd1 vssd1 vccd1 vccd1 _1422_ sky130_fd_sc_hd__xor2_2
XFILLER_114_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5346_ _0317_ _0318_ vssd1 vssd1 vccd1 vccd1 _0319_ sky130_fd_sc_hd__nand2_1
X_8134_ _3329_ _3330_ vssd1 vssd1 vccd1 vccd1 _3331_ sky130_fd_sc_hd__and2_1
XFILLER_0_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5277_ _0247_ _0249_ vssd1 vssd1 vccd1 vccd1 _0250_ sky130_fd_sc_hd__xor2_1
X_8065_ _3214_ _3220_ vssd1 vssd1 vccd1 vccd1 _3257_ sky130_fd_sc_hd__nor2_1
X_7016_ _2090_ _2098_ _2104_ vssd1 vssd1 vccd1 vccd1 _2105_ sky130_fd_sc_hd__o21ai_1
XFILLER_102_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4814__A _3815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7918_ _3096_ vssd1 vssd1 vccd1 vccd1 _3097_ sky130_fd_sc_hd__inv_2
XFILLER_102_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7849_ _3020_ vssd1 vssd1 vccd1 vccd1 _3021_ sky130_fd_sc_hd__clkbuf_4
XFILLER_23_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6476__A _4232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4724__A _3878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4950__B2 _3828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6180_ _1134_ _1185_ vssd1 vssd1 vccd1 vccd1 _1186_ sky130_fd_sc_hd__nand2_1
XFILLER_69_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5200_ _3988_ _0167_ _0171_ _0172_ vssd1 vssd1 vccd1 vccd1 _0173_ sky130_fd_sc_hd__o22a_1
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5131_ _4215_ _0103_ vssd1 vssd1 vccd1 vccd1 _0104_ sky130_fd_sc_hd__nor2_1
XFILLER_111_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5062_ _3855_ vssd1 vssd1 vccd1 vccd1 _4217_ sky130_fd_sc_hd__buf_6
XFILLER_111_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5964_ _0949_ _0955_ _0958_ vssd1 vssd1 vccd1 vccd1 _0959_ sky130_fd_sc_hd__o21a_1
X_7703_ _2858_ _2860_ vssd1 vssd1 vccd1 vccd1 _2861_ sky130_fd_sc_hd__nand2_1
X_5895_ _3892_ _0706_ _3832_ _0722_ vssd1 vssd1 vccd1 vccd1 _0887_ sky130_fd_sc_hd__a22o_1
XFILLER_80_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4915_ _4066_ _4069_ vssd1 vssd1 vccd1 vccd1 _4070_ sky130_fd_sc_hd__nand2_1
XFILLER_33_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4846_ _3763_ _3817_ vssd1 vssd1 vccd1 vccd1 _4001_ sky130_fd_sc_hd__nor2_1
X_7634_ _2774_ _2784_ _2708_ vssd1 vssd1 vccd1 vccd1 _2785_ sky130_fd_sc_hd__mux2_1
X_7565_ _2319_ _2706_ _2708_ vssd1 vssd1 vccd1 vccd1 _2709_ sky130_fd_sc_hd__and3_1
X_4777_ _3929_ _3931_ vssd1 vssd1 vccd1 vccd1 _3932_ sky130_fd_sc_hd__xnor2_1
X_6516_ _1551_ _1417_ _1553_ _1554_ vssd1 vssd1 vccd1 vccd1 _1555_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_107_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7496_ _2936_ _1836_ vssd1 vssd1 vccd1 vccd1 _2633_ sky130_fd_sc_hd__or2_1
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6447_ _1472_ _1478_ vssd1 vssd1 vccd1 vccd1 _1479_ sky130_fd_sc_hd__xor2_1
X_6378_ _1356_ _1386_ vssd1 vssd1 vccd1 vccd1 _1403_ sky130_fd_sc_hd__xor2_1
XFILLER_102_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5329_ _0285_ _0296_ vssd1 vssd1 vccd1 vccd1 _0302_ sky130_fd_sc_hd__xnor2_1
X_8117_ _3311_ _3312_ vssd1 vssd1 vccd1 vccd1 _3313_ sky130_fd_sc_hd__or2_1
XFILLER_87_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4457__B1 _1253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8048_ _3227_ _3228_ _3238_ vssd1 vssd1 vccd1 vccd1 _3239_ sky130_fd_sc_hd__or3_1
XFILLER_75_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7855__A _2993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5094__B _4232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4719__A _3793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6934__A _3615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8316__B1_N _1177_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5680_ _3813_ _0604_ _0619_ vssd1 vssd1 vccd1 vccd1 _0655_ sky130_fd_sc_hd__o21a_1
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4700_ _3772_ _3846_ _3851_ _3852_ vssd1 vssd1 vccd1 vccd1 _3855_ sky130_fd_sc_hd__o31ai_4
XANTENNA__7765__A _1253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5176__A1 _4222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4631_ _3339_ _3349_ _3424_ _2969_ _3360_ vssd1 vssd1 vccd1 vccd1 _3786_ sky130_fd_sc_hd__o2111a_1
XFILLER_8_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7484__B _0092_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5285__A _3800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4562_ _3690_ _3710_ _3711_ _3716_ vssd1 vssd1 vccd1 vccd1 _3717_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_8_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7350_ _2335_ _2471_ vssd1 vssd1 vccd1 vccd1 _2472_ sky130_fd_sc_hd__and2_1
X_6301_ _1315_ _1317_ vssd1 vssd1 vccd1 vccd1 _1318_ sky130_fd_sc_hd__nor2_1
X_4493_ _2969_ posit_add.in1\[1\] vssd1 vssd1 vccd1 vccd1 _3210_ sky130_fd_sc_hd__or2b_1
X_7281_ _2393_ _2395_ vssd1 vssd1 vccd1 vccd1 _2396_ sky130_fd_sc_hd__xnor2_1
XFILLER_116_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6232_ _1239_ _1240_ _1241_ vssd1 vssd1 vccd1 vccd1 _1243_ sky130_fd_sc_hd__a21bo_1
XFILLER_69_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6163_ _1167_ vssd1 vssd1 vccd1 vccd1 _1168_ sky130_fd_sc_hd__buf_2
XFILLER_69_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6094_ _0762_ _0722_ _0994_ vssd1 vssd1 vccd1 vccd1 _1096_ sky130_fd_sc_hd__and3_1
XFILLER_85_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5114_ _4240_ _4243_ _0077_ vssd1 vssd1 vccd1 vccd1 _0087_ sky130_fd_sc_hd__a21o_1
XFILLER_85_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5045_ _4031_ _4032_ vssd1 vssd1 vccd1 vccd1 _4200_ sky130_fd_sc_hd__nor2_1
XFILLER_84_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8050__B1 _0701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4364__A _1275_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6996_ _2047_ _2082_ vssd1 vssd1 vccd1 vccd1 _2083_ sky130_fd_sc_hd__nor2_1
XFILLER_25_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5947_ _0927_ _0939_ _0940_ vssd1 vssd1 vccd1 vccd1 _0941_ sky130_fd_sc_hd__a21bo_1
XFILLER_53_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5878_ _0833_ _0868_ vssd1 vssd1 vccd1 vccd1 _0869_ sky130_fd_sc_hd__and2_1
X_7617_ _2731_ _2745_ _2765_ vssd1 vssd1 vccd1 vccd1 _2766_ sky130_fd_sc_hd__o21ai_1
X_4829_ _3955_ _3983_ vssd1 vssd1 vccd1 vccd1 _3984_ sky130_fd_sc_hd__xnor2_1
XFILLER_107_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4914__A1 _2540_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7548_ _2654_ _2678_ _2674_ _0351_ vssd1 vssd1 vccd1 vccd1 _2690_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__6116__B1 _4017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7479_ _2612_ _2613_ _2494_ vssd1 vssd1 vccd1 vccd1 _2614_ sky130_fd_sc_hd__mux2_1
XFILLER_108_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7614__S _2652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6929__A _0218_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4449__A posit_add.in1\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6850_ _1482_ _1531_ _1915_ _1921_ vssd1 vssd1 vccd1 vccd1 _1922_ sky130_fd_sc_hd__a31oi_2
XFILLER_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5801_ _0760_ _0784_ vssd1 vssd1 vccd1 vccd1 _0785_ sky130_fd_sc_hd__xnor2_1
X_6781_ _0147_ _1413_ vssd1 vssd1 vccd1 vccd1 _1846_ sky130_fd_sc_hd__nand2_1
XFILLER_35_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5732_ _3866_ _0624_ vssd1 vssd1 vccd1 vccd1 _0713_ sky130_fd_sc_hd__nand2_1
X_8520_ clknet_3_4__leaf_clk _0006_ vssd1 vssd1 vccd1 vccd1 in_reg\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_62_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5663_ _0632_ _0636_ vssd1 vssd1 vccd1 vccd1 _0637_ sky130_fd_sc_hd__nand2_1
X_8451_ in_reg\[2\] posit_add.in1\[2\] _3655_ vssd1 vssd1 vccd1 vccd1 _3658_ sky130_fd_sc_hd__mux2_1
X_7402_ _2118_ _2120_ vssd1 vssd1 vccd1 vccd1 _2530_ sky130_fd_sc_hd__nand2_1
X_4614_ _3736_ _3768_ vssd1 vssd1 vccd1 vccd1 _3769_ sky130_fd_sc_hd__nor2_1
X_8382_ _3560_ _3593_ vssd1 vssd1 vccd1 vccd1 _3595_ sky130_fd_sc_hd__xnor2_1
X_5594_ _0507_ _0487_ _0515_ vssd1 vssd1 vccd1 vccd1 _0567_ sky130_fd_sc_hd__mux2_1
X_4545_ _3699_ vssd1 vssd1 vccd1 vccd1 _3700_ sky130_fd_sc_hd__clkbuf_4
X_7333_ _2409_ vssd1 vssd1 vccd1 vccd1 _2454_ sky130_fd_sc_hd__buf_2
XFILLER_116_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4476_ posit_add.in1\[12\] _3013_ _1253_ vssd1 vssd1 vccd1 vccd1 _3024_ sky130_fd_sc_hd__o21a_1
X_7264_ _2350_ _2376_ _2348_ vssd1 vssd1 vccd1 vccd1 _2378_ sky130_fd_sc_hd__o21ai_2
X_6215_ _1222_ _1223_ vssd1 vssd1 vccd1 vccd1 _1224_ sky130_fd_sc_hd__or2b_1
X_7195_ _1634_ _2301_ _2277_ vssd1 vssd1 vccd1 vccd1 _2302_ sky130_fd_sc_hd__o21bai_2
X_6146_ _1148_ _1149_ vssd1 vssd1 vccd1 vccd1 _1150_ sky130_fd_sc_hd__and2_1
XFILLER_85_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6077_ _1054_ _1076_ _1077_ _0971_ vssd1 vssd1 vccd1 vccd1 _1078_ sky130_fd_sc_hd__a211o_1
XFILLER_85_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5028_ _3828_ _3750_ _4182_ vssd1 vssd1 vccd1 vccd1 _4183_ sky130_fd_sc_hd__or3_1
XFILLER_72_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5918__A _3763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6979_ _1401_ _1537_ _2063_ vssd1 vssd1 vccd1 vccd1 _2064_ sky130_fd_sc_hd__or3_1
XFILLER_41_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6749__A _1384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4716__B _3838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4435__C posit_add.in1\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6931__B _1531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4330_ _1341_ _1374_ _1396_ _1407_ posit_add.in2\[15\] vssd1 vssd1 vccd1 vccd1 _1418_
+ sky130_fd_sc_hd__o41a_2
XFILLER_113_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4261_ counter\[4\] mode _0668_ counter\[3\] vssd1 vssd1 vccd1 vccd1 _0679_ sky130_fd_sc_hd__nor4b_2
XFILLER_113_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6000_ _0892_ _0702_ _0992_ _4016_ vssd1 vssd1 vccd1 vccd1 _0997_ sky130_fd_sc_hd__a211oi_2
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7951_ _3020_ _3132_ vssd1 vssd1 vccd1 vccd1 _3133_ sky130_fd_sc_hd__and2_1
X_6902_ _1911_ _1916_ vssd1 vssd1 vccd1 vccd1 _1980_ sky130_fd_sc_hd__xnor2_1
X_7882_ _3042_ _3056_ _3049_ _3048_ vssd1 vssd1 vccd1 vccd1 _3058_ sky130_fd_sc_hd__a22o_1
XANTENNA__8005__B1 _3192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6833_ _1866_ _1867_ vssd1 vssd1 vccd1 vccd1 _1904_ sky130_fd_sc_hd__xnor2_1
XANTENNA__4290__A1 in_reg\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6841__B _3703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6764_ _1802_ _1827_ vssd1 vssd1 vccd1 vccd1 _1828_ sky130_fd_sc_hd__xor2_1
XFILLER_11_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5715_ _0630_ _0622_ vssd1 vssd1 vccd1 vccd1 _0694_ sky130_fd_sc_hd__and2b_1
X_8503_ _3691_ vssd1 vssd1 vccd1 vccd1 _0069_ sky130_fd_sc_hd__clkbuf_1
X_6695_ _1750_ _1751_ vssd1 vssd1 vccd1 vccd1 _1752_ sky130_fd_sc_hd__nand2_1
X_5646_ _3811_ _3812_ _3775_ _2507_ vssd1 vssd1 vccd1 vccd1 _0619_ sky130_fd_sc_hd__a22o_2
X_8434_ _3644_ _3645_ _3641_ vssd1 vssd1 vccd1 vccd1 _3646_ sky130_fd_sc_hd__and3b_1
XFILLER_31_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5577_ _4119_ _4121_ _4123_ _4118_ vssd1 vssd1 vccd1 vccd1 _0550_ sky130_fd_sc_hd__o211a_1
XANTENNA__8479__A_N net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8365_ _3558_ _3576_ _3195_ vssd1 vssd1 vccd1 vccd1 _3577_ sky130_fd_sc_hd__a21oi_2
XFILLER_117_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4528_ _3134_ _2617_ _2804_ vssd1 vssd1 vccd1 vccd1 _3583_ sky130_fd_sc_hd__and3b_1
X_8296_ _3416_ _3500_ vssd1 vssd1 vccd1 vccd1 _3503_ sky130_fd_sc_hd__nor2_1
X_7316_ _2425_ _2426_ _2427_ _2434_ vssd1 vssd1 vccd1 vccd1 _2435_ sky130_fd_sc_hd__a31o_1
XFILLER_104_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5192__B _3838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4459_ _2661_ _2826_ vssd1 vssd1 vccd1 vccd1 _2837_ sky130_fd_sc_hd__xor2_1
X_7247_ _2354_ _2358_ vssd1 vssd1 vccd1 vccd1 _2359_ sky130_fd_sc_hd__and2_1
X_7178_ _2272_ _2281_ vssd1 vssd1 vccd1 vccd1 _2283_ sky130_fd_sc_hd__nor2_1
X_6129_ _1128_ _1131_ vssd1 vssd1 vccd1 vccd1 _1132_ sky130_fd_sc_hd__xor2_1
XANTENNA__5412__S _3729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5781__A1 _3866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6479__A _0303_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5500_ _0472_ _4147_ vssd1 vssd1 vccd1 vccd1 _0473_ sky130_fd_sc_hd__xnor2_1
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6480_ _1514_ _1485_ vssd1 vssd1 vccd1 vccd1 _1515_ sky130_fd_sc_hd__xnor2_1
XFILLER_9_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6389__A _4217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5431_ _3690_ _3830_ _3635_ _0347_ vssd1 vssd1 vccd1 vccd1 _0404_ sky130_fd_sc_hd__a31o_1
XFILLER_99_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8150_ out_reg\[4\] _1231_ _3346_ _3347_ vssd1 vssd1 vccd1 vccd1 _3348_ sky130_fd_sc_hd__o2bb2a_1
X_5362_ _0093_ _0096_ _0095_ vssd1 vssd1 vccd1 vccd1 _0335_ sky130_fd_sc_hd__or3_1
XFILLER_99_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7101_ _2174_ _2183_ _2196_ vssd1 vssd1 vccd1 vccd1 _2198_ sky130_fd_sc_hd__and3_1
X_4313_ _0786_ _0701_ vssd1 vssd1 vccd1 vccd1 _1231_ sky130_fd_sc_hd__nor2b_2
X_8081_ _3273_ vssd1 vssd1 vccd1 vccd1 _3274_ sky130_fd_sc_hd__clkinv_2
X_7032_ _1711_ _1355_ _1950_ vssd1 vssd1 vccd1 vccd1 _2123_ sky130_fd_sc_hd__and3_1
X_5293_ _0254_ _4187_ _0253_ vssd1 vssd1 vccd1 vccd1 _0266_ sky130_fd_sc_hd__nand3_1
XFILLER_114_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5740__B _3815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7013__A _1401_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7934_ _2901_ _2899_ _3034_ vssd1 vssd1 vccd1 vccd1 _3115_ sky130_fd_sc_hd__mux2_1
X_7865_ _2928_ _2948_ _2971_ vssd1 vssd1 vccd1 vccd1 _3039_ sky130_fd_sc_hd__mux2_1
XFILLER_42_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6816_ _1861_ _1883_ _1884_ vssd1 vssd1 vccd1 vccd1 _1885_ sky130_fd_sc_hd__a21boi_1
XFILLER_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7796_ _2928_ _2932_ vssd1 vssd1 vccd1 vccd1 _2963_ sky130_fd_sc_hd__nor2_1
XFILLER_23_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6747_ _1298_ _1299_ _1278_ vssd1 vssd1 vccd1 vccd1 _1809_ sky130_fd_sc_hd__o21ai_2
XFILLER_50_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6678_ _1691_ _1701_ vssd1 vssd1 vccd1 vccd1 _1733_ sky130_fd_sc_hd__nor2_1
XFILLER_109_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8417_ _1231_ vssd1 vssd1 vccd1 vccd1 _3631_ sky130_fd_sc_hd__inv_2
X_5629_ _0538_ _0594_ _0601_ vssd1 vssd1 vccd1 vccd1 _0602_ sky130_fd_sc_hd__and3b_1
X_8348_ _1330_ _3547_ _3556_ _3557_ _0600_ vssd1 vssd1 vccd1 vccd1 _3558_ sky130_fd_sc_hd__a311o_1
XFILLER_3_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5931__A _3735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5818__A2 _0702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8279_ _3419_ _3450_ _3482_ _3484_ vssd1 vssd1 vccd1 vccd1 _3485_ sky130_fd_sc_hd__a31oi_4
XFILLER_116_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6465__C _0105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8453__S _3655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5097__B _3925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5754__A1 _0687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5841__A _3770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5980_ _0881_ _0863_ _0880_ vssd1 vssd1 vccd1 vccd1 _0976_ sky130_fd_sc_hd__and3_1
XFILLER_92_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4931_ _4081_ _4085_ vssd1 vssd1 vccd1 vccd1 _4086_ sky130_fd_sc_hd__xnor2_1
XFILLER_45_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4862_ _4016_ vssd1 vssd1 vccd1 vccd1 _4017_ sky130_fd_sc_hd__buf_4
X_7650_ _3845_ _4126_ _2713_ vssd1 vssd1 vccd1 vccd1 _2802_ sky130_fd_sc_hd__mux2_1
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6601_ _1622_ _1647_ vssd1 vssd1 vccd1 vccd1 _1648_ sky130_fd_sc_hd__xnor2_1
XFILLER_33_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4793_ _3941_ _3946_ vssd1 vssd1 vccd1 vccd1 _3948_ sky130_fd_sc_hd__xnor2_1
X_7581_ _2723_ _2725_ vssd1 vssd1 vccd1 vccd1 _2726_ sky130_fd_sc_hd__nand2_1
XFILLER_119_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6532_ _1566_ _1567_ _1568_ _1570_ _1571_ vssd1 vssd1 vccd1 vccd1 _1573_ sky130_fd_sc_hd__a32oi_4
X_6463_ _1446_ _1428_ vssd1 vssd1 vccd1 vccd1 _1497_ sky130_fd_sc_hd__or2_1
XANTENNA__7498__B2 _2903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8202_ _2514_ _3250_ _3286_ vssd1 vssd1 vccd1 vccd1 _3404_ sky130_fd_sc_hd__a21bo_1
X_5414_ _0385_ vssd1 vssd1 vccd1 vccd1 _0387_ sky130_fd_sc_hd__inv_2
X_6394_ _1331_ _1333_ vssd1 vssd1 vccd1 vccd1 _1421_ sky130_fd_sc_hd__nand2_1
X_8133_ _3297_ _3300_ _3327_ vssd1 vssd1 vccd1 vccd1 _3330_ sky130_fd_sc_hd__a21o_1
XFILLER_114_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5345_ _0316_ _0314_ vssd1 vssd1 vccd1 vccd1 _0318_ sky130_fd_sc_hd__or2b_1
XFILLER_101_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5276_ _0205_ _0248_ vssd1 vssd1 vccd1 vccd1 _0249_ sky130_fd_sc_hd__and2_1
X_8064_ _3248_ _3254_ _3255_ vssd1 vssd1 vccd1 vccd1 _3256_ sky130_fd_sc_hd__a21oi_2
X_7015_ _2099_ _2103_ vssd1 vssd1 vccd1 vccd1 _2104_ sky130_fd_sc_hd__nand2_1
XFILLER_75_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4814__B _3702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7917_ _2998_ _3082_ _3095_ vssd1 vssd1 vccd1 vccd1 _3096_ sky130_fd_sc_hd__o21a_1
XFILLER_102_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4306__S _0819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7848_ _3014_ _3019_ vssd1 vssd1 vccd1 vccd1 _3020_ sky130_fd_sc_hd__xnor2_2
XFILLER_11_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7779_ _2938_ _2943_ vssd1 vssd1 vccd1 vccd1 _2944_ sky130_fd_sc_hd__and2_1
XFILLER_7_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6476__B _1510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4724__B _3855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5727__A1 _3866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4740__A _3893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4950__A2 _3795_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5130_ _3802_ _3838_ _4214_ vssd1 vssd1 vccd1 vccd1 _0103_ sky130_fd_sc_hd__a21oi_1
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5061_ _4211_ _4212_ _4215_ vssd1 vssd1 vccd1 vccd1 _4216_ sky130_fd_sc_hd__o21ba_1
XFILLER_111_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5963_ _0956_ _0957_ vssd1 vssd1 vccd1 vccd1 _0958_ sky130_fd_sc_hd__and2_1
XFILLER_65_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4634__B _3776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4914_ _2540_ _3817_ _4065_ vssd1 vssd1 vccd1 vccd1 _4069_ sky130_fd_sc_hd__o21ai_1
X_7702_ _2853_ _2857_ _2742_ _2778_ vssd1 vssd1 vccd1 vccd1 _2860_ sky130_fd_sc_hd__o2bb2a_1
X_5894_ _3792_ _0676_ vssd1 vssd1 vccd1 vccd1 _0886_ sky130_fd_sc_hd__nor2_1
XFILLER_80_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4845_ _3827_ _3771_ _3871_ vssd1 vssd1 vccd1 vccd1 _4000_ sky130_fd_sc_hd__o21ai_1
X_7633_ _3868_ _3893_ _2713_ vssd1 vssd1 vccd1 vccd1 _2784_ sky130_fd_sc_hd__mux2_1
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4776_ _3719_ _3930_ vssd1 vssd1 vccd1 vccd1 _3931_ sky130_fd_sc_hd__nor2_1
XANTENNA__4650__A _3802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7564_ _2707_ vssd1 vssd1 vccd1 vccd1 _2708_ sky130_fd_sc_hd__buf_2
XFILLER_119_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6515_ _1428_ _1423_ vssd1 vssd1 vccd1 vccd1 _1554_ sky130_fd_sc_hd__nor2_2
XANTENNA__8479__D net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7495_ _2936_ _1836_ _1803_ _3189_ vssd1 vssd1 vccd1 vccd1 _2632_ sky130_fd_sc_hd__a22o_1
X_6446_ _1466_ _1427_ _1474_ _1477_ vssd1 vssd1 vccd1 vccd1 _1478_ sky130_fd_sc_hd__a22oi_2
X_6377_ _1400_ _1401_ vssd1 vssd1 vccd1 vccd1 _1402_ sky130_fd_sc_hd__nor2_1
XFILLER_88_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5328_ _0299_ _0300_ vssd1 vssd1 vccd1 vccd1 _0301_ sky130_fd_sc_hd__nand2_1
XFILLER_0_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8116_ _0601_ _3305_ _3310_ _0600_ vssd1 vssd1 vccd1 vccd1 _3312_ sky130_fd_sc_hd__a31o_1
XFILLER_114_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8047_ _3236_ _3237_ vssd1 vssd1 vccd1 vccd1 _3238_ sky130_fd_sc_hd__nand2_1
XFILLER_102_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5259_ _0230_ _0231_ vssd1 vssd1 vccd1 vccd1 _0232_ sky130_fd_sc_hd__xor2_1
XFILLER_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8426__C_N _0701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5375__B _2452_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4719__B _3750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7398__B1 _2524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6950__A _1401_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_718 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7765__B _1275_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5176__A2 _0147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4630_ _3232_ _3307_ _3784_ _3477_ vssd1 vssd1 vccd1 vccd1 _3785_ sky130_fd_sc_hd__a211o_1
XANTENNA__8444__D_N net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7570__A0 _0218_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5285__B _3615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6300_ _1145_ _1148_ _1314_ vssd1 vssd1 vccd1 vccd1 _1317_ sky130_fd_sc_hd__and3_1
X_4561_ _3713_ _3715_ vssd1 vssd1 vccd1 vccd1 _3716_ sky130_fd_sc_hd__and2_1
XFILLER_116_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4492_ _2606_ _3189_ vssd1 vssd1 vccd1 vccd1 _3199_ sky130_fd_sc_hd__xor2_1
XFILLER_7_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7280_ _2369_ _2394_ vssd1 vssd1 vccd1 vccd1 _2395_ sky130_fd_sc_hd__xnor2_4
XFILLER_116_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6231_ _0802_ _1094_ _0787_ _1101_ vssd1 vssd1 vccd1 vccd1 _1241_ sky130_fd_sc_hd__or4b_1
XANTENNA__6397__A _1420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6162_ _1165_ _1166_ vssd1 vssd1 vccd1 vccd1 _1167_ sky130_fd_sc_hd__or2_1
XFILLER_103_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5113_ _0081_ _0085_ vssd1 vssd1 vccd1 vccd1 _0086_ sky130_fd_sc_hd__xnor2_1
XFILLER_111_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6093_ _1094_ vssd1 vssd1 vccd1 vccd1 _1095_ sky130_fd_sc_hd__buf_2
XFILLER_97_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5044_ _4154_ _4198_ vssd1 vssd1 vccd1 vccd1 _4199_ sky130_fd_sc_hd__xnor2_1
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4645__A _3719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6995_ _2075_ _2076_ _2081_ vssd1 vssd1 vccd1 vccd1 _2082_ sky130_fd_sc_hd__a21oi_1
XFILLER_80_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5946_ _0928_ _0938_ _0929_ vssd1 vssd1 vccd1 vccd1 _0940_ sky130_fd_sc_hd__nand3_1
XFILLER_40_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5877_ _3776_ _0624_ _0831_ _0832_ vssd1 vssd1 vccd1 vccd1 _0868_ sky130_fd_sc_hd__a22o_1
XFILLER_43_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4828_ _3963_ _3981_ _3982_ vssd1 vssd1 vccd1 vccd1 _3983_ sky130_fd_sc_hd__o21a_1
XFILLER_21_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7616_ _2712_ _2764_ vssd1 vssd1 vccd1 vccd1 _2765_ sky130_fd_sc_hd__or2_1
X_4759_ _3890_ _3913_ vssd1 vssd1 vccd1 vccd1 _3914_ sky130_fd_sc_hd__xor2_2
XANTENNA__4914__A2 _3817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7547_ _2682_ _2684_ vssd1 vssd1 vccd1 vccd1 _2689_ sky130_fd_sc_hd__xnor2_1
X_7478_ _2488_ _2392_ _2410_ vssd1 vssd1 vccd1 vccd1 _2613_ sky130_fd_sc_hd__mux2_1
X_6429_ _1435_ _1458_ vssd1 vssd1 vccd1 vccd1 _1459_ sky130_fd_sc_hd__xnor2_1
XFILLER_108_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4258__C in_reg\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8461__S _3655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4602__A1 _1682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7866__A _2954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6107__B2 _1097_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7304__B1 _2412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6929__B _1711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_692 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5800_ _0778_ _0783_ vssd1 vssd1 vccd1 vccd1 _0784_ sky130_fd_sc_hd__xnor2_1
XFILLER_90_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6780_ _1779_ _1844_ vssd1 vssd1 vccd1 vccd1 _1845_ sky130_fd_sc_hd__or2_1
XFILLER_50_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5731_ _0625_ _0637_ _0632_ vssd1 vssd1 vccd1 vccd1 _0711_ sky130_fd_sc_hd__o21ai_1
XFILLER_50_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5662_ _0633_ _3892_ _0634_ _3775_ vssd1 vssd1 vccd1 vccd1 _0636_ sky130_fd_sc_hd__a22o_1
X_8450_ _3657_ vssd1 vssd1 vccd1 vccd1 _0044_ sky130_fd_sc_hd__clkbuf_1
X_4613_ _3766_ _3767_ vssd1 vssd1 vccd1 vccd1 _3768_ sky130_fd_sc_hd__and2_1
X_8381_ _3437_ _3370_ _3438_ vssd1 vssd1 vccd1 vccd1 _3593_ sky130_fd_sc_hd__a21o_1
X_7401_ _2522_ _2523_ _2527_ vssd1 vssd1 vccd1 vccd1 _2528_ sky130_fd_sc_hd__a21o_1
X_5593_ _0519_ _0561_ _0563_ _0565_ vssd1 vssd1 vccd1 vccd1 _0566_ sky130_fd_sc_hd__or4_1
XFILLER_116_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4544_ _3625_ _3684_ _3698_ vssd1 vssd1 vccd1 vccd1 _3699_ sky130_fd_sc_hd__o21ai_4
X_7332_ _2436_ _2447_ _2451_ vssd1 vssd1 vccd1 vccd1 _2453_ sky130_fd_sc_hd__mux2_1
X_7263_ _2348_ _2350_ _2376_ vssd1 vssd1 vccd1 vccd1 _2377_ sky130_fd_sc_hd__or3_1
X_6214_ _1213_ _1214_ _1215_ _1164_ vssd1 vssd1 vccd1 vccd1 _1223_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_104_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4475_ posit_add.in1\[11\] posit_add.in1\[10\] _2573_ vssd1 vssd1 vccd1 vccd1 _3013_
+ sky130_fd_sc_hd__or3_2
X_7194_ _2274_ _2273_ _2300_ vssd1 vssd1 vccd1 vccd1 _2301_ sky130_fd_sc_hd__o21ai_1
X_6145_ _1144_ _1147_ vssd1 vssd1 vccd1 vccd1 _1149_ sky130_fd_sc_hd__or2_1
XFILLER_100_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6076_ _0977_ _0978_ vssd1 vssd1 vccd1 vccd1 _1077_ sky130_fd_sc_hd__nor2_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5027_ _3827_ _3816_ vssd1 vssd1 vccd1 vccd1 _4182_ sky130_fd_sc_hd__or2_1
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5388__A2 _3830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6978_ _1454_ _1718_ vssd1 vssd1 vccd1 vccd1 _2063_ sky130_fd_sc_hd__or2_1
XFILLER_80_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5929_ _0919_ _0920_ _0891_ vssd1 vssd1 vccd1 vccd1 _0922_ sky130_fd_sc_hd__a21o_1
XFILLER_110_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8579_ clknet_3_7__leaf_clk _0065_ vssd1 vssd1 vccd1 vccd1 posit_add.in2\[6\] sky130_fd_sc_hd__dfxtp_2
XFILLER_119_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6749__B _1510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_559 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5844__A _3776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4260_ counter\[2\] counter\[1\] counter\[0\] vssd1 vssd1 vccd1 vccd1 _0668_ sky130_fd_sc_hd__or3_1
XFILLER_79_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7950_ _3125_ _3131_ _3006_ vssd1 vssd1 vccd1 vccd1 _3132_ sky130_fd_sc_hd__mux2_1
XFILLER_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6901_ _1975_ _1977_ _1973_ vssd1 vssd1 vccd1 vccd1 _1978_ sky130_fd_sc_hd__a21oi_1
XFILLER_82_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7881_ _3055_ vssd1 vssd1 vccd1 vccd1 _3056_ sky130_fd_sc_hd__inv_2
XFILLER_35_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6832_ _1861_ _1883_ vssd1 vssd1 vccd1 vccd1 _1903_ sky130_fd_sc_hd__xnor2_1
XFILLER_63_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4923__A _3793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4578__B1 _3690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6763_ _1822_ _1824_ _1826_ vssd1 vssd1 vccd1 vccd1 _1827_ sky130_fd_sc_hd__a21oi_1
XFILLER_62_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5714_ _4222_ _0684_ _0692_ vssd1 vssd1 vccd1 vccd1 _0693_ sky130_fd_sc_hd__o21a_1
X_8502_ posit_add.in2\[10\] in_reg\[10\] _3676_ vssd1 vssd1 vccd1 vccd1 _3691_ sky130_fd_sc_hd__mux2_1
X_6694_ _1734_ _1745_ vssd1 vssd1 vccd1 vccd1 _1751_ sky130_fd_sc_hd__xor2_1
XFILLER_50_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7516__B1 _3830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5645_ _0612_ _0613_ _0615_ _0617_ _3801_ vssd1 vssd1 vccd1 vccd1 _0618_ sky130_fd_sc_hd__a2111o_1
X_8433_ counter\[0\] _3242_ counter\[1\] vssd1 vssd1 vccd1 vccd1 _3645_ sky130_fd_sc_hd__a21o_1
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5576_ _2540_ _0548_ _4130_ vssd1 vssd1 vccd1 vccd1 _0549_ sky130_fd_sc_hd__o21ai_1
X_8364_ _3565_ _3566_ _2621_ _3575_ vssd1 vssd1 vccd1 vccd1 _3576_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_117_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4527_ _3520_ _3541_ _3562_ vssd1 vssd1 vccd1 vccd1 _3573_ sky130_fd_sc_hd__and3_1
X_7315_ _1456_ _2412_ _2433_ vssd1 vssd1 vccd1 vccd1 _2434_ sky130_fd_sc_hd__a21oi_1
XFILLER_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8295_ _3419_ _3450_ _3482_ _3501_ vssd1 vssd1 vccd1 vccd1 _3502_ sky130_fd_sc_hd__and4_1
XFILLER_104_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4458_ posit_add.in1\[6\] _2815_ vssd1 vssd1 vccd1 vccd1 _2826_ sky130_fd_sc_hd__xor2_4
XFILLER_49_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7246_ _2356_ _2357_ vssd1 vssd1 vccd1 vccd1 _2358_ sky130_fd_sc_hd__nor2_2
XFILLER_77_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6585__A _1383_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7177_ _2272_ _2281_ vssd1 vssd1 vccd1 vccd1 _2282_ sky130_fd_sc_hd__and2_1
X_6128_ _1129_ _1130_ vssd1 vssd1 vccd1 vccd1 _1131_ sky130_fd_sc_hd__xnor2_1
XFILLER_86_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4389_ _1814_ _2034_ _2045_ _2056_ vssd1 vssd1 vccd1 vccd1 _2067_ sky130_fd_sc_hd__o22a_1
XFILLER_58_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6059_ _0956_ _0957_ _0955_ vssd1 vssd1 vccd1 vccd1 _1059_ sky130_fd_sc_hd__a21oi_1
XFILLER_100_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4309__S _1177_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_662 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4833__A _3853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5766__C1 _3924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5781__A2 _0762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6479__B _1423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5049__A1 _4045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5757__C1 _3866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7773__B _2937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5430_ _0347_ _0402_ _1748_ vssd1 vssd1 vccd1 vccd1 _0403_ sky130_fd_sc_hd__a21o_1
XFILLER_9_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6389__B _1414_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5361_ _0089_ _0132_ _0331_ _0333_ vssd1 vssd1 vccd1 vccd1 _0334_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_114_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7100_ _2174_ _2183_ _2196_ vssd1 vssd1 vccd1 vccd1 _2197_ sky130_fd_sc_hd__nand3_1
X_5292_ _0263_ _0264_ vssd1 vssd1 vccd1 vccd1 _0265_ sky130_fd_sc_hd__nand2_1
X_4312_ _0635_ vssd1 vssd1 vccd1 vccd1 _1220_ sky130_fd_sc_hd__buf_2
X_8080_ _3027_ _3272_ _3025_ vssd1 vssd1 vccd1 vccd1 _3273_ sky130_fd_sc_hd__mux2_1
XFILLER_99_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7031_ _2113_ _2114_ vssd1 vssd1 vccd1 vccd1 _2121_ sky130_fd_sc_hd__xor2_1
XFILLER_113_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4918__A _3739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5740__C _0702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7013__B _1782_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7933_ _3106_ _3113_ _2842_ vssd1 vssd1 vccd1 vccd1 _3114_ sky130_fd_sc_hd__mux2_1
XFILLER_27_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7864_ _2941_ vssd1 vssd1 vccd1 vccd1 _3038_ sky130_fd_sc_hd__buf_2
X_6815_ _1862_ _1882_ vssd1 vssd1 vccd1 vccd1 _1884_ sky130_fd_sc_hd__or2b_1
XANTENNA__5468__B _0440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7795_ _0388_ _2721_ _2667_ vssd1 vssd1 vccd1 vccd1 _2962_ sky130_fd_sc_hd__a21o_1
X_6746_ _1665_ _1511_ _1807_ vssd1 vssd1 vccd1 vccd1 _1808_ sky130_fd_sc_hd__a21o_1
XFILLER_51_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7683__B _2838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6677_ _1721_ _1731_ vssd1 vssd1 vccd1 vccd1 _1732_ sky130_fd_sc_hd__xnor2_1
X_5628_ _1319_ vssd1 vssd1 vccd1 vccd1 _0601_ sky130_fd_sc_hd__buf_2
X_8416_ _3624_ _3626_ _3629_ _1177_ vssd1 vssd1 vccd1 vccd1 _3630_ sky130_fd_sc_hd__a31o_1
XFILLER_117_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8347_ _1330_ _3547_ _3556_ vssd1 vssd1 vccd1 vccd1 _3557_ sky130_fd_sc_hd__a21oi_1
X_5559_ _0341_ _0489_ _0470_ vssd1 vssd1 vccd1 vccd1 _0532_ sky130_fd_sc_hd__mux2_1
XANTENNA__8465__A1 posit_add.in1\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8278_ _3419_ _3450_ _3483_ vssd1 vssd1 vccd1 vccd1 _3484_ sky130_fd_sc_hd__a21oi_1
XFILLER_116_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7229_ _3722_ _0373_ vssd1 vssd1 vccd1 vccd1 _2339_ sky130_fd_sc_hd__nand2_1
XFILLER_86_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5659__A _3792_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8035__A _1275_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5203__A1 _3800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7114__A _1711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4738__A _3892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4930_ _4083_ _4084_ vssd1 vssd1 vccd1 vccd1 _4085_ sky130_fd_sc_hd__and2b_1
XANTENNA__4473__A _2969_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4861_ posit_add.in2\[14\] _4015_ vssd1 vssd1 vccd1 vccd1 _4016_ sky130_fd_sc_hd__nor2_8
X_6600_ _1644_ _1646_ vssd1 vssd1 vccd1 vccd1 _1647_ sky130_fd_sc_hd__xor2_1
XFILLER_20_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4792_ _3780_ _3797_ vssd1 vssd1 vccd1 vccd1 _3947_ sky130_fd_sc_hd__xor2_1
XFILLER_60_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7580_ _2724_ vssd1 vssd1 vccd1 vccd1 _2725_ sky130_fd_sc_hd__inv_2
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6531_ _1549_ _1557_ vssd1 vssd1 vccd1 vccd1 _1571_ sky130_fd_sc_hd__xor2_2
X_6462_ _1481_ _1489_ _1494_ vssd1 vssd1 vccd1 vccd1 _1496_ sky130_fd_sc_hd__a21boi_1
XFILLER_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6393_ _3840_ vssd1 vssd1 vccd1 vccd1 _1420_ sky130_fd_sc_hd__buf_2
X_5413_ _0376_ _0379_ _0380_ _0385_ vssd1 vssd1 vccd1 vccd1 _0386_ sky130_fd_sc_hd__o211a_1
X_8201_ _3289_ _3401_ _3284_ vssd1 vssd1 vccd1 vccd1 _3402_ sky130_fd_sc_hd__or3b_1
X_5344_ _0314_ _0316_ vssd1 vssd1 vccd1 vccd1 _0317_ sky130_fd_sc_hd__or2b_1
XANTENNA__8447__A1 _2969_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8132_ _3297_ _3300_ _3327_ vssd1 vssd1 vccd1 vccd1 _3329_ sky130_fd_sc_hd__nand3_1
XFILLER_87_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5275_ _0204_ _0197_ _0202_ vssd1 vssd1 vccd1 vccd1 _0248_ sky130_fd_sc_hd__or3_1
X_8063_ _3248_ _3254_ _3212_ vssd1 vssd1 vccd1 vccd1 _3255_ sky130_fd_sc_hd__o21ai_1
X_7014_ _2032_ _2087_ _2101_ _2102_ vssd1 vssd1 vccd1 vccd1 _2103_ sky130_fd_sc_hd__o211a_1
XFILLER_87_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7916_ _2998_ _3094_ vssd1 vssd1 vccd1 vccd1 _3095_ sky130_fd_sc_hd__nand2_1
XFILLER_24_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7847_ _3016_ _3018_ vssd1 vssd1 vccd1 vccd1 _3019_ sky130_fd_sc_hd__xnor2_1
XFILLER_23_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7778_ _2654_ _2937_ vssd1 vssd1 vccd1 vccd1 _2943_ sky130_fd_sc_hd__nand2_1
X_6729_ _1668_ _1788_ vssd1 vssd1 vccd1 vccd1 _1789_ sky130_fd_sc_hd__xnor2_1
XFILLER_11_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6103__A _0795_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5389__A _1748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5727__A2 _0706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5060_ _3802_ _3838_ _4214_ vssd1 vssd1 vccd1 vccd1 _4215_ sky130_fd_sc_hd__and3_1
XFILLER_111_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5962_ _0937_ _0934_ _0936_ vssd1 vssd1 vccd1 vccd1 _0957_ sky130_fd_sc_hd__a21o_1
XFILLER_92_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4913_ _4047_ _4067_ vssd1 vssd1 vccd1 vccd1 _4068_ sky130_fd_sc_hd__xnor2_1
X_7701_ _2808_ _2857_ _2742_ _2767_ vssd1 vssd1 vccd1 vccd1 _2858_ sky130_fd_sc_hd__o2bb2a_1
X_5893_ _0693_ _3738_ _0855_ vssd1 vssd1 vccd1 vccd1 _0885_ sky130_fd_sc_hd__or3_1
XANTENNA__8365__B1 _3195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4844_ _3827_ _3771_ _3871_ vssd1 vssd1 vccd1 vccd1 _3999_ sky130_fd_sc_hd__or3_1
X_7632_ _2779_ _2781_ vssd1 vssd1 vccd1 vccd1 _2783_ sky130_fd_sc_hd__nand2_1
XFILLER_119_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4650__B _3804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4775_ _3722_ _3167_ _3746_ _3748_ vssd1 vssd1 vccd1 vccd1 _3930_ sky130_fd_sc_hd__nand4_4
XFILLER_20_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7563_ _2702_ _0390_ vssd1 vssd1 vccd1 vccd1 _2707_ sky130_fd_sc_hd__and2_1
XFILLER_119_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6514_ _1551_ _1417_ _1552_ vssd1 vssd1 vccd1 vccd1 _1553_ sky130_fd_sc_hd__o21a_2
XFILLER_119_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7494_ _3189_ _1803_ _2034_ _3232_ _2630_ vssd1 vssd1 vccd1 vccd1 _2631_ sky130_fd_sc_hd__o221a_1
XANTENNA__6858__A _1428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6445_ _1475_ _1476_ vssd1 vssd1 vccd1 vccd1 _1477_ sky130_fd_sc_hd__xnor2_1
X_6376_ _3817_ vssd1 vssd1 vccd1 vccd1 _1401_ sky130_fd_sc_hd__clkbuf_4
XFILLER_114_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5327_ _0298_ _0284_ vssd1 vssd1 vccd1 vccd1 _0300_ sky130_fd_sc_hd__or2b_1
XFILLER_0_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8115_ _1330_ _3305_ _3310_ vssd1 vssd1 vccd1 vccd1 _3311_ sky130_fd_sc_hd__a21oi_1
XANTENNA__5481__B _0440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8046_ _3229_ _3235_ vssd1 vssd1 vccd1 vccd1 _3237_ sky130_fd_sc_hd__or2_1
XFILLER_87_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5258_ _4157_ _4158_ _4160_ vssd1 vssd1 vccd1 vccd1 _0231_ sky130_fd_sc_hd__a21bo_1
XFILLER_68_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5189_ _0135_ _0156_ _0161_ vssd1 vssd1 vccd1 vccd1 _0162_ sky130_fd_sc_hd__o21ai_1
XFILLER_113_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5002__A _4016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5937__A _0762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8459__S _3655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7398__B2 _2335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6950__B _1718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4560_ _1858_ _2221_ _3714_ _2298_ vssd1 vssd1 vccd1 vccd1 _3715_ sky130_fd_sc_hd__a211o_1
XANTENNA__7570__A1 _4222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4491_ posit_add.in1\[2\] _3178_ vssd1 vssd1 vccd1 vccd1 _3189_ sky130_fd_sc_hd__xnor2_4
X_6230_ _0802_ _1095_ _1019_ _1102_ vssd1 vssd1 vccd1 vccd1 _1240_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__6397__B _1423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6161_ _1090_ _1089_ vssd1 vssd1 vccd1 vccd1 _1166_ sky130_fd_sc_hd__and2_1
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5112_ _4252_ _0084_ vssd1 vssd1 vccd1 vccd1 _0085_ sky130_fd_sc_hd__or2_1
X_6092_ _1091_ _1092_ vssd1 vssd1 vccd1 vccd1 _1094_ sky130_fd_sc_hd__xnor2_1
XFILLER_111_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5636__A1 _1748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5043_ _4194_ _4197_ vssd1 vssd1 vccd1 vccd1 _4198_ sky130_fd_sc_hd__xnor2_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6994_ _4217_ _2079_ _2080_ vssd1 vssd1 vccd1 vccd1 _2081_ sky130_fd_sc_hd__and3_1
XFILLER_53_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5945_ _0928_ _0929_ _0938_ vssd1 vssd1 vccd1 vccd1 _0939_ sky130_fd_sc_hd__a21o_1
XFILLER_80_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5876_ _3892_ _0634_ _0624_ _3832_ vssd1 vssd1 vccd1 vccd1 _0867_ sky130_fd_sc_hd__and4_1
XFILLER_80_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4661__A _3815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4827_ _3964_ _3980_ vssd1 vssd1 vccd1 vccd1 _3982_ sky130_fd_sc_hd__or2_1
XFILLER_21_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7615_ _2754_ _2763_ _2707_ vssd1 vssd1 vccd1 vccd1 _2764_ sky130_fd_sc_hd__mux2_1
X_4758_ _3891_ _3903_ _3912_ vssd1 vssd1 vccd1 vccd1 _3913_ sky130_fd_sc_hd__o21ai_2
XFILLER_5_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7546_ _2682_ _2685_ _2686_ vssd1 vssd1 vccd1 vccd1 _2688_ sky130_fd_sc_hd__o21ai_1
X_4689_ _3828_ _3750_ vssd1 vssd1 vccd1 vccd1 _3844_ sky130_fd_sc_hd__nor2_1
XANTENNA__6588__A _0080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7477_ _2381_ _2410_ _2589_ vssd1 vssd1 vccd1 vccd1 _2612_ sky130_fd_sc_hd__o21a_1
X_6428_ _1448_ _1453_ vssd1 vssd1 vccd1 vccd1 _1458_ sky130_fd_sc_hd__nand2_1
XFILLER_108_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6359_ _1375_ _1381_ vssd1 vssd1 vccd1 vccd1 _1382_ sky130_fd_sc_hd__xnor2_1
XFILLER_102_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4258__D in_reg\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8029_ _3217_ vssd1 vssd1 vccd1 vccd1 _3218_ sky130_fd_sc_hd__clkinv_2
XFILLER_17_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5667__A _4045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_498 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6929__C _1950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5866__A1 _2529_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8265__C1 _1177_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5730_ _0644_ _0708_ _0709_ vssd1 vssd1 vccd1 vccd1 _0710_ sky130_fd_sc_hd__nand3_1
XFILLER_95_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4481__A _2980_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5661_ _0631_ vssd1 vssd1 vccd1 vccd1 _0634_ sky130_fd_sc_hd__buf_2
X_7400_ _2454_ _2525_ _2526_ _2451_ vssd1 vssd1 vccd1 vccd1 _2527_ sky130_fd_sc_hd__o211a_1
X_4612_ _1803_ _3635_ _3712_ _2309_ vssd1 vssd1 vccd1 vccd1 _3767_ sky130_fd_sc_hd__a211o_1
X_8380_ _3590_ _0599_ _3591_ vssd1 vssd1 vccd1 vccd1 _3592_ sky130_fd_sc_hd__or3b_1
X_5592_ _0494_ _0564_ vssd1 vssd1 vccd1 vccd1 _0565_ sky130_fd_sc_hd__and2_1
X_4543_ _3690_ _2408_ _3696_ _1737_ vssd1 vssd1 vccd1 vccd1 _3698_ sky130_fd_sc_hd__a31o_1
X_7331_ _2450_ vssd1 vssd1 vccd1 vccd1 _2451_ sky130_fd_sc_hd__buf_2
X_7262_ _2347_ _2359_ _2370_ _2374_ vssd1 vssd1 vccd1 vccd1 _2376_ sky130_fd_sc_hd__a31oi_4
X_6213_ _1218_ _1219_ vssd1 vssd1 vccd1 vccd1 _1222_ sky130_fd_sc_hd__xnor2_1
X_4474_ _2881_ _2958_ _2991_ vssd1 vssd1 vccd1 vccd1 _3002_ sky130_fd_sc_hd__or3b_2
X_7193_ _0082_ _1446_ _0083_ vssd1 vssd1 vccd1 vccd1 _2300_ sky130_fd_sc_hd__o21ai_1
X_6144_ _1144_ _1147_ vssd1 vssd1 vccd1 vccd1 _1148_ sky130_fd_sc_hd__nand2_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6075_ _0942_ _1056_ _1074_ _0961_ _1075_ vssd1 vssd1 vccd1 vccd1 _1076_ sky130_fd_sc_hd__a311o_1
XFILLER_100_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7032__A _1711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5026_ _4179_ _4180_ vssd1 vssd1 vccd1 vccd1 _4181_ sky130_fd_sc_hd__xnor2_1
XFILLER_73_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6977_ _2060_ _2061_ vssd1 vssd1 vccd1 vccd1 _2062_ sky130_fd_sc_hd__xor2_1
XFILLER_53_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5928_ _0891_ _0919_ _0920_ vssd1 vssd1 vccd1 vccd1 _0921_ sky130_fd_sc_hd__nand3_1
XANTENNA__4596__A1 _2903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5859_ _0844_ _0847_ _0848_ _0759_ vssd1 vssd1 vccd1 vccd1 _0849_ sky130_fd_sc_hd__o211ai_2
XFILLER_21_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8578_ clknet_3_6__leaf_clk _0064_ vssd1 vssd1 vccd1 vccd1 posit_add.in2\[5\] sky130_fd_sc_hd__dfxtp_2
XFILLER_5_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7529_ _0369_ _2651_ vssd1 vssd1 vccd1 vccd1 _2669_ sky130_fd_sc_hd__xnor2_1
XFILLER_79_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4284__A0 in_reg\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6781__A _0147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5397__A _0369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6900_ _1976_ _1958_ vssd1 vssd1 vccd1 vccd1 _1977_ sky130_fd_sc_hd__xnor2_1
XFILLER_75_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7880_ _2941_ _3054_ vssd1 vssd1 vccd1 vccd1 _3055_ sky130_fd_sc_hd__or2_1
XANTENNA__8005__A2 _2621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6831_ _1890_ _1888_ vssd1 vssd1 vccd1 vccd1 _1901_ sky130_fd_sc_hd__xor2_1
XFILLER_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8501_ _3689_ vssd1 vssd1 vccd1 vccd1 _0068_ sky130_fd_sc_hd__clkbuf_1
X_6762_ _1804_ _1821_ vssd1 vssd1 vccd1 vccd1 _1826_ sky130_fd_sc_hd__nor2_1
XFILLER_50_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5713_ _3700_ _0686_ _0691_ _3923_ vssd1 vssd1 vccd1 vccd1 _0692_ sky130_fd_sc_hd__a211o_1
X_6693_ _1721_ _1747_ _1749_ vssd1 vssd1 vccd1 vccd1 _1750_ sky130_fd_sc_hd__a21o_1
X_5644_ _0616_ _0607_ _0614_ _3864_ _3718_ vssd1 vssd1 vccd1 vccd1 _0617_ sky130_fd_sc_hd__a221oi_1
X_8432_ counter\[1\] counter\[0\] _0786_ vssd1 vssd1 vccd1 vccd1 _3644_ sky130_fd_sc_hd__and3_1
XANTENNA__8411__A cmd\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8363_ _3571_ _3574_ vssd1 vssd1 vccd1 vccd1 _3575_ sky130_fd_sc_hd__xnor2_1
X_5575_ _4126_ vssd1 vssd1 vccd1 vccd1 _0548_ sky130_fd_sc_hd__clkbuf_4
X_7314_ _2432_ _2422_ _2416_ vssd1 vssd1 vccd1 vccd1 _2433_ sky130_fd_sc_hd__mux2_1
XFILLER_117_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4526_ _3232_ _3530_ _3552_ _3488_ vssd1 vssd1 vccd1 vccd1 _3562_ sky130_fd_sc_hd__o211ai_2
X_8294_ _3500_ vssd1 vssd1 vccd1 vccd1 _3501_ sky130_fd_sc_hd__clkinv_2
XFILLER_116_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4457_ posit_add.in1\[5\] posit_add.in1\[4\] _2551_ _1253_ vssd1 vssd1 vccd1 vccd1
+ _2815_ sky130_fd_sc_hd__o31a_1
X_7245_ _0430_ _0425_ vssd1 vssd1 vccd1 vccd1 _2357_ sky130_fd_sc_hd__nor2_1
XFILLER_104_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7176_ _2279_ _2280_ vssd1 vssd1 vccd1 vccd1 _2281_ sky130_fd_sc_hd__nor2_1
X_6127_ _0627_ _1095_ vssd1 vssd1 vccd1 vccd1 _1130_ sky130_fd_sc_hd__nor2_1
XFILLER_98_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4388_ posit_add.in2\[0\] _2034_ vssd1 vssd1 vccd1 vccd1 _2056_ sky130_fd_sc_hd__nor2_1
XFILLER_58_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6585__B _0082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6058_ _0956_ _0955_ _0957_ vssd1 vssd1 vccd1 vccd1 _1058_ sky130_fd_sc_hd__and3_1
XFILLER_46_619 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5009_ _4162_ _4163_ vssd1 vssd1 vccd1 vccd1 _4164_ sky130_fd_sc_hd__xnor2_1
XFILLER_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4569__A1 _2969_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8180__A1 _3378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8467__S _3654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5049__A2 _4153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5839__B _0754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5360_ _0079_ _0089_ _0132_ _0332_ vssd1 vssd1 vccd1 vccd1 _0333_ sky130_fd_sc_hd__a31oi_1
XFILLER_114_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5291_ _0260_ _0262_ vssd1 vssd1 vccd1 vccd1 _0264_ sky130_fd_sc_hd__nand2_1
X_4311_ _1199_ vssd1 vssd1 vccd1 vccd1 _0019_ sky130_fd_sc_hd__clkbuf_1
XFILLER_114_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7030_ _2119_ vssd1 vssd1 vccd1 vccd1 _2120_ sky130_fd_sc_hd__inv_2
XANTENNA__7682__A0 _3925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4918__B _3702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7013__C _1538_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4934__A _3883_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7932_ _2937_ _3041_ _3111_ vssd1 vssd1 vccd1 vccd1 _3113_ sky130_fd_sc_hd__a21o_1
X_7863_ _2948_ _3034_ _3036_ vssd1 vssd1 vccd1 vccd1 _3037_ sky130_fd_sc_hd__o21ai_1
XFILLER_23_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6814_ _1862_ _1882_ vssd1 vssd1 vccd1 vccd1 _1883_ sky130_fd_sc_hd__xnor2_1
XFILLER_50_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7794_ _2954_ _2955_ vssd1 vssd1 vccd1 vccd1 _2961_ sky130_fd_sc_hd__xor2_1
X_6745_ _1428_ _1510_ _1806_ vssd1 vssd1 vccd1 vccd1 _1807_ sky130_fd_sc_hd__o21ba_1
XFILLER_51_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6676_ _1724_ _1730_ vssd1 vssd1 vccd1 vccd1 _1731_ sky130_fd_sc_hd__xnor2_1
X_8415_ _1253_ _0082_ _2319_ _1330_ _3628_ vssd1 vssd1 vccd1 vccd1 _3629_ sky130_fd_sc_hd__a221o_1
X_5627_ _0599_ vssd1 vssd1 vccd1 vccd1 _0600_ sky130_fd_sc_hd__clkbuf_4
X_8346_ _0451_ _3259_ _3553_ _3554_ _3555_ vssd1 vssd1 vccd1 vccd1 _3556_ sky130_fd_sc_hd__a221oi_4
X_5558_ _0529_ _0530_ _0480_ vssd1 vssd1 vccd1 vccd1 _0531_ sky130_fd_sc_hd__mux2_1
XFILLER_117_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4509_ _2661_ _3232_ vssd1 vssd1 vccd1 vccd1 _3381_ sky130_fd_sc_hd__xor2_1
XFILLER_3_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8277_ _3416_ _3482_ vssd1 vssd1 vccd1 vccd1 _3483_ sky130_fd_sc_hd__and2b_1
X_5489_ _0461_ _0401_ vssd1 vssd1 vccd1 vccd1 _0462_ sky130_fd_sc_hd__or2_1
X_7228_ _0388_ _2336_ _2337_ vssd1 vssd1 vccd1 vccd1 _2338_ sky130_fd_sc_hd__a21oi_1
XFILLER_116_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5005__A _3701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7159_ _1765_ vssd1 vssd1 vccd1 vccd1 _2262_ sky130_fd_sc_hd__inv_2
XFILLER_100_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4844__A _3827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5659__B _0627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5203__A2 _3840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7874__B _2937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7114__B _4089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8226__A _0440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4860_ _1352_ _1374_ _1396_ _1407_ vssd1 vssd1 vccd1 vccd1 _4015_ sky130_fd_sc_hd__or4_2
XFILLER_60_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_644 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4791_ _3816_ _3702_ _3945_ vssd1 vssd1 vccd1 vccd1 _3946_ sky130_fd_sc_hd__or3_1
X_6530_ _1569_ _1568_ vssd1 vssd1 vccd1 vccd1 _1570_ sky130_fd_sc_hd__xnor2_2
XFILLER_13_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6461_ _1487_ _1488_ vssd1 vssd1 vccd1 vccd1 _1494_ sky130_fd_sc_hd__nand2_1
X_6392_ _1416_ _1417_ vssd1 vssd1 vccd1 vccd1 _1419_ sky130_fd_sc_hd__and2_1
X_5412_ _0384_ _3733_ _3729_ vssd1 vssd1 vccd1 vccd1 _0385_ sky130_fd_sc_hd__mux2_2
X_8200_ _3321_ _3354_ vssd1 vssd1 vccd1 vccd1 _3401_ sky130_fd_sc_hd__or2b_1
XFILLER_114_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5343_ _0315_ _0308_ vssd1 vssd1 vccd1 vccd1 _0316_ sky130_fd_sc_hd__xnor2_1
X_8131_ _3158_ _3326_ _3234_ vssd1 vssd1 vccd1 vccd1 _3327_ sky130_fd_sc_hd__mux2_1
XFILLER_114_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5274_ _0241_ _0245_ _0246_ vssd1 vssd1 vccd1 vccd1 _0247_ sky130_fd_sc_hd__o21ai_2
X_8062_ _3249_ _3252_ vssd1 vssd1 vccd1 vccd1 _3254_ sky130_fd_sc_hd__xor2_4
XFILLER_102_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7013_ _1401_ _1782_ _1538_ _2063_ vssd1 vssd1 vccd1 vccd1 _2102_ sky130_fd_sc_hd__or4_1
XANTENNA__5130__A1 _3802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7407__B1 _2534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4664__A posit_add.in1\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_419 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7915_ _3042_ _3081_ _3093_ vssd1 vssd1 vccd1 vccd1 _3094_ sky130_fd_sc_hd__o21ai_1
XFILLER_62_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7846_ _2987_ _3017_ vssd1 vssd1 vccd1 vccd1 _3018_ sky130_fd_sc_hd__and2_1
XANTENNA__7694__B _2802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8383__A1 _3182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7777_ _2673_ _2941_ vssd1 vssd1 vccd1 vccd1 _2942_ sky130_fd_sc_hd__or2_1
X_4989_ _4141_ _4142_ vssd1 vssd1 vccd1 vccd1 _4144_ sky130_fd_sc_hd__and2b_1
X_6728_ _1408_ _1409_ _0147_ vssd1 vssd1 vccd1 vccd1 _1788_ sky130_fd_sc_hd__and3_1
X_6659_ _1221_ _1224_ _1225_ vssd1 vssd1 vccd1 vccd1 _1712_ sky130_fd_sc_hd__a21oi_1
X_8329_ _3536_ _3537_ vssd1 vssd1 vccd1 vccd1 _3538_ sky130_fd_sc_hd__or2_1
XFILLER_117_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5121__A1 _0092_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5389__B _2507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5961_ _0937_ _0934_ _0936_ vssd1 vssd1 vccd1 vccd1 _0956_ sky130_fd_sc_hd__nand3_1
XFILLER_80_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4912_ _4048_ _4064_ _4066_ vssd1 vssd1 vccd1 vccd1 _4067_ sky130_fd_sc_hd__a21bo_1
X_7700_ _2676_ _2762_ vssd1 vssd1 vccd1 vccd1 _2857_ sky130_fd_sc_hd__nor2_1
X_5892_ _0853_ _0882_ vssd1 vssd1 vccd1 vccd1 _0884_ sky130_fd_sc_hd__xnor2_2
X_7631_ _2780_ vssd1 vssd1 vccd1 vccd1 _2781_ sky130_fd_sc_hd__inv_2
X_4843_ _3881_ _3883_ _3880_ _3997_ vssd1 vssd1 vccd1 vccd1 _3998_ sky130_fd_sc_hd__a31o_1
XFILLER_21_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4774_ _3926_ _3704_ _3928_ vssd1 vssd1 vccd1 vccd1 _3929_ sky130_fd_sc_hd__o21a_1
XFILLER_60_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7562_ _0375_ _2668_ vssd1 vssd1 vccd1 vccd1 _2706_ sky130_fd_sc_hd__xor2_2
X_6513_ _1420_ _1410_ _1415_ vssd1 vssd1 vccd1 vccd1 _1552_ sky130_fd_sc_hd__o21ai_1
X_7493_ posit_add.in1\[1\] _2034_ _3765_ _2969_ vssd1 vssd1 vccd1 vccd1 _2630_ sky130_fd_sc_hd__a211o_1
XFILLER_119_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6444_ _1383_ _3840_ vssd1 vssd1 vccd1 vccd1 _1476_ sky130_fd_sc_hd__or2_1
XANTENNA__6858__B _1718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6375_ _1399_ vssd1 vssd1 vccd1 vccd1 _1400_ sky130_fd_sc_hd__clkbuf_4
XFILLER_114_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5326_ _0284_ _0298_ vssd1 vssd1 vccd1 vccd1 _0299_ sky130_fd_sc_hd__or2b_1
XFILLER_0_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8114_ _3265_ _3309_ vssd1 vssd1 vccd1 vccd1 _3310_ sky130_fd_sc_hd__xor2_2
XFILLER_114_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5257_ _0183_ _0187_ vssd1 vssd1 vccd1 vccd1 _0230_ sky130_fd_sc_hd__xnor2_1
XFILLER_57_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8045_ _3229_ _3235_ vssd1 vssd1 vccd1 vccd1 _3236_ sky130_fd_sc_hd__nand2_1
XFILLER_88_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5188_ _0159_ _0160_ vssd1 vssd1 vccd1 vccd1 _0161_ sky130_fd_sc_hd__or2_1
XFILLER_28_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5002__B _3702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5937__B _3832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7829_ _2998_ vssd1 vssd1 vccd1 vccd1 _2999_ sky130_fd_sc_hd__clkbuf_4
XFILLER_24_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5953__A _3792_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4550__C1 _1682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8475__S _3654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8347__A1 _1330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_4__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_4__leaf_clk sky130_fd_sc_hd__clkbuf_16
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4490_ posit_add.in1\[0\] posit_add.in1\[1\] _1242_ vssd1 vssd1 vccd1 vccd1 _3178_
+ sky130_fd_sc_hd__o21ai_2
XFILLER_7_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4479__A _1253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6160_ _1090_ _1164_ vssd1 vssd1 vccd1 vccd1 _1165_ sky130_fd_sc_hd__nor2_1
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_411 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5111_ _3925_ _0082_ _0083_ vssd1 vssd1 vccd1 vccd1 _0084_ sky130_fd_sc_hd__o21a_1
X_6091_ _0884_ _0981_ vssd1 vssd1 vccd1 vccd1 _1092_ sky130_fd_sc_hd__xor2_2
XFILLER_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5636__A2 _2507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5042_ _4195_ _4027_ _4196_ vssd1 vssd1 vccd1 vccd1 _4197_ sky130_fd_sc_hd__o21ba_1
XFILLER_84_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6993_ _2075_ _2076_ vssd1 vssd1 vccd1 vccd1 _2080_ sky130_fd_sc_hd__xor2_1
XFILLER_65_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5944_ _0934_ _0936_ _0937_ vssd1 vssd1 vccd1 vccd1 _0938_ sky130_fd_sc_hd__a21bo_1
XFILLER_80_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4942__A _2540_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5875_ _0837_ _0838_ _0839_ vssd1 vssd1 vccd1 vccd1 _0866_ sky130_fd_sc_hd__nand3_1
X_4826_ _3964_ _3980_ vssd1 vssd1 vccd1 vccd1 _3981_ sky130_fd_sc_hd__xnor2_1
X_7614_ _0147_ _4045_ _2652_ vssd1 vssd1 vccd1 vccd1 _2763_ sky130_fd_sc_hd__mux2_1
XANTENNA__5021__B1 _3989_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7545_ _2682_ _2685_ _2686_ vssd1 vssd1 vccd1 vccd1 _2687_ sky130_fd_sc_hd__or3_1
XANTENNA__5773__A _3924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4757_ _3910_ _3911_ vssd1 vssd1 vccd1 vccd1 _3912_ sky130_fd_sc_hd__or2b_1
XFILLER_119_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4688_ _3818_ _3842_ vssd1 vssd1 vccd1 vccd1 _3843_ sky130_fd_sc_hd__xnor2_1
XANTENNA__6588__B _1400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7476_ _2520_ vssd1 vssd1 vccd1 vccd1 _2611_ sky130_fd_sc_hd__inv_2
X_6427_ _4250_ _0147_ _1455_ _1456_ vssd1 vssd1 vccd1 vccd1 _1457_ sky130_fd_sc_hd__or4_2
X_6358_ _1378_ _1380_ vssd1 vssd1 vccd1 vccd1 _1381_ sky130_fd_sc_hd__nand2_1
XANTENNA__7077__A1 _1456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5309_ _0280_ _0281_ vssd1 vssd1 vccd1 vccd1 _0282_ sky130_fd_sc_hd__nor2_1
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6289_ _1257_ _1302_ _1303_ _1304_ vssd1 vssd1 vccd1 vccd1 _1305_ sky130_fd_sc_hd__o211a_1
XFILLER_88_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4835__B1 _3989_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8028_ _0557_ _0569_ _3216_ vssd1 vssd1 vccd1 vccd1 _3217_ sky130_fd_sc_hd__o21ai_2
XFILLER_91_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8026__A0 _0451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7212__B _2319_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_588 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6779__A _1383_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5866__A2 _0773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7068__A1 _1676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6019__A _0779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4762__A _3736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8234__A _2993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5660_ _3700_ _0626_ _3923_ vssd1 vssd1 vccd1 vccd1 _0633_ sky130_fd_sc_hd__o21a_2
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4611_ _3765_ _2408_ _2452_ vssd1 vssd1 vccd1 vccd1 _3766_ sky130_fd_sc_hd__or3_1
X_5591_ _0530_ _0532_ _0480_ vssd1 vssd1 vccd1 vccd1 _0564_ sky130_fd_sc_hd__mux2_1
X_4542_ _2430_ _2452_ _2463_ vssd1 vssd1 vccd1 vccd1 _3696_ sky130_fd_sc_hd__o21a_1
X_7330_ _2449_ _2426_ _2427_ vssd1 vssd1 vccd1 vccd1 _2450_ sky130_fd_sc_hd__and3b_1
X_4473_ _2969_ posit_add.in1\[2\] posit_add.in1\[1\] _2980_ vssd1 vssd1 vccd1 vccd1
+ _2991_ sky130_fd_sc_hd__or4_1
X_7261_ _2361_ _2373_ _2368_ vssd1 vssd1 vccd1 vccd1 _2374_ sky130_fd_sc_hd__o21a_1
X_6212_ _1218_ _1219_ vssd1 vssd1 vccd1 vccd1 _1221_ sky130_fd_sc_hd__nand2_1
X_7192_ _2282_ _2283_ _2285_ vssd1 vssd1 vccd1 vccd1 _2299_ sky130_fd_sc_hd__or3b_1
XFILLER_112_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6143_ _1145_ _1146_ vssd1 vssd1 vccd1 vccd1 _1147_ sky130_fd_sc_hd__and2_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6074_ _0942_ _0960_ vssd1 vssd1 vccd1 vccd1 _1075_ sky130_fd_sc_hd__and2_1
XFILLER_100_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7032__B _1355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5025_ _4000_ _4001_ _3999_ vssd1 vssd1 vccd1 vccd1 _4180_ sky130_fd_sc_hd__a21bo_1
XANTENNA__8008__B1 _3194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6976_ _2011_ _2026_ vssd1 vssd1 vccd1 vccd1 _2061_ sky130_fd_sc_hd__xor2_1
XFILLER_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5927_ _0917_ _0918_ _0909_ vssd1 vssd1 vccd1 vccd1 _0920_ sky130_fd_sc_hd__a21o_1
XANTENNA__4391__B _1858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5858_ _0729_ _0730_ _0758_ vssd1 vssd1 vccd1 vccd1 _0848_ sky130_fd_sc_hd__o21ai_1
X_5789_ _0693_ vssd1 vssd1 vccd1 vccd1 _0773_ sky130_fd_sc_hd__clkbuf_4
X_8577_ clknet_3_6__leaf_clk _0063_ vssd1 vssd1 vccd1 vccd1 posit_add.in2\[4\] sky130_fd_sc_hd__dfxtp_2
X_4809_ _3939_ _3951_ vssd1 vssd1 vccd1 vccd1 _3964_ sky130_fd_sc_hd__xnor2_1
XFILLER_21_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7528_ _0388_ _2651_ _2667_ _0386_ vssd1 vssd1 vccd1 vccd1 _2668_ sky130_fd_sc_hd__a211o_1
X_7459_ _2587_ _2591_ _2569_ vssd1 vssd1 vccd1 vccd1 _2592_ sky130_fd_sc_hd__mux2_1
XFILLER_115_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4582__A _3736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6830_ _1896_ _1899_ vssd1 vssd1 vccd1 vccd1 _1900_ sky130_fd_sc_hd__nor2_1
XFILLER_90_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6761_ _1786_ _1823_ vssd1 vssd1 vccd1 vccd1 _1824_ sky130_fd_sc_hd__xnor2_1
X_8500_ posit_add.in2\[9\] in_reg\[9\] _3677_ vssd1 vssd1 vccd1 vccd1 _3689_ sky130_fd_sc_hd__mux2_1
X_5712_ _3718_ _0687_ _0688_ _0689_ _3801_ vssd1 vssd1 vccd1 vccd1 _0691_ sky130_fd_sc_hd__o311a_1
XFILLER_50_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6692_ _1724_ _1730_ vssd1 vssd1 vccd1 vccd1 _1749_ sky130_fd_sc_hd__nor2_1
XFILLER_31_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7516__A2 _3635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5643_ _2507_ _3775_ vssd1 vssd1 vccd1 vccd1 _0616_ sky130_fd_sc_hd__nand2_2
X_8431_ counter\[0\] _3242_ _3642_ vssd1 vssd1 vccd1 vccd1 _0038_ sky130_fd_sc_hd__a21oi_1
XANTENNA__8411__B cmd\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8362_ _3481_ _3532_ _3572_ vssd1 vssd1 vccd1 vccd1 _3574_ sky130_fd_sc_hd__or3b_1
X_5574_ _4140_ _0546_ vssd1 vssd1 vccd1 vccd1 _0547_ sky130_fd_sc_hd__nor2_1
XFILLER_116_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4525_ _3079_ _3296_ _3189_ _3046_ vssd1 vssd1 vccd1 vccd1 _3552_ sky130_fd_sc_hd__a211o_1
XANTENNA__8477__A0 in_reg\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7313_ _1899_ _2428_ _2429_ _2431_ vssd1 vssd1 vccd1 vccd1 _2432_ sky130_fd_sc_hd__o211a_1
X_8293_ _2611_ _3251_ vssd1 vssd1 vccd1 vccd1 _3500_ sky130_fd_sc_hd__and2_1
XANTENNA__5473__D _0445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4456_ _2793_ vssd1 vssd1 vccd1 vccd1 _2804_ sky130_fd_sc_hd__inv_2
X_7244_ _2355_ vssd1 vssd1 vccd1 vccd1 _2356_ sky130_fd_sc_hd__inv_2
X_4387_ _1506_ _1803_ vssd1 vssd1 vccd1 vccd1 _2045_ sky130_fd_sc_hd__or2_1
X_7175_ _1637_ _2278_ vssd1 vssd1 vccd1 vccd1 _2280_ sky130_fd_sc_hd__and2_1
X_6126_ _1096_ _1102_ _1120_ _1121_ vssd1 vssd1 vccd1 vccd1 _1129_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_98_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6057_ _0949_ _0958_ vssd1 vssd1 vccd1 vccd1 _1057_ sky130_fd_sc_hd__nand2_1
XFILLER_85_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5008_ _4017_ _3726_ _3927_ _4020_ vssd1 vssd1 vccd1 vccd1 _4163_ sky130_fd_sc_hd__o31a_1
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6959_ _2040_ _2041_ vssd1 vssd1 vccd1 vccd1 _2042_ sky130_fd_sc_hd__xor2_1
XFILLER_10_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5757__A1 _2507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6032__A _0773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8459__A0 in_reg\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6967__A _0147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5290_ _0260_ _0262_ vssd1 vssd1 vccd1 vccd1 _0263_ sky130_fd_sc_hd__or2_1
X_4310_ _0635_ _1188_ vssd1 vssd1 vccd1 vccd1 _1199_ sky130_fd_sc_hd__and2b_1
XFILLER_114_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7682__A1 _0080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4496__A1 _3232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7931_ _3110_ _3070_ _3038_ vssd1 vssd1 vccd1 vccd1 _3111_ sky130_fd_sc_hd__mux2_1
XFILLER_48_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7862_ _2950_ _3034_ vssd1 vssd1 vccd1 vccd1 _3036_ sky130_fd_sc_hd__or2b_1
XFILLER_35_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6813_ _1878_ _1881_ _1876_ vssd1 vssd1 vccd1 vccd1 _1882_ sky130_fd_sc_hd__a21o_1
XFILLER_51_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7793_ _2956_ _2959_ vssd1 vssd1 vccd1 vccd1 _2960_ sky130_fd_sc_hd__nor2_1
X_6744_ _4232_ _1664_ vssd1 vssd1 vccd1 vccd1 _1806_ sky130_fd_sc_hd__nor2_1
XFILLER_23_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6675_ _1727_ _1729_ vssd1 vssd1 vccd1 vccd1 _1730_ sky130_fd_sc_hd__xnor2_1
X_5626_ _0092_ cmd\[7\] cmd\[6\] vssd1 vssd1 vccd1 vccd1 _0599_ sky130_fd_sc_hd__or3b_4
X_8414_ cmd\[6\] _3186_ _3627_ cmd\[7\] vssd1 vssd1 vccd1 vccd1 _3628_ sky130_fd_sc_hd__a22oi_1
XFILLER_117_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8345_ _3553_ _3554_ vssd1 vssd1 vccd1 vccd1 _3555_ sky130_fd_sc_hd__nor2_1
X_5557_ _0490_ _0484_ _0470_ vssd1 vssd1 vccd1 vccd1 _0530_ sky130_fd_sc_hd__mux2_1
XFILLER_117_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4508_ _3339_ _3349_ _2826_ _3360_ vssd1 vssd1 vccd1 vccd1 _3371_ sky130_fd_sc_hd__o211a_1
X_8276_ _2514_ _3203_ _3205_ _2604_ vssd1 vssd1 vccd1 vccd1 _3482_ sky130_fd_sc_hd__a211o_2
X_5488_ _0092_ _0399_ vssd1 vssd1 vccd1 vccd1 _0461_ sky130_fd_sc_hd__nor2_1
XANTENNA__4397__A _1781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4439_ posit_add.in1\[7\] _2562_ vssd1 vssd1 vccd1 vccd1 _2617_ sky130_fd_sc_hd__or2_1
X_7227_ _0387_ _2335_ vssd1 vssd1 vccd1 vccd1 _2337_ sky130_fd_sc_hd__nor2_1
XFILLER_104_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7158_ _1773_ _2256_ _2260_ _1900_ vssd1 vssd1 vccd1 vccd1 _2261_ sky130_fd_sc_hd__or4bb_1
X_6109_ _1029_ _1110_ _1031_ vssd1 vssd1 vccd1 vccd1 _1111_ sky130_fd_sc_hd__a21oi_1
XFILLER_100_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7089_ _1664_ _1782_ _4126_ _2157_ vssd1 vssd1 vccd1 vccd1 _2185_ sky130_fd_sc_hd__or4_1
XANTENNA__5005__B _3795_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4844__B _3771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5659__C _3735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6787__A _1399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7114__C _1950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4473__C posit_add.in1\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4770__A _3924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4790_ _3942_ _3944_ _3756_ vssd1 vssd1 vccd1 vccd1 _3945_ sky130_fd_sc_hd__a21o_1
XFILLER_13_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6155__B2 _0762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6460_ _1480_ _1492_ vssd1 vssd1 vccd1 vccd1 _1493_ sky130_fd_sc_hd__xnor2_1
XFILLER_9_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6391_ _0303_ _1410_ vssd1 vssd1 vccd1 vccd1 _1417_ sky130_fd_sc_hd__or2_1
X_5411_ _3736_ _0382_ _0383_ vssd1 vssd1 vccd1 vccd1 _0384_ sky130_fd_sc_hd__o21ai_1
XFILLER_99_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5342_ _2540_ _3988_ vssd1 vssd1 vccd1 vccd1 _0315_ sky130_fd_sc_hd__nor2_1
X_8130_ _3021_ _3163_ _3028_ vssd1 vssd1 vccd1 vccd1 _3326_ sky130_fd_sc_hd__o21ba_1
XFILLER_99_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8061_ _2602_ _3251_ _2520_ vssd1 vssd1 vccd1 vccd1 _3252_ sky130_fd_sc_hd__mux2_2
XFILLER_114_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7012_ _2088_ vssd1 vssd1 vccd1 vccd1 _2101_ sky130_fd_sc_hd__inv_2
XFILLER_101_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5273_ _0201_ _0199_ vssd1 vssd1 vccd1 vccd1 _0246_ sky130_fd_sc_hd__xnor2_1
XFILLER_101_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5130__A2 _3838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7407__B2 _2416_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7914_ _3042_ _3092_ vssd1 vssd1 vccd1 vccd1 _3093_ sky130_fd_sc_hd__nand2_1
XFILLER_24_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7845_ _2986_ _2939_ _2985_ vssd1 vssd1 vccd1 vccd1 _3017_ sky130_fd_sc_hd__or3_1
XFILLER_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7776_ _2904_ _2940_ vssd1 vssd1 vccd1 vccd1 _2941_ sky130_fd_sc_hd__nor2_2
XFILLER_23_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5495__B1_N _0467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4988_ _4141_ _4142_ vssd1 vssd1 vccd1 vccd1 _4143_ sky130_fd_sc_hd__xnor2_1
XFILLER_109_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6727_ _1410_ _1401_ vssd1 vssd1 vccd1 vccd1 _1787_ sky130_fd_sc_hd__or2_1
XFILLER_109_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6658_ _1257_ _1302_ vssd1 vssd1 vccd1 vccd1 _1711_ sky130_fd_sc_hd__or2_2
X_5609_ _0510_ _0555_ _0575_ _0560_ _0557_ vssd1 vssd1 vccd1 vccd1 _0582_ sky130_fd_sc_hd__a32o_1
XANTENNA__6400__A _1353_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6589_ _0080_ _1400_ _1631_ vssd1 vssd1 vccd1 vccd1 _1635_ sky130_fd_sc_hd__o21ai_1
X_8328_ _3508_ _3535_ vssd1 vssd1 vccd1 vccd1 _3537_ sky130_fd_sc_hd__nor2_1
XFILLER_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8259_ _3259_ _0528_ vssd1 vssd1 vccd1 vccd1 _3464_ sky130_fd_sc_hd__nor2_1
XFILLER_78_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7231__A _0369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_387 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5960_ _0951_ _0954_ vssd1 vssd1 vccd1 vccd1 _0955_ sky130_fd_sc_hd__and2_1
XANTENNA__6980__A _1401_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5891_ _0863_ _0880_ _0881_ vssd1 vssd1 vccd1 vccd1 _0882_ sky130_fd_sc_hd__a21boi_1
X_4911_ _2540_ _3817_ _4065_ vssd1 vssd1 vccd1 vccd1 _4066_ sky130_fd_sc_hd__or3_1
X_7630_ _3793_ _3795_ _2713_ vssd1 vssd1 vccd1 vccd1 _2780_ sky130_fd_sc_hd__mux2_1
X_4842_ _3875_ _3879_ vssd1 vssd1 vccd1 vccd1 _3997_ sky130_fd_sc_hd__nor2_1
XFILLER_60_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4773_ _3927_ _3805_ vssd1 vssd1 vccd1 vccd1 _3928_ sky130_fd_sc_hd__or2_1
X_7561_ _2703_ vssd1 vssd1 vccd1 vccd1 _2704_ sky130_fd_sc_hd__buf_2
X_6512_ _4153_ _1414_ vssd1 vssd1 vccd1 vccd1 _1551_ sky130_fd_sc_hd__nand2_1
X_7492_ _1913_ vssd1 vssd1 vccd1 vccd1 _2629_ sky130_fd_sc_hd__inv_2
XFILLER_107_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6443_ _4217_ _1353_ _1354_ vssd1 vssd1 vccd1 vccd1 _1475_ sky130_fd_sc_hd__and3_1
XFILLER_106_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6220__A _0762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6374_ _1397_ _1398_ vssd1 vssd1 vccd1 vccd1 _1399_ sky130_fd_sc_hd__xor2_4
XFILLER_114_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5325_ _0285_ _0296_ _0297_ vssd1 vssd1 vccd1 vccd1 _0298_ sky130_fd_sc_hd__o21ai_1
X_8113_ _0586_ _3308_ _3259_ vssd1 vssd1 vccd1 vccd1 _3309_ sky130_fd_sc_hd__mux2_1
XFILLER_114_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5256_ _0227_ _0228_ vssd1 vssd1 vccd1 vccd1 _0229_ sky130_fd_sc_hd__nor2_1
X_8044_ _3124_ _3233_ _3234_ vssd1 vssd1 vccd1 vccd1 _3235_ sky130_fd_sc_hd__mux2_1
XFILLER_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7051__A _4089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5187_ _0135_ _0156_ vssd1 vssd1 vccd1 vccd1 _0160_ sky130_fd_sc_hd__xnor2_1
XANTENNA__8053__A1 _3213_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7828_ _2996_ _2997_ vssd1 vssd1 vccd1 vccd1 _2998_ sky130_fd_sc_hd__nand2_4
X_7759_ _2812_ _2872_ _1308_ vssd1 vssd1 vccd1 vccd1 _2922_ sky130_fd_sc_hd__mux2_1
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7226__A _0385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6784__B _4089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6090_ _1053_ _1078_ _1089_ _1090_ vssd1 vssd1 vccd1 vccd1 _1091_ sky130_fd_sc_hd__a211o_1
XFILLER_97_423 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5110_ _4228_ _4250_ vssd1 vssd1 vccd1 vccd1 _0083_ sky130_fd_sc_hd__or2_1
XFILLER_97_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5041_ _4009_ _4010_ vssd1 vssd1 vccd1 vccd1 _4196_ sky130_fd_sc_hd__and2b_1
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4495__A posit_add.in1\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6992_ _2077_ vssd1 vssd1 vccd1 vccd1 _2079_ sky130_fd_sc_hd__buf_2
XFILLER_53_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5943_ _0905_ _0930_ _0933_ vssd1 vssd1 vccd1 vccd1 _0937_ sky130_fd_sc_hd__or3b_1
XANTENNA__4942__B _3930_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5874_ _0844_ _0845_ _0846_ vssd1 vssd1 vccd1 vccd1 _0865_ sky130_fd_sc_hd__o21ai_1
XFILLER_61_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5021__A1 _3793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4825_ _3965_ _3978_ _3979_ vssd1 vssd1 vccd1 vccd1 _3980_ sky130_fd_sc_hd__a21oi_1
X_7613_ _2729_ _2702_ vssd1 vssd1 vccd1 vccd1 _2762_ sky130_fd_sc_hd__nand2_2
XANTENNA__5021__B2 _3771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7745__S _1297_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7544_ _0406_ _0403_ _2652_ vssd1 vssd1 vccd1 vccd1 _2686_ sky130_fd_sc_hd__mux2_1
X_4756_ _3891_ _3903_ vssd1 vssd1 vccd1 vccd1 _3911_ sky130_fd_sc_hd__xor2_1
XFILLER_119_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4687_ _3829_ _3839_ _3841_ vssd1 vssd1 vccd1 vccd1 _3842_ sky130_fd_sc_hd__o21ba_1
X_7475_ _2607_ _2609_ _1308_ vssd1 vssd1 vccd1 vccd1 _2610_ sky130_fd_sc_hd__a21o_1
X_6426_ _3930_ vssd1 vssd1 vccd1 vccd1 _1456_ sky130_fd_sc_hd__clkbuf_4
XFILLER_115_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6357_ _1350_ _1050_ _1377_ _1333_ _1379_ vssd1 vssd1 vccd1 vccd1 _1380_ sky130_fd_sc_hd__o221a_1
XANTENNA__7077__A2 _1538_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5308_ _0279_ _0275_ _0277_ vssd1 vssd1 vccd1 vccd1 _0281_ sky130_fd_sc_hd__and3_1
XFILLER_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6288_ _1227_ _1256_ vssd1 vssd1 vccd1 vccd1 _1304_ sky130_fd_sc_hd__or2_1
XFILLER_88_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4835__A1 _3828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5239_ _3881_ _3986_ _4177_ vssd1 vssd1 vccd1 vccd1 _0212_ sky130_fd_sc_hd__and3_1
XFILLER_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8027_ _0557_ _3215_ vssd1 vssd1 vccd1 vccd1 _3216_ sky130_fd_sc_hd__nand2_1
XFILLER_29_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5493__D1 _0440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6779__B _4126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7068__A2 _1537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4610_ posit_add.in2\[0\] vssd1 vssd1 vccd1 vccd1 _3765_ sky130_fd_sc_hd__inv_2
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5590_ _0535_ _0562_ vssd1 vssd1 vccd1 vccd1 _0563_ sky130_fd_sc_hd__and2_1
X_4541_ _1990_ vssd1 vssd1 vccd1 vccd1 _3690_ sky130_fd_sc_hd__clkbuf_4
XFILLER_116_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4472_ _2661_ vssd1 vssd1 vccd1 vccd1 _2980_ sky130_fd_sc_hd__inv_4
X_7260_ _2362_ _2372_ _2367_ vssd1 vssd1 vccd1 vccd1 _2373_ sky130_fd_sc_hd__o21ai_1
X_6211_ _1173_ _1182_ vssd1 vssd1 vccd1 vccd1 _1219_ sky130_fd_sc_hd__xor2_1
X_7191_ _2295_ _2296_ vssd1 vssd1 vccd1 vccd1 _2297_ sky130_fd_sc_hd__nand2_1
X_6142_ _1015_ _1031_ _1029_ vssd1 vssd1 vccd1 vccd1 _1146_ sky130_fd_sc_hd__or3_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6073_ _1067_ _1071_ _1073_ vssd1 vssd1 vccd1 vccd1 _1074_ sky130_fd_sc_hd__a21o_1
XANTENNA__4817__A1 _3739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7032__C _1950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5024_ _4172_ _4178_ vssd1 vssd1 vccd1 vccd1 _4179_ sky130_fd_sc_hd__xnor2_1
XANTENNA__4817__B2 _3735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8008__B2 _3195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6975_ _2048_ _2059_ vssd1 vssd1 vccd1 vccd1 _2060_ sky130_fd_sc_hd__or2b_1
XFILLER_81_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5926_ _0909_ _0917_ _0918_ vssd1 vssd1 vccd1 vccd1 _0919_ sky130_fd_sc_hd__nand3_1
XFILLER_81_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5857_ _0844_ _0845_ _0846_ vssd1 vssd1 vccd1 vccd1 _0847_ sky130_fd_sc_hd__nor3_1
XFILLER_70_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5788_ _3763_ _0702_ vssd1 vssd1 vccd1 vccd1 _0772_ sky130_fd_sc_hd__nor2_1
X_8576_ clknet_3_6__leaf_clk _0062_ vssd1 vssd1 vccd1 vccd1 posit_add.in2\[3\] sky130_fd_sc_hd__dfxtp_2
X_4808_ _3800_ _3726_ _3962_ vssd1 vssd1 vccd1 vccd1 _3963_ sky130_fd_sc_hd__or3_1
XFILLER_119_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4739_ _3167_ _3509_ _3573_ _3772_ vssd1 vssd1 vccd1 vccd1 _3894_ sky130_fd_sc_hd__a211oi_4
X_7527_ _0385_ _2651_ vssd1 vssd1 vccd1 vccd1 _2667_ sky130_fd_sc_hd__nor2_1
XFILLER_107_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7458_ _2451_ _2578_ _2590_ vssd1 vssd1 vccd1 vccd1 _2591_ sky130_fd_sc_hd__a21oi_1
X_6409_ _1371_ _1436_ _1394_ vssd1 vssd1 vccd1 vccd1 _1437_ sky130_fd_sc_hd__a21o_1
XFILLER_79_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7389_ _2495_ _2513_ _2514_ vssd1 vssd1 vccd1 vccd1 _2515_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7223__B _0687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4863__A _4017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5769__C1 _3924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8486__A1 in_reg\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7414__A _0548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5869__A _3719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4492__B _3189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6760_ _1793_ _1795_ vssd1 vssd1 vccd1 vccd1 _1823_ sky130_fd_sc_hd__xor2_1
XFILLER_23_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5711_ _3864_ _0619_ _0607_ _0112_ vssd1 vssd1 vccd1 vccd1 _0689_ sky130_fd_sc_hd__a211o_1
XFILLER_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6691_ _1724_ _1730_ vssd1 vssd1 vccd1 vccd1 _1747_ sky130_fd_sc_hd__nand2_1
XFILLER_31_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5642_ _3900_ _0609_ _0614_ _3864_ _3718_ vssd1 vssd1 vccd1 vccd1 _0615_ sky130_fd_sc_hd__o2111a_1
X_8430_ counter\[0\] _3242_ _3641_ vssd1 vssd1 vccd1 vccd1 _3642_ sky130_fd_sc_hd__o21ai_1
X_5573_ _4138_ _4125_ _4131_ vssd1 vssd1 vccd1 vccd1 _0546_ sky130_fd_sc_hd__and3_1
X_8361_ _3166_ _3416_ _3529_ vssd1 vssd1 vccd1 vccd1 _3572_ sky130_fd_sc_hd__or3_1
XANTENNA__5109__A _4232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4524_ _2969_ _3446_ _3530_ vssd1 vssd1 vccd1 vccd1 _3541_ sky130_fd_sc_hd__nand3_1
XANTENNA__8477__A1 _1253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7312_ _2333_ vssd1 vssd1 vccd1 vccd1 _2431_ sky130_fd_sc_hd__buf_2
XFILLER_116_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8292_ _1319_ _3485_ vssd1 vssd1 vccd1 vccd1 _3499_ sky130_fd_sc_hd__and2_1
XFILLER_116_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4455_ _2705_ _2782_ vssd1 vssd1 vccd1 vccd1 _2793_ sky130_fd_sc_hd__nand2_1
X_7243_ _0430_ _0425_ vssd1 vssd1 vccd1 vccd1 _2355_ sky130_fd_sc_hd__nand2_1
X_4386_ posit_add.in2\[1\] _2023_ vssd1 vssd1 vccd1 vccd1 _2034_ sky130_fd_sc_hd__xor2_4
X_7174_ _1637_ _2278_ vssd1 vssd1 vccd1 vccd1 _2279_ sky130_fd_sc_hd__nor2_1
XFILLER_112_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6125_ _1127_ vssd1 vssd1 vccd1 vccd1 _1128_ sky130_fd_sc_hd__buf_2
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6056_ _0960_ _1055_ vssd1 vssd1 vccd1 vccd1 _1056_ sky130_fd_sc_hd__nor2_1
XFILLER_105_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5007_ _4160_ _4161_ vssd1 vssd1 vccd1 vccd1 _4162_ sky130_fd_sc_hd__and2_1
XFILLER_73_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6958_ _1987_ _1989_ vssd1 vssd1 vccd1 vccd1 _2041_ sky130_fd_sc_hd__xor2_1
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5909_ _0898_ _0899_ _0894_ vssd1 vssd1 vccd1 vccd1 _0901_ sky130_fd_sc_hd__a21o_1
X_6889_ _1953_ _1954_ _1963_ _1964_ vssd1 vssd1 vccd1 vccd1 _1965_ sky130_fd_sc_hd__a31o_1
XFILLER_22_551 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8559_ clknet_3_0__leaf_clk _0045_ vssd1 vssd1 vccd1 vccd1 posit_add.in1\[2\] sky130_fd_sc_hd__dfxtp_2
XFILLER_108_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5019__A posit_add.in1\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_698 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5757__A2 _3815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4965__B1 _3804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7409__A _2534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7930_ _3109_ _3087_ _3044_ vssd1 vssd1 vccd1 vccd1 _3110_ sky130_fd_sc_hd__mux2_1
X_7861_ _2971_ vssd1 vssd1 vccd1 vccd1 _3034_ sky130_fd_sc_hd__buf_2
XFILLER_36_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6812_ _1845_ _1879_ vssd1 vssd1 vccd1 vccd1 _1881_ sky130_fd_sc_hd__xnor2_1
XFILLER_63_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7792_ _2942_ _2957_ vssd1 vssd1 vccd1 vccd1 _2959_ sky130_fd_sc_hd__nand2_1
XFILLER_36_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6743_ _1789_ _1790_ vssd1 vssd1 vccd1 vccd1 _1805_ sky130_fd_sc_hd__xor2_1
XANTENNA__6223__A _1097_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6674_ _1540_ _1728_ vssd1 vssd1 vccd1 vccd1 _1729_ sky130_fd_sc_hd__xnor2_1
X_5625_ _1330_ _0594_ _0597_ vssd1 vssd1 vccd1 vccd1 _0598_ sky130_fd_sc_hd__a21oi_1
X_8413_ _3225_ _4250_ vssd1 vssd1 vccd1 vccd1 _3627_ sky130_fd_sc_hd__nand2_1
XFILLER_3_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8344_ _3259_ _3337_ vssd1 vssd1 vccd1 vccd1 _3554_ sky130_fd_sc_hd__nor2_1
X_5556_ _0486_ _0505_ _0470_ vssd1 vssd1 vccd1 vccd1 _0529_ sky130_fd_sc_hd__mux2_1
X_4507_ _3328_ _3035_ vssd1 vssd1 vccd1 vccd1 _3360_ sky130_fd_sc_hd__xnor2_4
X_8275_ _3421_ _3415_ _3452_ _1308_ vssd1 vssd1 vccd1 vccd1 _3481_ sky130_fd_sc_hd__o31a_2
X_5487_ _0457_ _0459_ vssd1 vssd1 vccd1 vccd1 _0460_ sky130_fd_sc_hd__xnor2_1
XFILLER_117_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4438_ posit_add.in1\[14\] _2595_ vssd1 vssd1 vccd1 vccd1 _2606_ sky130_fd_sc_hd__xnor2_4
X_7226_ _0385_ _2335_ vssd1 vssd1 vccd1 vccd1 _2336_ sky130_fd_sc_hd__xnor2_1
XFILLER_98_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6893__A _1665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4369_ _1275_ _1352_ vssd1 vssd1 vccd1 vccd1 _1847_ sky130_fd_sc_hd__nand2_1
X_7157_ _2258_ _2259_ vssd1 vssd1 vccd1 vccd1 _2260_ sky130_fd_sc_hd__nor2_1
X_6108_ _1103_ _1109_ vssd1 vssd1 vccd1 vccd1 _1110_ sky130_fd_sc_hd__and2b_1
XFILLER_100_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7088_ _2163_ _2167_ vssd1 vssd1 vccd1 vccd1 _2184_ sky130_fd_sc_hd__xor2_1
XFILLER_86_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6039_ _0706_ _0993_ _0998_ _1005_ vssd1 vssd1 vccd1 vccd1 _1038_ sky130_fd_sc_hd__a22oi_1
XFILLER_100_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6787__B _4126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6624__B1 _1420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5212__A _4222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4473__D _2980_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6978__A _1454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5410_ _3757_ _3758_ _3690_ vssd1 vssd1 vccd1 vccd1 _0383_ sky130_fd_sc_hd__a21o_1
X_6390_ _0218_ _1414_ vssd1 vssd1 vccd1 vccd1 _1416_ sky130_fd_sc_hd__nand2_2
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5341_ _4199_ _4201_ _4203_ vssd1 vssd1 vccd1 vccd1 _0314_ sky130_fd_sc_hd__o21ba_1
X_8060_ _2597_ _3250_ _2486_ vssd1 vssd1 vccd1 vccd1 _3251_ sky130_fd_sc_hd__mux2_1
X_7011_ _2090_ _2098_ vssd1 vssd1 vccd1 vccd1 _2099_ sky130_fd_sc_hd__xor2_1
XANTENNA__5666__B2 _3892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5272_ _0243_ _0244_ vssd1 vssd1 vccd1 vccd1 _0245_ sky130_fd_sc_hd__and2b_1
XFILLER_114_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7407__A2 _2524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7913_ _3038_ _3054_ _3091_ vssd1 vssd1 vccd1 vccd1 _3092_ sky130_fd_sc_hd__a21oi_1
XFILLER_102_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7844_ _3012_ _3015_ _2993_ vssd1 vssd1 vccd1 vccd1 _3016_ sky130_fd_sc_hd__o21ai_1
XFILLER_51_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7775_ _2868_ _2935_ _2917_ vssd1 vssd1 vccd1 vccd1 _2940_ sky130_fd_sc_hd__a21oi_1
XFILLER_24_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6726_ _1677_ _1779_ _1780_ _1785_ vssd1 vssd1 vccd1 vccd1 _1786_ sky130_fd_sc_hd__a2bb2oi_2
XFILLER_51_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4987_ _4133_ _4117_ _4128_ _4136_ vssd1 vssd1 vccd1 vccd1 _4142_ sky130_fd_sc_hd__a31o_1
XFILLER_23_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6657_ _1706_ _1709_ vssd1 vssd1 vccd1 vccd1 _1710_ sky130_fd_sc_hd__xor2_1
XANTENNA__7343__A1 _0147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6588_ _0080_ _1400_ _1631_ vssd1 vssd1 vccd1 vccd1 _1634_ sky130_fd_sc_hd__or3_1
X_5608_ _0521_ _0570_ _0573_ _0580_ vssd1 vssd1 vccd1 vccd1 _0581_ sky130_fd_sc_hd__or4_1
XFILLER_117_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8327_ _3508_ _3535_ vssd1 vssd1 vccd1 vccd1 _3536_ sky130_fd_sc_hd__and2_1
XFILLER_3_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5539_ _0443_ _0510_ _0511_ vssd1 vssd1 vccd1 vccd1 _0512_ sky130_fd_sc_hd__o21ai_1
XANTENNA__6400__B _1354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8258_ _1319_ _3462_ vssd1 vssd1 vccd1 vccd1 _3463_ sky130_fd_sc_hd__nand2_1
X_8189_ _3023_ _3029_ vssd1 vssd1 vccd1 vccd1 _3389_ sky130_fd_sc_hd__nand2_1
X_7209_ _2292_ _2295_ _2314_ vssd1 vssd1 vccd1 vccd1 _2317_ sky130_fd_sc_hd__a21bo_1
XFILLER_59_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6798__A _3988_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6980__B _1538_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5890_ _0876_ _0879_ _0865_ _0864_ vssd1 vssd1 vccd1 vccd1 _0881_ sky130_fd_sc_hd__o211ai_1
XFILLER_93_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4910_ _4048_ _4064_ vssd1 vssd1 vccd1 vccd1 _4065_ sky130_fd_sc_hd__xnor2_1
XFILLER_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4841_ _3994_ _3995_ vssd1 vssd1 vccd1 vccd1 _3996_ sky130_fd_sc_hd__nand2_1
X_4772_ _3924_ _3702_ vssd1 vssd1 vccd1 vccd1 _3927_ sky130_fd_sc_hd__or2_1
X_7560_ _2676_ _2702_ vssd1 vssd1 vccd1 vccd1 _2703_ sky130_fd_sc_hd__nand2_1
X_6511_ _1544_ _1386_ _1547_ _1548_ vssd1 vssd1 vccd1 vccd1 _1549_ sky130_fd_sc_hd__a22oi_4
X_7491_ _2826_ _0402_ vssd1 vssd1 vccd1 vccd1 _2627_ sky130_fd_sc_hd__nor2_1
XANTENNA__6501__A _1537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6442_ _1399_ _1428_ vssd1 vssd1 vccd1 vccd1 _1474_ sky130_fd_sc_hd__nor2_1
XFILLER_115_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6220__B _1128_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6373_ _1375_ _1381_ _1371_ vssd1 vssd1 vccd1 vccd1 _1398_ sky130_fd_sc_hd__a21bo_1
X_8112_ _0535_ _0516_ _3306_ vssd1 vssd1 vccd1 vccd1 _3308_ sky130_fd_sc_hd__a21boi_1
XFILLER_114_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5324_ _0286_ _0295_ vssd1 vssd1 vccd1 vccd1 _0297_ sky130_fd_sc_hd__or2_1
X_5255_ _0215_ _0226_ vssd1 vssd1 vccd1 vccd1 _0228_ sky130_fd_sc_hd__and2_1
X_8043_ _3030_ vssd1 vssd1 vccd1 vccd1 _3234_ sky130_fd_sc_hd__buf_2
XANTENNA__7051__B _1676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5186_ _0157_ _0158_ vssd1 vssd1 vccd1 vccd1 _0159_ sky130_fd_sc_hd__and2_1
XFILLER_29_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8053__A2 _3224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5811__B2 _3866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5811__A1 _3901_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5787__A _3924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7827_ _2993_ _2995_ vssd1 vssd1 vccd1 vccd1 _2997_ sky130_fd_sc_hd__nand2_1
XFILLER_36_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7758_ _2849_ _2920_ vssd1 vssd1 vccd1 vccd1 _2921_ sky130_fd_sc_hd__xor2_2
X_6709_ _1765_ _1766_ vssd1 vssd1 vccd1 vccd1 _1767_ sky130_fd_sc_hd__and2_1
X_7689_ _2761_ _2822_ vssd1 vssd1 vccd1 vccd1 _2845_ sky130_fd_sc_hd__or2b_1
XFILLER_20_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7226__B _2335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5027__A _3827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4776__A _3719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5040_ _4009_ _3860_ _3888_ vssd1 vssd1 vccd1 vccd1 _4195_ sky130_fd_sc_hd__and3_1
XFILLER_69_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6991__A _1711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6991_ _1711_ _1950_ vssd1 vssd1 vccd1 vccd1 _2077_ sky130_fd_sc_hd__and2_1
XFILLER_65_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5942_ _0935_ _0926_ vssd1 vssd1 vccd1 vccd1 _0936_ sky130_fd_sc_hd__xnor2_1
XFILLER_93_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5873_ _0844_ _0845_ _0846_ vssd1 vssd1 vccd1 vccd1 _0864_ sky130_fd_sc_hd__or3_1
XFILLER_21_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4824_ _3967_ _3977_ vssd1 vssd1 vccd1 vccd1 _3979_ sky130_fd_sc_hd__and2b_1
XFILLER_21_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7612_ _2758_ _2759_ vssd1 vssd1 vccd1 vccd1 _2761_ sky130_fd_sc_hd__and2_1
XFILLER_33_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4755_ _3906_ _3909_ vssd1 vssd1 vccd1 vccd1 _3910_ sky130_fd_sc_hd__xor2_1
XANTENNA__5021__A2 _3988_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7543_ _2681_ _2684_ vssd1 vssd1 vccd1 vccd1 _2685_ sky130_fd_sc_hd__nor2_1
X_4686_ _3827_ _3739_ _3840_ _3828_ vssd1 vssd1 vccd1 vccd1 _3841_ sky130_fd_sc_hd__o22a_1
X_7474_ _2520_ _2569_ _2608_ vssd1 vssd1 vccd1 vccd1 _2609_ sky130_fd_sc_hd__a21oi_1
XFILLER_119_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6425_ _1445_ _1454_ vssd1 vssd1 vccd1 vccd1 _1455_ sky130_fd_sc_hd__or2_1
XANTENNA__6885__B _0548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6356_ _1349_ vssd1 vssd1 vccd1 vccd1 _1379_ sky130_fd_sc_hd__inv_2
XFILLER_115_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5307_ _0275_ _0277_ _0279_ vssd1 vssd1 vccd1 vccd1 _0280_ sky130_fd_sc_hd__a21oi_1
X_6287_ _1221_ _1224_ _1225_ vssd1 vssd1 vccd1 vccd1 _1303_ sky130_fd_sc_hd__a21o_1
XFILLER_102_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8026_ _0451_ _0512_ _0515_ vssd1 vssd1 vccd1 vccd1 _3215_ sky130_fd_sc_hd__mux2_1
XFILLER_75_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5238_ _3828_ _4037_ _4182_ _0210_ vssd1 vssd1 vccd1 vccd1 _0211_ sky130_fd_sc_hd__or4b_1
XANTENNA__4835__A2 _3988_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5169_ _0114_ _0115_ vssd1 vssd1 vccd1 vccd1 _0142_ sky130_fd_sc_hd__xnor2_1
XFILLER_56_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5796__B1 _0779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4540_ _1990_ _3659_ _3671_ _3678_ vssd1 vssd1 vccd1 vccd1 _3684_ sky130_fd_sc_hd__a31o_1
X_4471_ posit_add.in1\[0\] vssd1 vssd1 vccd1 vccd1 _2969_ sky130_fd_sc_hd__clkbuf_4
XFILLER_7_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6210_ _1211_ _1216_ _1217_ vssd1 vssd1 vccd1 vccd1 _1218_ sky130_fd_sc_hd__a21o_1
X_7190_ _2269_ _2294_ vssd1 vssd1 vccd1 vccd1 _2296_ sky130_fd_sc_hd__or2_1
XFILLER_112_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6141_ _1015_ _1031_ vssd1 vssd1 vccd1 vccd1 _1145_ sky130_fd_sc_hd__nand2_1
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6072_ _1057_ _1060_ _1066_ vssd1 vssd1 vccd1 vccd1 _1073_ sky130_fd_sc_hd__and3_1
XFILLER_112_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5023_ _4173_ _4177_ vssd1 vssd1 vccd1 vccd1 _4178_ sky130_fd_sc_hd__xnor2_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6974_ _2054_ _2058_ vssd1 vssd1 vccd1 vccd1 _2059_ sky130_fd_sc_hd__nand2_1
XFILLER_26_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5925_ _0915_ _0916_ _0912_ vssd1 vssd1 vccd1 vccd1 _0918_ sky130_fd_sc_hd__a21o_1
XFILLER_81_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5856_ _3770_ _0828_ vssd1 vssd1 vccd1 vccd1 _0846_ sky130_fd_sc_hd__xnor2_1
X_4807_ _3956_ _3957_ _3961_ vssd1 vssd1 vccd1 vccd1 _3962_ sky130_fd_sc_hd__o21a_1
XFILLER_21_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5787_ _3924_ _0660_ vssd1 vssd1 vccd1 vccd1 _0771_ sky130_fd_sc_hd__or2_1
X_8575_ clknet_3_6__leaf_clk _0061_ vssd1 vssd1 vccd1 vccd1 posit_add.in2\[2\] sky130_fd_sc_hd__dfxtp_2
XFILLER_119_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4738_ _3892_ vssd1 vssd1 vccd1 vccd1 _3893_ sky130_fd_sc_hd__clkbuf_4
X_7526_ _2662_ _2665_ vssd1 vssd1 vccd1 vccd1 _2666_ sky130_fd_sc_hd__nand2_1
XFILLER_119_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4669_ _3821_ _3823_ vssd1 vssd1 vccd1 vccd1 _3824_ sky130_fd_sc_hd__nand2_1
X_7457_ _2381_ _2454_ _2589_ _2493_ vssd1 vssd1 vccd1 vccd1 _2590_ sky130_fd_sc_hd__o211a_1
X_6408_ _1395_ vssd1 vssd1 vccd1 vccd1 _1436_ sky130_fd_sc_hd__inv_2
XFILLER_1_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7388_ _2481_ _2483_ vssd1 vssd1 vccd1 vccd1 _2514_ sky130_fd_sc_hd__nor2_4
XFILLER_103_532 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6339_ _0627_ _1338_ vssd1 vssd1 vccd1 vccd1 _1360_ sky130_fd_sc_hd__nand2_1
XFILLER_88_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4269__A0 in_reg\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8009_ _1220_ _3196_ vssd1 vssd1 vccd1 vccd1 _0020_ sky130_fd_sc_hd__nor2_1
XFILLER_91_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4582__C _3729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8266__B1_N _1177_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4265__S _0712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5710_ _3814_ _0604_ _3762_ vssd1 vssd1 vccd1 vccd1 _0688_ sky130_fd_sc_hd__a21oi_1
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6690_ _1734_ _1745_ vssd1 vssd1 vccd1 vccd1 _1746_ sky130_fd_sc_hd__or2_1
X_5641_ _4043_ _3898_ _3899_ vssd1 vssd1 vccd1 vccd1 _0614_ sky130_fd_sc_hd__or3_2
X_8360_ _3569_ _3570_ vssd1 vssd1 vccd1 vccd1 _3571_ sky130_fd_sc_hd__nor2_1
X_5572_ _0541_ _0544_ _0515_ vssd1 vssd1 vccd1 vccd1 _0545_ sky130_fd_sc_hd__o21ba_1
X_8291_ _1220_ _3497_ vssd1 vssd1 vccd1 vccd1 _0029_ sky130_fd_sc_hd__nor2_1
X_4523_ _3079_ _3296_ _3046_ vssd1 vssd1 vccd1 vccd1 _3530_ sky130_fd_sc_hd__a21oi_4
X_7311_ _1899_ _2428_ vssd1 vssd1 vccd1 vccd1 _2429_ sky130_fd_sc_hd__nand2_1
X_7242_ _0348_ _2351_ _2352_ vssd1 vssd1 vccd1 vccd1 _2354_ sky130_fd_sc_hd__o21a_2
X_4454_ _2738_ _2771_ vssd1 vssd1 vccd1 vccd1 _2782_ sky130_fd_sc_hd__nor2_1
XFILLER_98_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4385_ posit_add.in2\[0\] _1275_ vssd1 vssd1 vccd1 vccd1 _2023_ sky130_fd_sc_hd__nand2_2
X_7173_ _4251_ _2273_ _2275_ _2277_ vssd1 vssd1 vccd1 vccd1 _2278_ sky130_fd_sc_hd__a211o_1
XFILLER_112_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6124_ _1091_ _1126_ vssd1 vssd1 vccd1 vccd1 _1127_ sky130_fd_sc_hd__and2_1
XFILLER_105_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6055_ _0943_ _0944_ _0959_ vssd1 vssd1 vccd1 vccd1 _1055_ sky130_fd_sc_hd__a21oi_1
XANTENNA__4964__A _3771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5006_ _3802_ _3883_ _4159_ vssd1 vssd1 vccd1 vccd1 _4161_ sky130_fd_sc_hd__a21o_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5626__C_N cmd\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6957_ _2030_ _2038_ _2039_ vssd1 vssd1 vccd1 vccd1 _2040_ sky130_fd_sc_hd__a21o_1
XFILLER_81_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5795__A _4016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5908_ _0894_ _0898_ _0899_ vssd1 vssd1 vccd1 vccd1 _0900_ sky130_fd_sc_hd__nand3_1
X_6888_ _1961_ _1962_ vssd1 vssd1 vccd1 vccd1 _1964_ sky130_fd_sc_hd__and2b_1
X_5839_ _0826_ _0754_ vssd1 vssd1 vccd1 vccd1 _0827_ sky130_fd_sc_hd__and2b_1
XFILLER_10_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_563 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8558_ clknet_3_6__leaf_clk _0044_ vssd1 vssd1 vccd1 vccd1 posit_add.in1\[1\] sky130_fd_sc_hd__dfxtp_4
XFILLER_108_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7509_ _3068_ _1451_ _1539_ _2624_ _2646_ vssd1 vssd1 vccd1 vccd1 _2647_ sky130_fd_sc_hd__a221o_1
XFILLER_108_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8489_ _3682_ vssd1 vssd1 vccd1 vccd1 _0062_ sky130_fd_sc_hd__clkbuf_1
XFILLER_107_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7428__B1 _2557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4965__A1 _3832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4965__B2 _3893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7131__A2 _1676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7860_ _3032_ vssd1 vssd1 vccd1 vccd1 _3033_ sky130_fd_sc_hd__inv_2
X_6811_ _1852_ _1854_ vssd1 vssd1 vccd1 vccd1 _1879_ sky130_fd_sc_hd__xor2_1
XFILLER_36_666 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7791_ _2673_ _2941_ vssd1 vssd1 vccd1 vccd1 _2957_ sky130_fd_sc_hd__nand2_1
X_6742_ _1667_ _1673_ vssd1 vssd1 vccd1 vccd1 _1804_ sky130_fd_sc_hd__xnor2_1
XFILLER_51_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6223__B _1164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6673_ _4157_ _1533_ vssd1 vssd1 vccd1 vccd1 _1728_ sky130_fd_sc_hd__xor2_1
XANTENNA__5905__B1 _0706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5624_ _0595_ _0596_ vssd1 vssd1 vccd1 vccd1 _0597_ sky130_fd_sc_hd__and2_1
X_8412_ cmd\[7\] cmd\[6\] vssd1 vssd1 vccd1 vccd1 _3626_ sky130_fd_sc_hd__nand2_1
XFILLER_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8343_ _3518_ _3542_ vssd1 vssd1 vccd1 vccd1 _3553_ sky130_fd_sc_hd__or2_1
X_5555_ _0524_ _0527_ _0494_ vssd1 vssd1 vccd1 vccd1 _0528_ sky130_fd_sc_hd__mux2_1
X_4506_ _2738_ _3275_ _3285_ _3112_ vssd1 vssd1 vccd1 vccd1 _3349_ sky130_fd_sc_hd__o31a_4
X_8274_ _3227_ _3460_ _3478_ _3190_ vssd1 vssd1 vccd1 vccd1 _3480_ sky130_fd_sc_hd__o31a_1
XFILLER_2_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5486_ _0440_ _0458_ vssd1 vssd1 vccd1 vccd1 _0459_ sky130_fd_sc_hd__or2_1
X_4437_ posit_add.in1\[11\] posit_add.in1\[10\] _2573_ _2584_ _1242_ vssd1 vssd1 vccd1
+ vccd1 _2595_ sky130_fd_sc_hd__o41a_2
X_7225_ _2334_ vssd1 vssd1 vccd1 vccd1 _2335_ sky130_fd_sc_hd__clkbuf_4
X_7156_ _2003_ _1948_ vssd1 vssd1 vccd1 vccd1 _2259_ sky130_fd_sc_hd__xnor2_4
XFILLER_113_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6107_ _0996_ _0997_ _1102_ _1097_ vssd1 vssd1 vccd1 vccd1 _1109_ sky130_fd_sc_hd__a22o_1
XFILLER_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4368_ posit_add.in2\[3\] _1825_ vssd1 vssd1 vccd1 vccd1 _1836_ sky130_fd_sc_hd__xnor2_4
XFILLER_76_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7087_ _2170_ _2173_ _2172_ vssd1 vssd1 vccd1 vccd1 _2183_ sky130_fd_sc_hd__a21o_1
X_4299_ _1072_ vssd1 vssd1 vccd1 vccd1 _0014_ sky130_fd_sc_hd__clkbuf_1
XFILLER_58_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6038_ _1000_ _1036_ vssd1 vssd1 vccd1 vccd1 _1037_ sky130_fd_sc_hd__nor2_1
XFILLER_86_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8386__A1 _2621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7989_ _3150_ vssd1 vssd1 vccd1 vccd1 _3175_ sky130_fd_sc_hd__clkinv_2
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4947__A1 _3793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4869__A _3719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8076__A _0600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5212__B _3883_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6978__B _1718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5340_ _0311_ _0312_ vssd1 vssd1 vccd1 vccd1 _0313_ sky130_fd_sc_hd__nor2_1
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6994__A _4217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5271_ _0229_ _0234_ _0227_ vssd1 vssd1 vccd1 vccd1 _0244_ sky130_fd_sc_hd__a21o_1
X_7010_ _2058_ _2091_ _2097_ vssd1 vssd1 vccd1 vccd1 _2098_ sky130_fd_sc_hd__nand3_2
XANTENNA__5666__A2 _3878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7912_ _3038_ _3089_ vssd1 vssd1 vccd1 vccd1 _3091_ sky130_fd_sc_hd__and2b_1
XFILLER_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7843_ _3001_ vssd1 vssd1 vccd1 vccd1 _3015_ sky130_fd_sc_hd__inv_2
XFILLER_36_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4986_ _4097_ _4112_ vssd1 vssd1 vccd1 vccd1 _4141_ sky130_fd_sc_hd__xnor2_1
XFILLER_24_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7774_ _2665_ _2938_ vssd1 vssd1 vccd1 vccd1 _2939_ sky130_fd_sc_hd__nor2_1
X_6725_ _1783_ _1784_ vssd1 vssd1 vccd1 vccd1 _1785_ sky130_fd_sc_hd__xnor2_2
XANTENNA__5051__B1 _4033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6000__C1 _4016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6656_ _1707_ _1708_ vssd1 vssd1 vccd1 vccd1 _1709_ sky130_fd_sc_hd__xnor2_1
XANTENNA__4689__A _3828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6587_ _1598_ _1601_ vssd1 vssd1 vccd1 vccd1 _1633_ sky130_fd_sc_hd__or2_1
X_5607_ _0575_ _0576_ _0578_ _0579_ vssd1 vssd1 vccd1 vccd1 _0580_ sky130_fd_sc_hd__a22o_1
XFILLER_117_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7065__A _1454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8326_ _3437_ _3298_ _3438_ vssd1 vssd1 vccd1 vccd1 _3535_ sky130_fd_sc_hd__a21oi_1
X_5538_ _0440_ _0510_ vssd1 vssd1 vccd1 vccd1 _0511_ sky130_fd_sc_hd__nand2_1
XANTENNA__6400__C _4153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8257_ _3426_ _3433_ vssd1 vssd1 vccd1 vccd1 _3462_ sky130_fd_sc_hd__nand2_1
XFILLER_3_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7208_ _2008_ _2261_ _2268_ _2297_ _2315_ vssd1 vssd1 vccd1 vccd1 _2316_ sky130_fd_sc_hd__a311o_1
X_5469_ _0356_ _0363_ vssd1 vssd1 vccd1 vccd1 _0442_ sky130_fd_sc_hd__xor2_4
XFILLER_59_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8188_ _3329_ _3373_ vssd1 vssd1 vccd1 vccd1 _3388_ sky130_fd_sc_hd__and2b_1
X_7139_ _2197_ _2202_ _2182_ vssd1 vssd1 vccd1 vccd1 _2240_ sky130_fd_sc_hd__a21o_1
XFILLER_59_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_696 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6319__A _4210_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7270__A1 _0351_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4840_ _3992_ _3993_ vssd1 vssd1 vccd1 vccd1 _3995_ sky130_fd_sc_hd__or2_1
XFILLER_60_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4771_ _3925_ _3726_ vssd1 vssd1 vccd1 vccd1 _3926_ sky130_fd_sc_hd__nor2_1
X_6510_ _1400_ _1454_ vssd1 vssd1 vccd1 vccd1 _1548_ sky130_fd_sc_hd__nor2_1
XFILLER_60_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7490_ posit_add.in1\[7\] _2683_ vssd1 vssd1 vccd1 vccd1 _2626_ sky130_fd_sc_hd__xnor2_1
X_6441_ _1468_ _1471_ vssd1 vssd1 vccd1 vccd1 _1472_ sky130_fd_sc_hd__xnor2_1
X_6372_ _1394_ _1395_ vssd1 vssd1 vccd1 vccd1 _1397_ sky130_fd_sc_hd__or2_2
X_5323_ _0286_ _0295_ vssd1 vssd1 vccd1 vccd1 _0296_ sky130_fd_sc_hd__xnor2_1
X_8111_ _0451_ _0557_ vssd1 vssd1 vccd1 vccd1 _3306_ sky130_fd_sc_hd__nand2_1
X_5254_ _0215_ _0226_ vssd1 vssd1 vccd1 vccd1 _0227_ sky130_fd_sc_hd__nor2_1
X_8042_ _3151_ _3231_ _3021_ vssd1 vssd1 vccd1 vccd1 _3233_ sky130_fd_sc_hd__mux2_1
XANTENNA__6229__A _0706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5185_ _0154_ _0143_ vssd1 vssd1 vccd1 vccd1 _0158_ sky130_fd_sc_hd__or2b_1
XANTENNA__7051__C _1538_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5133__A _3925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7759__S _1308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8444__A net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5811__A2 _0795_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7826_ _2993_ _2995_ vssd1 vssd1 vccd1 vccd1 _2996_ sky130_fd_sc_hd__or2_1
XFILLER_24_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4969_ _4118_ _4123_ vssd1 vssd1 vccd1 vccd1 _4124_ sky130_fd_sc_hd__nor2_1
X_7757_ _1308_ _2874_ _2919_ vssd1 vssd1 vccd1 vccd1 _2920_ sky130_fd_sc_hd__a21oi_1
XFILLER_24_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6708_ _1762_ _1763_ _1764_ vssd1 vssd1 vccd1 vccd1 _1766_ sky130_fd_sc_hd__nand3_1
X_7688_ _2840_ _2839_ vssd1 vssd1 vccd1 vccd1 _2844_ sky130_fd_sc_hd__and2b_1
X_6639_ _1659_ _1674_ vssd1 vssd1 vccd1 vccd1 _1690_ sky130_fd_sc_hd__nor2_1
XFILLER_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5027__B _3816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8309_ _3259_ _3261_ vssd1 vssd1 vccd1 vccd1 _3517_ sky130_fd_sc_hd__or2_1
XFILLER_79_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_471 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4882__A _3750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7417__B _0548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4776__B _3930_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4264__C_N _0701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6991__B _1950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6990_ _2033_ _2042_ vssd1 vssd1 vccd1 vccd1 _2076_ sky130_fd_sc_hd__xor2_1
XFILLER_92_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5941_ _0923_ _0924_ vssd1 vssd1 vccd1 vccd1 _0935_ sky130_fd_sc_hd__nand2_1
XFILLER_93_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5872_ _3738_ _0860_ _0861_ vssd1 vssd1 vccd1 vccd1 _0863_ sky130_fd_sc_hd__o21ai_1
XFILLER_80_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4823_ _3967_ _3977_ vssd1 vssd1 vccd1 vccd1 _3978_ sky130_fd_sc_hd__xnor2_1
X_7611_ _3816_ _1384_ _2721_ vssd1 vssd1 vccd1 vccd1 _2759_ sky130_fd_sc_hd__mux2_1
XFILLER_21_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6512__A _4153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4754_ _3881_ _3907_ _3778_ _3908_ vssd1 vssd1 vccd1 vccd1 _3909_ sky130_fd_sc_hd__a31o_1
X_7542_ _0410_ _0420_ _2652_ vssd1 vssd1 vccd1 vccd1 _2684_ sky130_fd_sc_hd__mux2_1
XFILLER_119_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7473_ _2379_ _2448_ _2516_ vssd1 vssd1 vccd1 vccd1 _2608_ sky130_fd_sc_hd__and3_1
X_4685_ _3722_ _3835_ _3836_ _3837_ vssd1 vssd1 vccd1 vccd1 _3840_ sky130_fd_sc_hd__a31oi_4
XFILLER_108_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6424_ _3795_ vssd1 vssd1 vccd1 vccd1 _1454_ sky130_fd_sc_hd__clkbuf_4
XFILLER_115_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6355_ _1306_ _1310_ _1376_ _1377_ vssd1 vssd1 vccd1 vccd1 _1378_ sky130_fd_sc_hd__a211o_1
XFILLER_115_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6286_ _1277_ _1300_ _1301_ vssd1 vssd1 vccd1 vccd1 _1302_ sky130_fd_sc_hd__a21o_1
X_5306_ _0247_ _0278_ vssd1 vssd1 vccd1 vccd1 _0279_ sky130_fd_sc_hd__nand2_1
XANTENNA__7062__B _1456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5237_ _0165_ _0166_ vssd1 vssd1 vccd1 vccd1 _0210_ sky130_fd_sc_hd__xor2_1
X_8025_ _0594_ _0597_ vssd1 vssd1 vccd1 vccd1 _3214_ sky130_fd_sc_hd__or2_1
XFILLER_102_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5168_ _0125_ _0136_ _0140_ _4182_ vssd1 vssd1 vccd1 vccd1 _0141_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_56_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5099_ _4249_ _4253_ vssd1 vssd1 vccd1 vccd1 _4254_ sky130_fd_sc_hd__nand2_1
XFILLER_17_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7809_ _2956_ _2959_ vssd1 vssd1 vccd1 vccd1 _2977_ sky130_fd_sc_hd__and2_1
XFILLER_8_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5720__B2 _0698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4470_ _2914_ _2947_ vssd1 vssd1 vccd1 vccd1 _2958_ sky130_fd_sc_hd__or2_1
XFILLER_7_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4787__A _3739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6140_ _1002_ _1102_ vssd1 vssd1 vccd1 vccd1 _1144_ sky130_fd_sc_hd__xor2_1
XFILLER_98_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6071_ _0955_ _1061_ _1068_ _1070_ vssd1 vssd1 vccd1 vccd1 _1071_ sky130_fd_sc_hd__nor4_1
XFILLER_97_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4278__A1 in_reg\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5022_ _4175_ _4176_ vssd1 vssd1 vccd1 vccd1 _4177_ sky130_fd_sc_hd__nor2_1
XFILLER_66_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6507__A _1383_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6973_ _2055_ _2054_ _2057_ vssd1 vssd1 vccd1 vccd1 _2058_ sky130_fd_sc_hd__nand3_1
XFILLER_65_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5924_ _0912_ _0915_ _0916_ vssd1 vssd1 vccd1 vccd1 _0917_ sky130_fd_sc_hd__nand3_2
XFILLER_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5855_ _0710_ _0843_ _0842_ vssd1 vssd1 vccd1 vccd1 _0845_ sky130_fd_sc_hd__a21oi_1
XFILLER_21_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4806_ _3958_ _3960_ vssd1 vssd1 vccd1 vccd1 _3961_ sky130_fd_sc_hd__or2_1
XANTENNA__7338__A _2416_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5786_ _0764_ _0769_ vssd1 vssd1 vccd1 vccd1 _0770_ sky130_fd_sc_hd__xnor2_1
X_8574_ clknet_3_3__leaf_clk _0060_ vssd1 vssd1 vccd1 vccd1 posit_add.in2\[1\] sky130_fd_sc_hd__dfxtp_2
X_4737_ _3729_ _3733_ vssd1 vssd1 vccd1 vccd1 _3892_ sky130_fd_sc_hd__nor2_4
X_7525_ _2664_ vssd1 vssd1 vccd1 vccd1 _2665_ sky130_fd_sc_hd__inv_2
XFILLER_119_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4668_ _2760_ _3318_ _3822_ _3446_ vssd1 vssd1 vccd1 vccd1 _3823_ sky130_fd_sc_hd__a211o_1
X_7456_ _2425_ _2426_ _2427_ _2382_ vssd1 vssd1 vccd1 vccd1 _2589_ sky130_fd_sc_hd__a31o_1
X_6407_ _1404_ _1433_ _1434_ vssd1 vssd1 vccd1 vccd1 _1435_ sky130_fd_sc_hd__a21o_1
X_4599_ _3156_ _3751_ _3752_ _3753_ vssd1 vssd1 vccd1 vccd1 _3754_ sky130_fd_sc_hd__a31o_1
X_7387_ _2508_ _2512_ _2494_ vssd1 vssd1 vccd1 vccd1 _2513_ sky130_fd_sc_hd__mux2_1
XFILLER_115_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6338_ _0722_ _0993_ _0994_ _1097_ vssd1 vssd1 vccd1 vccd1 _1359_ sky130_fd_sc_hd__a22o_1
X_6269_ _1019_ _1128_ _1282_ vssd1 vssd1 vccd1 vccd1 _1283_ sky130_fd_sc_hd__a21o_1
XFILLER_95_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4269__A1 cmd\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8008_ out_reg\[0\] _1231_ _3194_ _3195_ vssd1 vssd1 vccd1 vccd1 _3196_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_29_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5769__A1 _0113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7682__S _2721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7997__A2 _3182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_675 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5640_ _0112_ _3864_ vssd1 vssd1 vccd1 vccd1 _0613_ sky130_fd_sc_hd__nor2_2
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5571_ _0543_ _0540_ _0470_ vssd1 vssd1 vccd1 vccd1 _0544_ sky130_fd_sc_hd__mux2_1
X_4522_ _2804_ _3002_ _3134_ vssd1 vssd1 vccd1 vccd1 _3520_ sky130_fd_sc_hd__a21oi_4
X_7310_ _1896_ _2418_ _2005_ vssd1 vssd1 vccd1 vccd1 _2428_ sky130_fd_sc_hd__o21ai_1
X_8290_ _3195_ _3495_ _3496_ vssd1 vssd1 vccd1 vccd1 _3497_ sky130_fd_sc_hd__o21ba_1
X_4453_ _2661_ _2760_ vssd1 vssd1 vccd1 vccd1 _2771_ sky130_fd_sc_hd__xnor2_1
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7241_ _0342_ _0349_ _0433_ vssd1 vssd1 vccd1 vccd1 _2352_ sky130_fd_sc_hd__a21o_1
XFILLER_98_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4384_ _2001_ vssd1 vssd1 vccd1 vccd1 _2012_ sky130_fd_sc_hd__clkbuf_2
X_7172_ _0080_ _1588_ _2274_ vssd1 vssd1 vccd1 vccd1 _2277_ sky130_fd_sc_hd__and3_1
X_6123_ _1090_ _1089_ _1078_ _1053_ vssd1 vssd1 vccd1 vccd1 _1126_ sky130_fd_sc_hd__o211ai_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6054_ _0971_ _0972_ vssd1 vssd1 vccd1 vccd1 _1054_ sky130_fd_sc_hd__nor2_1
XFILLER_112_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5005_ _3701_ _3795_ _4159_ vssd1 vssd1 vccd1 vccd1 _4160_ sky130_fd_sc_hd__or3b_1
XANTENNA__4964__B _3703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5141__A _0113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6956_ _2028_ _2029_ vssd1 vssd1 vccd1 vccd1 _2039_ sky130_fd_sc_hd__nor2_1
XFILLER_53_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5907_ _0896_ _0897_ _0895_ vssd1 vssd1 vccd1 vccd1 _0899_ sky130_fd_sc_hd__a21o_1
X_6887_ _1961_ _1962_ vssd1 vssd1 vccd1 vccd1 _1963_ sky130_fd_sc_hd__xnor2_1
XFILLER_22_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5838_ _0822_ _0824_ _0825_ vssd1 vssd1 vccd1 vccd1 _0826_ sky130_fd_sc_hd__a21boi_1
XFILLER_14_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5769_ _0113_ _0663_ _0751_ _0615_ _3924_ vssd1 vssd1 vccd1 vccd1 _0752_ sky130_fd_sc_hd__a221o_1
X_8557_ clknet_3_0__leaf_clk _0043_ vssd1 vssd1 vccd1 vccd1 posit_add.in1\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_108_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7508_ _3101_ _1484_ _2643_ _2644_ _2645_ vssd1 vssd1 vccd1 vccd1 _2646_ sky130_fd_sc_hd__o221a_1
XFILLER_108_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8488_ posit_add.in2\[3\] in_reg\[3\] _3677_ vssd1 vssd1 vccd1 vccd1 _3682_ sky130_fd_sc_hd__mux2_1
X_7439_ _2449_ _2541_ _2558_ _2569_ vssd1 vssd1 vccd1 vccd1 _2570_ sky130_fd_sc_hd__a211o_1
XFILLER_30_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4965__A2 _3868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6167__A1 _0795_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5390__A2 _1748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4653__A1 _1946_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4276__S _0830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6810_ _1876_ _1877_ vssd1 vssd1 vccd1 vccd1 _1878_ sky130_fd_sc_hd__nor2_1
XFILLER_51_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7587__S _2652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7790_ _2954_ _2955_ vssd1 vssd1 vccd1 vccd1 _2956_ sky130_fd_sc_hd__or2b_1
XFILLER_35_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6741_ _1675_ _1689_ vssd1 vssd1 vccd1 vccd1 _1802_ sky130_fd_sc_hd__xnor2_1
X_6672_ _1725_ _4157_ _1707_ _1708_ vssd1 vssd1 vccd1 vccd1 _1727_ sky130_fd_sc_hd__a22o_1
XANTENNA__5905__A1 _3878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5623_ _0593_ _0520_ _0538_ vssd1 vssd1 vccd1 vccd1 _0596_ sky130_fd_sc_hd__o21ai_1
X_8411_ cmd\[7\] cmd\[6\] _3623_ vssd1 vssd1 vccd1 vccd1 _3624_ sky130_fd_sc_hd__or3_1
XANTENNA__5905__B2 _3776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8342_ _3527_ _3551_ _0635_ vssd1 vssd1 vccd1 vccd1 _0031_ sky130_fd_sc_hd__a21oi_1
X_5554_ _0525_ _0526_ _0515_ vssd1 vssd1 vccd1 vccd1 _0527_ sky130_fd_sc_hd__mux2_1
XFILLER_105_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5136__A _3701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4505_ _3328_ _3068_ vssd1 vssd1 vccd1 vccd1 _3339_ sky130_fd_sc_hd__xnor2_4
X_8273_ _3227_ _3460_ _3478_ vssd1 vssd1 vccd1 vccd1 _3479_ sky130_fd_sc_hd__o21ai_1
X_5485_ _0446_ _0450_ _0449_ vssd1 vssd1 vccd1 vccd1 _0458_ sky130_fd_sc_hd__nor3_2
XFILLER_116_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4436_ posit_add.in1\[13\] posit_add.in1\[12\] vssd1 vssd1 vccd1 vccd1 _2584_ sky130_fd_sc_hd__or2_1
X_7224_ _2327_ _2330_ _2333_ vssd1 vssd1 vccd1 vccd1 _2334_ sky130_fd_sc_hd__and3_1
XFILLER_104_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4367_ posit_add.in2\[2\] _1770_ _1275_ vssd1 vssd1 vccd1 vccd1 _1825_ sky130_fd_sc_hd__o21a_2
X_7155_ _2000_ _2257_ vssd1 vssd1 vccd1 vccd1 _2258_ sky130_fd_sc_hd__or2_2
X_6106_ _1015_ _1029_ vssd1 vssd1 vccd1 vccd1 _1108_ sky130_fd_sc_hd__xnor2_1
XFILLER_98_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7086_ _2176_ _2178_ vssd1 vssd1 vccd1 vccd1 _2182_ sky130_fd_sc_hd__xor2_1
X_4298_ in_reg\[10\] in_reg\[11\] _0819_ vssd1 vssd1 vccd1 vccd1 _1072_ sky130_fd_sc_hd__mux2_1
XFILLER_86_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6037_ _1026_ _1034_ vssd1 vssd1 vccd1 vccd1 _1036_ sky130_fd_sc_hd__xnor2_1
XFILLER_86_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7988_ _3147_ vssd1 vssd1 vccd1 vccd1 _3174_ sky130_fd_sc_hd__clkinv_2
XFILLER_14_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6939_ _1414_ _1531_ vssd1 vssd1 vccd1 vccd1 _2020_ sky130_fd_sc_hd__nand2_1
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4869__B _3795_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6321__A1 _1097_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7900__A_N _2954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5270_ _0241_ _0242_ vssd1 vssd1 vccd1 vccd1 _0243_ sky130_fd_sc_hd__or2_1
XFILLER_99_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7911_ _3088_ _3067_ _3044_ vssd1 vssd1 vccd1 vccd1 _3089_ sky130_fd_sc_hd__mux2_1
XFILLER_83_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6515__A _1428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7842_ _2998_ _3006_ _3012_ vssd1 vssd1 vccd1 vccd1 _3014_ sky130_fd_sc_hd__or3b_1
XFILLER_63_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7773_ _2654_ _2937_ vssd1 vssd1 vccd1 vccd1 _2938_ sky130_fd_sc_hd__or2_1
X_4985_ _4139_ vssd1 vssd1 vccd1 vccd1 _4140_ sky130_fd_sc_hd__inv_2
X_6724_ _1383_ _3703_ vssd1 vssd1 vccd1 vccd1 _1784_ sky130_fd_sc_hd__or2_1
XFILLER_51_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6655_ _0080_ _1538_ vssd1 vssd1 vccd1 vccd1 _1708_ sky130_fd_sc_hd__nor2_1
XANTENNA__4689__B _3750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6586_ _1465_ _1631_ vssd1 vssd1 vccd1 vccd1 _1632_ sky130_fd_sc_hd__or2_1
X_5606_ _0535_ _0481_ _0534_ _0562_ vssd1 vssd1 vccd1 vccd1 _0579_ sky130_fd_sc_hd__or4_1
X_8325_ _3481_ _3531_ _3532_ _3533_ _3212_ vssd1 vssd1 vccd1 vccd1 _3534_ sky130_fd_sc_hd__o311a_1
X_5537_ _0470_ vssd1 vssd1 vccd1 vccd1 _0510_ sky130_fd_sc_hd__buf_2
X_8256_ _3458_ _3459_ _3303_ vssd1 vssd1 vccd1 vccd1 _3461_ sky130_fd_sc_hd__a21o_1
XFILLER_105_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5468_ _0398_ _0440_ vssd1 vssd1 vccd1 vccd1 _0441_ sky130_fd_sc_hd__xnor2_1
X_7207_ _2292_ _2314_ vssd1 vssd1 vccd1 vccd1 _2315_ sky130_fd_sc_hd__xor2_1
XFILLER_99_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7081__A _3986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4419_ _2012_ _2276_ _2287_ _1550_ vssd1 vssd1 vccd1 vccd1 _2397_ sky130_fd_sc_hd__a211o_1
X_5399_ _3101_ _3446_ _3145_ vssd1 vssd1 vccd1 vccd1 _0372_ sky130_fd_sc_hd__o21a_1
X_8187_ _3382_ _3386_ vssd1 vssd1 vccd1 vccd1 _3387_ sky130_fd_sc_hd__xor2_1
X_7138_ _2220_ _2238_ _2218_ vssd1 vssd1 vccd1 vccd1 _2239_ sky130_fd_sc_hd__a21o_1
X_7069_ _2161_ _2162_ vssd1 vssd1 vccd1 vccd1 _2163_ sky130_fd_sc_hd__nand2_1
XFILLER_100_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6319__B _0702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6335__A _1353_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4770_ _3924_ vssd1 vssd1 vccd1 vccd1 _3925_ sky130_fd_sc_hd__clkbuf_4
XFILLER_14_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6440_ _1469_ _1470_ vssd1 vssd1 vccd1 vccd1 _1471_ sky130_fd_sc_hd__and2b_1
X_6371_ _1365_ _1368_ _1393_ vssd1 vssd1 vccd1 vccd1 _1395_ sky130_fd_sc_hd__a21oi_1
X_5322_ _0291_ _0294_ vssd1 vssd1 vccd1 vccd1 _0295_ sky130_fd_sc_hd__and2_1
X_8110_ _3257_ _3267_ vssd1 vssd1 vccd1 vccd1 _3305_ sky130_fd_sc_hd__nand2_1
XFILLER_102_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5253_ _0179_ _0189_ vssd1 vssd1 vccd1 vccd1 _0226_ sky130_fd_sc_hd__xnor2_1
X_8041_ _3230_ vssd1 vssd1 vccd1 vccd1 _3231_ sky130_fd_sc_hd__clkinv_2
XANTENNA__7613__B _2702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5184_ _0138_ _0142_ vssd1 vssd1 vccd1 vccd1 _0157_ sky130_fd_sc_hd__or2b_1
XANTENNA__5414__A _0385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5133__B _3615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7825_ _2982_ _2994_ vssd1 vssd1 vccd1 vccd1 _2995_ sky130_fd_sc_hd__nor2_1
XFILLER_51_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6899__B _4126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4968_ _3845_ _3726_ _4119_ _4122_ vssd1 vssd1 vccd1 vccd1 _4123_ sky130_fd_sc_hd__or4b_1
XFILLER_11_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7756_ _1308_ _2814_ vssd1 vssd1 vccd1 vccd1 _2919_ sky130_fd_sc_hd__nor2_1
X_6707_ _1762_ _1763_ _1764_ vssd1 vssd1 vccd1 vccd1 _1765_ sky130_fd_sc_hd__a21o_1
X_4899_ _3878_ _3907_ _3789_ vssd1 vssd1 vccd1 vccd1 _4054_ sky130_fd_sc_hd__and3_1
XFILLER_11_139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7687_ _4250_ _0082_ _2710_ vssd1 vssd1 vccd1 vccd1 _2843_ sky130_fd_sc_hd__a21bo_1
XANTENNA__7076__A _1676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6638_ _1681_ _1688_ vssd1 vssd1 vccd1 vccd1 _1689_ sky130_fd_sc_hd__xnor2_1
XFILLER_106_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6569_ _1609_ _1611_ vssd1 vssd1 vccd1 vccd1 _1613_ sky130_fd_sc_hd__nand2_1
X_8308_ _3465_ _3490_ vssd1 vssd1 vccd1 vccd1 _3516_ sky130_fd_sc_hd__and2b_1
XFILLER_3_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8239_ _3182_ _3396_ _3442_ vssd1 vssd1 vccd1 vccd1 _3443_ sky130_fd_sc_hd__a21oi_1
XFILLER_87_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6065__A _3892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5940_ _0905_ _0930_ _0933_ vssd1 vssd1 vccd1 vccd1 _0934_ sky130_fd_sc_hd__o21bai_1
XFILLER_92_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6451__B1 _1414_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4284__S _0830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5871_ _0858_ _0859_ vssd1 vssd1 vccd1 vccd1 _0861_ sky130_fd_sc_hd__nand2_1
XANTENNA__5006__A1 _3802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7610_ _2743_ _2757_ vssd1 vssd1 vccd1 vccd1 _2758_ sky130_fd_sc_hd__nand2_1
X_4822_ _3968_ _3975_ _3976_ vssd1 vssd1 vccd1 vccd1 _3977_ sky130_fd_sc_hd__o21ai_1
XFILLER_21_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6512__B _1414_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4753_ _3773_ _3777_ vssd1 vssd1 vccd1 vccd1 _3908_ sky130_fd_sc_hd__and2_1
X_7541_ _2678_ _2680_ _2681_ vssd1 vssd1 vccd1 vccd1 _2682_ sky130_fd_sc_hd__o21ba_1
X_7472_ _2521_ _2571_ _2575_ _2605_ vssd1 vssd1 vccd1 vccd1 _2607_ sky130_fd_sc_hd__or4_1
X_4684_ _3832_ _3838_ vssd1 vssd1 vccd1 vccd1 _3839_ sky130_fd_sc_hd__nand2_1
X_6423_ _1450_ _1452_ vssd1 vssd1 vccd1 vccd1 _1453_ sky130_fd_sc_hd__nor2_1
XANTENNA__4517__B1 _2903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6354_ _1351_ _1335_ vssd1 vssd1 vccd1 vccd1 _1377_ sky130_fd_sc_hd__or2_1
XFILLER_115_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6285_ _1235_ _1254_ vssd1 vssd1 vccd1 vccd1 _1301_ sky130_fd_sc_hd__xnor2_1
X_5305_ _0246_ _0241_ _0245_ vssd1 vssd1 vccd1 vccd1 _0278_ sky130_fd_sc_hd__or3_1
XFILLER_115_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5236_ _0208_ vssd1 vssd1 vccd1 vccd1 _0209_ sky130_fd_sc_hd__inv_2
X_8024_ _3202_ _3208_ _3209_ _3212_ vssd1 vssd1 vccd1 vccd1 _3213_ sky130_fd_sc_hd__o211a_1
XFILLER_69_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5167_ _0138_ _0139_ vssd1 vssd1 vccd1 vccd1 _0140_ sky130_fd_sc_hd__nand2_1
XFILLER_56_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5098_ _4251_ _4252_ vssd1 vssd1 vccd1 vccd1 _4253_ sky130_fd_sc_hd__xnor2_1
XFILLER_29_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6745__A1 _1428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7808_ _2961_ _2972_ _2974_ _2975_ vssd1 vssd1 vccd1 vccd1 _2976_ sky130_fd_sc_hd__o22a_1
XFILLER_40_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7739_ _2833_ _2885_ _1297_ vssd1 vssd1 vccd1 vccd1 _2900_ sky130_fd_sc_hd__mux2_1
XFILLER_116_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4787__B _3750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6070_ _1065_ _1069_ vssd1 vssd1 vccd1 vccd1 _1070_ sky130_fd_sc_hd__or2_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5021_ _3793_ _3988_ _3989_ _3771_ vssd1 vssd1 vccd1 vccd1 _4176_ sky130_fd_sc_hd__o22a_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6507__B _1401_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6972_ _2017_ _2049_ _2053_ vssd1 vssd1 vccd1 vccd1 _2057_ sky130_fd_sc_hd__a21o_1
XFILLER_65_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4308__A _0701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5923_ _0914_ _0913_ _0900_ vssd1 vssd1 vccd1 vccd1 _0916_ sky130_fd_sc_hd__a21bo_1
X_5854_ _0710_ _0842_ _0843_ vssd1 vssd1 vccd1 vccd1 _0844_ sky130_fd_sc_hd__and3_1
XFILLER_22_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8573_ clknet_3_6__leaf_clk _0059_ vssd1 vssd1 vccd1 vccd1 posit_add.in2\[0\] sky130_fd_sc_hd__dfxtp_2
X_4805_ _3793_ _3817_ _3959_ vssd1 vssd1 vccd1 vccd1 _3960_ sky130_fd_sc_hd__or3_1
X_5785_ _0766_ _0768_ vssd1 vssd1 vccd1 vccd1 _0769_ sky130_fd_sc_hd__xnor2_2
XFILLER_21_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7524_ _2657_ _2663_ vssd1 vssd1 vccd1 vccd1 _2664_ sky130_fd_sc_hd__xnor2_1
XFILLER_119_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4736_ _3857_ _3858_ vssd1 vssd1 vccd1 vccd1 _3891_ sky130_fd_sc_hd__xnor2_1
X_4667_ _3339_ _3349_ _2727_ _3360_ vssd1 vssd1 vccd1 vccd1 _3822_ sky130_fd_sc_hd__o211a_1
X_7455_ _2565_ _2587_ _2486_ vssd1 vssd1 vccd1 vccd1 _2588_ sky130_fd_sc_hd__mux2_1
X_6406_ _1425_ _1432_ vssd1 vssd1 vccd1 vccd1 _1434_ sky130_fd_sc_hd__and2b_1
X_7386_ _2511_ _2381_ _2409_ vssd1 vssd1 vccd1 vccd1 _2512_ sky130_fd_sc_hd__mux2_1
XFILLER_115_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6337_ _1004_ _1342_ vssd1 vssd1 vccd1 vccd1 _1358_ sky130_fd_sc_hd__or2_1
X_4598_ _2969_ _3530_ _3723_ _3520_ _3488_ vssd1 vssd1 vccd1 vccd1 _3753_ sky130_fd_sc_hd__o2111a_1
XFILLER_1_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6268_ _0802_ _1168_ vssd1 vssd1 vccd1 vccd1 _1282_ sky130_fd_sc_hd__nor2_1
X_6199_ _1203_ _1205_ vssd1 vssd1 vccd1 vccd1 _1207_ sky130_fd_sc_hd__and2_1
XFILLER_88_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5219_ _0178_ _0191_ vssd1 vssd1 vccd1 vccd1 _0192_ sky130_fd_sc_hd__xnor2_1
X_8007_ _1177_ vssd1 vssd1 vccd1 vccd1 _3195_ sky130_fd_sc_hd__clkbuf_4
XFILLER_29_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6966__A1 _3817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6433__A _1420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7529__A _0369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8159__B1 _2621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5570_ _0542_ _0539_ _0338_ vssd1 vssd1 vccd1 vccd1 _0543_ sky130_fd_sc_hd__mux2_1
XFILLER_117_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4521_ _3456_ _3498_ vssd1 vssd1 vccd1 vccd1 _3509_ sky130_fd_sc_hd__nand2_2
X_4452_ posit_add.in1\[9\] _2749_ vssd1 vssd1 vccd1 vccd1 _2760_ sky130_fd_sc_hd__xor2_4
X_7240_ _0349_ _0433_ vssd1 vssd1 vccd1 vccd1 _2351_ sky130_fd_sc_hd__nand2_1
XFILLER_104_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4383_ _1561_ _1638_ _1715_ vssd1 vssd1 vccd1 vccd1 _2001_ sky130_fd_sc_hd__and3_1
X_7171_ _2273_ _1624_ _2274_ vssd1 vssd1 vccd1 vccd1 _2275_ sky130_fd_sc_hd__and3b_1
X_6122_ _1123_ _1124_ vssd1 vssd1 vccd1 vccd1 _1125_ sky130_fd_sc_hd__or2b_1
XFILLER_98_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6053_ _0962_ _0973_ _0979_ _1052_ vssd1 vssd1 vccd1 vccd1 _1053_ sky130_fd_sc_hd__o31a_1
XFILLER_105_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5004_ _4157_ _4158_ vssd1 vssd1 vccd1 vccd1 _4159_ sky130_fd_sc_hd__xor2_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5141__B _4217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6955_ _2033_ _2037_ vssd1 vssd1 vccd1 vccd1 _2038_ sky130_fd_sc_hd__nor2_1
X_5906_ _0895_ _0896_ _0897_ vssd1 vssd1 vccd1 vccd1 _0898_ sky130_fd_sc_hd__nand3_1
XANTENNA__6253__A _0773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6886_ _1842_ _1953_ vssd1 vssd1 vccd1 vccd1 _1962_ sky130_fd_sc_hd__xnor2_1
XFILLER_22_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5837_ _3815_ _0693_ _0823_ vssd1 vssd1 vccd1 vccd1 _0825_ sky130_fd_sc_hd__or3_1
XFILLER_22_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5768_ _3814_ _0665_ vssd1 vssd1 vccd1 vccd1 _0751_ sky130_fd_sc_hd__nand2_1
X_8556_ clknet_3_1__leaf_clk _0042_ vssd1 vssd1 vccd1 vccd1 counter\[4\] sky130_fd_sc_hd__dfxtp_1
X_8487_ _3681_ vssd1 vssd1 vccd1 vccd1 _0061_ sky130_fd_sc_hd__clkbuf_1
X_4719_ _3793_ _3750_ vssd1 vssd1 vccd1 vccd1 _3874_ sky130_fd_sc_hd__or2_1
X_7507_ _3068_ _1451_ vssd1 vssd1 vccd1 vccd1 _2645_ sky130_fd_sc_hd__or2_1
XFILLER_108_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5699_ _0675_ vssd1 vssd1 vccd1 vccd1 _0676_ sky130_fd_sc_hd__buf_2
X_7438_ _2486_ vssd1 vssd1 vccd1 vccd1 _2569_ sky130_fd_sc_hd__buf_2
XFILLER_107_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7369_ _2396_ _2407_ _2449_ vssd1 vssd1 vccd1 vccd1 _2493_ sky130_fd_sc_hd__or3_1
XFILLER_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7958__S _2999_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6167__A2 _1128_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4653__A2 _3635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4292__S _0830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6740_ _1778_ _1800_ vssd1 vssd1 vccd1 vccd1 _1801_ sky130_fd_sc_hd__xor2_1
XANTENNA__7169__A _0080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6671_ _1446_ _0548_ vssd1 vssd1 vccd1 vccd1 _1725_ sky130_fd_sc_hd__nor2_1
XFILLER_50_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5905__A2 _0722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5622_ _0592_ _0538_ _0520_ vssd1 vssd1 vccd1 vccd1 _0595_ sky130_fd_sc_hd__or3_1
X_8410_ _3227_ _3188_ _3187_ vssd1 vssd1 vccd1 vccd1 _3623_ sky130_fd_sc_hd__o21ai_1
X_5553_ _0444_ _0443_ _0510_ vssd1 vssd1 vccd1 vccd1 _0526_ sky130_fd_sc_hd__mux2_1
X_8341_ _3534_ _3549_ _3550_ _3195_ vssd1 vssd1 vccd1 vccd1 _3551_ sky130_fd_sc_hd__a2bb2o_1
X_4504_ _2661_ vssd1 vssd1 vccd1 vccd1 _3328_ sky130_fd_sc_hd__clkbuf_8
X_8272_ _3475_ _3476_ vssd1 vssd1 vccd1 vccd1 _3478_ sky130_fd_sc_hd__nand2_1
XANTENNA__4321__A _1308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5484_ _0416_ _0438_ vssd1 vssd1 vccd1 vccd1 _0457_ sky130_fd_sc_hd__xnor2_2
XFILLER_105_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7223_ _0698_ _0687_ _2332_ vssd1 vssd1 vccd1 vccd1 _2333_ sky130_fd_sc_hd__nand3b_2
XANTENNA__5136__B _3750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4435_ posit_add.in1\[9\] posit_add.in1\[8\] posit_add.in1\[7\] _2562_ vssd1 vssd1
+ vccd1 vccd1 _2573_ sky130_fd_sc_hd__or4_2
XFILLER_116_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4366_ _1781_ _1803_ vssd1 vssd1 vccd1 vccd1 _1814_ sky130_fd_sc_hd__nand2_1
X_7154_ _1999_ _1949_ vssd1 vssd1 vccd1 vccd1 _2257_ sky130_fd_sc_hd__and2b_1
XFILLER_113_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6105_ _1095_ _1106_ vssd1 vssd1 vccd1 vccd1 _1107_ sky130_fd_sc_hd__xnor2_1
XANTENNA__6618__A0 _1420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7085_ _2152_ _2180_ vssd1 vssd1 vccd1 vccd1 _2181_ sky130_fd_sc_hd__nand2_1
X_4297_ _1051_ vssd1 vssd1 vccd1 vccd1 _0013_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5152__A _3816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6036_ _1026_ _1034_ vssd1 vssd1 vccd1 vccd1 _1035_ sky130_fd_sc_hd__and2_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7987_ _3154_ vssd1 vssd1 vccd1 vccd1 _3173_ sky130_fd_sc_hd__clkinv_2
XFILLER_14_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6938_ _2013_ _2018_ vssd1 vssd1 vccd1 vccd1 _2019_ sky130_fd_sc_hd__xnor2_1
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6869_ _1932_ _1937_ vssd1 vssd1 vccd1 vccd1 _1943_ sky130_fd_sc_hd__or2b_1
XFILLER_41_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8539_ clknet_3_1__leaf_clk _0025_ vssd1 vssd1 vccd1 vccd1 out_reg\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_10_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5062__A _3855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5997__A _4016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4406__A posit_add.in2\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7910_ _3087_ vssd1 vssd1 vccd1 vccd1 _3088_ sky130_fd_sc_hd__clkinv_2
XANTENNA__5700__A _3719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7841_ _2995_ _3008_ _3009_ _3011_ vssd1 vssd1 vccd1 vccd1 _3012_ sky130_fd_sc_hd__or4_1
XFILLER_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6515__B _1423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4984_ _4125_ _4131_ _4138_ vssd1 vssd1 vccd1 vccd1 _4139_ sky130_fd_sc_hd__a21o_1
X_7772_ _2918_ _2935_ vssd1 vssd1 vccd1 vccd1 _2937_ sky130_fd_sc_hd__nor2_4
XFILLER_36_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6723_ _1353_ _1354_ _1782_ vssd1 vssd1 vccd1 vccd1 _1783_ sky130_fd_sc_hd__and3_1
XFILLER_23_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6654_ _4018_ _1532_ vssd1 vssd1 vccd1 vccd1 _1707_ sky130_fd_sc_hd__xor2_1
XFILLER_32_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5605_ _0574_ _0577_ _0545_ vssd1 vssd1 vccd1 vccd1 _0578_ sky130_fd_sc_hd__a21o_1
X_6585_ _1383_ _0082_ vssd1 vssd1 vccd1 vccd1 _1631_ sky130_fd_sc_hd__or2_1
XFILLER_11_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8324_ _3481_ _3532_ _3531_ vssd1 vssd1 vccd1 vccd1 _3533_ sky130_fd_sc_hd__o21ai_1
X_5536_ _0508_ vssd1 vssd1 vccd1 vccd1 _0509_ sky130_fd_sc_hd__inv_2
X_8255_ _3458_ _3459_ vssd1 vssd1 vccd1 vccd1 _3460_ sky130_fd_sc_hd__nor2_2
X_5467_ _4250_ _0082_ _0399_ _0401_ _0439_ vssd1 vssd1 vccd1 vccd1 _0440_ sky130_fd_sc_hd__o32a_4
X_4418_ _1726_ _2353_ _2364_ _2375_ vssd1 vssd1 vccd1 vccd1 _2386_ sky130_fd_sc_hd__o211a_1
X_7206_ _2312_ _2313_ vssd1 vssd1 vccd1 vccd1 _2314_ sky130_fd_sc_hd__and2_1
XFILLER_99_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5398_ _2760_ _3307_ _3822_ _3477_ vssd1 vssd1 vccd1 vccd1 _0371_ sky130_fd_sc_hd__a211o_1
X_8186_ _3365_ _3385_ vssd1 vssd1 vccd1 vccd1 _3386_ sky130_fd_sc_hd__xnor2_1
XFILLER_113_470 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7137_ _2223_ _2237_ vssd1 vssd1 vccd1 vccd1 _2238_ sky130_fd_sc_hd__nor2_1
X_4349_ _1506_ _1583_ _1605_ vssd1 vssd1 vccd1 vccd1 _1627_ sky130_fd_sc_hd__a21oi_1
X_7068_ _1676_ _1537_ _2160_ _2086_ vssd1 vssd1 vccd1 vccd1 _2162_ sky130_fd_sc_hd__o31ai_1
XFILLER_86_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6019_ _0779_ _0803_ _0992_ vssd1 vssd1 vccd1 vccd1 _1017_ sky130_fd_sc_hd__or3_2
XFILLER_101_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6425__B _1454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6160__B _1164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5057__A _3925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4553__A1 _1946_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6616__A _4037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6335__B _1354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6370_ _1365_ _1368_ _1393_ vssd1 vssd1 vccd1 vccd1 _1394_ sky130_fd_sc_hd__and3_1
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5321_ _0292_ _0293_ vssd1 vssd1 vccd1 vccd1 _0294_ sky130_fd_sc_hd__or2b_1
XFILLER_114_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8040_ _3176_ _2993_ _3065_ vssd1 vssd1 vccd1 vccd1 _3230_ sky130_fd_sc_hd__mux2_1
XFILLER_102_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5252_ _0211_ _0222_ _0224_ vssd1 vssd1 vccd1 vccd1 _0225_ sky130_fd_sc_hd__a21o_1
X_5183_ _0141_ _0155_ vssd1 vssd1 vccd1 vccd1 _0156_ sky130_fd_sc_hd__or2b_1
XFILLER_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5133__C _0105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7824_ _2981_ _2960_ _2979_ vssd1 vssd1 vccd1 vccd1 _2994_ sky130_fd_sc_hd__nor3_1
XFILLER_51_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4967_ _4119_ _4121_ vssd1 vssd1 vccd1 vccd1 _4122_ sky130_fd_sc_hd__xor2_1
X_7755_ _2904_ _2917_ vssd1 vssd1 vccd1 vccd1 _2918_ sky130_fd_sc_hd__or2_2
X_6706_ _1565_ _1580_ vssd1 vssd1 vccd1 vccd1 _1764_ sky130_fd_sc_hd__xnor2_1
X_4898_ _4051_ _4052_ vssd1 vssd1 vccd1 vccd1 _4053_ sky130_fd_sc_hd__xor2_1
X_7686_ _2710_ _2841_ _1297_ vssd1 vssd1 vccd1 vccd1 _2842_ sky130_fd_sc_hd__a21oi_4
XANTENNA__7076__B _1718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6637_ _1683_ _1687_ vssd1 vssd1 vccd1 vccd1 _1688_ sky130_fd_sc_hd__xor2_1
X_6568_ _1609_ _1611_ vssd1 vssd1 vccd1 vccd1 _1612_ sky130_fd_sc_hd__nor2_1
XFILLER_22_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8307_ _3462_ _3468_ _3491_ _1319_ vssd1 vssd1 vccd1 vccd1 _3515_ sky130_fd_sc_hd__o31a_1
XFILLER_3_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5519_ _0487_ _0491_ _0480_ vssd1 vssd1 vccd1 vccd1 _0492_ sky130_fd_sc_hd__mux2_1
X_6499_ _1226_ _1305_ _1191_ vssd1 vssd1 vccd1 vccd1 _1536_ sky130_fd_sc_hd__o21ai_1
XFILLER_105_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8238_ _3440_ _3441_ vssd1 vssd1 vccd1 vccd1 _3442_ sky130_fd_sc_hd__nor2_1
XFILLER_59_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8169_ _1330_ _3359_ _3367_ vssd1 vssd1 vccd1 vccd1 _3368_ sky130_fd_sc_hd__a21oi_1
XFILLER_87_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7966__S _2999_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6171__A _0706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4526__A1 _3232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6451__B2 _0121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6451__A1 _0218_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5870_ _0858_ _0859_ vssd1 vssd1 vccd1 vccd1 _0860_ sky130_fd_sc_hd__xnor2_1
XFILLER_80_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7876__S _2999_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5006__A2 _3883_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4821_ _3970_ _3974_ vssd1 vssd1 vccd1 vccd1 _3976_ sky130_fd_sc_hd__nand2_1
X_4752_ _3772_ _3826_ vssd1 vssd1 vccd1 vccd1 _3907_ sky130_fd_sc_hd__nor2_2
XFILLER_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7540_ _3328_ _1781_ vssd1 vssd1 vccd1 vccd1 _2681_ sky130_fd_sc_hd__nor2_1
XFILLER_119_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4683_ _3721_ _3835_ _3836_ _3837_ vssd1 vssd1 vccd1 vccd1 _3838_ sky130_fd_sc_hd__a31o_4
X_7471_ _2487_ _2576_ _2599_ _2603_ _2604_ vssd1 vssd1 vccd1 vccd1 _2605_ sky130_fd_sc_hd__o41a_1
X_6422_ _0148_ _1449_ _4213_ vssd1 vssd1 vccd1 vccd1 _1452_ sky130_fd_sc_hd__and3b_1
X_6353_ _1323_ _1329_ vssd1 vssd1 vccd1 vccd1 _1376_ sky130_fd_sc_hd__or2_1
X_6284_ _1278_ _1298_ _1299_ vssd1 vssd1 vccd1 vccd1 _1300_ sky130_fd_sc_hd__or3_2
X_5304_ _2540_ _4232_ _0276_ vssd1 vssd1 vccd1 vccd1 _0277_ sky130_fd_sc_hd__or3b_1
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5235_ _0206_ _0207_ vssd1 vssd1 vccd1 vccd1 _0208_ sky130_fd_sc_hd__or2_1
X_8023_ _3211_ vssd1 vssd1 vccd1 vccd1 _3212_ sky130_fd_sc_hd__buf_2
XFILLER_96_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5166_ _3881_ _3855_ _0137_ vssd1 vssd1 vccd1 vccd1 _0139_ sky130_fd_sc_hd__a21o_1
XFILLER_56_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5097_ _4228_ _3925_ vssd1 vssd1 vccd1 vccd1 _4252_ sky130_fd_sc_hd__nor2_1
XFILLER_84_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5999_ _4016_ _0892_ _0702_ _0991_ vssd1 vssd1 vccd1 vccd1 _0996_ sky130_fd_sc_hd__or4_2
XANTENNA__6745__A2 _1510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7807_ _2961_ _2972_ vssd1 vssd1 vccd1 vccd1 _2975_ sky130_fd_sc_hd__xnor2_1
XFILLER_40_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7738_ _2898_ vssd1 vssd1 vccd1 vccd1 _2899_ sky130_fd_sc_hd__inv_2
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7669_ _2761_ _2821_ _2822_ vssd1 vssd1 vccd1 vccd1 _2823_ sky130_fd_sc_hd__o21a_1
XFILLER_109_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7630__A0 _3793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5245__A _4228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5020_ _3776_ _3878_ _3855_ _4174_ vssd1 vssd1 vccd1 vccd1 _4175_ sky130_fd_sc_hd__and4_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6971_ _1414_ _3804_ vssd1 vssd1 vccd1 vccd1 _2055_ sky130_fd_sc_hd__and2_1
XFILLER_81_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5922_ _0900_ _0913_ _0914_ vssd1 vssd1 vccd1 vccd1 _0915_ sky130_fd_sc_hd__nand3b_2
XFILLER_81_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5853_ _0708_ _0709_ _0644_ vssd1 vssd1 vccd1 vccd1 _0843_ sky130_fd_sc_hd__a21o_1
XFILLER_22_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5784_ _0715_ _0767_ vssd1 vssd1 vccd1 vccd1 _0768_ sky130_fd_sc_hd__xor2_1
X_8572_ clknet_3_2__leaf_clk _0058_ vssd1 vssd1 vccd1 vccd1 posit_add.in1\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4804_ _3878_ _3868_ vssd1 vssd1 vccd1 vccd1 _3959_ sky130_fd_sc_hd__nand2_1
XFILLER_21_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4735_ _3888_ _3889_ vssd1 vssd1 vccd1 vccd1 _3890_ sky130_fd_sc_hd__nand2_1
XFILLER_21_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7523_ _0399_ _2654_ vssd1 vssd1 vccd1 vccd1 _2663_ sky130_fd_sc_hd__or2_1
XFILLER_119_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4666_ _2694_ _3318_ _3820_ _3488_ vssd1 vssd1 vccd1 vccd1 _3821_ sky130_fd_sc_hd__a211o_1
X_7454_ _2522_ _2577_ _2586_ vssd1 vssd1 vccd1 vccd1 _2587_ sky130_fd_sc_hd__a21oi_1
X_6405_ _1425_ _1432_ vssd1 vssd1 vccd1 vccd1 _1433_ sky130_fd_sc_hd__xnor2_1
XANTENNA__5163__A1 _3816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4597_ _3189_ _3318_ _3745_ _3488_ vssd1 vssd1 vccd1 vccd1 _3752_ sky130_fd_sc_hd__a211o_1
X_7385_ _0218_ _2431_ _2442_ _2503_ _2510_ vssd1 vssd1 vccd1 vccd1 _2511_ sky130_fd_sc_hd__o221a_1
X_6336_ _1344_ _1343_ vssd1 vssd1 vccd1 vccd1 _1357_ sky130_fd_sc_hd__and2b_1
XFILLER_103_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6267_ _1279_ _1280_ vssd1 vssd1 vccd1 vccd1 _1281_ sky130_fd_sc_hd__nor2_1
X_6198_ _1203_ _1205_ vssd1 vssd1 vccd1 vccd1 _1206_ sky130_fd_sc_hd__xor2_1
XFILLER_88_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5218_ _0179_ _0189_ _0190_ vssd1 vssd1 vccd1 vccd1 _0191_ sky130_fd_sc_hd__a21bo_1
X_8006_ _0598_ _0600_ _0602_ _3193_ vssd1 vssd1 vccd1 vccd1 _3194_ sky130_fd_sc_hd__o31a_1
X_5149_ _3881_ _0121_ _4182_ vssd1 vssd1 vccd1 vccd1 _0122_ sky130_fd_sc_hd__and3_1
XFILLER_29_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6433__B _1399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5065__A _4210_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4520_ _2936_ _3318_ _3467_ _3488_ vssd1 vssd1 vccd1 vccd1 _3498_ sky130_fd_sc_hd__a211o_1
XFILLER_11_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4451_ posit_add.in1\[8\] _2617_ _1242_ vssd1 vssd1 vccd1 vccd1 _2749_ sky130_fd_sc_hd__o21a_1
XFILLER_7_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7170_ _4250_ _0303_ vssd1 vssd1 vccd1 vccd1 _2274_ sky130_fd_sc_hd__nor2_1
X_6121_ _1117_ _1110_ vssd1 vssd1 vccd1 vccd1 _1124_ sky130_fd_sc_hd__xnor2_1
XFILLER_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4382_ _1759_ _1979_ _1561_ vssd1 vssd1 vccd1 vccd1 _1990_ sky130_fd_sc_hd__o21ai_4
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6052_ _0978_ _0971_ vssd1 vssd1 vccd1 vccd1 _1052_ sky130_fd_sc_hd__or2b_1
XFILLER_112_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_387 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5003_ _3924_ _3930_ vssd1 vssd1 vccd1 vccd1 _4158_ sky130_fd_sc_hd__nor2_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6954_ _1988_ _2035_ _2036_ vssd1 vssd1 vccd1 vccd1 _2037_ sky130_fd_sc_hd__a21boi_1
XFILLER_19_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5905_ _3878_ _0722_ _0706_ _3776_ vssd1 vssd1 vccd1 vccd1 _0897_ sky130_fd_sc_hd__a22o_1
XFILLER_81_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6885_ _1599_ _0548_ _1960_ vssd1 vssd1 vccd1 vccd1 _1961_ sky130_fd_sc_hd__or3_1
XFILLER_14_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5836_ _3815_ _0693_ _0823_ vssd1 vssd1 vccd1 vccd1 _0824_ sky130_fd_sc_hd__o21ai_1
X_5767_ _2507_ _3815_ _3792_ _0732_ vssd1 vssd1 vccd1 vccd1 _0750_ sky130_fd_sc_hd__a22o_1
X_8555_ clknet_3_0__leaf_clk _0041_ vssd1 vssd1 vccd1 vccd1 counter\[3\] sky130_fd_sc_hd__dfxtp_1
X_5698_ _0660_ _0674_ _3924_ vssd1 vssd1 vccd1 vccd1 _0675_ sky130_fd_sc_hd__mux2_1
X_8486_ posit_add.in2\[2\] in_reg\[2\] _3677_ vssd1 vssd1 vccd1 vccd1 _3681_ sky130_fd_sc_hd__mux2_1
X_4718_ _3869_ _3870_ _3872_ vssd1 vssd1 vccd1 vccd1 _3873_ sky130_fd_sc_hd__o21ai_1
X_7506_ _3101_ _1484_ _1583_ _2727_ vssd1 vssd1 vccd1 vccd1 _2644_ sky130_fd_sc_hd__a22o_1
X_4649_ _3803_ vssd1 vssd1 vccd1 vccd1 _3804_ sky130_fd_sc_hd__buf_4
X_7437_ _2565_ _2567_ vssd1 vssd1 vccd1 vccd1 _2568_ sky130_fd_sc_hd__nand2_1
XANTENNA__6884__A1 _1423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4895__B1 _3868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7368_ _2378_ _2481_ _2410_ _2491_ vssd1 vssd1 vccd1 vccd1 _2492_ sky130_fd_sc_hd__a2bb2o_1
X_6319_ _4210_ _0702_ _0993_ _1097_ vssd1 vssd1 vccd1 vccd1 _1338_ sky130_fd_sc_hd__or4b_2
XFILLER_89_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8086__B1 _0701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7299_ _2415_ vssd1 vssd1 vccd1 vccd1 _2416_ sky130_fd_sc_hd__clkbuf_4
XFILLER_91_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6444__A _1383_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4899__A _3878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6619__A _3986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7169__B _1446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6670_ _1681_ _1722_ _1723_ vssd1 vssd1 vccd1 vccd1 _1724_ sky130_fd_sc_hd__o21a_1
XFILLER_31_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5621_ _0520_ _0593_ vssd1 vssd1 vccd1 vccd1 _0594_ sky130_fd_sc_hd__and2b_1
X_5552_ _0397_ _0440_ _0468_ _0511_ vssd1 vssd1 vccd1 vccd1 _0525_ sky130_fd_sc_hd__o31ai_1
X_8340_ out_reg\[10\] _3242_ vssd1 vssd1 vccd1 vccd1 _3550_ sky130_fd_sc_hd__nand2_1
X_4503_ _3307_ vssd1 vssd1 vccd1 vccd1 _3318_ sky130_fd_sc_hd__buf_2
XFILLER_8_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8271_ _3455_ _3474_ vssd1 vssd1 vccd1 vccd1 _3476_ sky130_fd_sc_hd__or2_1
XFILLER_105_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5483_ _0447_ _0453_ _0441_ _0455_ vssd1 vssd1 vccd1 vccd1 _0456_ sky130_fd_sc_hd__or4b_1
X_7222_ _3925_ _3828_ _3771_ _3845_ vssd1 vssd1 vccd1 vccd1 _2332_ sky130_fd_sc_hd__and4_1
X_4434_ posit_add.in1\[6\] posit_add.in1\[5\] posit_add.in1\[4\] _2551_ vssd1 vssd1
+ vccd1 vccd1 _2562_ sky130_fd_sc_hd__or4_1
XFILLER_6_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8068__A0 _0440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4365_ posit_add.in2\[2\] _1792_ vssd1 vssd1 vccd1 vccd1 _1803_ sky130_fd_sc_hd__xor2_4
X_7153_ _2085_ _2247_ _2253_ _2255_ vssd1 vssd1 vccd1 vccd1 _2256_ sky130_fd_sc_hd__a31oi_4
XFILLER_113_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6104_ _1104_ _1105_ vssd1 vssd1 vccd1 vccd1 _1106_ sky130_fd_sc_hd__xnor2_1
XFILLER_98_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7084_ _2153_ _2175_ _2179_ vssd1 vssd1 vccd1 vccd1 _2180_ sky130_fd_sc_hd__o21a_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6035_ _1004_ _1027_ _1032_ _1033_ vssd1 vssd1 vccd1 vccd1 _1034_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_100_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4296_ in_reg\[9\] in_reg\[10\] _0819_ vssd1 vssd1 vccd1 vccd1 _1051_ sky130_fd_sc_hd__mux2_1
XANTENNA__5152__B _3989_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4629__B1 _3189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7043__A1 _1456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7986_ _3102_ _3162_ _3165_ _3171_ vssd1 vssd1 vccd1 vccd1 _3172_ sky130_fd_sc_hd__or4b_1
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6937_ _1665_ _2014_ _2017_ vssd1 vssd1 vccd1 vccd1 _2018_ sky130_fd_sc_hd__a21bo_1
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6868_ _1936_ vssd1 vssd1 vccd1 vccd1 _1942_ sky130_fd_sc_hd__inv_2
XFILLER_22_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5819_ _4222_ _3700_ _0113_ _0706_ _0804_ vssd1 vssd1 vccd1 vccd1 _0805_ sky130_fd_sc_hd__a41o_1
XFILLER_50_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6799_ _1401_ _1510_ vssd1 vssd1 vccd1 vccd1 _1866_ sky130_fd_sc_hd__nor2_1
X_8538_ clknet_3_1__leaf_clk _0024_ vssd1 vssd1 vccd1 vccd1 out_reg\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_10_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8469_ in_reg\[11\] posit_add.in1\[11\] _3654_ vssd1 vssd1 vccd1 vccd1 _3669_ sky130_fd_sc_hd__mux2_1
XFILLER_2_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6439__A _0080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8231__B1 _0600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4406__B _1781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6068__B _3739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7879__S _2954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7840_ _2974_ _3010_ vssd1 vssd1 vccd1 vccd1 _3011_ sky130_fd_sc_hd__and2_1
XFILLER_91_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4983_ _4136_ _4137_ vssd1 vssd1 vccd1 vccd1 _4138_ sky130_fd_sc_hd__or2_1
X_7771_ _2926_ _2934_ vssd1 vssd1 vccd1 vccd1 _2935_ sky130_fd_sc_hd__nor2_1
XFILLER_23_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6722_ _3868_ vssd1 vssd1 vccd1 vccd1 _1782_ sky130_fd_sc_hd__clkbuf_4
XFILLER_16_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6653_ _1625_ _1705_ vssd1 vssd1 vccd1 vccd1 _1706_ sky130_fd_sc_hd__nand2_1
XANTENNA__6000__A2 _0702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5604_ _0494_ _0556_ vssd1 vssd1 vccd1 vccd1 _0577_ sky130_fd_sc_hd__or2_1
X_6584_ _1623_ _1629_ vssd1 vssd1 vccd1 vccd1 _1630_ sky130_fd_sc_hd__xor2_1
XFILLER_11_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8323_ _3485_ _3505_ _1308_ vssd1 vssd1 vccd1 vccd1 _3532_ sky130_fd_sc_hd__o21a_1
X_5535_ _0503_ _0507_ _0480_ vssd1 vssd1 vccd1 vccd1 _0508_ sky130_fd_sc_hd__mux2_1
XFILLER_105_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8254_ _3394_ _3395_ _3442_ _3182_ vssd1 vssd1 vccd1 vccd1 _3459_ sky130_fd_sc_hd__o31a_1
X_5466_ _0416_ _0438_ _0413_ vssd1 vssd1 vccd1 vccd1 _0439_ sky130_fd_sc_hd__a21o_1
XFILLER_105_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4417_ posit_add.in2\[2\] _1792_ vssd1 vssd1 vccd1 vccd1 _2375_ sky130_fd_sc_hd__xnor2_1
X_7205_ _2308_ _2311_ vssd1 vssd1 vccd1 vccd1 _2313_ sky130_fd_sc_hd__nand2_1
XFILLER_101_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8185_ _3383_ _3384_ _3259_ vssd1 vssd1 vccd1 vccd1 _3385_ sky130_fd_sc_hd__mux2_1
X_5397_ _0369_ vssd1 vssd1 vccd1 vccd1 _0370_ sky130_fd_sc_hd__clkinv_2
XFILLER_113_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7136_ _2226_ _2235_ _2236_ vssd1 vssd1 vccd1 vccd1 _2237_ sky130_fd_sc_hd__o21ba_1
XFILLER_86_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4348_ _1429_ _1583_ _1605_ vssd1 vssd1 vccd1 vccd1 _1616_ sky130_fd_sc_hd__o21a_1
XANTENNA_input3_A io_in[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7789__S _2721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7067_ _1676_ _1537_ _2086_ _2160_ vssd1 vssd1 vccd1 vccd1 _2161_ sky130_fd_sc_hd__or4_1
XFILLER_100_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8461__A0 in_reg\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4279_ _0862_ vssd1 vssd1 vccd1 vccd1 _0004_ sky130_fd_sc_hd__clkbuf_1
XFILLER_74_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6018_ _0779_ _0803_ _0992_ vssd1 vssd1 vccd1 vccd1 _1016_ sky130_fd_sc_hd__a21o_1
XFILLER_100_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7969_ _3051_ _3064_ _3065_ vssd1 vssd1 vccd1 vccd1 _3153_ sky130_fd_sc_hd__mux2_1
XFILLER_14_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6722__A _3868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_447 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_609 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5057__B _4037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5073__A _3827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_720 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6335__C _1355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_414 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5320_ _0290_ _0288_ vssd1 vssd1 vccd1 vccd1 _0293_ sky130_fd_sc_hd__xnor2_1
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4298__S _0819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5251_ _0171_ _0223_ vssd1 vssd1 vccd1 vccd1 _0224_ sky130_fd_sc_hd__xor2_1
XANTENNA__7494__A1 _3189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7494__B2 _3232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5182_ _0143_ _0154_ vssd1 vssd1 vccd1 vccd1 _0155_ sky130_fd_sc_hd__xnor2_1
XFILLER_110_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7823_ _2658_ _2659_ _2989_ _2992_ vssd1 vssd1 vccd1 vccd1 _2993_ sky130_fd_sc_hd__o22ai_4
XFILLER_36_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7754_ _2906_ _2908_ _2916_ vssd1 vssd1 vccd1 vccd1 _2917_ sky130_fd_sc_hd__or3_1
X_4966_ _4101_ _4120_ vssd1 vssd1 vccd1 vccd1 _4121_ sky130_fd_sc_hd__nand2_1
X_6705_ _1758_ _1754_ vssd1 vssd1 vccd1 vccd1 _1763_ sky130_fd_sc_hd__or2b_1
XFILLER_51_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4897_ _3892_ _3832_ _3943_ _3868_ vssd1 vssd1 vccd1 vccd1 _4052_ sky130_fd_sc_hd__and4_1
XFILLER_51_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7685_ _2835_ _2839_ _2840_ vssd1 vssd1 vccd1 vccd1 _2841_ sky130_fd_sc_hd__a21oi_2
X_6636_ _1685_ _1686_ vssd1 vssd1 vccd1 vccd1 _1687_ sky130_fd_sc_hd__xor2_2
X_6567_ _1493_ _1504_ _1610_ vssd1 vssd1 vccd1 vccd1 _1611_ sky130_fd_sc_hd__a21oi_1
XFILLER_106_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8306_ _3511_ _3512_ _3190_ vssd1 vssd1 vccd1 vccd1 _3514_ sky130_fd_sc_hd__o21a_1
X_5518_ _0489_ _0490_ _0469_ vssd1 vssd1 vccd1 vccd1 _0491_ sky130_fd_sc_hd__mux2_1
X_6498_ _1191_ _1226_ _1305_ vssd1 vssd1 vccd1 vccd1 _1535_ sky130_fd_sc_hd__or3_1
XFILLER_3_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8237_ _3391_ _3439_ vssd1 vssd1 vccd1 vccd1 _3441_ sky130_fd_sc_hd__nor2_1
X_5449_ _3736_ _0420_ _0421_ vssd1 vssd1 vccd1 vccd1 _0422_ sky130_fd_sc_hd__mux2_1
XFILLER_87_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8168_ _3365_ _3366_ vssd1 vssd1 vccd1 vccd1 _3367_ sky130_fd_sc_hd__nor2_1
XFILLER_113_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7119_ _2202_ _2204_ _2217_ vssd1 vssd1 vccd1 vccd1 _2218_ sky130_fd_sc_hd__and3_1
XFILLER_87_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6717__A _0303_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7237__A1 _0351_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8099_ _3290_ _3291_ _3292_ vssd1 vssd1 vccd1 vccd1 _3293_ sky130_fd_sc_hd__o21ai_1
XFILLER_101_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7945__C1 _2941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5068__A _4222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6362__A _1383_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4820_ _3970_ _3974_ vssd1 vssd1 vccd1 vccd1 _3975_ sky130_fd_sc_hd__xnor2_1
XFILLER_33_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4751_ _3896_ _3905_ vssd1 vssd1 vccd1 vccd1 _3906_ sky130_fd_sc_hd__xnor2_1
XFILLER_119_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4682_ _3594_ _3156_ _3786_ vssd1 vssd1 vccd1 vccd1 _3837_ sky130_fd_sc_hd__and3_1
X_7470_ _2520_ vssd1 vssd1 vccd1 vccd1 _2604_ sky130_fd_sc_hd__buf_2
XFILLER_119_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5714__A1 _4222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6421_ _4211_ _1449_ _0148_ vssd1 vssd1 vccd1 vccd1 _1450_ sky130_fd_sc_hd__and3_1
XFILLER_108_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6352_ _1373_ vssd1 vssd1 vccd1 vccd1 _1375_ sky130_fd_sc_hd__inv_2
XANTENNA__4610__A posit_add.in2\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6283_ _1260_ _1273_ vssd1 vssd1 vccd1 vccd1 _1299_ sky130_fd_sc_hd__xnor2_1
X_5303_ _0274_ _0273_ vssd1 vssd1 vccd1 vccd1 _0276_ sky130_fd_sc_hd__xnor2_1
XFILLER_102_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5234_ _0164_ _0205_ vssd1 vssd1 vccd1 vccd1 _0207_ sky130_fd_sc_hd__and2_1
X_8022_ cmd\[6\] _2319_ cmd\[7\] vssd1 vssd1 vccd1 vccd1 _3211_ sky130_fd_sc_hd__and3b_1
X_5165_ _3855_ _0137_ vssd1 vssd1 vccd1 vccd1 _0138_ sky130_fd_sc_hd__nand2_1
XANTENNA__8416__B1 _1177_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5096_ _4250_ _3988_ vssd1 vssd1 vccd1 vccd1 _4251_ sky130_fd_sc_hd__or2_2
XFILLER_83_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7806_ _2842_ _2973_ vssd1 vssd1 vccd1 vccd1 _2974_ sky130_fd_sc_hd__nand2_1
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5998_ _0795_ _0994_ vssd1 vssd1 vccd1 vccd1 _0995_ sky130_fd_sc_hd__nand2_1
XFILLER_52_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4949_ _4101_ _4103_ vssd1 vssd1 vccd1 vccd1 _4104_ sky130_fd_sc_hd__or2b_1
X_7737_ _2741_ _2897_ vssd1 vssd1 vccd1 vccd1 _2898_ sky130_fd_sc_hd__xnor2_1
X_7668_ _2758_ _2759_ vssd1 vssd1 vccd1 vccd1 _2822_ sky130_fd_sc_hd__or2_1
XFILLER_33_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6619_ _3986_ _1414_ vssd1 vssd1 vccd1 vccd1 _1668_ sky130_fd_sc_hd__nand2_2
XFILLER_20_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7599_ _2712_ _2745_ vssd1 vssd1 vccd1 vccd1 _2746_ sky130_fd_sc_hd__nor2_1
XFILLER_106_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7630__A1 _3795_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4430__A _1748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6672__A2 _4157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6970_ _2017_ _2049_ _2053_ vssd1 vssd1 vccd1 vccd1 _2054_ sky130_fd_sc_hd__nand3_1
XFILLER_81_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5921_ _0870_ _0871_ _0872_ vssd1 vssd1 vccd1 vccd1 _0914_ sky130_fd_sc_hd__nand3_1
XFILLER_81_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5852_ _0837_ _0838_ _0839_ _0840_ vssd1 vssd1 vccd1 vccd1 _0842_ sky130_fd_sc_hd__a31o_1
XFILLER_61_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5783_ _3901_ _0634_ vssd1 vssd1 vccd1 vccd1 _0767_ sky130_fd_sc_hd__nand2_1
X_8571_ clknet_3_5__leaf_clk _0057_ vssd1 vssd1 vccd1 vccd1 posit_add.in1\[14\] sky130_fd_sc_hd__dfxtp_4
XFILLER_61_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4803_ _3956_ _3957_ vssd1 vssd1 vccd1 vccd1 _3958_ sky130_fd_sc_hd__xnor2_1
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4734_ _3862_ _3887_ vssd1 vssd1 vccd1 vccd1 _3889_ sky130_fd_sc_hd__or2_1
X_7522_ _2653_ _2660_ vssd1 vssd1 vccd1 vccd1 _2662_ sky130_fd_sc_hd__xnor2_4
XFILLER_119_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4665_ _3339_ _3349_ _3819_ _3360_ vssd1 vssd1 vccd1 vccd1 _3820_ sky130_fd_sc_hd__o211a_1
X_7453_ _2454_ _2465_ _2580_ _2451_ vssd1 vssd1 vccd1 vccd1 _2586_ sky130_fd_sc_hd__o211a_1
X_6404_ _1426_ _1431_ vssd1 vssd1 vccd1 vccd1 _1432_ sky130_fd_sc_hd__xor2_1
XANTENNA__5163__A2 _4232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4596_ _2903_ _3318_ _3742_ _3446_ vssd1 vssd1 vccd1 vccd1 _3751_ sky130_fd_sc_hd__a211o_1
X_7384_ _2504_ _2509_ _2444_ vssd1 vssd1 vccd1 vccd1 _2510_ sky130_fd_sc_hd__o21ai_1
XFILLER_89_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6335_ _1353_ _1354_ _1355_ vssd1 vssd1 vccd1 vccd1 _1356_ sky130_fd_sc_hd__and3_1
XFILLER_89_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6266_ _1268_ _1267_ _1266_ vssd1 vssd1 vccd1 vccd1 _1280_ sky130_fd_sc_hd__a21oi_1
X_8005_ _2619_ _2621_ _2622_ _3192_ vssd1 vssd1 vccd1 vccd1 _3193_ sky130_fd_sc_hd__o31a_1
X_6197_ _1176_ _1204_ vssd1 vssd1 vccd1 vccd1 _1205_ sky130_fd_sc_hd__and2b_1
XFILLER_103_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5217_ _0188_ _0182_ vssd1 vssd1 vccd1 vccd1 _0190_ sky130_fd_sc_hd__or2b_1
XFILLER_57_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5148_ _4174_ vssd1 vssd1 vccd1 vccd1 _0121_ sky130_fd_sc_hd__buf_4
XFILLER_84_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5079_ _3988_ _4223_ vssd1 vssd1 vccd1 vccd1 _4234_ sky130_fd_sc_hd__nor2_1
XFILLER_84_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6730__A _1423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8421__S _0819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7826__A _2993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5065__B _4037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4450_ _2606_ _2727_ vssd1 vssd1 vccd1 vccd1 _2738_ sky130_fd_sc_hd__xnor2_2
XFILLER_7_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4381_ _1770_ _1814_ _1968_ vssd1 vssd1 vccd1 vccd1 _1979_ sky130_fd_sc_hd__o21ba_1
X_6120_ _1117_ _1122_ _1031_ vssd1 vssd1 vccd1 vccd1 _1123_ sky130_fd_sc_hd__o21ba_1
XFILLER_112_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6051_ _1035_ _1037_ _1049_ vssd1 vssd1 vccd1 vccd1 _1050_ sky130_fd_sc_hd__o21ai_2
XFILLER_86_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5002_ _4016_ _3702_ vssd1 vssd1 vccd1 vccd1 _4157_ sky130_fd_sc_hd__nor2_2
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8506__S _3676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6953_ _2031_ _2032_ vssd1 vssd1 vccd1 vccd1 _2036_ sky130_fd_sc_hd__nand2_1
XFILLER_81_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5081__A1 _4222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5904_ _3770_ _0773_ _0823_ vssd1 vssd1 vccd1 vccd1 _0896_ sky130_fd_sc_hd__or3_1
X_6884_ _1423_ _0548_ _1958_ _1959_ vssd1 vssd1 vccd1 vccd1 _1960_ sky130_fd_sc_hd__o31a_1
XFILLER_81_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_3_5__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_5__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5835_ _3792_ _0700_ vssd1 vssd1 vccd1 vccd1 _0823_ sky130_fd_sc_hd__or2_1
XFILLER_62_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5766_ _3718_ _3775_ _0746_ _0748_ _3924_ vssd1 vssd1 vccd1 vccd1 _0749_ sky130_fd_sc_hd__o221a_1
X_8554_ clknet_3_0__leaf_clk _0040_ vssd1 vssd1 vccd1 vccd1 counter\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5697_ _3700_ _0662_ _0664_ _0669_ _0673_ vssd1 vssd1 vccd1 vccd1 _0674_ sky130_fd_sc_hd__o32a_1
X_4717_ _3871_ _3782_ vssd1 vssd1 vccd1 vccd1 _3872_ sky130_fd_sc_hd__or2_1
X_8485_ _3680_ vssd1 vssd1 vccd1 vccd1 _0060_ sky130_fd_sc_hd__clkbuf_1
X_7505_ _2640_ _2641_ _2642_ vssd1 vssd1 vccd1 vccd1 _2643_ sky130_fd_sc_hd__a21oi_1
XANTENNA__4592__B1 _3232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4648_ _3722_ _3724_ vssd1 vssd1 vccd1 vccd1 _3803_ sky130_fd_sc_hd__and2_1
X_7436_ _2566_ _2467_ _2494_ vssd1 vssd1 vccd1 vccd1 _2567_ sky130_fd_sc_hd__mux2_1
XFILLER_30_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6884__A2 _0548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4579_ _3729_ _3733_ vssd1 vssd1 vccd1 vccd1 _3734_ sky130_fd_sc_hd__or2_1
XANTENNA__4895__B2 _3776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7367_ _2350_ _2376_ vssd1 vssd1 vccd1 vccd1 _2491_ sky130_fd_sc_hd__nor2_1
X_6318_ _1045_ _1042_ vssd1 vssd1 vccd1 vccd1 _1337_ sky130_fd_sc_hd__and2b_1
XFILLER_1_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7298_ _2327_ _2330_ vssd1 vssd1 vccd1 vccd1 _2415_ sky130_fd_sc_hd__and2_1
X_6249_ _1238_ _1245_ vssd1 vssd1 vccd1 vccd1 _1261_ sky130_fd_sc_hd__xor2_1
XFILLER_89_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7597__A0 _1355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6444__B _3840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6021__B1 _0754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6619__B _1414_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6635__A _1400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5620_ _0538_ _0558_ _0591_ _0592_ vssd1 vssd1 vccd1 vccd1 _0593_ sky130_fd_sc_hd__a31o_1
X_5551_ _0522_ _0523_ _0515_ vssd1 vssd1 vccd1 vccd1 _0524_ sky130_fd_sc_hd__mux2_1
X_4502_ _3079_ _3296_ _3046_ vssd1 vssd1 vccd1 vccd1 _3307_ sky130_fd_sc_hd__a21o_2
X_8270_ _3455_ _3474_ vssd1 vssd1 vccd1 vccd1 _3475_ sky130_fd_sc_hd__nand2_1
XFILLER_117_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5482_ _0450_ _0454_ vssd1 vssd1 vccd1 vccd1 _0455_ sky130_fd_sc_hd__xnor2_2
X_7221_ _2312_ _2325_ _2329_ vssd1 vssd1 vccd1 vccd1 _2330_ sky130_fd_sc_hd__o21a_1
X_4433_ posit_add.in1\[0\] posit_add.in1\[3\] posit_add.in1\[2\] posit_add.in1\[1\]
+ vssd1 vssd1 vccd1 vccd1 _2551_ sky130_fd_sc_hd__or4_2
XFILLER_116_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4364_ _1275_ _1770_ vssd1 vssd1 vccd1 vccd1 _1792_ sky130_fd_sc_hd__nand2_2
X_7152_ _2251_ _2083_ _2252_ vssd1 vssd1 vccd1 vccd1 _2255_ sky130_fd_sc_hd__o21a_1
XFILLER_113_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6103_ _0795_ _1102_ vssd1 vssd1 vccd1 vccd1 _1105_ sky130_fd_sc_hd__nand2_1
X_7083_ _2176_ _2178_ vssd1 vssd1 vccd1 vccd1 _2179_ sky130_fd_sc_hd__or2b_1
X_4295_ _1030_ vssd1 vssd1 vccd1 vccd1 _0012_ sky130_fd_sc_hd__clkbuf_1
XFILLER_86_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6034_ _1015_ _1022_ vssd1 vssd1 vccd1 vccd1 _1033_ sky130_fd_sc_hd__nand2_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7043__A2 _1537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7985_ _2950_ _3034_ _3170_ vssd1 vssd1 vccd1 vccd1 _3171_ sky130_fd_sc_hd__o21ba_1
XANTENNA__8240__A1 _3182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6936_ _1509_ _3703_ _2016_ vssd1 vssd1 vccd1 vccd1 _2017_ sky130_fd_sc_hd__or3b_1
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6867_ _1903_ _1940_ vssd1 vssd1 vccd1 vccd1 _1941_ sky130_fd_sc_hd__xnor2_1
X_5818_ _3719_ _0702_ _0692_ vssd1 vssd1 vccd1 vccd1 _0804_ sky130_fd_sc_hd__o21a_1
X_6798_ _3988_ _1664_ vssd1 vssd1 vccd1 vccd1 _1865_ sky130_fd_sc_hd__nor2_1
X_5749_ _0677_ _0707_ _0704_ vssd1 vssd1 vccd1 vccd1 _0731_ sky130_fd_sc_hd__a21boi_1
XANTENNA__5762__C1 _3924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8537_ clknet_3_0__leaf_clk _0023_ vssd1 vssd1 vccd1 vccd1 out_reg\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_41_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8468_ _3668_ vssd1 vssd1 vccd1 vccd1 _0053_ sky130_fd_sc_hd__clkbuf_1
X_7419_ _2223_ _2226_ vssd1 vssd1 vccd1 vccd1 _2548_ sky130_fd_sc_hd__and2_1
X_8399_ _2993_ _3610_ _3611_ vssd1 vssd1 vccd1 vccd1 _3612_ sky130_fd_sc_hd__a21oi_1
XFILLER_89_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6439__B _1423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4406__C _1803_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6190__A _0773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4703__A _3816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_607 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4982_ _4132_ _4135_ vssd1 vssd1 vccd1 vccd1 _4137_ sky130_fd_sc_hd__and2_1
X_7770_ _2928_ _2933_ vssd1 vssd1 vccd1 vccd1 _2934_ sky130_fd_sc_hd__nand2_1
XFILLER_23_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4493__B_N posit_add.in1\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6721_ _1400_ _0548_ vssd1 vssd1 vccd1 vccd1 _1780_ sky130_fd_sc_hd__nor2_1
XFILLER_32_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6652_ _1703_ vssd1 vssd1 vccd1 vccd1 _1705_ sky130_fd_sc_hd__inv_2
X_5603_ _0555_ _0543_ _0510_ vssd1 vssd1 vccd1 vccd1 _0576_ sky130_fd_sc_hd__mux2_1
XFILLER_31_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6583_ _1603_ _1628_ vssd1 vssd1 vccd1 vccd1 _1629_ sky130_fd_sc_hd__xnor2_1
X_8322_ _3416_ _3529_ vssd1 vssd1 vccd1 vccd1 _3531_ sky130_fd_sc_hd__nor2_1
XFILLER_11_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5534_ _0505_ _0506_ _0469_ vssd1 vssd1 vccd1 vccd1 _0507_ sky130_fd_sc_hd__mux2_1
X_8253_ _3455_ _3457_ vssd1 vssd1 vccd1 vccd1 _3458_ sky130_fd_sc_hd__nor2_1
X_5465_ _0425_ _0437_ _0423_ vssd1 vssd1 vccd1 vccd1 _0438_ sky130_fd_sc_hd__a21o_1
XFILLER_117_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4416_ _2122_ _2166_ _2199_ vssd1 vssd1 vccd1 vccd1 _2364_ sky130_fd_sc_hd__o21a_2
X_8184_ _0557_ _3260_ _3306_ vssd1 vssd1 vccd1 vccd1 _3384_ sky130_fd_sc_hd__o21ai_1
X_7204_ _2308_ _2311_ vssd1 vssd1 vccd1 vccd1 _2312_ sky130_fd_sc_hd__or2_1
XFILLER_99_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7135_ _1782_ _2079_ _2225_ vssd1 vssd1 vccd1 vccd1 _2236_ sky130_fd_sc_hd__and3_1
X_5396_ _3729_ _0365_ _0366_ _3736_ _0368_ vssd1 vssd1 vccd1 vccd1 _0369_ sky130_fd_sc_hd__a221oi_4
X_4347_ posit_add.in2\[9\] _1594_ vssd1 vssd1 vccd1 vccd1 _1605_ sky130_fd_sc_hd__xor2_2
XFILLER_113_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7066_ _4126_ _1718_ vssd1 vssd1 vccd1 vccd1 _2160_ sky130_fd_sc_hd__nor2_1
XANTENNA__8461__A1 posit_add.in1\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4278_ in_reg\[0\] in_reg\[1\] _0830_ vssd1 vssd1 vccd1 vccd1 _0862_ sky130_fd_sc_hd__mux2_1
X_6017_ _1014_ vssd1 vssd1 vccd1 vccd1 _1015_ sky130_fd_sc_hd__clkbuf_2
XFILLER_100_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7968_ _3121_ _3151_ _3021_ vssd1 vssd1 vccd1 vccd1 _3152_ sky130_fd_sc_hd__mux2_1
XFILLER_15_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6919_ _1952_ _1996_ vssd1 vssd1 vccd1 vccd1 _1998_ sky130_fd_sc_hd__nor2_1
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7899_ _2965_ _3066_ _2971_ vssd1 vssd1 vccd1 vccd1 _3076_ sky130_fd_sc_hd__mux2_1
XFILLER_52_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5250_ _3988_ _0167_ _0172_ vssd1 vssd1 vccd1 vccd1 _0223_ sky130_fd_sc_hd__o21ba_1
XANTENNA__7494__A2 _1803_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5181_ _0145_ _0151_ _0153_ vssd1 vssd1 vccd1 vccd1 _0154_ sky130_fd_sc_hd__o21ba_1
XFILLER_110_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4608__A _3762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7822_ _2990_ _2659_ _2677_ _2662_ vssd1 vssd1 vccd1 vccd1 _2992_ sky130_fd_sc_hd__o22ai_2
X_4965_ _3832_ _3868_ _3804_ _3893_ vssd1 vssd1 vccd1 vccd1 _4120_ sky130_fd_sc_hd__a22o_1
XFILLER_51_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7753_ _2911_ _2915_ vssd1 vssd1 vccd1 vccd1 _2916_ sky130_fd_sc_hd__or2_1
X_6704_ _1756_ _1757_ vssd1 vssd1 vccd1 vccd1 _1762_ sky130_fd_sc_hd__nand2_1
XFILLER_11_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4896_ _3792_ _3755_ _3959_ _4050_ vssd1 vssd1 vccd1 vccd1 _4051_ sky130_fd_sc_hd__o31a_1
X_7684_ _2836_ _2838_ vssd1 vssd1 vccd1 vccd1 _2840_ sky130_fd_sc_hd__nor2_1
X_6635_ _1400_ _1456_ vssd1 vssd1 vccd1 vccd1 _1686_ sky130_fd_sc_hd__nor2_1
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6566_ _1480_ _1492_ vssd1 vssd1 vccd1 vccd1 _1610_ sky130_fd_sc_hd__and2b_1
X_8305_ _3511_ _3512_ vssd1 vssd1 vccd1 vccd1 _3513_ sky130_fd_sc_hd__nand2_1
X_5517_ _0488_ _0482_ _0337_ vssd1 vssd1 vccd1 vccd1 _0490_ sky130_fd_sc_hd__mux2_1
XFILLER_105_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6497_ _4157_ _1533_ vssd1 vssd1 vccd1 vccd1 _1534_ sky130_fd_sc_hd__nor2_1
X_8236_ _3391_ _3439_ vssd1 vssd1 vccd1 vccd1 _3440_ sky130_fd_sc_hd__and2_1
XFILLER_105_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5448_ _1781_ _0418_ vssd1 vssd1 vccd1 vccd1 _0421_ sky130_fd_sc_hd__nand2_1
XFILLER_87_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5379_ _3079_ _3296_ _3101_ _3046_ vssd1 vssd1 vccd1 vccd1 _0352_ sky130_fd_sc_hd__a211o_1
X_8167_ _3340_ _3364_ vssd1 vssd1 vccd1 vccd1 _3366_ sky130_fd_sc_hd__and2_1
X_7118_ _2206_ _2212_ _2216_ vssd1 vssd1 vccd1 vccd1 _2217_ sky130_fd_sc_hd__o21ai_1
XFILLER_59_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8098_ _3290_ _3291_ _2621_ vssd1 vssd1 vccd1 vccd1 _3292_ sky130_fd_sc_hd__a21oi_1
X_7049_ _2104_ _2140_ vssd1 vssd1 vccd1 vccd1 _2141_ sky130_fd_sc_hd__nand2_1
XANTENNA__6717__B _1537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6733__A _1399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5068__B _3838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5812__A _3763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6627__B _1456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6362__B _1384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5411__A1 _3736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4750_ _3869_ _3904_ vssd1 vssd1 vccd1 vccd1 _3905_ sky130_fd_sc_hd__xnor2_1
XFILLER_61_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4681_ _3783_ _3785_ _3156_ vssd1 vssd1 vccd1 vccd1 _3836_ sky130_fd_sc_hd__a21o_1
X_6420_ _1446_ _1401_ vssd1 vssd1 vccd1 vccd1 _1449_ sky130_fd_sc_hd__nor2_1
X_6351_ _1371_ _1372_ vssd1 vssd1 vccd1 vccd1 _1373_ sky130_fd_sc_hd__nand2_1
X_5302_ _0273_ _0274_ vssd1 vssd1 vccd1 vccd1 _0275_ sky130_fd_sc_hd__or2b_1
X_6282_ _1287_ _1290_ _1293_ _1296_ vssd1 vssd1 vccd1 vccd1 _1298_ sky130_fd_sc_hd__a31o_1
XFILLER_103_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5233_ _0164_ _0205_ vssd1 vssd1 vccd1 vccd1 _0206_ sky130_fd_sc_hd__nor2_1
X_8021_ _3202_ _3207_ vssd1 vssd1 vccd1 vccd1 _3209_ sky130_fd_sc_hd__nand2_1
XFILLER_69_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5164_ _3881_ _3776_ _3838_ _0121_ vssd1 vssd1 vccd1 vccd1 _0137_ sky130_fd_sc_hd__and4_1
XFILLER_69_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5095_ _4210_ vssd1 vssd1 vccd1 vccd1 _4250_ sky130_fd_sc_hd__buf_4
XFILLER_84_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6553__A _1400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7805_ _2962_ _2971_ vssd1 vssd1 vccd1 vccd1 _2973_ sky130_fd_sc_hd__xor2_1
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5997_ _4016_ _0992_ vssd1 vssd1 vccd1 vccd1 _0994_ sky130_fd_sc_hd__nor2_4
XFILLER_12_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4948_ _4078_ _4102_ vssd1 vssd1 vccd1 vccd1 _4103_ sky130_fd_sc_hd__and2_1
X_7736_ _2831_ _2896_ _1286_ vssd1 vssd1 vccd1 vccd1 _2897_ sky130_fd_sc_hd__mux2_1
XFILLER_24_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4879_ _3937_ _3953_ vssd1 vssd1 vccd1 vccd1 _4034_ sky130_fd_sc_hd__or2b_1
X_7667_ _2773_ _2819_ _2820_ vssd1 vssd1 vccd1 vccd1 _2821_ sky130_fd_sc_hd__a21oi_1
X_6618_ _1420_ _1661_ _1666_ vssd1 vssd1 vccd1 vccd1 _1667_ sky130_fd_sc_hd__mux2_1
XANTENNA__4801__A _3735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7598_ _2733_ _2744_ _2708_ vssd1 vssd1 vccd1 vccd1 _2745_ sky130_fd_sc_hd__mux2_1
X_6549_ _1587_ _1590_ vssd1 vssd1 vccd1 vccd1 _1591_ sky130_fd_sc_hd__xor2_1
XFILLER_106_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8219_ _3419_ _3420_ vssd1 vssd1 vccd1 vccd1 _3421_ sky130_fd_sc_hd__nor2_1
XFILLER_58_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8407__B2 _3195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8407__A1 _3608_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6969__A1 _1510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6463__A _1446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5079__A _3988_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4430__B _2507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5920_ _0871_ _0872_ _0870_ vssd1 vssd1 vccd1 vccd1 _0913_ sky130_fd_sc_hd__a21o_1
XFILLER_0_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5851_ _0641_ _0834_ _0835_ vssd1 vssd1 vccd1 vccd1 _0840_ sky130_fd_sc_hd__and3_1
XANTENNA__7385__A1 _0218_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5782_ _0113_ _0762_ vssd1 vssd1 vccd1 vccd1 _0766_ sky130_fd_sc_hd__nand2_1
X_8570_ clknet_3_5__leaf_clk _0056_ vssd1 vssd1 vccd1 vccd1 posit_add.in1\[13\] sky130_fd_sc_hd__dfxtp_2
X_4802_ _3781_ _3790_ vssd1 vssd1 vccd1 vccd1 _3957_ sky130_fd_sc_hd__xnor2_1
XFILLER_21_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4733_ _3862_ _3887_ vssd1 vssd1 vccd1 vccd1 _3888_ sky130_fd_sc_hd__nand2_1
X_7521_ _2654_ _2657_ _0399_ vssd1 vssd1 vccd1 vccd1 _2660_ sky130_fd_sc_hd__a21o_1
XFILLER_119_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7452_ _2514_ _2579_ _2583_ vssd1 vssd1 vccd1 vccd1 _2585_ sky130_fd_sc_hd__o21ai_1
XFILLER_119_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6403_ _1427_ _1430_ vssd1 vssd1 vccd1 vccd1 _1431_ sky130_fd_sc_hd__xor2_1
X_4664_ posit_add.in1\[8\] _2628_ vssd1 vssd1 vccd1 vccd1 _3819_ sky130_fd_sc_hd__xnor2_1
X_4595_ _3167_ _3744_ _3749_ _3594_ vssd1 vssd1 vccd1 vccd1 _3750_ sky130_fd_sc_hd__a211o_4
X_7383_ _2316_ _2317_ _2326_ vssd1 vssd1 vccd1 vccd1 _2509_ sky130_fd_sc_hd__and3_1
X_6334_ _4037_ vssd1 vssd1 vccd1 vccd1 _1355_ sky130_fd_sc_hd__inv_2
XFILLER_115_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6265_ _1268_ _1266_ _1267_ vssd1 vssd1 vccd1 vccd1 _1279_ sky130_fd_sc_hd__and3_1
XFILLER_1_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5216_ _0182_ _0188_ vssd1 vssd1 vccd1 vccd1 _0189_ sky130_fd_sc_hd__xnor2_1
X_8004_ _3184_ _3191_ vssd1 vssd1 vccd1 vccd1 _3192_ sky130_fd_sc_hd__nand2_1
X_6196_ _1017_ _1028_ _1102_ _0706_ vssd1 vssd1 vccd1 vccd1 _1204_ sky130_fd_sc_hd__a22o_1
XFILLER_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5147_ _0118_ _0119_ vssd1 vssd1 vccd1 vccd1 _0120_ sky130_fd_sc_hd__or2_1
XFILLER_28_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5078_ _4228_ _3701_ vssd1 vssd1 vccd1 vccd1 _4233_ sky130_fd_sc_hd__nor2_1
XFILLER_84_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7376__B2 _2416_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7376__A1 _4153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7719_ _2847_ _2876_ _2877_ vssd1 vssd1 vccd1 vccd1 _2878_ sky130_fd_sc_hd__o21ai_1
XFILLER_100_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6730__B _1454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4441__A posit_add.in1\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4380_ _1836_ _1869_ _1891_ _1924_ _1957_ vssd1 vssd1 vccd1 vccd1 _1968_ sky130_fd_sc_hd__a2111o_1
XFILLER_50_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6050_ _1047_ _1048_ vssd1 vssd1 vccd1 vccd1 _1049_ sky130_fd_sc_hd__nor2_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5001_ _3719_ _3817_ vssd1 vssd1 vccd1 vccd1 _4156_ sky130_fd_sc_hd__nor2_1
XFILLER_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6952_ _1384_ _1538_ _1931_ vssd1 vssd1 vccd1 vccd1 _2035_ sky130_fd_sc_hd__o21ai_1
XFILLER_93_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4616__A _3770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5081__A2 _3855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5903_ _2529_ _0676_ vssd1 vssd1 vccd1 vccd1 _0895_ sky130_fd_sc_hd__nor2_1
X_6883_ _1955_ _1956_ vssd1 vssd1 vccd1 vccd1 _1959_ sky130_fd_sc_hd__or2_1
XFILLER_53_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5834_ _3763_ _0676_ vssd1 vssd1 vccd1 vccd1 _0822_ sky130_fd_sc_hd__nor2_1
XFILLER_62_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6030__A1 _0779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5765_ _3865_ _0747_ _0112_ vssd1 vssd1 vccd1 vccd1 _0748_ sky130_fd_sc_hd__a21o_1
X_8553_ clknet_3_0__leaf_clk _0039_ vssd1 vssd1 vccd1 vccd1 counter\[1\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__5447__A _3690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5696_ _3865_ _0670_ _0671_ _0672_ _3801_ vssd1 vssd1 vccd1 vccd1 _0673_ sky130_fd_sc_hd__a311o_1
X_4716_ _3776_ _3838_ vssd1 vssd1 vccd1 vccd1 _3871_ sky130_fd_sc_hd__nand2_1
X_8484_ posit_add.in2\[1\] in_reg\[1\] _3677_ vssd1 vssd1 vccd1 vccd1 _3680_ sky130_fd_sc_hd__mux2_1
X_7504_ _2727_ _1583_ _3919_ _2760_ vssd1 vssd1 vccd1 vccd1 _2642_ sky130_fd_sc_hd__o22ai_1
X_4647_ _3801_ vssd1 vssd1 vccd1 vccd1 _3802_ sky130_fd_sc_hd__buf_4
X_7435_ _2454_ _2424_ _2435_ vssd1 vssd1 vccd1 vccd1 _2566_ sky130_fd_sc_hd__o21ai_1
XFILLER_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7366_ _2382_ _2410_ _2489_ vssd1 vssd1 vccd1 vccd1 _2490_ sky130_fd_sc_hd__o21a_1
X_6317_ _1331_ _1333_ _1335_ vssd1 vssd1 vccd1 vccd1 _1336_ sky130_fd_sc_hd__a21o_1
XFILLER_89_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4578_ _3730_ _3732_ _3690_ vssd1 vssd1 vccd1 vccd1 _3733_ sky130_fd_sc_hd__o21ai_2
XFILLER_1_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7297_ _2259_ _2413_ vssd1 vssd1 vccd1 vccd1 _2414_ sky130_fd_sc_hd__xor2_4
X_6248_ _1228_ _1259_ vssd1 vssd1 vccd1 vccd1 _1260_ sky130_fd_sc_hd__nor2_1
X_6179_ _1132_ _1133_ vssd1 vssd1 vccd1 vccd1 _1185_ sky130_fd_sc_hd__or2_1
XFILLER_103_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5910__A _3770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7597__A1 _3881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4280__A0 in_reg\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6021__A1 _3701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_590 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6635__B _1456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4436__A posit_add.in1\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6651__A _0548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7747__A _1297_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5771__B1 _3802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5550_ _0506_ _0500_ _0510_ vssd1 vssd1 vccd1 vccd1 _0523_ sky130_fd_sc_hd__mux2_1
X_4501_ _2738_ _3275_ _3285_ _3112_ vssd1 vssd1 vccd1 vccd1 _3296_ sky130_fd_sc_hd__o31ai_4
X_5481_ _0447_ _0440_ vssd1 vssd1 vccd1 vccd1 _0454_ sky130_fd_sc_hd__or2_1
X_4432_ _2529_ vssd1 vssd1 vccd1 vccd1 _2540_ sky130_fd_sc_hd__buf_2
X_7220_ _2328_ _0092_ _2323_ _2273_ vssd1 vssd1 vccd1 vccd1 _2329_ sky130_fd_sc_hd__o211a_1
XFILLER_104_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7151_ _2251_ _2252_ vssd1 vssd1 vccd1 vccd1 _2253_ sky130_fd_sc_hd__and2b_2
X_4363_ _1429_ vssd1 vssd1 vccd1 vccd1 _1781_ sky130_fd_sc_hd__clkbuf_4
XFILLER_113_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6102_ _1096_ _1103_ vssd1 vssd1 vccd1 vccd1 _1104_ sky130_fd_sc_hd__or2_1
XFILLER_98_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7082_ _2153_ _2175_ vssd1 vssd1 vccd1 vccd1 _2178_ sky130_fd_sc_hd__xor2_1
X_4294_ in_reg\[8\] in_reg\[9\] _0830_ vssd1 vssd1 vccd1 vccd1 _1030_ sky130_fd_sc_hd__mux2_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6033_ _1015_ _1029_ _1031_ vssd1 vssd1 vccd1 vccd1 _1032_ sky130_fd_sc_hd__a21o_1
XFILLER_86_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7984_ _3042_ _3037_ _3043_ _2999_ _3169_ vssd1 vssd1 vccd1 vccd1 _3170_ sky130_fd_sc_hd__a221o_1
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6935_ _1969_ _2015_ vssd1 vssd1 vccd1 vccd1 _2016_ sky130_fd_sc_hd__xnor2_1
XFILLER_42_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6866_ _1929_ _1938_ _1939_ vssd1 vssd1 vccd1 vccd1 _1940_ sky130_fd_sc_hd__a21oi_1
XFILLER_50_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5817_ _4016_ _0802_ vssd1 vssd1 vccd1 vccd1 _0803_ sky130_fd_sc_hd__or2_2
X_6797_ _1811_ _1816_ vssd1 vssd1 vccd1 vccd1 _1864_ sky130_fd_sc_hd__xnor2_1
XANTENNA__5177__A _3925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5748_ _0727_ _0728_ _0643_ _0710_ vssd1 vssd1 vccd1 vccd1 _0730_ sky130_fd_sc_hd__o211a_1
X_8536_ clknet_3_1__leaf_clk _0022_ vssd1 vssd1 vccd1 vccd1 out_reg\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_41_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5679_ _3718_ _0645_ _0653_ _3699_ vssd1 vssd1 vccd1 vccd1 _0654_ sky130_fd_sc_hd__o31ai_1
X_8467_ in_reg\[10\] posit_add.in1\[10\] _3654_ vssd1 vssd1 vccd1 vccd1 _3668_ sky130_fd_sc_hd__mux2_1
X_7418_ _1531_ _3804_ _1813_ _2546_ vssd1 vssd1 vccd1 vccd1 _2547_ sky130_fd_sc_hd__o22a_1
X_8398_ _3182_ _3596_ vssd1 vssd1 vccd1 vccd1 _3611_ sky130_fd_sc_hd__nand2_1
XFILLER_104_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7349_ _1619_ _2468_ vssd1 vssd1 vccd1 vccd1 _2471_ sky130_fd_sc_hd__xnor2_1
XFILLER_104_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_700 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7567__A _2319_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4703__B _3795_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5753__B1 _3762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8398__A _3182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_619 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4981_ _4132_ _4135_ vssd1 vssd1 vccd1 vccd1 _4136_ sky130_fd_sc_hd__nor2_1
XFILLER_17_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6720_ _1599_ _1676_ vssd1 vssd1 vccd1 vccd1 _1779_ sky130_fd_sc_hd__or2_1
XFILLER_51_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6651_ _0548_ _1537_ vssd1 vssd1 vccd1 vccd1 _1703_ sky130_fd_sc_hd__or2_1
X_6582_ _1624_ _4251_ _1498_ _1626_ vssd1 vssd1 vccd1 vccd1 _1628_ sky130_fd_sc_hd__o31a_1
X_5602_ _0574_ vssd1 vssd1 vccd1 vccd1 _0575_ sky130_fd_sc_hd__inv_2
XFILLER_118_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8321_ _3502_ _3528_ vssd1 vssd1 vccd1 vccd1 _3529_ sky130_fd_sc_hd__xnor2_1
X_5533_ _0504_ _0498_ _0337_ vssd1 vssd1 vccd1 vccd1 _0506_ sky130_fd_sc_hd__mux2_1
XFILLER_117_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8252_ _3440_ _3454_ _3438_ vssd1 vssd1 vccd1 vccd1 _3457_ sky130_fd_sc_hd__o21bai_1
X_5464_ _0433_ _0435_ _0436_ vssd1 vssd1 vccd1 vccd1 _0437_ sky130_fd_sc_hd__o21bai_2
X_4415_ _2331_ _2342_ _1968_ vssd1 vssd1 vccd1 vccd1 _2353_ sky130_fd_sc_hd__mux2_2
X_5395_ _2309_ _3920_ _0367_ vssd1 vssd1 vccd1 vccd1 _0368_ sky130_fd_sc_hd__a21oi_1
X_8183_ _0573_ vssd1 vssd1 vccd1 vccd1 _3383_ sky130_fd_sc_hd__clkinv_2
X_7203_ _2271_ _2288_ _2310_ vssd1 vssd1 vccd1 vccd1 _2311_ sky130_fd_sc_hd__a21oi_1
X_7134_ _2228_ _2229_ _2234_ vssd1 vssd1 vccd1 vccd1 _2235_ sky130_fd_sc_hd__o21ba_1
X_4346_ posit_add.in2\[8\] _1352_ _1374_ _1264_ vssd1 vssd1 vccd1 vccd1 _1594_ sky130_fd_sc_hd__o31a_1
XFILLER_98_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7065_ _1454_ _2158_ vssd1 vssd1 vccd1 vccd1 _2159_ sky130_fd_sc_hd__nand2_1
XANTENNA__6556__A _1353_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4277_ _0841_ vssd1 vssd1 vccd1 vccd1 _0003_ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6016_ _0998_ _1005_ vssd1 vssd1 vccd1 vccd1 _1014_ sky130_fd_sc_hd__and2_1
XFILLER_100_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7967_ _3146_ _3150_ _3006_ vssd1 vssd1 vccd1 vccd1 _3151_ sky130_fd_sc_hd__mux2_1
X_6918_ _1952_ _1996_ vssd1 vssd1 vccd1 vccd1 _1997_ sky130_fd_sc_hd__xor2_1
XFILLER_54_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4804__A _3878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7898_ _3072_ vssd1 vssd1 vccd1 vccd1 _3075_ sky130_fd_sc_hd__clkinv_2
XFILLER_14_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6849_ _1414_ _1782_ _1848_ vssd1 vssd1 vccd1 vccd1 _1921_ sky130_fd_sc_hd__and3_1
XFILLER_50_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4538__A1 _1682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8519_ clknet_3_4__leaf_clk _0005_ vssd1 vssd1 vccd1 vccd1 in_reg\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_108_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4714__A _3866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5180_ _0152_ _3838_ _0113_ vssd1 vssd1 vccd1 vccd1 _0153_ sky130_fd_sc_hd__and3b_1
XFILLER_110_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6376__A _3817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6454__A1 _4217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7821_ _2980_ _0347_ vssd1 vssd1 vccd1 vccd1 _2990_ sky130_fd_sc_hd__nor2_1
XANTENNA__4768__B2 _3729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4964_ _3771_ _3703_ vssd1 vssd1 vccd1 vccd1 _4119_ sky130_fd_sc_hd__or2_1
X_7752_ _2846_ _2913_ vssd1 vssd1 vccd1 vccd1 _2915_ sky130_fd_sc_hd__xnor2_2
XANTENNA__7000__A _1454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6703_ _1746_ _1752_ _1760_ vssd1 vssd1 vccd1 vccd1 _1761_ sky130_fd_sc_hd__a21o_1
XFILLER_51_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4895_ _3722_ _3754_ _3878_ _3868_ _3776_ vssd1 vssd1 vccd1 vccd1 _4050_ sky130_fd_sc_hd__a32o_1
X_7683_ _2836_ _2838_ vssd1 vssd1 vccd1 vccd1 _2839_ sky130_fd_sc_hd__nand2_1
X_6634_ _1684_ _1544_ vssd1 vssd1 vccd1 vccd1 _1685_ sky130_fd_sc_hd__xnor2_1
X_6565_ _1592_ _1608_ vssd1 vssd1 vccd1 vccd1 _1609_ sky130_fd_sc_hd__xnor2_1
XFILLER_20_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6496_ _1446_ _1456_ vssd1 vssd1 vccd1 vccd1 _1533_ sky130_fd_sc_hd__nor2_1
X_8304_ _3460_ _3478_ _3227_ vssd1 vssd1 vccd1 vccd1 _3512_ sky130_fd_sc_hd__a21o_1
X_5516_ _0340_ _0488_ _0337_ vssd1 vssd1 vccd1 vccd1 _0489_ sky130_fd_sc_hd__mux2_1
XFILLER_118_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8235_ _3437_ _3179_ _3438_ vssd1 vssd1 vccd1 vccd1 _3439_ sky130_fd_sc_hd__a21oi_1
X_5447_ _3690_ _0419_ vssd1 vssd1 vccd1 vccd1 _0420_ sky130_fd_sc_hd__xnor2_1
XFILLER_87_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8166_ _3340_ _3364_ vssd1 vssd1 vccd1 vccd1 _3365_ sky130_fd_sc_hd__nor2_1
X_5378_ _0346_ _0350_ vssd1 vssd1 vccd1 vccd1 _0351_ sky130_fd_sc_hd__or2_2
XFILLER_113_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7117_ _2213_ _2215_ vssd1 vssd1 vccd1 vccd1 _2216_ sky130_fd_sc_hd__nand2_1
X_4329_ posit_add.in2\[13\] posit_add.in2\[12\] vssd1 vssd1 vccd1 vccd1 _1407_ sky130_fd_sc_hd__or2_1
X_8097_ _3247_ _3254_ _0601_ vssd1 vssd1 vccd1 vccd1 _3291_ sky130_fd_sc_hd__o21a_1
X_7048_ _2099_ _2103_ vssd1 vssd1 vccd1 vccd1 _2140_ sky130_fd_sc_hd__or2_1
XFILLER_101_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6733__B _1676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8122__A1 _3314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5812__B _3815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7633__A0 _3868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4680_ _3833_ _3834_ _3520_ vssd1 vssd1 vccd1 vccd1 _3835_ sky130_fd_sc_hd__a21o_1
X_6350_ _1370_ _1357_ _1346_ vssd1 vssd1 vccd1 vccd1 _1372_ sky130_fd_sc_hd__or3_1
XFILLER_115_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5301_ _0244_ _0243_ vssd1 vssd1 vccd1 vccd1 _0274_ sky130_fd_sc_hd__xnor2_1
XFILLER_6_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6281_ _1287_ _1293_ _1295_ vssd1 vssd1 vccd1 vccd1 _1296_ sky130_fd_sc_hd__o21a_1
XANTENNA__7490__A posit_add.in1\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4686__B1 _3840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5232_ _0197_ _0202_ _0204_ vssd1 vssd1 vccd1 vccd1 _0205_ sky130_fd_sc_hd__o21ai_1
X_8020_ _3200_ _3207_ vssd1 vssd1 vccd1 vccd1 _3208_ sky130_fd_sc_hd__xnor2_1
X_5163_ _3816_ _4232_ _0124_ vssd1 vssd1 vccd1 vccd1 _0136_ sky130_fd_sc_hd__o21ai_1
XFILLER_96_441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7624__A0 _3883_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5094_ _3701_ _4232_ vssd1 vssd1 vccd1 vccd1 _4249_ sky130_fd_sc_hd__nor2_1
XFILLER_110_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7649__B _2800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7804_ _2962_ _2971_ vssd1 vssd1 vccd1 vccd1 _2972_ sky130_fd_sc_hd__and2b_1
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5996_ _0992_ vssd1 vssd1 vccd1 vccd1 _0993_ sky130_fd_sc_hd__buf_2
X_4947_ _3793_ _3726_ _3959_ vssd1 vssd1 vccd1 vccd1 _4102_ sky130_fd_sc_hd__o21ai_1
X_7735_ _2825_ _2883_ _2827_ vssd1 vssd1 vccd1 vccd1 _2896_ sky130_fd_sc_hd__a21oi_1
XFILLER_33_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4878_ _4031_ _4032_ vssd1 vssd1 vccd1 vccd1 _4033_ sky130_fd_sc_hd__xnor2_2
X_7666_ _2768_ _2769_ vssd1 vssd1 vccd1 vccd1 _2820_ sky130_fd_sc_hd__and2b_1
X_6617_ _1665_ _1511_ vssd1 vssd1 vccd1 vccd1 _1666_ sky130_fd_sc_hd__nand2_1
XANTENNA__5166__A1 _3881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4801__B _3739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7597_ _1355_ _3881_ _2713_ vssd1 vssd1 vccd1 vccd1 _2744_ sky130_fd_sc_hd__mux2_1
X_6548_ _4219_ _1497_ _4213_ _1589_ vssd1 vssd1 vccd1 vccd1 _1590_ sky130_fd_sc_hd__o31a_1
XFILLER_106_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6479_ _0303_ _1423_ vssd1 vssd1 vccd1 vccd1 _1514_ sky130_fd_sc_hd__or2_1
XANTENNA__7604__S _2721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8218_ _3407_ _3417_ vssd1 vssd1 vccd1 vccd1 _3420_ sky130_fd_sc_hd__nor2_1
XFILLER_58_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8149_ out_reg\[3\] _3242_ _1177_ vssd1 vssd1 vccd1 vccd1 _3347_ sky130_fd_sc_hd__a21boi_1
XFILLER_87_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6969__A2 _4126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7091__A1 _4089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6744__A _4232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6463__B _1428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7294__B _0687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5095__A _4210_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7514__S _2652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4439__A posit_add.in1\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7606__A0 _3986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6654__A _4018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5850_ _0825_ _0824_ _0822_ vssd1 vssd1 vccd1 vccd1 _0839_ sky130_fd_sc_hd__a21o_1
X_5781_ _3866_ _0762_ _0716_ _0763_ vssd1 vssd1 vccd1 vccd1 _0764_ sky130_fd_sc_hd__a31o_1
XANTENNA__5396__A1 _3729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5396__B2 _3736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4801_ _3735_ _3739_ _3604_ _3794_ vssd1 vssd1 vccd1 vccd1 _3956_ sky130_fd_sc_hd__or4_1
X_4732_ _3873_ _3886_ vssd1 vssd1 vccd1 vccd1 _3887_ sky130_fd_sc_hd__xnor2_1
X_7520_ _0403_ _0406_ _2652_ vssd1 vssd1 vccd1 vccd1 _2659_ sky130_fd_sc_hd__mux2_2
X_4663_ _3816_ _3817_ vssd1 vssd1 vccd1 vccd1 _3818_ sky130_fd_sc_hd__nor2_1
XFILLER_9_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7451_ _2522_ _2581_ _2582_ _2569_ vssd1 vssd1 vccd1 vccd1 _2583_ sky130_fd_sc_hd__a211o_1
XFILLER_119_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6402_ _1383_ _1428_ vssd1 vssd1 vccd1 vccd1 _1430_ sky130_fd_sc_hd__nor2_1
X_4594_ _3746_ _3748_ _3167_ vssd1 vssd1 vccd1 vccd1 _3749_ sky130_fd_sc_hd__a21oi_1
X_7382_ _2501_ _2506_ _2410_ vssd1 vssd1 vccd1 vccd1 _2508_ sky130_fd_sc_hd__mux2_1
X_6333_ _1351_ _1050_ _1336_ vssd1 vssd1 vccd1 vccd1 _1354_ sky130_fd_sc_hd__nand3_4
XANTENNA__8098__B1 _2621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6264_ _1258_ _1276_ vssd1 vssd1 vccd1 vccd1 _1278_ sky130_fd_sc_hd__xnor2_1
XFILLER_103_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5215_ _0183_ _0187_ _0185_ vssd1 vssd1 vccd1 vccd1 _0188_ sky130_fd_sc_hd__a21oi_1
X_8003_ _3165_ _3181_ _3182_ _3190_ vssd1 vssd1 vccd1 vccd1 _3191_ sky130_fd_sc_hd__o31a_1
X_6195_ _1197_ _1201_ _1202_ vssd1 vssd1 vccd1 vccd1 _1203_ sky130_fd_sc_hd__a21o_1
X_5146_ _0102_ _0117_ vssd1 vssd1 vccd1 vccd1 _0119_ sky130_fd_sc_hd__and2_1
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5077_ _3989_ vssd1 vssd1 vccd1 vccd1 _4232_ sky130_fd_sc_hd__buf_4
XFILLER_56_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5979_ _0881_ _0880_ _0863_ vssd1 vssd1 vccd1 vccd1 _0975_ sky130_fd_sc_hd__a21oi_1
XFILLER_80_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7718_ _2779_ _2780_ vssd1 vssd1 vccd1 vccd1 _2877_ sky130_fd_sc_hd__or2_1
XFILLER_100_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7649_ _2799_ _2800_ vssd1 vssd1 vccd1 vccd1 _2801_ sky130_fd_sc_hd__nor2_1
XFILLER_4_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8089__B1 _3282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_448 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5643__A _2507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4259__A in_reg\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6921__B _1999_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4722__A _3729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5000_ _3998_ _4007_ vssd1 vssd1 vccd1 vccd1 _4155_ sky130_fd_sc_hd__nand2_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6951_ _1931_ _2031_ _2032_ vssd1 vssd1 vccd1 vccd1 _2033_ sky130_fd_sc_hd__and3_1
XFILLER_93_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5902_ _0867_ _0893_ vssd1 vssd1 vccd1 vccd1 _0894_ sky130_fd_sc_hd__nor2_1
X_6882_ _1955_ _1956_ vssd1 vssd1 vccd1 vccd1 _1958_ sky130_fd_sc_hd__xnor2_1
XFILLER_81_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5833_ _0791_ _0820_ vssd1 vssd1 vccd1 vccd1 _0821_ sky130_fd_sc_hd__xnor2_1
XFILLER_22_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8552_ clknet_3_1__leaf_clk _0038_ vssd1 vssd1 vccd1 vccd1 counter\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5764_ _3814_ _2518_ _0365_ vssd1 vssd1 vccd1 vccd1 _0747_ sky130_fd_sc_hd__a21o_1
X_7503_ _2760_ _3919_ _3643_ _2639_ vssd1 vssd1 vccd1 vccd1 _2641_ sky130_fd_sc_hd__o2bb2a_1
X_5695_ _3900_ _4044_ _0647_ _3717_ _3761_ vssd1 vssd1 vccd1 vccd1 _0672_ sky130_fd_sc_hd__o2111a_1
X_8483_ _3679_ vssd1 vssd1 vccd1 vccd1 _0059_ sky130_fd_sc_hd__clkbuf_1
X_4715_ _3771_ _3840_ _3615_ _3793_ vssd1 vssd1 vccd1 vccd1 _3870_ sky130_fd_sc_hd__o22a_1
X_4646_ _3625_ _3684_ _3698_ vssd1 vssd1 vccd1 vccd1 _3801_ sky130_fd_sc_hd__o21a_2
X_7434_ _2451_ _2523_ _2564_ vssd1 vssd1 vccd1 vccd1 _2565_ sky130_fd_sc_hd__a21oi_1
X_4577_ _1880_ _2452_ _3731_ _2397_ vssd1 vssd1 vccd1 vccd1 _3732_ sky130_fd_sc_hd__o211a_1
XANTENNA__5541__A1 _0445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7365_ _2425_ _2426_ _2427_ _2488_ vssd1 vssd1 vccd1 vccd1 _2489_ sky130_fd_sc_hd__a31o_1
X_6316_ _1050_ _1334_ vssd1 vssd1 vccd1 vccd1 _1335_ sky130_fd_sc_hd__nand2_1
XANTENNA__4895__A3 _3878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7296_ _2256_ _2258_ _2000_ vssd1 vssd1 vccd1 vccd1 _2413_ sky130_fd_sc_hd__o21bai_2
XFILLER_1_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6247_ _0722_ _1164_ vssd1 vssd1 vccd1 vccd1 _1259_ sky130_fd_sc_hd__nand2_1
XFILLER_89_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6178_ _1173_ _1182_ _1183_ vssd1 vssd1 vccd1 vccd1 _1184_ sky130_fd_sc_hd__a21oi_1
XFILLER_111_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5129_ _4229_ _4230_ vssd1 vssd1 vccd1 vccd1 _0102_ sky130_fd_sc_hd__xnor2_1
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4280__A1 in_reg\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7853__A _2993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8482__A0 posit_add.in2\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_720 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_672 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6651__B _1537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4452__A posit_add.in1\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4500_ _2650_ _2672_ _2771_ vssd1 vssd1 vccd1 vccd1 _3285_ sky130_fd_sc_hd__nor3_2
XANTENNA__7763__A _1308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5480_ _0449_ _0452_ vssd1 vssd1 vccd1 vccd1 _0453_ sky130_fd_sc_hd__xnor2_1
XFILLER_117_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4431_ _2518_ vssd1 vssd1 vccd1 vccd1 _2529_ sky130_fd_sc_hd__buf_4
XANTENNA__8170__C1 _0600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5283__A _3893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7150_ _2248_ _2249_ _2250_ vssd1 vssd1 vccd1 vccd1 _2252_ sky130_fd_sc_hd__or3_1
X_4362_ posit_add.in2\[0\] posit_add.in2\[1\] vssd1 vssd1 vccd1 vccd1 _1770_ sky130_fd_sc_hd__or2_1
XFILLER_6_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6101_ _1097_ _0996_ _0997_ _1102_ vssd1 vssd1 vccd1 vccd1 _1103_ sky130_fd_sc_hd__and4_1
X_7081_ _3986_ _2079_ vssd1 vssd1 vccd1 vccd1 _2176_ sky130_fd_sc_hd__nand2_1
X_4293_ _1009_ vssd1 vssd1 vccd1 vccd1 _0011_ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6032_ _0773_ _1017_ vssd1 vssd1 vccd1 vccd1 _1031_ sky130_fd_sc_hd__nor2_2
XFILLER_98_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7983_ _2858_ _3168_ vssd1 vssd1 vccd1 vccd1 _3169_ sky130_fd_sc_hd__xnor2_1
XFILLER_39_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6934_ _3615_ _1663_ vssd1 vssd1 vccd1 vccd1 _2015_ sky130_fd_sc_hd__or2_1
XFILLER_54_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6865_ _1928_ _1927_ vssd1 vssd1 vccd1 vccd1 _1939_ sky130_fd_sc_hd__and2b_1
XFILLER_34_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5816_ _0676_ vssd1 vssd1 vccd1 vccd1 _0802_ sky130_fd_sc_hd__buf_2
X_6796_ _1805_ _1820_ vssd1 vssd1 vccd1 vccd1 _1863_ sky130_fd_sc_hd__xnor2_1
XANTENNA__4362__A posit_add.in2\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5747_ _0643_ _0710_ _0727_ _0728_ vssd1 vssd1 vccd1 vccd1 _0729_ sky130_fd_sc_hd__a211oi_1
XANTENNA__5762__A1 _3719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8535_ clknet_3_2__leaf_clk _0021_ vssd1 vssd1 vccd1 vccd1 out_reg\[1\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__5177__B _0105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8466_ _3667_ vssd1 vssd1 vccd1 vccd1 _0052_ sky130_fd_sc_hd__clkbuf_1
XFILLER_108_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5678_ _3813_ _0604_ _0619_ _3761_ vssd1 vssd1 vccd1 vccd1 _0653_ sky130_fd_sc_hd__o211a_1
X_7417_ _1664_ _0548_ vssd1 vssd1 vccd1 vccd1 _2546_ sky130_fd_sc_hd__nor2_1
XANTENNA__5193__A _3893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4629_ _3339_ _3349_ _3189_ _3360_ vssd1 vssd1 vccd1 vccd1 _3784_ sky130_fd_sc_hd__o211a_1
X_8397_ _3609_ _3593_ vssd1 vssd1 vccd1 vccd1 _3610_ sky130_fd_sc_hd__or2_1
X_7348_ _1652_ _2469_ vssd1 vssd1 vccd1 vccd1 _2470_ sky130_fd_sc_hd__xnor2_2
XFILLER_104_666 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7279_ _2362_ _2389_ _2361_ vssd1 vssd1 vccd1 vccd1 _2394_ sky130_fd_sc_hd__o21ba_1
XFILLER_106_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4272__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7258__A1 _2352_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8207__B1 _2621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4980_ _4133_ _4134_ vssd1 vssd1 vccd1 vccd1 _4135_ sky130_fd_sc_hd__xor2_1
XFILLER_16_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6650_ _1691_ _1701_ vssd1 vssd1 vccd1 vccd1 _1702_ sky130_fd_sc_hd__xor2_1
X_6581_ _4235_ _1497_ _1625_ vssd1 vssd1 vccd1 vccd1 _1626_ sky130_fd_sc_hd__a21o_1
X_5601_ _0535_ _0479_ vssd1 vssd1 vccd1 vccd1 _0574_ sky130_fd_sc_hd__nand2_1
XFILLER_118_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8320_ _2604_ _3287_ vssd1 vssd1 vccd1 vccd1 _3528_ sky130_fd_sc_hd__or2_1
X_5532_ _0485_ _0504_ _0338_ vssd1 vssd1 vccd1 vccd1 _0505_ sky130_fd_sc_hd__mux2_1
XANTENNA__7497__A1 _2903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8251_ _3391_ _3439_ _3454_ vssd1 vssd1 vccd1 vccd1 _3455_ sky130_fd_sc_hd__and3_1
X_5463_ _0426_ _0429_ vssd1 vssd1 vccd1 vccd1 _0436_ sky130_fd_sc_hd__and2b_1
XFILLER_105_419 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4414_ _2078_ _2089_ _1869_ _1957_ vssd1 vssd1 vccd1 vccd1 _2342_ sky130_fd_sc_hd__a31oi_1
X_5394_ _1484_ _3830_ _3729_ _3736_ vssd1 vssd1 vccd1 vccd1 _0367_ sky130_fd_sc_hd__a211o_1
X_7202_ _1630_ _1641_ _2286_ vssd1 vssd1 vccd1 vccd1 _2310_ sky130_fd_sc_hd__and3_1
X_8182_ _0601_ _3380_ vssd1 vssd1 vccd1 vccd1 _3382_ sky130_fd_sc_hd__nand2_1
XFILLER_99_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7133_ _2230_ _2233_ vssd1 vssd1 vccd1 vccd1 _2234_ sky130_fd_sc_hd__and2_1
X_4345_ posit_add.in2\[10\] _1572_ vssd1 vssd1 vccd1 vccd1 _1583_ sky130_fd_sc_hd__xnor2_4
XFILLER_98_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7064_ _2156_ _2157_ vssd1 vssd1 vccd1 vccd1 _2158_ sky130_fd_sc_hd__nor2_1
XANTENNA__6556__B _1354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4276_ net3 in_reg\[0\] _0830_ vssd1 vssd1 vccd1 vccd1 _0841_ sky130_fd_sc_hd__mux2_1
X_6015_ _1011_ _1012_ vssd1 vssd1 vccd1 vccd1 _1013_ sky130_fd_sc_hd__nand2_1
XFILLER_67_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7966_ _3011_ _3009_ _2999_ vssd1 vssd1 vccd1 vccd1 _3150_ sky130_fd_sc_hd__mux2_1
XANTENNA__5432__A0 _3729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6917_ _1965_ _1994_ _1995_ vssd1 vssd1 vccd1 vccd1 _1996_ sky130_fd_sc_hd__a21boi_1
XANTENNA__4804__B _3868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7897_ _3073_ vssd1 vssd1 vccd1 vccd1 _3074_ sky130_fd_sc_hd__clkinv_2
X_6848_ _1918_ _1919_ vssd1 vssd1 vccd1 vccd1 _1920_ sky130_fd_sc_hd__xor2_1
XFILLER_52_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4538__A2 _3635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6779_ _1383_ _4126_ vssd1 vssd1 vccd1 vccd1 _1844_ sky130_fd_sc_hd__or2_1
X_8518_ clknet_3_4__leaf_clk _0004_ vssd1 vssd1 vccd1 vccd1 in_reg\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8449_ in_reg\[1\] posit_add.in1\[1\] _3655_ vssd1 vssd1 vccd1 vccd1 _3657_ sky130_fd_sc_hd__mux2_1
XFILLER_2_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4714__B _3868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5826__A _2529_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7820_ _2666_ _2987_ _2988_ vssd1 vssd1 vccd1 vccd1 _2989_ sky130_fd_sc_hd__a21oi_2
XFILLER_91_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4963_ _4106_ _4107_ vssd1 vssd1 vccd1 vccd1 _4118_ sky130_fd_sc_hd__xnor2_1
XFILLER_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7751_ _2912_ _2876_ _1297_ vssd1 vssd1 vccd1 vccd1 _2913_ sky130_fd_sc_hd__mux2_1
XANTENNA__7000__B _1537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6702_ _1754_ _1758_ vssd1 vssd1 vccd1 vccd1 _1760_ sky130_fd_sc_hd__xor2_1
X_7682_ _3925_ _0080_ _2721_ vssd1 vssd1 vccd1 vccd1 _2838_ sky130_fd_sc_hd__mux2_1
X_6633_ _1383_ _1454_ vssd1 vssd1 vccd1 vccd1 _1684_ sky130_fd_sc_hd__or2_1
X_4894_ _3965_ _3978_ vssd1 vssd1 vccd1 vccd1 _4049_ sky130_fd_sc_hd__xnor2_1
XFILLER_20_612 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6564_ _1606_ _1607_ vssd1 vssd1 vccd1 vccd1 _1608_ sky130_fd_sc_hd__xor2_1
X_6495_ _1443_ _1444_ _1531_ vssd1 vssd1 vccd1 vccd1 _1532_ sky130_fd_sc_hd__o21a_1
X_5515_ _0313_ _0322_ vssd1 vssd1 vccd1 vccd1 _0488_ sky130_fd_sc_hd__xor2_1
X_8303_ _3508_ _3510_ vssd1 vssd1 vccd1 vccd1 _3511_ sky130_fd_sc_hd__or2_1
X_5446_ _1781_ _0418_ vssd1 vssd1 vccd1 vccd1 _0419_ sky130_fd_sc_hd__or2_1
X_8234_ _2993_ _3234_ vssd1 vssd1 vccd1 vccd1 _3438_ sky130_fd_sc_hd__and2_1
XFILLER_99_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8165_ _3361_ _3363_ _3259_ vssd1 vssd1 vccd1 vccd1 _3364_ sky130_fd_sc_hd__mux2_1
X_5377_ _0348_ _0349_ vssd1 vssd1 vccd1 vccd1 _0350_ sky130_fd_sc_hd__nor2_2
X_7116_ _2206_ _2214_ vssd1 vssd1 vccd1 vccd1 _2215_ sky130_fd_sc_hd__xnor2_1
X_4328_ posit_add.in2\[11\] posit_add.in2\[9\] posit_add.in2\[8\] posit_add.in2\[10\]
+ vssd1 vssd1 vccd1 vccd1 _1396_ sky130_fd_sc_hd__or4_1
X_8096_ _3284_ _3289_ vssd1 vssd1 vccd1 vccd1 _3290_ sky130_fd_sc_hd__xnor2_2
X_7047_ _2098_ _2124_ _2130_ _2138_ vssd1 vssd1 vccd1 vccd1 _2139_ sky130_fd_sc_hd__a31o_1
XFILLER_74_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4259_ in_reg\[1\] in_reg\[0\] in_reg\[3\] in_reg\[2\] vssd1 vssd1 vccd1 vccd1 _0657_
+ sky130_fd_sc_hd__or4_1
XFILLER_59_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input1_A io_in[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7949_ _3119_ _3130_ _2998_ vssd1 vssd1 vccd1 vccd1 _3131_ sky130_fd_sc_hd__mux2_1
XFILLER_27_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_522 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5812__C _0627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7633__A1 _3893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5300_ _0252_ _0269_ _0272_ vssd1 vssd1 vccd1 vccd1 _0273_ sky130_fd_sc_hd__o21ba_1
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6280_ _1262_ _1294_ vssd1 vssd1 vccd1 vccd1 _1295_ sky130_fd_sc_hd__xnor2_1
XFILLER_6_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4686__A1 _3827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5231_ _0161_ _0203_ vssd1 vssd1 vccd1 vccd1 _0204_ sky130_fd_sc_hd__and2_1
XANTENNA__4686__B2 _3828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5162_ _0120_ _0122_ vssd1 vssd1 vccd1 vccd1 _0135_ sky130_fd_sc_hd__xor2_1
XFILLER_110_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5093_ _4233_ _4237_ vssd1 vssd1 vccd1 vccd1 _4248_ sky130_fd_sc_hd__and2_1
XANTENNA__7624__A1 _3776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6834__B _4153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7803_ _2970_ vssd1 vssd1 vccd1 vccd1 _2971_ sky130_fd_sc_hd__clkbuf_4
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5995_ _0991_ vssd1 vssd1 vccd1 vccd1 _0992_ sky130_fd_sc_hd__buf_2
XFILLER_52_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7734_ _2891_ _2894_ vssd1 vssd1 vccd1 vccd1 _2895_ sky130_fd_sc_hd__or2b_1
X_4946_ _3828_ _3845_ _3930_ _3726_ vssd1 vssd1 vccd1 vccd1 _4101_ sky130_fd_sc_hd__or4_1
XFILLER_52_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4877_ _3935_ _3728_ _3933_ vssd1 vssd1 vccd1 vccd1 _4032_ sky130_fd_sc_hd__o21ba_1
XFILLER_20_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7665_ _2783_ _2817_ _2818_ vssd1 vssd1 vccd1 vccd1 _2819_ sky130_fd_sc_hd__a21boi_1
X_6616_ _4037_ _1664_ vssd1 vssd1 vccd1 vccd1 _1665_ sky130_fd_sc_hd__nor2_2
XANTENNA__5166__A2 _3855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7596_ _2742_ vssd1 vssd1 vccd1 vccd1 _2743_ sky130_fd_sc_hd__clkbuf_4
X_6547_ _1498_ _1447_ _1588_ vssd1 vssd1 vccd1 vccd1 _1589_ sky130_fd_sc_hd__a21o_1
XFILLER_118_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6478_ _1512_ _1424_ vssd1 vssd1 vccd1 vccd1 _1513_ sky130_fd_sc_hd__xnor2_4
XFILLER_106_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5429_ _1946_ vssd1 vssd1 vccd1 vccd1 _0402_ sky130_fd_sc_hd__inv_2
X_8217_ _3418_ vssd1 vssd1 vccd1 vccd1 _3419_ sky130_fd_sc_hd__buf_2
XANTENNA__6728__C _0147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8148_ _3212_ _3325_ _3335_ _3345_ _1177_ vssd1 vssd1 vccd1 vccd1 _3346_ sky130_fd_sc_hd__a2111oi_4
XFILLER_99_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8079_ _3142_ vssd1 vssd1 vccd1 vccd1 _3272_ sky130_fd_sc_hd__clkinv_2
XANTENNA__7620__S _2721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8040__A1 _2993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8451__S _3655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6620__A2_N _1414_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7606__A1 _3901_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4800_ _3807_ _3954_ vssd1 vssd1 vccd1 vccd1 _3955_ sky130_fd_sc_hd__xnor2_1
XFILLER_61_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5780_ _0714_ _0715_ vssd1 vssd1 vccd1 vccd1 _0763_ sky130_fd_sc_hd__nor2_1
XFILLER_61_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4731_ _3856_ _3885_ vssd1 vssd1 vccd1 vccd1 _3886_ sky130_fd_sc_hd__xnor2_1
X_4662_ _3755_ vssd1 vssd1 vccd1 vccd1 _3817_ sky130_fd_sc_hd__buf_4
XFILLER_9_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7450_ _2450_ _2561_ _2563_ vssd1 vssd1 vccd1 vccd1 _2582_ sky130_fd_sc_hd__and3_1
X_6401_ _4037_ vssd1 vssd1 vccd1 vccd1 _1428_ sky130_fd_sc_hd__buf_4
XANTENNA__4356__B1 _1682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4593_ _2969_ _3318_ _3747_ _3488_ vssd1 vssd1 vccd1 vccd1 _3748_ sky130_fd_sc_hd__a211o_2
X_7381_ _4217_ _2431_ _2437_ _2503_ _2505_ vssd1 vssd1 vccd1 vccd1 _2506_ sky130_fd_sc_hd__o221a_1
X_6332_ _1050_ _1336_ _1351_ vssd1 vssd1 vccd1 vccd1 _1353_ sky130_fd_sc_hd__a21o_2
X_6263_ _1258_ _1276_ vssd1 vssd1 vccd1 vccd1 _1277_ sky130_fd_sc_hd__or2_1
XFILLER_89_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5214_ _0185_ _0186_ vssd1 vssd1 vccd1 vccd1 _0187_ sky130_fd_sc_hd__nor2_1
X_8002_ cmd\[7\] cmd\[6\] _3188_ vssd1 vssd1 vccd1 vccd1 _3190_ sky130_fd_sc_hd__nor3_4
X_6194_ _1007_ _1198_ _1101_ vssd1 vssd1 vccd1 vccd1 _1202_ sky130_fd_sc_hd__and3_1
XFILLER_111_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5145_ _0102_ _0117_ vssd1 vssd1 vccd1 vccd1 _0118_ sky130_fd_sc_hd__nor2_1
XFILLER_84_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5076_ _4229_ _4230_ vssd1 vssd1 vccd1 vccd1 _4231_ sky130_fd_sc_hd__and2_1
XFILLER_72_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5978_ _0915_ _0917_ _0964_ _0879_ vssd1 vssd1 vccd1 vccd1 _0974_ sky130_fd_sc_hd__a211o_1
XANTENNA__6580__A _0303_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4929_ _4077_ _4078_ vssd1 vssd1 vccd1 vccd1 _4084_ sky130_fd_sc_hd__xor2_1
X_7717_ _2849_ _2874_ _2875_ vssd1 vssd1 vccd1 vccd1 _2876_ sky130_fd_sc_hd__a21oi_1
XFILLER_40_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4304__S _0819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7648_ _3771_ _3703_ _2713_ vssd1 vssd1 vccd1 vccd1 _2800_ sky130_fd_sc_hd__mux2_1
XFILLER_20_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7579_ _2675_ _2720_ _2722_ vssd1 vssd1 vccd1 vccd1 _2724_ sky130_fd_sc_hd__o21a_1
XFILLER_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4275__A _0819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5834__A _3763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6665__A _0082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6950_ _1401_ _1718_ vssd1 vssd1 vccd1 vccd1 _2032_ sky130_fd_sc_hd__nor2_1
XANTENNA__5066__B2 _1748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5901_ _0634_ _3832_ _0892_ _3735_ vssd1 vssd1 vccd1 vccd1 _0893_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_81_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6881_ _1408_ _1409_ _1531_ vssd1 vssd1 vccd1 vccd1 _1956_ sky130_fd_sc_hd__nand3_1
X_5832_ _0814_ _0818_ vssd1 vssd1 vccd1 vccd1 _0820_ sky130_fd_sc_hd__xnor2_1
XFILLER_34_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5763_ _3866_ _0670_ vssd1 vssd1 vccd1 vccd1 _0746_ sky130_fd_sc_hd__nor2_1
X_8551_ clknet_3_0__leaf_clk _0037_ vssd1 vssd1 vccd1 vccd1 mode sky130_fd_sc_hd__dfxtp_1
X_4714_ _3866_ _3868_ vssd1 vssd1 vccd1 vccd1 _3869_ sky130_fd_sc_hd__nand2_1
X_7502_ _2626_ _1682_ _3643_ _2639_ _2638_ vssd1 vssd1 vccd1 vccd1 _2640_ sky130_fd_sc_hd__a221o_1
X_5694_ _0616_ _0609_ _3717_ vssd1 vssd1 vccd1 vccd1 _0671_ sky130_fd_sc_hd__a21o_1
X_8482_ posit_add.in2\[0\] in_reg\[0\] _3677_ vssd1 vssd1 vccd1 vccd1 _3679_ sky130_fd_sc_hd__mux2_1
X_4645_ _3719_ vssd1 vssd1 vccd1 vccd1 _3800_ sky130_fd_sc_hd__clkbuf_4
X_7433_ _2494_ _2561_ _2563_ vssd1 vssd1 vccd1 vccd1 _2564_ sky130_fd_sc_hd__and3_1
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4576_ _2012_ _2111_ _2210_ _2375_ vssd1 vssd1 vccd1 vccd1 _3731_ sky130_fd_sc_hd__a211o_1
X_7364_ _2343_ _0442_ vssd1 vssd1 vccd1 vccd1 _2488_ sky130_fd_sc_hd__xor2_2
X_6315_ _1049_ _1035_ _1037_ vssd1 vssd1 vccd1 vccd1 _1334_ sky130_fd_sc_hd__or3_1
XANTENNA__7154__A_N _1999_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7295_ _2411_ vssd1 vssd1 vccd1 vccd1 _2412_ sky130_fd_sc_hd__buf_4
X_6246_ _1237_ _1249_ vssd1 vssd1 vccd1 vccd1 _1258_ sky130_fd_sc_hd__xnor2_1
XFILLER_39_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6177_ _1180_ _1181_ vssd1 vssd1 vccd1 vccd1 _1183_ sky130_fd_sc_hd__and2b_1
XFILLER_85_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8243__A1 _3445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5128_ _0079_ _0100_ vssd1 vssd1 vccd1 vccd1 _0101_ sky130_fd_sc_hd__and2_1
XANTENNA__6254__B1 _1128_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5059_ _4213_ _4212_ vssd1 vssd1 vccd1 vccd1 _4214_ sky130_fd_sc_hd__xnor2_1
XFILLER_55_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_695 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4568__B1 _3232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5548__B _0467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4430_ _1748_ _2507_ vssd1 vssd1 vccd1 vccd1 _2518_ sky130_fd_sc_hd__nand2_1
XFILLER_6_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6100_ _1101_ vssd1 vssd1 vccd1 vccd1 _1102_ sky130_fd_sc_hd__buf_2
X_4361_ _1638_ _1715_ vssd1 vssd1 vccd1 vccd1 _1759_ sky130_fd_sc_hd__nand2_1
XFILLER_112_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7080_ _2170_ _2174_ vssd1 vssd1 vccd1 vccd1 _2175_ sky130_fd_sc_hd__and2_1
X_4292_ in_reg\[7\] in_reg\[8\] _0830_ vssd1 vssd1 vccd1 vccd1 _1009_ sky130_fd_sc_hd__mux2_1
XANTENNA__8473__A1 posit_add.in1\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6031_ _1017_ _1028_ _1008_ vssd1 vssd1 vccd1 vccd1 _1029_ sky130_fd_sc_hd__mux2_2
XFILLER_100_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7982_ _3166_ _2860_ vssd1 vssd1 vccd1 vccd1 _3168_ sky130_fd_sc_hd__nor2_1
XFILLER_26_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6933_ _1300_ _3986_ _1809_ vssd1 vssd1 vccd1 vccd1 _2014_ sky130_fd_sc_hd__and3_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6864_ _1932_ _1937_ vssd1 vssd1 vccd1 vccd1 _1938_ sky130_fd_sc_hd__xnor2_1
XFILLER_81_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5815_ _0793_ _0800_ vssd1 vssd1 vccd1 vccd1 _0801_ sky130_fd_sc_hd__xnor2_1
XFILLER_34_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6795_ _1822_ _1824_ vssd1 vssd1 vccd1 vccd1 _1862_ sky130_fd_sc_hd__xnor2_1
X_5746_ _0725_ _0726_ _0719_ vssd1 vssd1 vccd1 vccd1 _0728_ sky130_fd_sc_hd__a21oi_1
X_8534_ clknet_3_2__leaf_clk _0020_ vssd1 vssd1 vccd1 vccd1 out_reg\[0\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__5177__C _3795_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5677_ _0112_ _0645_ _0649_ _0650_ _0651_ vssd1 vssd1 vccd1 vccd1 _0652_ sky130_fd_sc_hd__o32a_1
X_8465_ in_reg\[9\] posit_add.in1\[9\] _3655_ vssd1 vssd1 vccd1 vccd1 _3667_ sky130_fd_sc_hd__mux2_1
X_7416_ _2230_ _2544_ _2234_ vssd1 vssd1 vccd1 vccd1 _2545_ sky130_fd_sc_hd__o21ba_1
X_4628_ _2936_ _3307_ _3467_ _3435_ vssd1 vssd1 vccd1 vccd1 _3783_ sky130_fd_sc_hd__a211o_1
XANTENNA__5193__B _0121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8396_ _3560_ vssd1 vssd1 vccd1 vccd1 _3609_ sky130_fd_sc_hd__clkinv_2
X_4559_ _1726_ _2353_ _2364_ _1836_ vssd1 vssd1 vccd1 vccd1 _3714_ sky130_fd_sc_hd__o211a_1
X_7347_ _1619_ _2468_ _2266_ vssd1 vssd1 vccd1 vccd1 _2469_ sky130_fd_sc_hd__o21a_1
XFILLER_1_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7278_ _2385_ _2388_ _2390_ _2392_ vssd1 vssd1 vccd1 vccd1 _2393_ sky130_fd_sc_hd__o31a_2
XFILLER_104_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6229_ _0706_ _1127_ vssd1 vssd1 vccd1 vccd1 _1239_ sky130_fd_sc_hd__and2_1
XFILLER_106_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_607 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7727__B1 _2838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7864__A _2941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5384__A _3736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6662__B _1711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6580_ _0303_ _1446_ vssd1 vssd1 vccd1 vccd1 _1625_ sky130_fd_sc_hd__nor2_1
X_5600_ _0571_ _0572_ _0557_ vssd1 vssd1 vccd1 vccd1 _0573_ sky130_fd_sc_hd__mux2_1
XFILLER_31_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5531_ _0208_ _0327_ vssd1 vssd1 vccd1 vccd1 _0504_ sky130_fd_sc_hd__xnor2_1
XFILLER_117_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8250_ _3234_ _3164_ vssd1 vssd1 vccd1 vccd1 _3454_ sky130_fd_sc_hd__or2_1
XANTENNA__7497__A2 _1858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5462_ _0434_ _0396_ _0350_ vssd1 vssd1 vccd1 vccd1 _0435_ sky130_fd_sc_hd__a21oi_4
X_7201_ _2306_ _2307_ vssd1 vssd1 vccd1 vccd1 _2308_ sky130_fd_sc_hd__nand2_1
X_4413_ _1814_ _2034_ _2045_ _2056_ vssd1 vssd1 vccd1 vccd1 _2331_ sky130_fd_sc_hd__o22ai_1
X_5393_ _1748_ _3706_ _3708_ vssd1 vssd1 vccd1 vccd1 _0366_ sky130_fd_sc_hd__and3_1
X_8181_ _3359_ _3367_ vssd1 vssd1 vccd1 vccd1 _3380_ sky130_fd_sc_hd__or2_1
X_7132_ _3804_ _2079_ _2185_ _2231_ vssd1 vssd1 vccd1 vccd1 _2233_ sky130_fd_sc_hd__and4_1
X_4344_ posit_add.in2\[9\] posit_add.in2\[8\] _1352_ _1374_ _1264_ vssd1 vssd1 vccd1
+ vccd1 _1572_ sky130_fd_sc_hd__o41a_2
XFILLER_113_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7063_ _1531_ _1813_ vssd1 vssd1 vccd1 vccd1 _2157_ sky130_fd_sc_hd__nand2_1
X_6014_ _0998_ _1005_ _1006_ _1010_ vssd1 vssd1 vccd1 vccd1 _1012_ sky130_fd_sc_hd__a22o_1
XFILLER_98_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4275_ _0819_ vssd1 vssd1 vccd1 vccd1 _0830_ sky130_fd_sc_hd__buf_4
XANTENNA__4638__A _3792_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7965_ _3124_ _3135_ _3143_ _3148_ vssd1 vssd1 vccd1 vccd1 _3149_ sky130_fd_sc_hd__or4_1
X_6916_ _1993_ _1992_ vssd1 vssd1 vccd1 vccd1 _1995_ sky130_fd_sc_hd__or2b_1
XFILLER_42_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7896_ _3062_ _3072_ _2842_ vssd1 vssd1 vccd1 vccd1 _3073_ sky130_fd_sc_hd__mux2_1
XFILLER_23_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6847_ _1872_ _1874_ vssd1 vssd1 vccd1 vccd1 _1919_ sky130_fd_sc_hd__xor2_1
XFILLER_23_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6778_ _1776_ _1842_ vssd1 vssd1 vccd1 vccd1 _1843_ sky130_fd_sc_hd__or2_1
X_5729_ _0704_ _0707_ _0677_ vssd1 vssd1 vccd1 vccd1 _0709_ sky130_fd_sc_hd__a21o_1
X_8517_ clknet_3_1__leaf_clk _0003_ vssd1 vssd1 vccd1 vccd1 in_reg\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_10_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8448_ _3656_ vssd1 vssd1 vccd1 vccd1 _0043_ sky130_fd_sc_hd__clkbuf_1
X_8379_ _3588_ _3589_ vssd1 vssd1 vccd1 vccd1 _3591_ sky130_fd_sc_hd__nand2_1
XANTENNA__5932__A _2529_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4548__A _3702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4631__C1 _2969_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4433__D posit_add.in1\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5842__A _0627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6673__A _4157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4962_ _4104_ _4116_ vssd1 vssd1 vccd1 vccd1 _4117_ sky130_fd_sc_hd__xnor2_2
X_7750_ _2817_ vssd1 vssd1 vccd1 vccd1 _2912_ sky130_fd_sc_hd__clkinv_2
X_4893_ _3963_ _3981_ vssd1 vssd1 vccd1 vccd1 _4048_ sky130_fd_sc_hd__xor2_2
X_6701_ _1756_ _1757_ vssd1 vssd1 vccd1 vccd1 _1758_ sky130_fd_sc_hd__xnor2_1
X_7681_ _2743_ _2797_ vssd1 vssd1 vccd1 vccd1 _2836_ sky130_fd_sc_hd__nand2_1
XFILLER_32_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6632_ _1655_ _1668_ _1672_ _1669_ vssd1 vssd1 vccd1 vccd1 _1683_ sky130_fd_sc_hd__o22ai_2
XANTENNA__8364__B1 _2621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6563_ _1463_ _1479_ vssd1 vssd1 vccd1 vccd1 _1607_ sky130_fd_sc_hd__nand2_1
XANTENNA__8116__B1 _0600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6494_ _3907_ vssd1 vssd1 vccd1 vccd1 _1531_ sky130_fd_sc_hd__buf_4
X_8302_ _3437_ _3273_ _3475_ _3438_ vssd1 vssd1 vccd1 vccd1 _3510_ sky130_fd_sc_hd__a31o_1
X_5514_ _0484_ _0486_ _0470_ vssd1 vssd1 vccd1 vccd1 _0487_ sky130_fd_sc_hd__mux2_1
XFILLER_118_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8233_ _3234_ vssd1 vssd1 vccd1 vccd1 _3437_ sky130_fd_sc_hd__inv_2
X_5445_ _3830_ _3635_ vssd1 vssd1 vccd1 vccd1 _0418_ sky130_fd_sc_hd__nand2_1
X_8164_ _3362_ vssd1 vssd1 vccd1 vccd1 _3363_ sky130_fd_sc_hd__inv_2
X_7115_ _2207_ _2211_ vssd1 vssd1 vccd1 vccd1 _2214_ sky130_fd_sc_hd__and2_1
XFILLER_59_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5376_ _0343_ _0344_ vssd1 vssd1 vccd1 vccd1 _0349_ sky130_fd_sc_hd__and2_1
XFILLER_113_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4327_ _1352_ _1374_ vssd1 vssd1 vccd1 vccd1 _1385_ sky130_fd_sc_hd__nor2_1
XFILLER_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8095_ _2585_ _3288_ _2604_ vssd1 vssd1 vccd1 vccd1 _3289_ sky130_fd_sc_hd__mux2_2
XFILLER_113_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7046_ _2131_ _2132_ _2137_ vssd1 vssd1 vccd1 vccd1 _2138_ sky130_fd_sc_hd__and3_1
XFILLER_101_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4258_ in_reg\[5\] in_reg\[4\] in_reg\[7\] in_reg\[6\] vssd1 vssd1 vccd1 vccd1 _0646_
+ sky130_fd_sc_hd__or4_1
XFILLER_74_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7948_ _3118_ _3129_ _2842_ vssd1 vssd1 vccd1 vccd1 _3130_ sky130_fd_sc_hd__mux2_1
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7879_ _3053_ _3039_ _2954_ vssd1 vssd1 vccd1 vccd1 _3054_ sky130_fd_sc_hd__mux2_1
XFILLER_10_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8022__B _2319_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_534 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8449__S _3655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5837__A _3815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4741__A _3893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5230_ _0159_ _0160_ vssd1 vssd1 vccd1 vccd1 _0203_ sky130_fd_sc_hd__nand2_1
XANTENNA__4686__A2 _3739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5161_ _0118_ _0130_ vssd1 vssd1 vccd1 vccd1 _0134_ sky130_fd_sc_hd__xnor2_1
XFILLER_69_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5092_ _4240_ _4243_ vssd1 vssd1 vccd1 vccd1 _4247_ sky130_fd_sc_hd__nand2_1
XFILLER_110_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5994_ _0821_ _0990_ vssd1 vssd1 vccd1 vccd1 _0991_ sky130_fd_sc_hd__xnor2_1
XFILLER_64_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7802_ _2964_ _2968_ _2918_ vssd1 vssd1 vccd1 vccd1 _2970_ sky130_fd_sc_hd__mux2_1
XFILLER_25_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4945_ _4080_ _4086_ vssd1 vssd1 vccd1 vccd1 _4100_ sky130_fd_sc_hd__xnor2_1
X_7733_ _2844_ _2893_ vssd1 vssd1 vccd1 vccd1 _2894_ sky130_fd_sc_hd__xnor2_1
XFILLER_24_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4876_ _4028_ _4030_ vssd1 vssd1 vccd1 vccd1 _4031_ sky130_fd_sc_hd__xnor2_2
XFILLER_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7664_ _2779_ _2781_ vssd1 vssd1 vccd1 vccd1 _2818_ sky130_fd_sc_hd__or2_1
XFILLER_32_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6615_ _1663_ vssd1 vssd1 vccd1 vccd1 _1664_ sky130_fd_sc_hd__buf_2
X_7595_ _2729_ _2702_ vssd1 vssd1 vccd1 vccd1 _2742_ sky130_fd_sc_hd__and2_1
X_6546_ _1420_ _1446_ vssd1 vssd1 vccd1 vccd1 _1588_ sky130_fd_sc_hd__nor2_1
X_6477_ _1416_ _1417_ vssd1 vssd1 vccd1 vccd1 _1512_ sky130_fd_sc_hd__xor2_2
X_8216_ _3289_ _3406_ _3417_ _3284_ vssd1 vssd1 vccd1 vccd1 _3418_ sky130_fd_sc_hd__and4b_1
X_5428_ _3328_ _0121_ _0400_ vssd1 vssd1 vccd1 vccd1 _0401_ sky130_fd_sc_hd__a21oi_1
XFILLER_114_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8147_ _3166_ _3336_ _3342_ _3344_ vssd1 vssd1 vccd1 vccd1 _3345_ sky130_fd_sc_hd__o31a_1
X_5359_ _0079_ _0132_ _0089_ vssd1 vssd1 vccd1 vccd1 _0332_ sky130_fd_sc_hd__a21oi_1
XFILLER_59_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8078_ _3228_ _3238_ vssd1 vssd1 vccd1 vccd1 _3271_ sky130_fd_sc_hd__and2_1
XFILLER_101_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7029_ _2112_ _2115_ _2117_ vssd1 vssd1 vccd1 vccd1 _2119_ sky130_fd_sc_hd__and3_1
XFILLER_114_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4730_ _3880_ _3884_ vssd1 vssd1 vccd1 vccd1 _3885_ sky130_fd_sc_hd__xnor2_1
XFILLER_9_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4661_ _3815_ vssd1 vssd1 vccd1 vccd1 _3816_ sky130_fd_sc_hd__clkbuf_4
XFILLER_9_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6400_ _1353_ _1354_ _4153_ vssd1 vssd1 vccd1 vccd1 _1427_ sky130_fd_sc_hd__and3_1
X_7380_ _2499_ _2504_ _2330_ vssd1 vssd1 vccd1 vccd1 _2505_ sky130_fd_sc_hd__or3b_1
X_6331_ _1349_ _1350_ vssd1 vssd1 vccd1 vccd1 _1351_ sky130_fd_sc_hd__or2_1
X_4592_ _3339_ _3349_ _3232_ _3360_ vssd1 vssd1 vccd1 vccd1 _3747_ sky130_fd_sc_hd__o211a_1
XFILLER_115_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6262_ _1260_ _1273_ _1274_ vssd1 vssd1 vccd1 vccd1 _1276_ sky130_fd_sc_hd__a21oi_1
XFILLER_89_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6193_ _1198_ _1200_ vssd1 vssd1 vccd1 vccd1 _1201_ sky130_fd_sc_hd__xnor2_1
X_5213_ _4222_ _3883_ _0184_ vssd1 vssd1 vccd1 vccd1 _0186_ sky130_fd_sc_hd__a21oi_1
XFILLER_69_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8001_ _3042_ _3138_ _3187_ vssd1 vssd1 vccd1 vccd1 _3188_ sky130_fd_sc_hd__o21ai_2
X_5144_ _0104_ _0110_ _0114_ _0116_ vssd1 vssd1 vccd1 vccd1 _0117_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_111_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5075_ _4226_ _4216_ vssd1 vssd1 vccd1 vccd1 _4230_ sky130_fd_sc_hd__xnor2_1
XANTENNA__4292__A0 in_reg\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5977_ _0971_ _0972_ vssd1 vssd1 vccd1 vccd1 _0973_ sky130_fd_sc_hd__or2_2
XANTENNA__6580__B _1446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4928_ _4052_ _4082_ vssd1 vssd1 vccd1 vccd1 _4083_ sky130_fd_sc_hd__or2_1
X_7716_ _2788_ _2789_ vssd1 vssd1 vccd1 vccd1 _2875_ sky130_fd_sc_hd__and2b_1
X_7647_ _2796_ _2798_ vssd1 vssd1 vccd1 vccd1 _2799_ sky130_fd_sc_hd__nand2_1
X_4859_ _3856_ _3885_ _4013_ vssd1 vssd1 vccd1 vccd1 _4014_ sky130_fd_sc_hd__a21o_1
XFILLER_119_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_0__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_20_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7578_ _2675_ _2720_ _2722_ vssd1 vssd1 vccd1 vccd1 _2723_ sky130_fd_sc_hd__or3_1
XFILLER_69_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6529_ _1566_ _1567_ vssd1 vssd1 vccd1 vccd1 _1569_ sky130_fd_sc_hd__nand2_1
XANTENNA__6101__A _1097_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4259__C in_reg\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5387__A _3830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6011__A _4017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6665__B _1718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4510__A1 _2969_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5900_ _0762_ vssd1 vssd1 vccd1 vccd1 _0892_ sky130_fd_sc_hd__clkinv_2
XFILLER_81_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6880_ _1413_ _1782_ vssd1 vssd1 vccd1 vccd1 _1955_ sky130_fd_sc_hd__nand2_1
XFILLER_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5831_ _0815_ _0817_ vssd1 vssd1 vccd1 vccd1 _0818_ sky130_fd_sc_hd__xnor2_1
XFILLER_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5762_ _3719_ _0740_ _0743_ _3924_ vssd1 vssd1 vccd1 vccd1 _0745_ sky130_fd_sc_hd__a211o_1
X_8550_ clknet_3_1__leaf_clk _0036_ vssd1 vssd1 vccd1 vccd1 io_out[3] sky130_fd_sc_hd__dfxtp_2
XFILLER_61_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7501_ _2626_ _1682_ _2627_ _2637_ vssd1 vssd1 vccd1 vccd1 _2638_ sky130_fd_sc_hd__o22a_1
X_4713_ _3867_ vssd1 vssd1 vccd1 vccd1 _3868_ sky130_fd_sc_hd__clkbuf_4
X_5693_ _0365_ _3791_ _3813_ vssd1 vssd1 vccd1 vccd1 _0670_ sky130_fd_sc_hd__mux2_1
X_8481_ _3676_ vssd1 vssd1 vccd1 vccd1 _3677_ sky130_fd_sc_hd__clkbuf_4
X_4644_ _3756_ _3779_ _3798_ vssd1 vssd1 vccd1 vccd1 _3799_ sky130_fd_sc_hd__a21o_1
X_7432_ _2379_ _2396_ _2407_ _2434_ vssd1 vssd1 vccd1 vccd1 _2563_ sky130_fd_sc_hd__or4_1
X_4575_ _2430_ _2441_ _2463_ _2298_ vssd1 vssd1 vccd1 vccd1 _3730_ sky130_fd_sc_hd__o211a_1
X_7363_ _2453_ _2480_ _2486_ vssd1 vssd1 vccd1 vccd1 _2487_ sky130_fd_sc_hd__mux2_1
XFILLER_116_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6314_ _1332_ _1327_ _1321_ vssd1 vssd1 vccd1 vccd1 _1333_ sky130_fd_sc_hd__o21bai_1
XFILLER_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7294_ _0698_ _0687_ _2332_ vssd1 vssd1 vccd1 vccd1 _2411_ sky130_fd_sc_hd__and3b_1
XANTENNA__8341__A1_N _3534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6245_ _1227_ _1256_ vssd1 vssd1 vccd1 vccd1 _1257_ sky130_fd_sc_hd__xnor2_1
XFILLER_103_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6176_ _1180_ _1181_ vssd1 vssd1 vccd1 vccd1 _1182_ sky130_fd_sc_hd__xnor2_1
XFILLER_69_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5127_ _4246_ _0078_ vssd1 vssd1 vccd1 vccd1 _0100_ sky130_fd_sc_hd__or2_1
XFILLER_84_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5058_ _4210_ _3615_ vssd1 vssd1 vccd1 vccd1 _4213_ sky130_fd_sc_hd__nor2_1
XFILLER_72_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8457__S _3655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6006__A _4210_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8170__A1 _1330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4360_ _1737_ vssd1 vssd1 vccd1 vccd1 _1748_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__4313__B_N _0701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4291_ _0988_ vssd1 vssd1 vccd1 vccd1 _0010_ sky130_fd_sc_hd__clkbuf_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6030_ _0779_ _0803_ _0992_ vssd1 vssd1 vccd1 vccd1 _1028_ sky130_fd_sc_hd__a21oi_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7984__B2 _2999_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7981_ _2929_ vssd1 vssd1 vccd1 vccd1 _3166_ sky130_fd_sc_hd__buf_2
X_6932_ _1967_ _1971_ vssd1 vssd1 vccd1 vccd1 _2013_ sky130_fd_sc_hd__xnor2_1
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6842__C _1782_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6863_ _1933_ _1936_ vssd1 vssd1 vccd1 vccd1 _1937_ sky130_fd_sc_hd__xnor2_1
X_5814_ _0794_ _0799_ vssd1 vssd1 vccd1 vccd1 _0800_ sky130_fd_sc_hd__xnor2_1
XFILLER_62_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_611 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6794_ _1843_ _1860_ vssd1 vssd1 vccd1 vccd1 _1861_ sky130_fd_sc_hd__xnor2_1
XFILLER_22_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5745_ _0719_ _0725_ _0726_ vssd1 vssd1 vccd1 vccd1 _0727_ sky130_fd_sc_hd__and3_1
X_8533_ clknet_3_0__leaf_clk _0019_ vssd1 vssd1 vccd1 vccd1 last_SCLK sky130_fd_sc_hd__dfxtp_1
X_5676_ _3900_ _0609_ vssd1 vssd1 vccd1 vccd1 _0651_ sky130_fd_sc_hd__nor2_1
X_8464_ _3666_ vssd1 vssd1 vccd1 vccd1 _0051_ sky130_fd_sc_hd__clkbuf_1
XFILLER_108_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7415_ _2185_ _2543_ _2231_ _2079_ _3804_ vssd1 vssd1 vccd1 vccd1 _2544_ sky130_fd_sc_hd__a32o_1
X_4627_ _3167_ _3509_ _3771_ _3573_ _3594_ vssd1 vssd1 vccd1 vccd1 _3782_ sky130_fd_sc_hd__a2111o_2
X_8395_ _3606_ _3607_ vssd1 vssd1 vccd1 vccd1 _3608_ sky130_fd_sc_hd__or2_1
XFILLER_104_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4558_ _1803_ _2221_ _3712_ _2408_ vssd1 vssd1 vccd1 vccd1 _3713_ sky130_fd_sc_hd__a211o_1
X_7346_ _1771_ _2456_ _2264_ vssd1 vssd1 vccd1 vccd1 _2468_ sky130_fd_sc_hd__a21boi_1
XFILLER_89_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4489_ _3156_ vssd1 vssd1 vccd1 vccd1 _3167_ sky130_fd_sc_hd__buf_4
XFILLER_9_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7277_ _2349_ _2391_ vssd1 vssd1 vccd1 vccd1 _2392_ sky130_fd_sc_hd__nand2_2
X_6228_ _1232_ _1233_ vssd1 vssd1 vccd1 vccd1 _1238_ sky130_fd_sc_hd__xnor2_1
X_6159_ _1089_ vssd1 vssd1 vccd1 vccd1 _1164_ sky130_fd_sc_hd__clkbuf_4
XFILLER_106_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_619 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4834__A posit_add.in1\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4562__A1_N _3690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5665__A _0627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7880__A _2941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6496__A _1446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5575__A _4126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7294__A_N _0698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5530_ _0500_ _0502_ _0470_ vssd1 vssd1 vccd1 vccd1 _0503_ sky130_fd_sc_hd__mux2_1
X_5461_ _0348_ _0349_ vssd1 vssd1 vccd1 vccd1 _0434_ sky130_fd_sc_hd__nand2_1
X_4412_ _1913_ _2221_ _2232_ _2309_ vssd1 vssd1 vccd1 vccd1 _2320_ sky130_fd_sc_hd__a211o_1
XANTENNA__7790__A _2954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7200_ _2279_ _2282_ _2305_ vssd1 vssd1 vccd1 vccd1 _2307_ sky130_fd_sc_hd__or3_1
X_5392_ _3690_ _3716_ _3774_ vssd1 vssd1 vccd1 vccd1 _0365_ sky130_fd_sc_hd__a21oi_4
X_8180_ _3378_ _3379_ _0635_ vssd1 vssd1 vccd1 vccd1 _0025_ sky130_fd_sc_hd__a21oi_1
XFILLER_99_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7131_ _1664_ _1676_ _2125_ vssd1 vssd1 vccd1 vccd1 _2231_ sky130_fd_sc_hd__o21ai_1
X_4343_ _1495_ _1517_ _1550_ vssd1 vssd1 vccd1 vccd1 _1561_ sky130_fd_sc_hd__a21oi_4
XANTENNA__4919__A _3892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7062_ _1664_ _1456_ vssd1 vssd1 vccd1 vccd1 _2156_ sky130_fd_sc_hd__or2_1
XFILLER_86_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4274_ _0808_ vssd1 vssd1 vccd1 vccd1 _0819_ sky130_fd_sc_hd__clkbuf_4
XFILLER_101_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6013_ _0998_ _1005_ _1006_ _1010_ vssd1 vssd1 vccd1 vccd1 _1011_ sky130_fd_sc_hd__nand4_1
XFILLER_98_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7964_ _3144_ _3147_ _3021_ vssd1 vssd1 vccd1 vccd1 _3148_ sky130_fd_sc_hd__mux2_1
XFILLER_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6915_ _1992_ _1993_ vssd1 vssd1 vccd1 vccd1 _1994_ sky130_fd_sc_hd__xnor2_1
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7895_ _3070_ _3071_ _3038_ vssd1 vssd1 vccd1 vccd1 _3072_ sky130_fd_sc_hd__mux2_1
XFILLER_35_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6846_ _1911_ _1916_ _1917_ vssd1 vssd1 vccd1 vccd1 _1918_ sky130_fd_sc_hd__a21o_1
XFILLER_52_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6777_ _1420_ _1718_ vssd1 vssd1 vccd1 vccd1 _1842_ sky130_fd_sc_hd__or2_1
XFILLER_22_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7684__B _2838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5728_ _0677_ _0704_ _0707_ vssd1 vssd1 vccd1 vccd1 _0708_ sky130_fd_sc_hd__nand3_1
X_8516_ clknet_3_6__leaf_clk _0002_ vssd1 vssd1 vccd1 vccd1 cmd\[7\] sky130_fd_sc_hd__dfxtp_4
XFILLER_50_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5659_ _3792_ _0627_ _3735_ _0631_ vssd1 vssd1 vccd1 vccd1 _0632_ sky130_fd_sc_hd__or4b_1
X_8447_ in_reg\[0\] _2969_ _3655_ vssd1 vssd1 vccd1 vccd1 _3656_ sky130_fd_sc_hd__mux2_1
X_8378_ _3588_ _3589_ vssd1 vssd1 vccd1 vccd1 _3590_ sky130_fd_sc_hd__nor2_1
XFILLER_104_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7329_ _2402_ _2448_ vssd1 vssd1 vccd1 vccd1 _2449_ sky130_fd_sc_hd__xnor2_1
XFILLER_104_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5408__C1 _3830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6620__B2 _1384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5842__B _3770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5111__A1 _3925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5662__A2 _3892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4961_ _4109_ _4108_ vssd1 vssd1 vccd1 vccd1 _4116_ sky130_fd_sc_hd__xnor2_1
X_6700_ _1575_ _1576_ vssd1 vssd1 vccd1 vccd1 _1757_ sky130_fd_sc_hd__xor2_1
XFILLER_51_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4892_ _3984_ _4046_ vssd1 vssd1 vccd1 vccd1 _4047_ sky130_fd_sc_hd__xnor2_1
X_7680_ _2728_ _2833_ _2834_ vssd1 vssd1 vccd1 vccd1 _2835_ sky130_fd_sc_hd__o21ai_1
X_6631_ _1400_ _1676_ _1679_ _1680_ vssd1 vssd1 vccd1 vccd1 _1681_ sky130_fd_sc_hd__o31a_1
XFILLER_32_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6562_ _1603_ _1604_ vssd1 vssd1 vccd1 vccd1 _1606_ sky130_fd_sc_hd__nand2_1
X_8301_ _3437_ _3273_ _3475_ vssd1 vssd1 vccd1 vccd1 _3508_ sky130_fd_sc_hd__a21oi_1
XFILLER_20_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6493_ _1461_ _1529_ vssd1 vssd1 vccd1 vccd1 _1530_ sky130_fd_sc_hd__xnor2_1
X_5513_ _0483_ _0485_ _0338_ vssd1 vssd1 vccd1 vccd1 _0486_ sky130_fd_sc_hd__mux2_1
X_8232_ _3427_ _3433_ _3434_ vssd1 vssd1 vccd1 vccd1 _3436_ sky130_fd_sc_hd__o21ai_1
X_5444_ _0407_ _0410_ vssd1 vssd1 vccd1 vccd1 _0417_ sky130_fd_sc_hd__xnor2_1
XFILLER_105_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8163_ _0535_ _3215_ _3306_ vssd1 vssd1 vccd1 vccd1 _3362_ sky130_fd_sc_hd__a21boi_1
X_7114_ _1711_ _4089_ _1950_ vssd1 vssd1 vccd1 vccd1 _2213_ sky130_fd_sc_hd__and3_1
X_5375_ _0347_ _2452_ vssd1 vssd1 vccd1 vccd1 _0348_ sky130_fd_sc_hd__xnor2_2
X_4326_ _1363_ vssd1 vssd1 vccd1 vccd1 _1374_ sky130_fd_sc_hd__clkbuf_2
X_8094_ _3287_ vssd1 vssd1 vccd1 vccd1 _3288_ sky130_fd_sc_hd__clkinv_2
X_7045_ _2134_ _2135_ _2136_ vssd1 vssd1 vccd1 vccd1 _2137_ sky130_fd_sc_hd__and3_1
XFILLER_86_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4257_ net4 vssd1 vssd1 vccd1 vccd1 _0635_ sky130_fd_sc_hd__buf_2
XFILLER_47_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7947_ _2937_ _3056_ _3128_ vssd1 vssd1 vccd1 vccd1 _3129_ sky130_fd_sc_hd__a21bo_1
XFILLER_42_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7878_ _3052_ vssd1 vssd1 vccd1 vccd1 _3053_ sky130_fd_sc_hd__clkinv_2
X_6829_ _1838_ _1898_ vssd1 vssd1 vccd1 vccd1 _1899_ sky130_fd_sc_hd__xnor2_1
XFILLER_23_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8022__C cmd\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8465__S _3655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8346__A1 _0451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4741__B _3832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6949__A _1384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7544__S _2652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5160_ _0101_ _0131_ vssd1 vssd1 vccd1 vccd1 _0133_ sky130_fd_sc_hd__xnor2_1
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5091_ _4227_ _4231_ _4245_ vssd1 vssd1 vccd1 vccd1 _4246_ sky130_fd_sc_hd__o21a_1
XFILLER_110_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5993_ _0884_ _0981_ _0986_ _0989_ vssd1 vssd1 vccd1 vccd1 _0990_ sky130_fd_sc_hd__a31o_1
XFILLER_64_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7801_ _2904_ _2906_ _2966_ _2967_ _2891_ vssd1 vssd1 vccd1 vccd1 _2968_ sky130_fd_sc_hd__o32ai_1
XFILLER_24_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4944_ _4091_ _4098_ vssd1 vssd1 vccd1 vccd1 _4099_ sky130_fd_sc_hd__or2_1
X_7732_ _2835_ _2886_ _1297_ vssd1 vssd1 vccd1 vccd1 _2893_ sky130_fd_sc_hd__mux2_1
XANTENNA__8337__A1 _1308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4875_ _3914_ _3936_ _4029_ vssd1 vssd1 vccd1 vccd1 _4030_ sky130_fd_sc_hd__o21bai_2
X_7663_ _2790_ _2814_ _2816_ vssd1 vssd1 vccd1 vccd1 _2817_ sky130_fd_sc_hd__o21bai_1
X_6614_ _1277_ _1662_ _1302_ vssd1 vssd1 vccd1 vccd1 _1663_ sky130_fd_sc_hd__a21bo_1
X_7594_ _2739_ _2740_ vssd1 vssd1 vccd1 vccd1 _2741_ sky130_fd_sc_hd__xnor2_1
X_6545_ _1472_ _1478_ _1586_ vssd1 vssd1 vccd1 vccd1 _1587_ sky130_fd_sc_hd__o21ai_1
XFILLER_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5763__A _3866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6476_ _4232_ _1510_ vssd1 vssd1 vccd1 vccd1 _1511_ sky130_fd_sc_hd__nor2_4
X_8215_ _2604_ _2615_ _3416_ vssd1 vssd1 vccd1 vccd1 _3417_ sky130_fd_sc_hd__o21ba_1
X_5427_ _0347_ _4210_ vssd1 vssd1 vccd1 vccd1 _0400_ sky130_fd_sc_hd__nor2_1
XFILLER_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8146_ _0599_ _3343_ vssd1 vssd1 vccd1 vccd1 _3344_ sky130_fd_sc_hd__nor2_1
X_5358_ _0133_ _0163_ _0330_ vssd1 vssd1 vccd1 vccd1 _0331_ sky130_fd_sc_hd__o21bai_1
XFILLER_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4309_ last_SCLK net2 _1177_ vssd1 vssd1 vccd1 vccd1 _1188_ sky130_fd_sc_hd__mux2_1
X_8077_ _3166_ _3257_ _3267_ _3269_ vssd1 vssd1 vccd1 vccd1 _3270_ sky130_fd_sc_hd__o31a_1
XFILLER_101_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7028_ _2112_ _2115_ _2117_ vssd1 vssd1 vccd1 vccd1 _2118_ sky130_fd_sc_hd__a21o_1
X_5289_ _4156_ _4164_ _0261_ vssd1 vssd1 vccd1 vccd1 _0262_ sky130_fd_sc_hd__a21oi_1
XFILLER_75_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5003__A _3924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6009__A _4017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4660_ _3814_ vssd1 vssd1 vccd1 vccd1 _3815_ sky130_fd_sc_hd__clkbuf_4
XFILLER_14_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6330_ _1348_ _1337_ _1047_ vssd1 vssd1 vccd1 vccd1 _1350_ sky130_fd_sc_hd__nor3_1
X_4591_ _3189_ _3318_ _3745_ _3446_ vssd1 vssd1 vccd1 vccd1 _3746_ sky130_fd_sc_hd__a211o_2
X_6261_ _1272_ _1261_ vssd1 vssd1 vccd1 vccd1 _1274_ sky130_fd_sc_hd__and2b_1
XFILLER_115_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6192_ _1098_ _1100_ _4016_ _0802_ vssd1 vssd1 vccd1 vccd1 _1200_ sky130_fd_sc_hd__a211o_1
X_5212_ _4222_ _3883_ _0184_ vssd1 vssd1 vccd1 vccd1 _0185_ sky130_fd_sc_hd__and3_1
X_8000_ _3185_ _0121_ _3186_ vssd1 vssd1 vccd1 vccd1 _3187_ sky130_fd_sc_hd__o21a_1
X_5143_ _0115_ vssd1 vssd1 vccd1 vccd1 _0116_ sky130_fd_sc_hd__clkinv_2
XFILLER_111_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5074_ _4228_ _3800_ vssd1 vssd1 vccd1 vccd1 _4229_ sky130_fd_sc_hd__nor2_1
XFILLER_84_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5976_ _0968_ _0969_ _0970_ vssd1 vssd1 vccd1 vccd1 _0972_ sky130_fd_sc_hd__a21oi_1
XFILLER_80_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4927_ _3845_ _3817_ _3930_ _3828_ vssd1 vssd1 vccd1 vccd1 _4082_ sky130_fd_sc_hd__o22a_1
X_7715_ _2850_ _2872_ _2873_ vssd1 vssd1 vccd1 vccd1 _2874_ sky130_fd_sc_hd__o21ai_1
X_4858_ _3886_ _3873_ vssd1 vssd1 vccd1 vccd1 _4013_ sky130_fd_sc_hd__and2b_1
XFILLER_60_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7646_ _2742_ _2797_ vssd1 vssd1 vccd1 vccd1 _2798_ sky130_fd_sc_hd__or2_1
XFILLER_60_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4789_ _3893_ _3943_ vssd1 vssd1 vccd1 vccd1 _3944_ sky130_fd_sc_hd__nand2_1
X_7577_ _3802_ _4217_ _2721_ vssd1 vssd1 vccd1 vccd1 _2722_ sky130_fd_sc_hd__mux2_1
XFILLER_119_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6528_ _1511_ _1513_ vssd1 vssd1 vccd1 vccd1 _1568_ sky130_fd_sc_hd__xor2_4
XFILLER_4_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6459_ _1490_ _1491_ vssd1 vssd1 vccd1 vccd1 _1492_ sky130_fd_sc_hd__and2_1
XFILLER_79_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4259__D in_reg\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8129_ _3322_ _3324_ vssd1 vssd1 vccd1 vccd1 _3325_ sky130_fd_sc_hd__xnor2_2
XFILLER_48_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4572__A _3719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7883__A _2937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6011__B _0773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4747__A _3901_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4510__A2 _2980_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4466__B _2903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7777__B _2941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5830_ _0778_ _0783_ _0816_ vssd1 vssd1 vccd1 vccd1 _0817_ sky130_fd_sc_hd__o21a_1
X_5761_ _0113_ _0741_ _0742_ vssd1 vssd1 vccd1 vccd1 _0743_ sky130_fd_sc_hd__and3_1
XANTENNA__4577__A2 _2452_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7500_ _2826_ _0402_ _2636_ vssd1 vssd1 vccd1 vccd1 _2637_ sky130_fd_sc_hd__a21oi_1
X_8480_ _3675_ vssd1 vssd1 vccd1 vccd1 _3676_ sky130_fd_sc_hd__clkbuf_4
X_4712_ _3721_ _3156_ _3746_ _3748_ vssd1 vssd1 vccd1 vccd1 _3867_ sky130_fd_sc_hd__and4_1
X_5692_ _0666_ _0667_ _3718_ _3865_ vssd1 vssd1 vccd1 vccd1 _0669_ sky130_fd_sc_hd__a211oi_1
XFILLER_30_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7431_ _2425_ _2426_ _2427_ _2460_ vssd1 vssd1 vccd1 vccd1 _2561_ sky130_fd_sc_hd__a31o_1
X_4643_ _3780_ _3797_ vssd1 vssd1 vccd1 vccd1 _3798_ sky130_fd_sc_hd__and2b_1
X_4574_ _3678_ vssd1 vssd1 vccd1 vccd1 _3729_ sky130_fd_sc_hd__buf_4
X_7362_ _2484_ vssd1 vssd1 vccd1 vccd1 _2486_ sky130_fd_sc_hd__clkbuf_4
X_6313_ _1322_ vssd1 vssd1 vccd1 vccd1 _1332_ sky130_fd_sc_hd__inv_2
X_7293_ _2409_ vssd1 vssd1 vccd1 vccd1 _2410_ sky130_fd_sc_hd__buf_2
XFILLER_116_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6244_ _1235_ _1254_ _1255_ vssd1 vssd1 vccd1 vccd1 _1256_ sky130_fd_sc_hd__a21oi_1
XANTENNA__7732__S _1297_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6175_ _1029_ _1122_ vssd1 vssd1 vccd1 vccd1 _1181_ sky130_fd_sc_hd__xnor2_1
XFILLER_97_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4376__B _1913_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5126_ _0090_ _0098_ vssd1 vssd1 vccd1 vccd1 _0099_ sky130_fd_sc_hd__xor2_1
XFILLER_111_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5057_ _3925_ _4037_ vssd1 vssd1 vccd1 vccd1 _4212_ sky130_fd_sc_hd__or2_1
XFILLER_29_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5488__A _0092_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5959_ _0949_ _0953_ vssd1 vssd1 vccd1 vccd1 _0954_ sky130_fd_sc_hd__nor2_1
XFILLER_80_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7629_ _2762_ _2778_ vssd1 vssd1 vccd1 vccd1 _2779_ sky130_fd_sc_hd__nor2_1
XFILLER_5_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_644 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5951__A _0773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_704 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8473__S _3654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4290_ in_reg\[6\] in_reg\[7\] _0830_ vssd1 vssd1 vccd1 vccd1 _0988_ sky130_fd_sc_hd__mux2_1
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4477__A posit_add.in1\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7980_ _3160_ _3164_ _3030_ vssd1 vssd1 vccd1 vccd1 _3165_ sky130_fd_sc_hd__mux2_1
XFILLER_26_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6931_ _1414_ _1531_ _2010_ vssd1 vssd1 vccd1 vccd1 _2011_ sky130_fd_sc_hd__and3_1
XFILLER_81_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6862_ _1843_ _1934_ vssd1 vssd1 vccd1 vccd1 _1936_ sky130_fd_sc_hd__and2_1
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5813_ _0796_ _0798_ vssd1 vssd1 vccd1 vccd1 _0799_ sky130_fd_sc_hd__nand2_1
XFILLER_50_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8532_ clknet_3_5__leaf_clk _0018_ vssd1 vssd1 vccd1 vccd1 in_reg\[15\] sky130_fd_sc_hd__dfxtp_1
X_6793_ _1857_ _1859_ vssd1 vssd1 vccd1 vccd1 _1860_ sky130_fd_sc_hd__xor2_1
XFILLER_50_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5744_ _0721_ _0724_ _0720_ vssd1 vssd1 vccd1 vccd1 _0726_ sky130_fd_sc_hd__a21o_1
XANTENNA__8412__A cmd\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5675_ _3900_ _0609_ _3717_ vssd1 vssd1 vccd1 vccd1 _0650_ sky130_fd_sc_hd__a21o_1
X_8463_ in_reg\[8\] posit_add.in1\[8\] _3655_ vssd1 vssd1 vccd1 vccd1 _3666_ sky130_fd_sc_hd__mux2_1
XFILLER_30_391 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7414_ _0548_ _2158_ vssd1 vssd1 vccd1 vccd1 _2543_ sky130_fd_sc_hd__nand2_1
X_4626_ _3763_ _3725_ vssd1 vssd1 vccd1 vccd1 _3781_ sky130_fd_sc_hd__nor2_1
X_8394_ _3585_ _3602_ _3605_ _2621_ vssd1 vssd1 vccd1 vccd1 _3607_ sky130_fd_sc_hd__a31o_1
XANTENNA__8449__A0 in_reg\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7345_ _2454_ _2460_ _2466_ vssd1 vssd1 vccd1 vccd1 _2467_ sky130_fd_sc_hd__o21ai_1
X_4557_ _1726_ _2353_ _2364_ _2034_ vssd1 vssd1 vccd1 vccd1 _3712_ sky130_fd_sc_hd__o211a_1
XFILLER_103_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4488_ _3145_ vssd1 vssd1 vccd1 vccd1 _3156_ sky130_fd_sc_hd__buf_2
X_7276_ _2347_ _2359_ _2370_ _2374_ vssd1 vssd1 vccd1 vccd1 _2391_ sky130_fd_sc_hd__a31o_1
X_6227_ _1235_ _1236_ vssd1 vssd1 vccd1 vccd1 _1237_ sky130_fd_sc_hd__nor2_1
XFILLER_58_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6158_ _1159_ _1162_ vssd1 vssd1 vccd1 vccd1 _1163_ sky130_fd_sc_hd__nand2_1
XFILLER_103_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5109_ _4232_ vssd1 vssd1 vccd1 vccd1 _0082_ sky130_fd_sc_hd__buf_4
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6089_ _0973_ _1076_ vssd1 vssd1 vccd1 vccd1 _1090_ sky130_fd_sc_hd__xnor2_2
XFILLER_57_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5681__A _2507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6777__A _1420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6496__B _1456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7415__B2 _3804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5856__A _3770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5460_ _0432_ vssd1 vssd1 vccd1 vccd1 _0433_ sky130_fd_sc_hd__clkbuf_4
X_4411_ _2298_ vssd1 vssd1 vccd1 vccd1 _2309_ sky130_fd_sc_hd__buf_2
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5901__B2 _3735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5391_ _0356_ _0363_ vssd1 vssd1 vccd1 vccd1 _0364_ sky130_fd_sc_hd__or2b_1
XFILLER_98_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7130_ _2228_ _2229_ vssd1 vssd1 vccd1 vccd1 _2230_ sky130_fd_sc_hd__xor2_1
X_4342_ _1429_ _1539_ vssd1 vssd1 vccd1 vccd1 _1550_ sky130_fd_sc_hd__xor2_4
XANTENNA__4919__B _3883_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7061_ _2131_ _2132_ _2137_ vssd1 vssd1 vccd1 vccd1 _2154_ sky130_fd_sc_hd__a21oi_1
XFILLER_99_689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4273_ net4 _0797_ vssd1 vssd1 vccd1 vccd1 _0808_ sky130_fd_sc_hd__or2_1
XFILLER_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6012_ _1007_ _0993_ _1008_ vssd1 vssd1 vccd1 vccd1 _1010_ sky130_fd_sc_hd__a21bo_1
.ends

