VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tholin_nand_scaled
  CLASS BLOCK ;
  FOREIGN tholin_nand_scaled ;
  ORIGIN 0.000 0.000 ;
  SIZE 87.300 BY 97.300 ;
  OBS
      LAYER nwell ;
        RECT 4.000 77.800 85.900 97.300 ;
        RECT 4.000 54.700 38.600 77.800 ;
        RECT 51.300 54.700 85.900 77.800 ;
      LAYER li1 ;
        RECT 0.100 84.500 87.300 97.300 ;
        RECT 9.300 64.500 14.700 84.500 ;
        RECT 56.700 70.100 62.000 70.200 ;
        RECT 26.900 64.500 62.100 70.100 ;
        RECT 74.800 64.600 80.200 84.500 ;
        RECT 12.600 40.300 17.800 45.600 ;
        RECT 56.700 37.500 62.000 64.500 ;
        RECT 71.900 43.200 77.200 48.500 ;
        RECT 56.700 32.600 78.600 37.500 ;
        RECT 10.200 12.200 16.000 26.000 ;
        RECT 73.500 25.500 78.600 32.600 ;
        RECT 25.600 20.100 63.500 25.500 ;
        RECT 73.500 20.100 78.700 25.500 ;
        RECT 0.000 0.000 87.300 12.200 ;
      LAYER met4 ;
        RECT 0.970 85.240 86.480 96.220 ;
        RECT 0.520 1.070 85.870 11.130 ;
  END
END tholin_nand_scaled
END LIBRARY

