magic
tech sky130B
magscale 1 2
timestamp 1682095681
<< viali >>
rect 12817 22049 12851 22083
rect 10517 21981 10551 22015
rect 21465 21981 21499 22015
rect 22661 21981 22695 22015
rect 7113 21913 7147 21947
rect 7665 21913 7699 21947
rect 10272 21913 10306 21947
rect 12633 21913 12667 21947
rect 17049 21913 17083 21947
rect 17601 21913 17635 21947
rect 7757 21845 7791 21879
rect 9137 21845 9171 21879
rect 11069 21845 11103 21879
rect 12081 21845 12115 21879
rect 14289 21845 14323 21879
rect 14933 21845 14967 21879
rect 15669 21845 15703 21879
rect 17693 21845 17727 21879
rect 22569 21845 22603 21879
rect 17693 21641 17727 21675
rect 19993 21641 20027 21675
rect 16129 21573 16163 21607
rect 18337 21573 18371 21607
rect 22201 21573 22235 21607
rect 2780 21505 2814 21539
rect 4629 21505 4663 21539
rect 4896 21505 4930 21539
rect 10077 21505 10111 21539
rect 10333 21505 10367 21539
rect 12081 21505 12115 21539
rect 13093 21505 13127 21539
rect 14197 21505 14231 21539
rect 15117 21505 15151 21539
rect 17969 21505 18003 21539
rect 20283 21505 20317 21539
rect 21097 21505 21131 21539
rect 21281 21505 21315 21539
rect 22385 21505 22419 21539
rect 2513 21437 2547 21471
rect 13921 21437 13955 21471
rect 14933 21437 14967 21471
rect 15025 21437 15059 21471
rect 15209 21437 15243 21471
rect 17877 21437 17911 21471
rect 20453 21437 20487 21471
rect 21189 21437 21223 21471
rect 12173 21369 12207 21403
rect 14749 21369 14783 21403
rect 15761 21369 15795 21403
rect 16313 21369 16347 21403
rect 22017 21369 22051 21403
rect 3893 21301 3927 21335
rect 6009 21301 6043 21335
rect 8953 21301 8987 21335
rect 11161 21301 11195 21335
rect 13001 21301 13035 21335
rect 16129 21301 16163 21335
rect 11713 21097 11747 21131
rect 14289 21097 14323 21131
rect 21281 21097 21315 21131
rect 12265 21029 12299 21063
rect 13461 21029 13495 21063
rect 14565 21029 14599 21063
rect 16221 21029 16255 21063
rect 5365 20961 5399 20995
rect 5825 20961 5859 20995
rect 9137 20961 9171 20995
rect 11345 20961 11379 20995
rect 14656 20961 14690 20995
rect 14749 20961 14783 20995
rect 2053 20893 2087 20927
rect 6092 20893 6126 20927
rect 11529 20893 11563 20927
rect 11805 20893 11839 20927
rect 12449 20893 12483 20927
rect 12817 20893 12851 20927
rect 13737 20893 13771 20927
rect 14473 20893 14507 20927
rect 15393 20893 15427 20927
rect 15577 20893 15611 20927
rect 16405 20893 16439 20927
rect 16681 20893 16715 20927
rect 16957 20893 16991 20927
rect 17601 20893 17635 20927
rect 21189 20893 21223 20927
rect 21373 20893 21407 20927
rect 14933 20859 14967 20893
rect 2298 20825 2332 20859
rect 5098 20825 5132 20859
rect 9404 20825 9438 20859
rect 12541 20825 12575 20859
rect 12633 20825 12667 20859
rect 13461 20825 13495 20859
rect 3433 20757 3467 20791
rect 3985 20757 4019 20791
rect 7205 20757 7239 20791
rect 10517 20757 10551 20791
rect 13645 20757 13679 20791
rect 15393 20757 15427 20791
rect 10333 20553 10367 20587
rect 12265 20553 12299 20587
rect 14841 20553 14875 20587
rect 15669 20553 15703 20587
rect 18429 20553 18463 20587
rect 22109 20553 22143 20587
rect 19533 20485 19567 20519
rect 4353 20417 4387 20451
rect 8953 20417 8987 20451
rect 9220 20417 9254 20451
rect 12173 20417 12207 20451
rect 13185 20417 13219 20451
rect 13553 20417 13587 20451
rect 13921 20417 13955 20451
rect 14197 20417 14231 20451
rect 15025 20417 15059 20451
rect 15209 20417 15243 20451
rect 15853 20417 15887 20451
rect 16037 20417 16071 20451
rect 16129 20417 16163 20451
rect 16313 20417 16347 20451
rect 17279 20417 17313 20451
rect 17417 20417 17451 20451
rect 17509 20417 17543 20451
rect 17693 20417 17727 20451
rect 18613 20417 18647 20451
rect 18705 20417 18739 20451
rect 18889 20417 18923 20451
rect 18981 20417 19015 20451
rect 19441 20417 19475 20451
rect 19625 20417 19659 20451
rect 22017 20417 22051 20451
rect 22201 20417 22235 20451
rect 2605 20349 2639 20383
rect 17049 20349 17083 20383
rect 13553 20281 13587 20315
rect 15945 20281 15979 20315
rect 11161 20213 11195 20247
rect 15209 20213 15243 20247
rect 12173 20009 12207 20043
rect 14749 20009 14783 20043
rect 18245 20009 18279 20043
rect 15945 19941 15979 19975
rect 16497 19941 16531 19975
rect 2053 19873 2087 19907
rect 6653 19873 6687 19907
rect 9137 19873 9171 19907
rect 12817 19873 12851 19907
rect 15393 19873 15427 19907
rect 16681 19873 16715 19907
rect 20269 19873 20303 19907
rect 9404 19805 9438 19839
rect 10977 19805 11011 19839
rect 12633 19805 12667 19839
rect 14657 19805 14691 19839
rect 14841 19805 14875 19839
rect 16405 19805 16439 19839
rect 17417 19805 17451 19839
rect 17601 19805 17635 19839
rect 20545 19805 20579 19839
rect 2298 19737 2332 19771
rect 6386 19737 6420 19771
rect 16681 19737 16715 19771
rect 3433 19669 3467 19703
rect 5273 19669 5307 19703
rect 10517 19669 10551 19703
rect 11621 19669 11655 19703
rect 12541 19669 12575 19703
rect 17233 19669 17267 19703
rect 4261 19465 4295 19499
rect 6653 19465 6687 19499
rect 10333 19465 10367 19499
rect 17509 19465 17543 19499
rect 7766 19397 7800 19431
rect 17417 19397 17451 19431
rect 20453 19397 20487 19431
rect 3148 19329 3182 19363
rect 8033 19329 8067 19363
rect 8953 19329 8987 19363
rect 9220 19329 9254 19363
rect 14657 19329 14691 19363
rect 14841 19329 14875 19363
rect 15301 19329 15335 19363
rect 17325 19329 17359 19363
rect 17785 19329 17819 19363
rect 19349 19329 19383 19363
rect 19533 19329 19567 19363
rect 19625 19329 19659 19363
rect 20269 19329 20303 19363
rect 20545 19329 20579 19363
rect 21281 19329 21315 19363
rect 2881 19261 2915 19295
rect 15485 19261 15519 19295
rect 19165 19261 19199 19295
rect 20085 19261 20119 19295
rect 21005 19261 21039 19295
rect 14749 19125 14783 19159
rect 5825 18921 5859 18955
rect 7665 18921 7699 18955
rect 14289 18921 14323 18955
rect 16037 18921 16071 18955
rect 18337 18921 18371 18955
rect 19441 18921 19475 18955
rect 22385 18921 22419 18955
rect 16865 18853 16899 18887
rect 9137 18785 9171 18819
rect 13185 18785 13219 18819
rect 13277 18785 13311 18819
rect 13553 18785 13587 18819
rect 15393 18785 15427 18819
rect 18613 18785 18647 18819
rect 3433 18717 3467 18751
rect 6377 18717 6411 18751
rect 13093 18717 13127 18751
rect 13369 18717 13403 18751
rect 14473 18717 14507 18751
rect 14933 18717 14967 18751
rect 15761 18717 15795 18751
rect 15853 18717 15887 18751
rect 16681 18717 16715 18751
rect 16957 18717 16991 18751
rect 18521 18717 18555 18751
rect 18705 18717 18739 18751
rect 18797 18717 18831 18751
rect 19579 18717 19613 18751
rect 19717 18717 19751 18751
rect 19937 18717 19971 18751
rect 20085 18717 20119 18751
rect 20729 18717 20763 18751
rect 21005 18717 21039 18751
rect 22109 18717 22143 18751
rect 3188 18649 3222 18683
rect 9404 18649 9438 18683
rect 14565 18649 14599 18683
rect 14657 18649 14691 18683
rect 14775 18649 14809 18683
rect 15485 18649 15519 18683
rect 19809 18649 19843 18683
rect 22293 18649 22327 18683
rect 2053 18581 2087 18615
rect 10517 18581 10551 18615
rect 16497 18581 16531 18615
rect 20545 18581 20579 18615
rect 20913 18581 20947 18615
rect 9137 18377 9171 18411
rect 13553 18377 13587 18411
rect 14657 18377 14691 18411
rect 19809 18377 19843 18411
rect 20913 18377 20947 18411
rect 22017 18377 22051 18411
rect 7849 18309 7883 18343
rect 14289 18309 14323 18343
rect 2881 18241 2915 18275
rect 13093 18241 13127 18275
rect 13377 18241 13411 18275
rect 14197 18241 14231 18275
rect 14473 18241 14507 18275
rect 16957 18241 16991 18275
rect 17141 18241 17175 18275
rect 20065 18241 20099 18275
rect 20158 18241 20192 18275
rect 20274 18241 20308 18275
rect 20453 18241 20487 18275
rect 22293 18241 22327 18275
rect 22382 18244 22416 18278
rect 22477 18241 22511 18275
rect 22661 18241 22695 18275
rect 2605 18173 2639 18207
rect 13185 18173 13219 18207
rect 13299 18173 13333 18207
rect 15669 18105 15703 18139
rect 4169 18037 4203 18071
rect 15209 18037 15243 18071
rect 16221 18037 16255 18071
rect 16957 18037 16991 18071
rect 17601 18037 17635 18071
rect 19349 18037 19383 18071
rect 13277 17833 13311 17867
rect 19441 17833 19475 17867
rect 19809 17833 19843 17867
rect 22661 17833 22695 17867
rect 7113 17697 7147 17731
rect 9137 17697 9171 17731
rect 17693 17697 17727 17731
rect 19717 17697 19751 17731
rect 2053 17629 2087 17663
rect 9404 17629 9438 17663
rect 12817 17629 12851 17663
rect 13093 17629 13127 17663
rect 14473 17629 14507 17663
rect 16221 17629 16255 17663
rect 16497 17629 16531 17663
rect 17417 17629 17451 17663
rect 17601 17629 17635 17663
rect 18153 17629 18187 17663
rect 18245 17629 18279 17663
rect 18889 17629 18923 17663
rect 19809 17629 19843 17663
rect 21833 17629 21867 17663
rect 22109 17629 22143 17663
rect 2320 17561 2354 17595
rect 6846 17561 6880 17595
rect 14933 17561 14967 17595
rect 15485 17561 15519 17595
rect 3433 17493 3467 17527
rect 5733 17493 5767 17527
rect 10517 17493 10551 17527
rect 12909 17493 12943 17527
rect 14381 17493 14415 17527
rect 16037 17493 16071 17527
rect 16405 17493 16439 17527
rect 17233 17493 17267 17527
rect 21649 17493 21683 17527
rect 22017 17493 22051 17527
rect 12173 17289 12207 17323
rect 12633 17289 12667 17323
rect 14013 17289 14047 17323
rect 19073 17289 19107 17323
rect 19717 17289 19751 17323
rect 20729 17289 20763 17323
rect 16957 17221 16991 17255
rect 8861 17153 8895 17187
rect 12817 17153 12851 17187
rect 12909 17153 12943 17187
rect 13185 17153 13219 17187
rect 14289 17153 14323 17187
rect 15485 17153 15519 17187
rect 16865 17153 16899 17187
rect 17141 17153 17175 17187
rect 17877 17153 17911 17187
rect 18981 17153 19015 17187
rect 19349 17153 19383 17187
rect 20913 17153 20947 17187
rect 21005 17153 21039 17187
rect 2697 17085 2731 17119
rect 2973 17085 3007 17119
rect 9137 17085 9171 17119
rect 14197 17085 14231 17119
rect 14381 17085 14415 17119
rect 14473 17085 14507 17119
rect 15301 17085 15335 17119
rect 18153 17085 18187 17119
rect 20729 17085 20763 17119
rect 11069 17017 11103 17051
rect 13093 17017 13127 17051
rect 17141 17017 17175 17051
rect 19441 17017 19475 17051
rect 20269 17017 20303 17051
rect 4261 16949 4295 16983
rect 8401 16949 8435 16983
rect 10425 16949 10459 16983
rect 16037 16949 16071 16983
rect 17693 16949 17727 16983
rect 18061 16949 18095 16983
rect 19257 16949 19291 16983
rect 15485 16745 15519 16779
rect 22017 16745 22051 16779
rect 22201 16745 22235 16779
rect 15025 16677 15059 16711
rect 16497 16677 16531 16711
rect 20177 16677 20211 16711
rect 6653 16609 6687 16643
rect 7113 16609 7147 16643
rect 9137 16609 9171 16643
rect 9413 16609 9447 16643
rect 12633 16609 12667 16643
rect 15945 16609 15979 16643
rect 17141 16609 17175 16643
rect 17785 16609 17819 16643
rect 20361 16609 20395 16643
rect 2053 16541 2087 16575
rect 7380 16541 7414 16575
rect 11897 16541 11931 16575
rect 12081 16541 12115 16575
rect 12831 16551 12865 16585
rect 12982 16541 13016 16575
rect 13105 16541 13139 16575
rect 13195 16541 13229 16575
rect 14381 16541 14415 16575
rect 14529 16541 14563 16575
rect 14846 16541 14880 16575
rect 15669 16541 15703 16575
rect 15761 16541 15795 16575
rect 16037 16541 16071 16575
rect 17325 16541 17359 16575
rect 20085 16541 20119 16575
rect 20269 16541 20303 16575
rect 20545 16541 20579 16575
rect 2320 16473 2354 16507
rect 6386 16473 6420 16507
rect 14657 16473 14691 16507
rect 14749 16473 14783 16507
rect 17417 16473 17451 16507
rect 17509 16473 17543 16507
rect 17647 16473 17681 16507
rect 22385 16473 22419 16507
rect 3433 16405 3467 16439
rect 5273 16405 5307 16439
rect 8493 16405 8527 16439
rect 10701 16405 10735 16439
rect 12081 16405 12115 16439
rect 13737 16405 13771 16439
rect 18889 16405 18923 16439
rect 19901 16405 19935 16439
rect 21005 16405 21039 16439
rect 22185 16405 22219 16439
rect 9137 16201 9171 16235
rect 18337 16201 18371 16235
rect 20453 16201 20487 16235
rect 4353 16133 4387 16167
rect 7849 16133 7883 16167
rect 20821 16133 20855 16167
rect 11713 16065 11747 16099
rect 11989 16065 12023 16099
rect 12725 16065 12759 16099
rect 13093 16065 13127 16099
rect 17049 16065 17083 16099
rect 17325 16065 17359 16099
rect 18705 16065 18739 16099
rect 19625 16065 19659 16099
rect 19809 16065 19843 16099
rect 20637 16065 20671 16099
rect 20729 16065 20763 16099
rect 21005 16065 21039 16099
rect 21097 16065 21131 16099
rect 11805 15997 11839 16031
rect 14197 15997 14231 16031
rect 16129 15997 16163 16031
rect 16957 15997 16991 16031
rect 17233 15997 17267 16031
rect 18613 15997 18647 16031
rect 22109 15997 22143 16031
rect 19901 15929 19935 15963
rect 3065 15861 3099 15895
rect 12173 15861 12207 15895
rect 15025 15861 15059 15895
rect 15669 15861 15703 15895
rect 17141 15861 17175 15895
rect 18705 15861 18739 15895
rect 22661 15861 22695 15895
rect 14289 15657 14323 15691
rect 15117 15657 15151 15691
rect 19993 15657 20027 15691
rect 22109 15657 22143 15691
rect 22753 15657 22787 15691
rect 16681 15589 16715 15623
rect 18153 15589 18187 15623
rect 4997 15521 5031 15555
rect 9137 15521 9171 15555
rect 11989 15521 12023 15555
rect 15301 15521 15335 15555
rect 15393 15521 15427 15555
rect 19441 15521 19475 15555
rect 2237 15453 2271 15487
rect 2513 15453 2547 15487
rect 3985 15453 4019 15487
rect 11253 15453 11287 15487
rect 11345 15453 11379 15487
rect 11529 15453 11563 15487
rect 12541 15453 12575 15487
rect 13645 15453 13679 15487
rect 14289 15453 14323 15487
rect 14473 15453 14507 15487
rect 15485 15453 15519 15487
rect 15577 15453 15611 15487
rect 16681 15453 16715 15487
rect 18705 15453 18739 15487
rect 18889 15453 18923 15487
rect 21097 15453 21131 15487
rect 22293 15453 22327 15487
rect 3341 15385 3375 15419
rect 4261 15385 4295 15419
rect 5264 15385 5298 15419
rect 9404 15385 9438 15419
rect 12909 15385 12943 15419
rect 16773 15385 16807 15419
rect 16957 15385 16991 15419
rect 18797 15385 18831 15419
rect 20821 15385 20855 15419
rect 2053 15317 2087 15351
rect 2421 15317 2455 15351
rect 3065 15317 3099 15351
rect 6377 15317 6411 15351
rect 10517 15317 10551 15351
rect 16221 15317 16255 15351
rect 4813 15113 4847 15147
rect 11713 15113 11747 15147
rect 20361 15113 20395 15147
rect 22661 15113 22695 15147
rect 1869 15045 1903 15079
rect 5181 15045 5215 15079
rect 6561 15045 6595 15079
rect 19349 15045 19383 15079
rect 1593 14977 1627 15011
rect 1777 14977 1811 15011
rect 1961 14977 1995 15011
rect 4997 14977 5031 15011
rect 5089 14977 5123 15011
rect 5365 14977 5399 15011
rect 6009 14977 6043 15011
rect 6745 14977 6779 15011
rect 6837 14977 6871 15011
rect 9689 14977 9723 15011
rect 12541 14977 12575 15011
rect 13093 14977 13127 15011
rect 13277 14977 13311 15011
rect 13369 14977 13403 15011
rect 13829 14977 13863 15011
rect 14749 14977 14783 15011
rect 15577 14977 15611 15011
rect 15853 14977 15887 15011
rect 19525 14977 19559 15011
rect 19625 14977 19659 15011
rect 19809 14977 19843 15011
rect 19901 14977 19935 15011
rect 20913 14977 20947 15011
rect 21097 14977 21131 15011
rect 22017 14977 22051 15011
rect 22110 14977 22144 15011
rect 22293 14977 22327 15011
rect 22385 14977 22419 15011
rect 22523 14977 22557 15011
rect 2697 14909 2731 14943
rect 2973 14909 3007 14943
rect 9413 14909 9447 14943
rect 10241 14909 10275 14943
rect 14105 14909 14139 14943
rect 15025 14909 15059 14943
rect 18889 14909 18923 14943
rect 20637 14909 20671 14943
rect 11161 14841 11195 14875
rect 14841 14841 14875 14875
rect 20729 14841 20763 14875
rect 2145 14773 2179 14807
rect 4261 14773 4295 14807
rect 6561 14773 6595 14807
rect 8125 14773 8159 14807
rect 14749 14773 14783 14807
rect 16865 14773 16899 14807
rect 20821 14773 20855 14807
rect 23121 14773 23155 14807
rect 2053 14569 2087 14603
rect 4721 14569 4755 14603
rect 5825 14569 5859 14603
rect 6837 14569 6871 14603
rect 9137 14569 9171 14603
rect 12633 14569 12667 14603
rect 15025 14569 15059 14603
rect 19441 14569 19475 14603
rect 20453 14569 20487 14603
rect 22385 14569 22419 14603
rect 10701 14501 10735 14535
rect 2421 14433 2455 14467
rect 4169 14433 4203 14467
rect 11069 14433 11103 14467
rect 12173 14433 12207 14467
rect 12357 14433 12391 14467
rect 12449 14433 12483 14467
rect 16221 14433 16255 14467
rect 17509 14433 17543 14467
rect 2237 14365 2271 14399
rect 3065 14365 3099 14399
rect 3157 14365 3191 14399
rect 3433 14365 3467 14399
rect 4261 14365 4295 14399
rect 4353 14365 4387 14399
rect 6009 14365 6043 14399
rect 6377 14365 6411 14399
rect 7021 14365 7055 14399
rect 7389 14365 7423 14399
rect 7941 14365 7975 14399
rect 9321 14365 9355 14399
rect 9689 14365 9723 14399
rect 12265 14365 12299 14399
rect 14289 14365 14323 14399
rect 14381 14365 14415 14399
rect 14565 14365 14599 14399
rect 14749 14365 14783 14399
rect 17325 14365 17359 14399
rect 17417 14365 17451 14399
rect 17601 14365 17635 14399
rect 19625 14365 19659 14399
rect 19717 14365 19751 14399
rect 19901 14365 19935 14399
rect 19993 14365 20027 14399
rect 21097 14365 21131 14399
rect 21741 14365 21775 14399
rect 22569 14365 22603 14399
rect 22845 14365 22879 14399
rect 3249 14297 3283 14331
rect 6101 14297 6135 14331
rect 6193 14297 6227 14331
rect 7113 14297 7147 14331
rect 7205 14297 7239 14331
rect 8401 14297 8435 14331
rect 9413 14297 9447 14331
rect 9505 14297 9539 14331
rect 11161 14297 11195 14331
rect 11253 14297 11287 14331
rect 13461 14297 13495 14331
rect 14657 14297 14691 14331
rect 16037 14297 16071 14331
rect 2881 14229 2915 14263
rect 15669 14229 15703 14263
rect 16129 14229 16163 14263
rect 17141 14229 17175 14263
rect 21833 14229 21867 14263
rect 22753 14229 22787 14263
rect 3985 14025 4019 14059
rect 5089 14025 5123 14059
rect 9597 14025 9631 14059
rect 12817 14025 12851 14059
rect 15577 14025 15611 14059
rect 20361 14025 20395 14059
rect 2872 13957 2906 13991
rect 8484 13957 8518 13991
rect 15853 13957 15887 13991
rect 22661 13957 22695 13991
rect 2145 13889 2179 13923
rect 2605 13889 2639 13923
rect 5457 13889 5491 13923
rect 5549 13889 5583 13923
rect 8217 13889 8251 13923
rect 10057 13889 10091 13923
rect 10241 13889 10275 13923
rect 10915 13889 10949 13923
rect 11069 13889 11103 13923
rect 14565 13889 14599 13923
rect 14657 13889 14691 13923
rect 14841 13889 14875 13923
rect 14933 13889 14967 13923
rect 15761 13889 15795 13923
rect 15945 13889 15979 13923
rect 16129 13889 16163 13923
rect 17877 13889 17911 13923
rect 17969 13889 18003 13923
rect 18153 13889 18187 13923
rect 18245 13889 18279 13923
rect 19257 13889 19291 13923
rect 20637 13889 20671 13923
rect 20729 13889 20763 13923
rect 20821 13889 20855 13923
rect 20999 13889 21033 13923
rect 22293 13889 22327 13923
rect 22569 13889 22603 13923
rect 22845 13889 22879 13923
rect 1869 13821 1903 13855
rect 5641 13821 5675 13855
rect 11805 13821 11839 13855
rect 19073 13821 19107 13855
rect 19349 13821 19383 13855
rect 19441 13821 19475 13855
rect 19533 13821 19567 13855
rect 23029 13821 23063 13855
rect 1961 13753 1995 13787
rect 17693 13753 17727 13787
rect 2053 13685 2087 13719
rect 7481 13685 7515 13719
rect 10241 13685 10275 13719
rect 10885 13685 10919 13719
rect 14105 13685 14139 13719
rect 15117 13685 15151 13719
rect 16957 13685 16991 13719
rect 4445 13481 4479 13515
rect 4629 13481 4663 13515
rect 5273 13481 5307 13515
rect 6653 13481 6687 13515
rect 9689 13481 9723 13515
rect 15669 13481 15703 13515
rect 16589 13481 16623 13515
rect 19441 13481 19475 13515
rect 20637 13481 20671 13515
rect 21465 13481 21499 13515
rect 2697 13413 2731 13447
rect 6561 13413 6595 13447
rect 11253 13413 11287 13447
rect 14841 13413 14875 13447
rect 6193 13345 6227 13379
rect 10333 13345 10367 13379
rect 19625 13345 19659 13379
rect 19901 13345 19935 13379
rect 21005 13345 21039 13379
rect 2145 13277 2179 13311
rect 2329 13277 2363 13311
rect 2513 13277 2547 13311
rect 3433 13277 3467 13311
rect 5181 13277 5215 13311
rect 7205 13277 7239 13311
rect 7849 13277 7883 13311
rect 10241 13277 10275 13311
rect 10609 13277 10643 13311
rect 10701 13277 10735 13311
rect 11897 13277 11931 13311
rect 12449 13277 12483 13311
rect 14289 13277 14323 13311
rect 14565 13277 14599 13311
rect 15301 13277 15335 13311
rect 15485 13277 15519 13311
rect 16129 13277 16163 13311
rect 16405 13277 16439 13311
rect 17049 13277 17083 13311
rect 17141 13277 17175 13311
rect 17325 13277 17359 13311
rect 17417 13277 17451 13311
rect 19718 13277 19752 13311
rect 19809 13277 19843 13311
rect 20821 13277 20855 13311
rect 21649 13277 21683 13311
rect 21925 13277 21959 13311
rect 22753 13277 22787 13311
rect 2421 13209 2455 13243
rect 4261 13209 4295 13243
rect 4461 13209 4495 13243
rect 16221 13209 16255 13243
rect 23029 13209 23063 13243
rect 3249 13141 3283 13175
rect 7205 13141 7239 13175
rect 14473 13141 14507 13175
rect 14657 13141 14691 13175
rect 17601 13141 17635 13175
rect 18889 13141 18923 13175
rect 21833 13141 21867 13175
rect 3334 12937 3368 12971
rect 4195 12937 4229 12971
rect 8217 12937 8251 12971
rect 19441 12937 19475 12971
rect 22293 12937 22327 12971
rect 2605 12869 2639 12903
rect 3433 12869 3467 12903
rect 3985 12869 4019 12903
rect 12541 12869 12575 12903
rect 14657 12869 14691 12903
rect 15301 12869 15335 12903
rect 17233 12869 17267 12903
rect 21465 12869 21499 12903
rect 22779 12869 22813 12903
rect 3157 12801 3191 12835
rect 3249 12801 3283 12835
rect 5273 12801 5307 12835
rect 5365 12801 5399 12835
rect 7297 12801 7331 12835
rect 7389 12801 7423 12835
rect 7573 12801 7607 12835
rect 7665 12801 7699 12835
rect 8125 12801 8159 12835
rect 8309 12801 8343 12835
rect 8953 12801 8987 12835
rect 9045 12801 9079 12835
rect 9321 12801 9355 12835
rect 10425 12801 10459 12835
rect 10517 12801 10551 12835
rect 10701 12801 10735 12835
rect 11897 12801 11931 12835
rect 12173 12801 12207 12835
rect 12357 12801 12391 12835
rect 13645 12801 13679 12835
rect 14013 12801 14047 12835
rect 15853 12801 15887 12835
rect 16865 12801 16899 12835
rect 16958 12801 16992 12835
rect 17141 12801 17175 12835
rect 17349 12801 17383 12835
rect 19625 12801 19659 12835
rect 19717 12801 19751 12835
rect 19901 12801 19935 12835
rect 20085 12801 20119 12835
rect 21097 12801 21131 12835
rect 22477 12801 22511 12835
rect 22569 12801 22603 12835
rect 22661 12801 22695 12835
rect 22937 12801 22971 12835
rect 9229 12733 9263 12767
rect 11161 12733 11195 12767
rect 13737 12733 13771 12767
rect 14197 12733 14231 12767
rect 15945 12733 15979 12767
rect 16037 12733 16071 12767
rect 16129 12733 16163 12767
rect 4353 12665 4387 12699
rect 7113 12665 7147 12699
rect 18061 12665 18095 12699
rect 19809 12665 19843 12699
rect 1777 12597 1811 12631
rect 2513 12597 2547 12631
rect 4169 12597 4203 12631
rect 6561 12597 6595 12631
rect 8769 12597 8803 12631
rect 16313 12597 16347 12631
rect 17509 12597 17543 12631
rect 18613 12597 18647 12631
rect 4077 12393 4111 12427
rect 6009 12393 6043 12427
rect 7389 12393 7423 12427
rect 8125 12393 8159 12427
rect 11529 12393 11563 12427
rect 11989 12393 12023 12427
rect 13645 12393 13679 12427
rect 15393 12393 15427 12427
rect 16313 12393 16347 12427
rect 19441 12393 19475 12427
rect 20729 12393 20763 12427
rect 6745 12325 6779 12359
rect 12541 12325 12575 12359
rect 16497 12325 16531 12359
rect 21097 12325 21131 12359
rect 2237 12257 2271 12291
rect 11805 12257 11839 12291
rect 2053 12189 2087 12223
rect 2421 12189 2455 12223
rect 2973 12189 3007 12223
rect 3157 12189 3191 12223
rect 3985 12189 4019 12223
rect 4169 12189 4203 12223
rect 6561 12189 6595 12223
rect 6745 12189 6779 12223
rect 7205 12189 7239 12223
rect 7389 12189 7423 12223
rect 8401 12189 8435 12223
rect 10057 12189 10091 12223
rect 10425 12189 10459 12223
rect 10701 12189 10735 12223
rect 11713 12189 11747 12223
rect 13553 12189 13587 12223
rect 13737 12189 13771 12223
rect 14289 12189 14323 12223
rect 14473 12189 14507 12223
rect 14841 12189 14875 12223
rect 17509 12189 17543 12223
rect 17601 12189 17635 12223
rect 17693 12189 17727 12223
rect 17877 12189 17911 12223
rect 20729 12189 20763 12223
rect 20821 12189 20855 12223
rect 21741 12189 21775 12223
rect 21833 12189 21867 12223
rect 22017 12189 22051 12223
rect 22109 12189 22143 12223
rect 23121 12189 23155 12223
rect 2881 12121 2915 12155
rect 8125 12121 8159 12155
rect 9229 12121 9263 12155
rect 11989 12121 12023 12155
rect 16129 12121 16163 12155
rect 21557 12121 21591 12155
rect 22845 12121 22879 12155
rect 2145 12053 2179 12087
rect 2329 12053 2363 12087
rect 4629 12053 4663 12087
rect 8309 12053 8343 12087
rect 9781 12053 9815 12087
rect 13093 12053 13127 12087
rect 16329 12053 16363 12087
rect 17233 12053 17267 12087
rect 18429 12053 18463 12087
rect 20085 12053 20119 12087
rect 1869 11849 1903 11883
rect 2513 11849 2547 11883
rect 2697 11849 2731 11883
rect 4813 11849 4847 11883
rect 5917 11849 5951 11883
rect 7941 11849 7975 11883
rect 11897 11849 11931 11883
rect 12081 11849 12115 11883
rect 17877 11849 17911 11883
rect 19717 11849 19751 11883
rect 19993 11849 20027 11883
rect 21373 11849 21407 11883
rect 23029 11849 23063 11883
rect 2881 11781 2915 11815
rect 5181 11781 5215 11815
rect 9413 11781 9447 11815
rect 11713 11781 11747 11815
rect 13461 11781 13495 11815
rect 14289 11781 14323 11815
rect 19625 11781 19659 11815
rect 1593 11713 1627 11747
rect 1685 11713 1719 11747
rect 3985 11713 4019 11747
rect 4078 11713 4112 11747
rect 4997 11713 5031 11747
rect 5089 11713 5123 11747
rect 5299 11713 5333 11747
rect 5457 11713 5491 11747
rect 7297 11713 7331 11747
rect 7849 11713 7883 11747
rect 8125 11713 8159 11747
rect 8677 11713 8711 11747
rect 9229 11713 9263 11747
rect 10333 11713 10367 11747
rect 10977 11713 11011 11747
rect 11161 11713 11195 11747
rect 13369 11713 13403 11747
rect 13829 11713 13863 11747
rect 17417 11713 17451 11747
rect 17601 11713 17635 11747
rect 17693 11713 17727 11747
rect 19441 11713 19475 11747
rect 19809 11713 19843 11747
rect 21281 11713 21315 11747
rect 21465 11713 21499 11747
rect 22109 11713 22143 11747
rect 23029 11713 23063 11747
rect 23213 11713 23247 11747
rect 1869 11645 1903 11679
rect 3341 11645 3375 11679
rect 7021 11645 7055 11679
rect 7113 11645 7147 11679
rect 7205 11645 7239 11679
rect 10057 11645 10091 11679
rect 13553 11645 13587 11679
rect 17509 11645 17543 11679
rect 22385 11645 22419 11679
rect 20453 11577 20487 11611
rect 2697 11509 2731 11543
rect 4169 11509 4203 11543
rect 6837 11509 6871 11543
rect 10793 11509 10827 11543
rect 11897 11509 11931 11543
rect 14749 11509 14783 11543
rect 15393 11509 15427 11543
rect 15945 11509 15979 11543
rect 18429 11509 18463 11543
rect 18981 11509 19015 11543
rect 4629 11305 4663 11339
rect 9137 11305 9171 11339
rect 13645 11305 13679 11339
rect 19533 11305 19567 11339
rect 19625 11305 19659 11339
rect 22293 11305 22327 11339
rect 3157 11237 3191 11271
rect 14933 11237 14967 11271
rect 20821 11237 20855 11271
rect 4077 11169 4111 11203
rect 4445 11169 4479 11203
rect 5549 11169 5583 11203
rect 8493 11169 8527 11203
rect 15761 11169 15795 11203
rect 18429 11169 18463 11203
rect 19441 11169 19475 11203
rect 22845 11169 22879 11203
rect 1593 11101 1627 11135
rect 2421 11101 2455 11135
rect 2789 11101 2823 11135
rect 2973 11101 3007 11135
rect 3985 11101 4019 11135
rect 4353 11101 4387 11135
rect 6653 11101 6687 11135
rect 7389 11101 7423 11135
rect 9321 11101 9355 11135
rect 9505 11101 9539 11135
rect 9781 11101 9815 11135
rect 10609 11101 10643 11135
rect 10793 11101 10827 11135
rect 11897 11101 11931 11135
rect 12081 11101 12115 11135
rect 12173 11101 12207 11135
rect 12633 11101 12667 11135
rect 13093 11101 13127 11135
rect 13461 11101 13495 11135
rect 14289 11101 14323 11135
rect 14382 11101 14416 11135
rect 14754 11101 14788 11135
rect 15485 11101 15519 11135
rect 15669 11101 15703 11135
rect 16865 11101 16899 11135
rect 17417 11101 17451 11135
rect 18337 11101 18371 11135
rect 18613 11101 18647 11135
rect 18705 11101 18739 11135
rect 19717 11101 19751 11135
rect 22109 11101 22143 11135
rect 22385 11101 22419 11135
rect 9413 11033 9447 11067
rect 9643 11033 9677 11067
rect 10701 11033 10735 11067
rect 13277 11033 13311 11067
rect 13369 11033 13403 11067
rect 14565 11033 14599 11067
rect 14657 11033 14691 11067
rect 16313 11033 16347 11067
rect 18889 11033 18923 11067
rect 20269 11033 20303 11067
rect 4169 10965 4203 10999
rect 11437 10965 11471 10999
rect 21373 10965 21407 10999
rect 1777 10761 1811 10795
rect 5289 10761 5323 10795
rect 6653 10761 6687 10795
rect 11161 10761 11195 10795
rect 13645 10761 13679 10795
rect 14473 10761 14507 10795
rect 15761 10761 15795 10795
rect 15945 10761 15979 10795
rect 19349 10761 19383 10795
rect 2237 10693 2271 10727
rect 4537 10693 4571 10727
rect 5089 10693 5123 10727
rect 7021 10693 7055 10727
rect 7159 10693 7193 10727
rect 9229 10693 9263 10727
rect 11989 10693 12023 10727
rect 13813 10693 13847 10727
rect 14013 10693 14047 10727
rect 15577 10693 15611 10727
rect 16129 10693 16163 10727
rect 17049 10693 17083 10727
rect 21281 10693 21315 10727
rect 23029 10693 23063 10727
rect 1961 10625 1995 10659
rect 2697 10625 2731 10659
rect 2881 10625 2915 10659
rect 3617 10625 3651 10659
rect 6837 10625 6871 10659
rect 6929 10625 6963 10659
rect 7941 10625 7975 10659
rect 8033 10625 8067 10659
rect 8125 10625 8159 10659
rect 9045 10625 9079 10659
rect 12449 10625 12483 10659
rect 12725 10625 12759 10659
rect 14749 10625 14783 10659
rect 14841 10625 14875 10659
rect 14933 10625 14967 10659
rect 15117 10625 15151 10659
rect 15853 10625 15887 10659
rect 17693 10625 17727 10659
rect 18061 10625 18095 10659
rect 18705 10625 18739 10659
rect 18889 10625 18923 10659
rect 19187 10625 19221 10659
rect 19901 10625 19935 10659
rect 20085 10625 20119 10659
rect 22293 10625 22327 10659
rect 2145 10557 2179 10591
rect 3525 10557 3559 10591
rect 7297 10557 7331 10591
rect 17601 10557 17635 10591
rect 18245 10557 18279 10591
rect 18981 10557 19015 10591
rect 22109 10557 22143 10591
rect 22201 10557 22235 10591
rect 22385 10557 22419 10591
rect 3985 10489 4019 10523
rect 9413 10489 9447 10523
rect 12633 10489 12667 10523
rect 19073 10489 19107 10523
rect 19993 10489 20027 10523
rect 2145 10421 2179 10455
rect 2881 10421 2915 10455
rect 5273 10421 5307 10455
rect 5457 10421 5491 10455
rect 6009 10421 6043 10455
rect 7757 10421 7791 10455
rect 10425 10421 10459 10455
rect 13829 10421 13863 10455
rect 20821 10421 20855 10455
rect 22569 10421 22603 10455
rect 4813 10217 4847 10251
rect 6193 10217 6227 10251
rect 8585 10217 8619 10251
rect 13553 10217 13587 10251
rect 14933 10217 14967 10251
rect 17693 10217 17727 10251
rect 21649 10217 21683 10251
rect 2237 10149 2271 10183
rect 4353 10149 4387 10183
rect 10517 10149 10551 10183
rect 12265 10149 12299 10183
rect 14381 10149 14415 10183
rect 19441 10149 19475 10183
rect 20637 10149 20671 10183
rect 6377 10081 6411 10115
rect 6653 10081 6687 10115
rect 7941 10081 7975 10115
rect 8125 10081 8159 10115
rect 12909 10081 12943 10115
rect 22661 10081 22695 10115
rect 2329 10013 2363 10047
rect 2513 10013 2547 10047
rect 3433 10013 3467 10047
rect 4997 10013 5031 10047
rect 5089 10013 5123 10047
rect 5319 10013 5353 10047
rect 5457 10013 5491 10047
rect 6469 10013 6503 10047
rect 6561 10013 6595 10047
rect 9137 10013 9171 10047
rect 9781 10013 9815 10047
rect 10701 10013 10735 10047
rect 11069 10013 11103 10047
rect 12449 10013 12483 10047
rect 12817 10013 12851 10047
rect 15117 10013 15151 10047
rect 15209 10013 15243 10047
rect 15393 10013 15427 10047
rect 15485 10013 15519 10047
rect 16129 10013 16163 10047
rect 16313 10013 16347 10047
rect 17141 10013 17175 10047
rect 17233 10013 17267 10047
rect 17417 10013 17451 10047
rect 17509 10013 17543 10047
rect 18153 10013 18187 10047
rect 18245 10013 18279 10047
rect 18429 10013 18463 10047
rect 19993 10013 20027 10047
rect 20177 10013 20211 10047
rect 20269 10013 20303 10047
rect 20361 10013 20395 10047
rect 21557 10013 21591 10047
rect 22385 10013 22419 10047
rect 22477 10013 22511 10047
rect 22569 10013 22603 10047
rect 3157 9945 3191 9979
rect 5181 9945 5215 9979
rect 9597 9945 9631 9979
rect 10793 9945 10827 9979
rect 10885 9945 10919 9979
rect 16681 9945 16715 9979
rect 1685 9877 1719 9911
rect 7389 9877 7423 9911
rect 8217 9877 8251 9911
rect 22201 9877 22235 9911
rect 23213 9877 23247 9911
rect 9045 9673 9079 9707
rect 14473 9673 14507 9707
rect 1685 9605 1719 9639
rect 2881 9605 2915 9639
rect 4629 9605 4663 9639
rect 5917 9605 5951 9639
rect 8309 9605 8343 9639
rect 12173 9605 12207 9639
rect 16129 9605 16163 9639
rect 18521 9605 18555 9639
rect 18705 9605 18739 9639
rect 22201 9605 22235 9639
rect 23121 9605 23155 9639
rect 1869 9537 1903 9571
rect 2053 9537 2087 9571
rect 3709 9537 3743 9571
rect 3801 9537 3835 9571
rect 4813 9537 4847 9571
rect 4905 9537 4939 9571
rect 5457 9537 5491 9571
rect 7665 9537 7699 9571
rect 7849 9537 7883 9571
rect 7941 9537 7975 9571
rect 8033 9537 8067 9571
rect 8861 9537 8895 9571
rect 10057 9537 10091 9571
rect 10977 9537 11011 9571
rect 13645 9537 13679 9571
rect 13921 9537 13955 9571
rect 15577 9537 15611 9571
rect 16865 9537 16899 9571
rect 17601 9537 17635 9571
rect 18245 9537 18279 9571
rect 19257 9537 19291 9571
rect 19533 9537 19567 9571
rect 20361 9537 20395 9571
rect 20453 9537 20487 9571
rect 20637 9537 20671 9571
rect 20729 9537 20763 9571
rect 22109 9537 22143 9571
rect 22385 9537 22419 9571
rect 3524 9469 3558 9503
rect 3617 9469 3651 9503
rect 5825 9469 5859 9503
rect 9321 9469 9355 9503
rect 10241 9469 10275 9503
rect 12541 9469 12575 9503
rect 17233 9469 17267 9503
rect 20177 9469 20211 9503
rect 2697 9401 2731 9435
rect 13093 9401 13127 9435
rect 13645 9401 13679 9435
rect 17141 9401 17175 9435
rect 19349 9401 19383 9435
rect 3985 9333 4019 9367
rect 4721 9333 4755 9367
rect 6653 9333 6687 9367
rect 7205 9333 7239 9367
rect 9873 9333 9907 9367
rect 11069 9333 11103 9367
rect 12633 9333 12667 9367
rect 12725 9333 12759 9367
rect 14933 9333 14967 9367
rect 17003 9333 17037 9367
rect 18521 9333 18555 9367
rect 19717 9333 19751 9367
rect 21189 9333 21223 9367
rect 22569 9333 22603 9367
rect 2145 9129 2179 9163
rect 6837 9129 6871 9163
rect 9873 9129 9907 9163
rect 14289 9129 14323 9163
rect 17233 9129 17267 9163
rect 22753 9129 22787 9163
rect 9689 9061 9723 9095
rect 11805 9061 11839 9095
rect 13277 9061 13311 9095
rect 14657 9061 14691 9095
rect 16865 9061 16899 9095
rect 21281 9061 21315 9095
rect 2605 8993 2639 9027
rect 6468 8993 6502 9027
rect 9229 8993 9263 9027
rect 16736 8993 16770 9027
rect 16957 8993 16991 9027
rect 18889 8993 18923 9027
rect 2329 8925 2363 8959
rect 3249 8925 3283 8959
rect 3433 8925 3467 8959
rect 3985 8925 4019 8959
rect 5365 8925 5399 8959
rect 6383 8925 6417 8959
rect 6560 8925 6594 8959
rect 6653 8925 6687 8959
rect 9873 8925 9907 8959
rect 10057 8925 10091 8959
rect 11069 8925 11103 8959
rect 11529 8925 11563 8959
rect 11621 8925 11655 8959
rect 12725 8925 12759 8959
rect 12817 8925 12851 8959
rect 13001 8925 13035 8959
rect 13093 8925 13127 8959
rect 14289 8925 14323 8959
rect 14381 8925 14415 8959
rect 15525 8925 15559 8959
rect 18245 8925 18279 8959
rect 19901 8925 19935 8959
rect 21189 8925 21223 8959
rect 21373 8925 21407 8959
rect 21465 8925 21499 8959
rect 21649 8925 21683 8959
rect 2421 8857 2455 8891
rect 3065 8857 3099 8891
rect 4261 8857 4295 8891
rect 5089 8857 5123 8891
rect 11805 8857 11839 8891
rect 15117 8857 15151 8891
rect 15301 8857 15335 8891
rect 15669 8857 15703 8891
rect 16589 8857 16623 8891
rect 20269 8857 20303 8891
rect 10977 8789 11011 8823
rect 15393 8789 15427 8823
rect 17969 8789 18003 8823
rect 21005 8789 21039 8823
rect 22201 8789 22235 8823
rect 23213 8789 23247 8823
rect 3801 8585 3835 8619
rect 9137 8585 9171 8619
rect 9597 8585 9631 8619
rect 11713 8585 11747 8619
rect 16313 8585 16347 8619
rect 7021 8517 7055 8551
rect 13093 8517 13127 8551
rect 15945 8517 15979 8551
rect 16145 8517 16179 8551
rect 19625 8517 19659 8551
rect 20361 8517 20395 8551
rect 21097 8517 21131 8551
rect 21281 8517 21315 8551
rect 1685 8449 1719 8483
rect 1869 8449 1903 8483
rect 2789 8449 2823 8483
rect 3341 8449 3375 8483
rect 3617 8449 3651 8483
rect 4905 8449 4939 8483
rect 6561 8449 6595 8483
rect 7481 8449 7515 8483
rect 8125 8449 8159 8483
rect 8585 8449 8619 8483
rect 10149 8449 10183 8483
rect 10333 8449 10367 8483
rect 11069 8449 11103 8483
rect 11897 8449 11931 8483
rect 11989 8449 12023 8483
rect 12173 8449 12207 8483
rect 12265 8449 12299 8483
rect 14197 8449 14231 8483
rect 14473 8449 14507 8483
rect 17509 8449 17543 8483
rect 18337 8449 18371 8483
rect 18797 8449 18831 8483
rect 21373 8449 21407 8483
rect 22477 8449 22511 8483
rect 22569 8449 22603 8483
rect 22845 8449 22879 8483
rect 2329 8381 2363 8415
rect 2881 8381 2915 8415
rect 3525 8381 3559 8415
rect 5181 8381 5215 8415
rect 8309 8381 8343 8415
rect 14105 8381 14139 8415
rect 14657 8381 14691 8415
rect 15209 8381 15243 8415
rect 17325 8381 17359 8415
rect 17785 8381 17819 8415
rect 22753 8381 22787 8415
rect 1869 8313 1903 8347
rect 10333 8313 10367 8347
rect 21097 8313 21131 8347
rect 22293 8313 22327 8347
rect 3341 8245 3375 8279
rect 7941 8245 7975 8279
rect 8125 8245 8159 8279
rect 16129 8245 16163 8279
rect 2421 8041 2455 8075
rect 4537 8041 4571 8075
rect 5733 8041 5767 8075
rect 7757 8041 7791 8075
rect 8125 8041 8159 8075
rect 10517 8041 10551 8075
rect 13645 8041 13679 8075
rect 18521 8041 18555 8075
rect 21005 8041 21039 8075
rect 22385 8041 22419 8075
rect 19625 7973 19659 8007
rect 3157 7905 3191 7939
rect 9413 7905 9447 7939
rect 10425 7905 10459 7939
rect 11805 7905 11839 7939
rect 14381 7905 14415 7939
rect 1961 7837 1995 7871
rect 2237 7837 2271 7871
rect 3341 7837 3375 7871
rect 4353 7837 4387 7871
rect 4445 7837 4479 7871
rect 5549 7837 5583 7871
rect 5733 7837 5767 7871
rect 6561 7837 6595 7871
rect 6837 7837 6871 7871
rect 8033 7837 8067 7871
rect 8125 7837 8159 7871
rect 9597 7837 9631 7871
rect 9965 7837 9999 7871
rect 10885 7837 10919 7871
rect 11897 7837 11931 7871
rect 13553 7837 13587 7871
rect 13737 7837 13771 7871
rect 14473 7837 14507 7871
rect 14749 7837 14783 7871
rect 14841 7837 14875 7871
rect 15945 7837 15979 7871
rect 16589 7837 16623 7871
rect 16957 7837 16991 7871
rect 17141 7837 17175 7871
rect 17325 7837 17359 7871
rect 17601 7837 17635 7871
rect 18061 7837 18095 7871
rect 19441 7837 19475 7871
rect 19625 7837 19659 7871
rect 20545 7837 20579 7871
rect 20821 7837 20855 7871
rect 22661 7837 22695 7871
rect 22753 7837 22787 7871
rect 22845 7837 22879 7871
rect 23029 7837 23063 7871
rect 5273 7769 5307 7803
rect 6745 7769 6779 7803
rect 7297 7769 7331 7803
rect 15485 7769 15519 7803
rect 20637 7769 20671 7803
rect 2053 7701 2087 7735
rect 4721 7701 4755 7735
rect 5917 7701 5951 7735
rect 9873 7701 9907 7735
rect 10701 7701 10735 7735
rect 10793 7701 10827 7735
rect 11161 7701 11195 7735
rect 12449 7701 12483 7735
rect 16037 7701 16071 7735
rect 21465 7701 21499 7735
rect 9965 7497 9999 7531
rect 11713 7497 11747 7531
rect 12725 7497 12759 7531
rect 14933 7497 14967 7531
rect 15025 7497 15059 7531
rect 23029 7497 23063 7531
rect 9137 7429 9171 7463
rect 9229 7429 9263 7463
rect 11069 7429 11103 7463
rect 14749 7429 14783 7463
rect 15301 7429 15335 7463
rect 20269 7429 20303 7463
rect 1777 7361 1811 7395
rect 1931 7361 1965 7395
rect 2881 7361 2915 7395
rect 3893 7361 3927 7395
rect 4353 7361 4387 7395
rect 5549 7361 5583 7395
rect 6653 7361 6687 7395
rect 8125 7361 8159 7395
rect 8217 7361 8251 7395
rect 8953 7361 8987 7395
rect 9321 7361 9355 7395
rect 10333 7361 10367 7395
rect 12081 7361 12115 7395
rect 12909 7361 12943 7395
rect 13185 7361 13219 7395
rect 15117 7361 15151 7395
rect 15945 7361 15979 7395
rect 17325 7361 17359 7395
rect 17509 7361 17543 7395
rect 18061 7361 18095 7395
rect 18245 7361 18279 7395
rect 19533 7361 19567 7395
rect 19809 7361 19843 7395
rect 20821 7361 20855 7395
rect 21005 7361 21039 7395
rect 22385 7361 22419 7395
rect 22569 7361 22603 7395
rect 22661 7361 22695 7395
rect 22799 7361 22833 7395
rect 4629 7293 4663 7327
rect 5365 7293 5399 7327
rect 6837 7293 6871 7327
rect 8033 7293 8067 7327
rect 8309 7293 8343 7327
rect 8493 7293 8527 7327
rect 10241 7293 10275 7327
rect 11889 7293 11923 7327
rect 11989 7293 12023 7327
rect 12173 7293 12207 7327
rect 13093 7293 13127 7327
rect 2145 7225 2179 7259
rect 4537 7225 4571 7259
rect 9505 7225 9539 7259
rect 19625 7225 19659 7259
rect 21005 7225 21039 7259
rect 2973 7157 3007 7191
rect 3801 7157 3835 7191
rect 4445 7157 4479 7191
rect 10333 7157 10367 7191
rect 12909 7157 12943 7191
rect 13829 7157 13863 7191
rect 15945 7157 15979 7191
rect 18521 7157 18555 7191
rect 2421 6953 2455 6987
rect 8493 6953 8527 6987
rect 15669 6953 15703 6987
rect 16405 6953 16439 6987
rect 22477 6953 22511 6987
rect 10517 6885 10551 6919
rect 11345 6885 11379 6919
rect 13277 6885 13311 6919
rect 14473 6885 14507 6919
rect 22385 6885 22419 6919
rect 3433 6817 3467 6851
rect 5365 6817 5399 6851
rect 5825 6817 5859 6851
rect 9597 6817 9631 6851
rect 9689 6817 9723 6851
rect 9965 6817 9999 6851
rect 17049 6817 17083 6851
rect 17601 6817 17635 6851
rect 18245 6817 18279 6851
rect 20361 6817 20395 6851
rect 22293 6817 22327 6851
rect 23213 6817 23247 6851
rect 2053 6749 2087 6783
rect 2421 6749 2455 6783
rect 3065 6749 3099 6783
rect 3249 6749 3283 6783
rect 4629 6749 4663 6783
rect 5733 6749 5767 6783
rect 6101 6749 6135 6783
rect 6285 6749 6319 6783
rect 7205 6749 7239 6783
rect 7389 6749 7423 6783
rect 7665 6749 7699 6783
rect 7757 6749 7791 6783
rect 8309 6749 8343 6783
rect 9505 6749 9539 6783
rect 9781 6749 9815 6783
rect 14933 6749 14967 6783
rect 15117 6749 15151 6783
rect 18337 6749 18371 6783
rect 18889 6749 18923 6783
rect 19441 6749 19475 6783
rect 19625 6749 19659 6783
rect 19993 6749 20027 6783
rect 20177 6749 20211 6783
rect 21373 6749 21407 6783
rect 22661 6749 22695 6783
rect 4353 6681 4387 6715
rect 15025 6681 15059 6715
rect 21649 6681 21683 6715
rect 2605 6613 2639 6647
rect 11805 6613 11839 6647
rect 22569 6613 22603 6647
rect 3433 6409 3467 6443
rect 6745 6409 6779 6443
rect 6837 6409 6871 6443
rect 9781 6409 9815 6443
rect 11069 6409 11103 6443
rect 13737 6409 13771 6443
rect 18337 6409 18371 6443
rect 22017 6409 22051 6443
rect 23029 6409 23063 6443
rect 4169 6341 4203 6375
rect 4629 6341 4663 6375
rect 6009 6341 6043 6375
rect 6929 6341 6963 6375
rect 7113 6341 7147 6375
rect 8309 6341 8343 6375
rect 12909 6341 12943 6375
rect 15117 6341 15151 6375
rect 15669 6341 15703 6375
rect 21281 6341 21315 6375
rect 2237 6273 2271 6307
rect 2421 6273 2455 6307
rect 2697 6273 2731 6307
rect 2789 6273 2823 6307
rect 3065 6273 3099 6307
rect 4261 6273 4295 6307
rect 5273 6273 5307 6307
rect 5549 6273 5583 6307
rect 6561 6273 6595 6307
rect 8033 6273 8067 6307
rect 8126 6273 8160 6307
rect 8398 6273 8432 6307
rect 8498 6273 8532 6307
rect 9137 6273 9171 6307
rect 9321 6273 9355 6307
rect 9413 6273 9447 6307
rect 9505 6273 9539 6307
rect 10885 6273 10919 6307
rect 11161 6273 11195 6307
rect 11713 6273 11747 6307
rect 11897 6273 11931 6307
rect 12081 6273 12115 6307
rect 12173 6273 12207 6307
rect 12817 6273 12851 6307
rect 13001 6273 13035 6307
rect 13139 6273 13173 6307
rect 13921 6273 13955 6307
rect 14197 6273 14231 6307
rect 15209 6273 15243 6307
rect 17877 6273 17911 6307
rect 17969 6273 18003 6307
rect 18153 6273 18187 6307
rect 19257 6273 19291 6307
rect 19809 6273 19843 6307
rect 20913 6273 20947 6307
rect 21189 6273 21223 6307
rect 22201 6273 22235 6307
rect 22385 6273 22419 6307
rect 22937 6273 22971 6307
rect 23121 6273 23155 6307
rect 4721 6205 4755 6239
rect 5365 6205 5399 6239
rect 13277 6205 13311 6239
rect 14105 6205 14139 6239
rect 20361 6205 20395 6239
rect 22477 6205 22511 6239
rect 8677 6137 8711 6171
rect 12633 6137 12667 6171
rect 14933 6137 14967 6171
rect 10701 6069 10735 6103
rect 16129 6069 16163 6103
rect 16865 6069 16899 6103
rect 2053 5865 2087 5899
rect 3985 5865 4019 5899
rect 9229 5865 9263 5899
rect 12357 5865 12391 5899
rect 18429 5865 18463 5899
rect 18613 5865 18647 5899
rect 21649 5865 21683 5899
rect 22569 5865 22603 5899
rect 2329 5797 2363 5831
rect 6285 5797 6319 5831
rect 11253 5797 11287 5831
rect 12817 5797 12851 5831
rect 14657 5797 14691 5831
rect 15209 5797 15243 5831
rect 19901 5797 19935 5831
rect 8033 5729 8067 5763
rect 10701 5729 10735 5763
rect 13001 5729 13035 5763
rect 13093 5729 13127 5763
rect 15853 5729 15887 5763
rect 16773 5729 16807 5763
rect 17233 5729 17267 5763
rect 17969 5729 18003 5763
rect 20545 5729 20579 5763
rect 22937 5729 22971 5763
rect 1869 5661 1903 5695
rect 2053 5661 2087 5695
rect 2145 5661 2179 5695
rect 3157 5661 3191 5695
rect 3341 5661 3375 5695
rect 5089 5661 5123 5695
rect 5273 5661 5307 5695
rect 6101 5661 6135 5695
rect 7021 5661 7055 5695
rect 7205 5661 7239 5695
rect 7757 5661 7791 5695
rect 7941 5661 7975 5695
rect 8125 5661 8159 5695
rect 8309 5661 8343 5695
rect 10149 5661 10183 5695
rect 10241 5661 10275 5695
rect 10425 5661 10459 5695
rect 10517 5661 10551 5695
rect 11713 5661 11747 5695
rect 11897 5661 11931 5695
rect 11989 5661 12023 5695
rect 12081 5661 12115 5695
rect 13185 5661 13219 5695
rect 13277 5661 13311 5695
rect 14289 5661 14323 5695
rect 14473 5661 14507 5695
rect 14749 5661 14783 5695
rect 15209 5661 15243 5695
rect 15393 5661 15427 5695
rect 16037 5661 16071 5695
rect 16221 5661 16255 5695
rect 16957 5661 16991 5695
rect 17325 5661 17359 5695
rect 19809 5661 19843 5695
rect 20085 5661 20119 5695
rect 21005 5661 21039 5695
rect 21189 5661 21223 5695
rect 21281 5661 21315 5695
rect 21419 5661 21453 5695
rect 22753 5661 22787 5695
rect 2881 5593 2915 5627
rect 4169 5593 4203 5627
rect 4353 5593 4387 5627
rect 7113 5593 7147 5627
rect 18797 5593 18831 5627
rect 2973 5525 3007 5559
rect 8493 5525 8527 5559
rect 18587 5525 18621 5559
rect 2513 5321 2547 5355
rect 5825 5321 5859 5355
rect 6837 5321 6871 5355
rect 14749 5321 14783 5355
rect 15669 5321 15703 5355
rect 21373 5321 21407 5355
rect 22109 5321 22143 5355
rect 4353 5253 4387 5287
rect 12449 5253 12483 5287
rect 13645 5253 13679 5287
rect 14657 5253 14691 5287
rect 15117 5253 15151 5287
rect 16313 5253 16347 5287
rect 19533 5253 19567 5287
rect 20729 5253 20763 5287
rect 22569 5253 22603 5287
rect 1961 5185 1995 5219
rect 2053 5185 2087 5219
rect 2237 5185 2271 5219
rect 2329 5185 2363 5219
rect 3433 5185 3467 5219
rect 5733 5185 5767 5219
rect 6561 5185 6595 5219
rect 6745 5185 6779 5219
rect 7665 5185 7699 5219
rect 7941 5185 7975 5219
rect 8585 5185 8619 5219
rect 14933 5185 14967 5219
rect 15945 5185 15979 5219
rect 16221 5185 16255 5219
rect 17417 5185 17451 5219
rect 17785 5185 17819 5219
rect 19441 5185 19475 5219
rect 20545 5185 20579 5219
rect 22753 5185 22787 5219
rect 22845 5185 22879 5219
rect 3157 5117 3191 5151
rect 5089 5117 5123 5151
rect 9689 5117 9723 5151
rect 15854 5117 15888 5151
rect 17233 5117 17267 5151
rect 17693 5117 17727 5151
rect 18337 5117 18371 5151
rect 19533 5117 19567 5151
rect 8585 5049 8619 5083
rect 9137 4981 9171 5015
rect 13093 4981 13127 5015
rect 14197 4981 14231 5015
rect 19993 4981 20027 5015
rect 20913 4981 20947 5015
rect 1869 4777 1903 4811
rect 2697 4777 2731 4811
rect 9597 4777 9631 4811
rect 11253 4777 11287 4811
rect 12725 4777 12759 4811
rect 16865 4777 16899 4811
rect 20545 4777 20579 4811
rect 10057 4709 10091 4743
rect 21097 4709 21131 4743
rect 6837 4641 6871 4675
rect 9137 4641 9171 4675
rect 9229 4641 9263 4675
rect 10701 4641 10735 4675
rect 22109 4641 22143 4675
rect 2329 4573 2363 4607
rect 2789 4573 2823 4607
rect 4445 4573 4479 4607
rect 4537 4573 4571 4607
rect 4997 4573 5031 4607
rect 5733 4573 5767 4607
rect 5917 4573 5951 4607
rect 6377 4573 6411 4607
rect 6561 4573 6595 4607
rect 6929 4573 6963 4607
rect 8033 4573 8067 4607
rect 9413 4573 9447 4607
rect 10241 4573 10275 4607
rect 10333 4573 10367 4607
rect 10609 4573 10643 4607
rect 12265 4573 12299 4607
rect 12541 4573 12575 4607
rect 13369 4573 13403 4607
rect 13737 4573 13771 4607
rect 14381 4573 14415 4607
rect 15485 4573 15519 4607
rect 16221 4573 16255 4607
rect 16314 4573 16348 4607
rect 16497 4573 16531 4607
rect 16727 4573 16761 4607
rect 17877 4573 17911 4607
rect 19441 4573 19475 4607
rect 19717 4573 19751 4607
rect 20453 4573 20487 4607
rect 22661 4573 22695 4607
rect 23029 4573 23063 4607
rect 4261 4505 4295 4539
rect 4629 4505 4663 4539
rect 7573 4505 7607 4539
rect 12357 4505 12391 4539
rect 13461 4505 13495 4539
rect 13553 4505 13587 4539
rect 16589 4505 16623 4539
rect 19533 4505 19567 4539
rect 19901 4505 19935 4539
rect 3433 4437 3467 4471
rect 5825 4437 5859 4471
rect 13185 4437 13219 4471
rect 14933 4437 14967 4471
rect 17417 4437 17451 4471
rect 18889 4437 18923 4471
rect 6745 4233 6779 4267
rect 8493 4233 8527 4267
rect 10885 4233 10919 4267
rect 12081 4233 12115 4267
rect 14013 4233 14047 4267
rect 14565 4233 14599 4267
rect 17969 4233 18003 4267
rect 18521 4233 18555 4267
rect 5733 4165 5767 4199
rect 6653 4165 6687 4199
rect 18889 4165 18923 4199
rect 1869 4097 1903 4131
rect 2145 4097 2179 4131
rect 2605 4097 2639 4131
rect 2697 4097 2731 4131
rect 4629 4097 4663 4131
rect 5181 4097 5215 4131
rect 5365 4097 5399 4131
rect 6837 4097 6871 4131
rect 7389 4097 7423 4131
rect 8401 4097 8435 4131
rect 8585 4097 8619 4131
rect 10701 4097 10735 4131
rect 10793 4097 10827 4131
rect 11713 4097 11747 4131
rect 11989 4097 12023 4131
rect 12909 4097 12943 4131
rect 15761 4097 15795 4131
rect 15853 4097 15887 4131
rect 15945 4097 15979 4131
rect 16129 4097 16163 4131
rect 16865 4097 16899 4131
rect 17417 4097 17451 4131
rect 18705 4097 18739 4131
rect 18797 4097 18831 4131
rect 19073 4097 19107 4131
rect 19993 4097 20027 4131
rect 20177 4097 20211 4131
rect 20361 4097 20395 4131
rect 20545 4097 20579 4131
rect 20821 4097 20855 4131
rect 22753 4097 22787 4131
rect 4353 4029 4387 4063
rect 7205 4029 7239 4063
rect 11161 4029 11195 4063
rect 11885 4029 11919 4063
rect 12265 4029 12299 4063
rect 12357 4029 12391 4063
rect 15485 4029 15519 4063
rect 19533 4029 19567 4063
rect 2053 3961 2087 3995
rect 9045 3961 9079 3995
rect 1685 3893 1719 3927
rect 2881 3893 2915 3927
rect 3709 3893 3743 3927
rect 7849 3893 7883 3927
rect 9689 3893 9723 3927
rect 13461 3893 13495 3927
rect 22293 3893 22327 3927
rect 4077 3689 4111 3723
rect 7389 3689 7423 3723
rect 9413 3689 9447 3723
rect 13737 3689 13771 3723
rect 15209 3689 15243 3723
rect 18061 3689 18095 3723
rect 21833 3689 21867 3723
rect 22385 3689 22419 3723
rect 5733 3621 5767 3655
rect 9505 3621 9539 3655
rect 14289 3621 14323 3655
rect 19533 3621 19567 3655
rect 4997 3553 5031 3587
rect 10333 3553 10367 3587
rect 12081 3553 12115 3587
rect 12173 3553 12207 3587
rect 12265 3553 12299 3587
rect 18705 3553 18739 3587
rect 2053 3485 2087 3519
rect 2421 3485 2455 3519
rect 2513 3485 2547 3519
rect 2697 3485 2731 3519
rect 2861 3485 2895 3519
rect 4813 3485 4847 3519
rect 6285 3485 6319 3519
rect 6929 3485 6963 3519
rect 7113 3485 7147 3519
rect 8309 3485 8343 3519
rect 8493 3485 8527 3519
rect 8585 3485 8619 3519
rect 9137 3485 9171 3519
rect 9321 3485 9355 3519
rect 9597 3485 9631 3519
rect 11713 3485 11747 3519
rect 13461 3485 13495 3519
rect 13553 3485 13587 3519
rect 14565 3485 14599 3519
rect 14749 3485 14783 3519
rect 15853 3485 15887 3519
rect 16129 3485 16163 3519
rect 16589 3485 16623 3519
rect 16957 3485 16991 3519
rect 17325 3485 17359 3519
rect 18245 3485 18279 3519
rect 18547 3485 18581 3519
rect 19441 3485 19475 3519
rect 20177 3485 20211 3519
rect 20361 3485 20395 3519
rect 20729 3485 20763 3519
rect 21189 3485 21223 3519
rect 23305 3485 23339 3519
rect 3341 3417 3375 3451
rect 4905 3417 4939 3451
rect 5273 3417 5307 3451
rect 9873 3417 9907 3451
rect 13093 3417 13127 3451
rect 15761 3417 15795 3451
rect 18337 3417 18371 3451
rect 18429 3417 18463 3451
rect 11161 3349 11195 3383
rect 14473 3349 14507 3383
rect 2605 3145 2639 3179
rect 8401 3145 8435 3179
rect 9873 3145 9907 3179
rect 11713 3145 11747 3179
rect 12817 3145 12851 3179
rect 13645 3145 13679 3179
rect 14197 3145 14231 3179
rect 14749 3145 14783 3179
rect 16865 3145 16899 3179
rect 18245 3145 18279 3179
rect 20361 3145 20395 3179
rect 6745 3077 6779 3111
rect 9229 3077 9263 3111
rect 10333 3077 10367 3111
rect 18613 3077 18647 3111
rect 20177 3077 20211 3111
rect 2237 3009 2271 3043
rect 2329 3009 2363 3043
rect 2421 3009 2455 3043
rect 3525 3009 3559 3043
rect 3985 3009 4019 3043
rect 4169 3009 4203 3043
rect 4445 3009 4479 3043
rect 4629 3009 4663 3043
rect 5273 3009 5307 3043
rect 5825 3009 5859 3043
rect 7021 3009 7055 3043
rect 8309 3009 8343 3043
rect 8493 3009 8527 3043
rect 9597 3009 9631 3043
rect 10609 3009 10643 3043
rect 12449 3009 12483 3043
rect 12633 3009 12667 3043
rect 14657 3009 14691 3043
rect 14841 3009 14875 3043
rect 15761 3009 15795 3043
rect 15945 3009 15979 3043
rect 17049 3009 17083 3043
rect 17325 3009 17359 3043
rect 18429 3009 18463 3043
rect 18705 3009 18739 3043
rect 19993 3009 20027 3043
rect 3341 2941 3375 2975
rect 5365 2941 5399 2975
rect 5641 2941 5675 2975
rect 9689 2941 9723 2975
rect 10333 2941 10367 2975
rect 4261 2873 4295 2907
rect 4353 2873 4387 2907
rect 7849 2873 7883 2907
rect 10517 2873 10551 2907
rect 11161 2873 11195 2907
rect 20821 2873 20855 2907
rect 1685 2805 1719 2839
rect 15853 2805 15887 2839
rect 17233 2805 17267 2839
rect 19165 2805 19199 2839
rect 22017 2805 22051 2839
rect 22845 2805 22879 2839
rect 5365 2601 5399 2635
rect 6009 2601 6043 2635
rect 16313 2601 16347 2635
rect 18797 2601 18831 2635
rect 19441 2601 19475 2635
rect 21373 2601 21407 2635
rect 4997 2533 5031 2567
rect 5085 2533 5119 2567
rect 4077 2465 4111 2499
rect 7665 2465 7699 2499
rect 17509 2465 17543 2499
rect 20085 2465 20119 2499
rect 2513 2397 2547 2431
rect 3433 2397 3467 2431
rect 4261 2397 4295 2431
rect 4905 2397 4939 2431
rect 5181 2397 5215 2431
rect 7021 2397 7055 2431
rect 7481 2397 7515 2431
rect 8585 2397 8619 2431
rect 9873 2397 9907 2431
rect 10517 2397 10551 2431
rect 11161 2397 11195 2431
rect 11897 2397 11931 2431
rect 12541 2397 12575 2431
rect 13185 2397 13219 2431
rect 14289 2397 14323 2431
rect 14933 2397 14967 2431
rect 15577 2397 15611 2431
rect 16865 2397 16899 2431
rect 18153 2397 18187 2431
rect 20729 2397 20763 2431
rect 22017 2397 22051 2431
rect 22661 2397 22695 2431
rect 2237 2329 2271 2363
rect 3157 2329 3191 2363
rect 6745 2329 6779 2363
rect 9137 2329 9171 2363
<< metal1 >>
rect 1104 22330 23828 22352
rect 1104 22278 3790 22330
rect 3842 22278 3854 22330
rect 3906 22278 3918 22330
rect 3970 22278 3982 22330
rect 4034 22278 4046 22330
rect 4098 22278 9471 22330
rect 9523 22278 9535 22330
rect 9587 22278 9599 22330
rect 9651 22278 9663 22330
rect 9715 22278 9727 22330
rect 9779 22278 15152 22330
rect 15204 22278 15216 22330
rect 15268 22278 15280 22330
rect 15332 22278 15344 22330
rect 15396 22278 15408 22330
rect 15460 22278 20833 22330
rect 20885 22278 20897 22330
rect 20949 22278 20961 22330
rect 21013 22278 21025 22330
rect 21077 22278 21089 22330
rect 21141 22278 23828 22330
rect 1104 22256 23828 22278
rect 12805 22083 12863 22089
rect 12805 22049 12817 22083
rect 12851 22080 12863 22083
rect 21174 22080 21180 22092
rect 12851 22052 21180 22080
rect 12851 22049 12863 22052
rect 12805 22043 12863 22049
rect 21174 22040 21180 22052
rect 21232 22040 21238 22092
rect 10502 22012 10508 22024
rect 10463 21984 10508 22012
rect 10502 21972 10508 21984
rect 10560 21972 10566 22024
rect 19978 22012 19984 22024
rect 12406 21984 19984 22012
rect 7101 21947 7159 21953
rect 7101 21913 7113 21947
rect 7147 21944 7159 21947
rect 7466 21944 7472 21956
rect 7147 21916 7472 21944
rect 7147 21913 7159 21916
rect 7101 21907 7159 21913
rect 7466 21904 7472 21916
rect 7524 21944 7530 21956
rect 7653 21947 7711 21953
rect 7653 21944 7665 21947
rect 7524 21916 7665 21944
rect 7524 21904 7530 21916
rect 7653 21913 7665 21916
rect 7699 21913 7711 21947
rect 7653 21907 7711 21913
rect 10260 21947 10318 21953
rect 10260 21913 10272 21947
rect 10306 21944 10318 21947
rect 12406 21944 12434 21984
rect 19978 21972 19984 21984
rect 20036 21972 20042 22024
rect 21453 22015 21511 22021
rect 21453 21981 21465 22015
rect 21499 22012 21511 22015
rect 22370 22012 22376 22024
rect 21499 21984 22376 22012
rect 21499 21981 21511 21984
rect 21453 21975 21511 21981
rect 22370 21972 22376 21984
rect 22428 22012 22434 22024
rect 22649 22015 22707 22021
rect 22649 22012 22661 22015
rect 22428 21984 22661 22012
rect 22428 21972 22434 21984
rect 22649 21981 22661 21984
rect 22695 21981 22707 22015
rect 22649 21975 22707 21981
rect 10306 21916 12434 21944
rect 12621 21947 12679 21953
rect 10306 21913 10318 21916
rect 10260 21907 10318 21913
rect 12621 21913 12633 21947
rect 12667 21913 12679 21947
rect 12621 21907 12679 21913
rect 17037 21947 17095 21953
rect 17037 21913 17049 21947
rect 17083 21944 17095 21947
rect 17402 21944 17408 21956
rect 17083 21916 17408 21944
rect 17083 21913 17095 21916
rect 17037 21907 17095 21913
rect 6270 21836 6276 21888
rect 6328 21876 6334 21888
rect 7745 21879 7803 21885
rect 7745 21876 7757 21879
rect 6328 21848 7757 21876
rect 6328 21836 6334 21848
rect 7745 21845 7757 21848
rect 7791 21845 7803 21879
rect 7745 21839 7803 21845
rect 8938 21836 8944 21888
rect 8996 21876 9002 21888
rect 9125 21879 9183 21885
rect 9125 21876 9137 21879
rect 8996 21848 9137 21876
rect 8996 21836 9002 21848
rect 9125 21845 9137 21848
rect 9171 21845 9183 21879
rect 9125 21839 9183 21845
rect 11057 21879 11115 21885
rect 11057 21845 11069 21879
rect 11103 21876 11115 21879
rect 11330 21876 11336 21888
rect 11103 21848 11336 21876
rect 11103 21845 11115 21848
rect 11057 21839 11115 21845
rect 11330 21836 11336 21848
rect 11388 21836 11394 21888
rect 12069 21879 12127 21885
rect 12069 21845 12081 21879
rect 12115 21876 12127 21879
rect 12434 21876 12440 21888
rect 12115 21848 12440 21876
rect 12115 21845 12127 21848
rect 12069 21839 12127 21845
rect 12434 21836 12440 21848
rect 12492 21876 12498 21888
rect 12636 21876 12664 21907
rect 17402 21904 17408 21916
rect 17460 21944 17466 21956
rect 17589 21947 17647 21953
rect 17589 21944 17601 21947
rect 17460 21916 17601 21944
rect 17460 21904 17466 21916
rect 17589 21913 17601 21916
rect 17635 21913 17647 21947
rect 17589 21907 17647 21913
rect 12492 21848 12664 21876
rect 12492 21836 12498 21848
rect 13998 21836 14004 21888
rect 14056 21876 14062 21888
rect 14277 21879 14335 21885
rect 14277 21876 14289 21879
rect 14056 21848 14289 21876
rect 14056 21836 14062 21848
rect 14277 21845 14289 21848
rect 14323 21845 14335 21879
rect 14277 21839 14335 21845
rect 14921 21879 14979 21885
rect 14921 21845 14933 21879
rect 14967 21876 14979 21879
rect 15102 21876 15108 21888
rect 14967 21848 15108 21876
rect 14967 21845 14979 21848
rect 14921 21839 14979 21845
rect 15102 21836 15108 21848
rect 15160 21836 15166 21888
rect 15654 21876 15660 21888
rect 15615 21848 15660 21876
rect 15654 21836 15660 21848
rect 15712 21836 15718 21888
rect 17678 21876 17684 21888
rect 17639 21848 17684 21876
rect 17678 21836 17684 21848
rect 17736 21836 17742 21888
rect 22370 21836 22376 21888
rect 22428 21876 22434 21888
rect 22557 21879 22615 21885
rect 22557 21876 22569 21879
rect 22428 21848 22569 21876
rect 22428 21836 22434 21848
rect 22557 21845 22569 21848
rect 22603 21845 22615 21879
rect 22557 21839 22615 21845
rect 1104 21786 23987 21808
rect 1104 21734 6630 21786
rect 6682 21734 6694 21786
rect 6746 21734 6758 21786
rect 6810 21734 6822 21786
rect 6874 21734 6886 21786
rect 6938 21734 12311 21786
rect 12363 21734 12375 21786
rect 12427 21734 12439 21786
rect 12491 21734 12503 21786
rect 12555 21734 12567 21786
rect 12619 21734 17992 21786
rect 18044 21734 18056 21786
rect 18108 21734 18120 21786
rect 18172 21734 18184 21786
rect 18236 21734 18248 21786
rect 18300 21734 23673 21786
rect 23725 21734 23737 21786
rect 23789 21734 23801 21786
rect 23853 21734 23865 21786
rect 23917 21734 23929 21786
rect 23981 21734 23987 21786
rect 1104 21712 23987 21734
rect 2498 21632 2504 21684
rect 2556 21672 2562 21684
rect 5810 21672 5816 21684
rect 2556 21644 5816 21672
rect 2556 21632 2562 21644
rect 5810 21632 5816 21644
rect 5868 21632 5874 21684
rect 17681 21675 17739 21681
rect 17681 21672 17693 21675
rect 11992 21644 17693 21672
rect 5350 21604 5356 21616
rect 2516 21576 5356 21604
rect 2038 21428 2044 21480
rect 2096 21468 2102 21480
rect 2516 21477 2544 21576
rect 2774 21545 2780 21548
rect 2768 21499 2780 21545
rect 2832 21536 2838 21548
rect 4632 21545 4660 21576
rect 5350 21564 5356 21576
rect 5408 21564 5414 21616
rect 9122 21564 9128 21616
rect 9180 21604 9186 21616
rect 11992 21604 12020 21644
rect 17681 21641 17693 21644
rect 17727 21641 17739 21675
rect 19150 21672 19156 21684
rect 17681 21635 17739 21641
rect 18248 21644 19156 21672
rect 13814 21604 13820 21616
rect 9180 21576 10364 21604
rect 9180 21564 9186 21576
rect 4617 21539 4675 21545
rect 2832 21508 2868 21536
rect 2774 21496 2780 21499
rect 2832 21496 2838 21508
rect 4617 21505 4629 21539
rect 4663 21505 4675 21539
rect 4617 21499 4675 21505
rect 4884 21539 4942 21545
rect 4884 21505 4896 21539
rect 4930 21536 4942 21539
rect 5442 21536 5448 21548
rect 4930 21508 5448 21536
rect 4930 21505 4942 21508
rect 4884 21499 4942 21505
rect 5442 21496 5448 21508
rect 5500 21496 5506 21548
rect 10336 21545 10364 21576
rect 10612 21576 12020 21604
rect 12820 21576 13820 21604
rect 10065 21539 10123 21545
rect 10065 21505 10077 21539
rect 10111 21536 10123 21539
rect 10321 21539 10379 21545
rect 10111 21508 10272 21536
rect 10111 21505 10123 21508
rect 10065 21499 10123 21505
rect 2501 21471 2559 21477
rect 2501 21468 2513 21471
rect 2096 21440 2513 21468
rect 2096 21428 2102 21440
rect 2501 21437 2513 21440
rect 2547 21437 2559 21471
rect 10244 21468 10272 21508
rect 10321 21505 10333 21539
rect 10367 21536 10379 21539
rect 10502 21536 10508 21548
rect 10367 21508 10508 21536
rect 10367 21505 10379 21508
rect 10321 21499 10379 21505
rect 10502 21496 10508 21508
rect 10560 21496 10566 21548
rect 10612 21468 10640 21576
rect 12069 21539 12127 21545
rect 12069 21505 12081 21539
rect 12115 21505 12127 21539
rect 12069 21499 12127 21505
rect 10244 21440 10640 21468
rect 2501 21431 2559 21437
rect 1854 21292 1860 21344
rect 1912 21332 1918 21344
rect 3881 21335 3939 21341
rect 3881 21332 3893 21335
rect 1912 21304 3893 21332
rect 1912 21292 1918 21304
rect 3881 21301 3893 21304
rect 3927 21301 3939 21335
rect 3881 21295 3939 21301
rect 5997 21335 6055 21341
rect 5997 21301 6009 21335
rect 6043 21332 6055 21335
rect 6178 21332 6184 21344
rect 6043 21304 6184 21332
rect 6043 21301 6055 21304
rect 5997 21295 6055 21301
rect 6178 21292 6184 21304
rect 6236 21292 6242 21344
rect 8846 21292 8852 21344
rect 8904 21332 8910 21344
rect 8941 21335 8999 21341
rect 8941 21332 8953 21335
rect 8904 21304 8953 21332
rect 8904 21292 8910 21304
rect 8941 21301 8953 21304
rect 8987 21301 8999 21335
rect 8941 21295 8999 21301
rect 11149 21335 11207 21341
rect 11149 21301 11161 21335
rect 11195 21332 11207 21335
rect 11330 21332 11336 21344
rect 11195 21304 11336 21332
rect 11195 21301 11207 21304
rect 11149 21295 11207 21301
rect 11330 21292 11336 21304
rect 11388 21292 11394 21344
rect 11790 21292 11796 21344
rect 11848 21332 11854 21344
rect 12084 21332 12112 21499
rect 12161 21403 12219 21409
rect 12161 21369 12173 21403
rect 12207 21400 12219 21403
rect 12820 21400 12848 21576
rect 13814 21564 13820 21576
rect 13872 21564 13878 21616
rect 14550 21564 14556 21616
rect 14608 21604 14614 21616
rect 16117 21607 16175 21613
rect 14608 21576 15240 21604
rect 14608 21564 14614 21576
rect 13078 21536 13084 21548
rect 13039 21508 13084 21536
rect 13078 21496 13084 21508
rect 13136 21496 13142 21548
rect 13998 21496 14004 21548
rect 14056 21496 14062 21548
rect 14090 21496 14096 21548
rect 14148 21536 14154 21548
rect 14185 21539 14243 21545
rect 14185 21536 14197 21539
rect 14148 21508 14197 21536
rect 14148 21496 14154 21508
rect 14185 21505 14197 21508
rect 14231 21505 14243 21539
rect 15102 21536 15108 21548
rect 14185 21499 14243 21505
rect 14292 21508 15108 21536
rect 13262 21428 13268 21480
rect 13320 21468 13326 21480
rect 13909 21471 13967 21477
rect 13909 21468 13921 21471
rect 13320 21440 13921 21468
rect 13320 21428 13326 21440
rect 13909 21437 13921 21440
rect 13955 21468 13967 21471
rect 14016 21468 14044 21496
rect 13955 21440 14044 21468
rect 13955 21437 13967 21440
rect 13909 21431 13967 21437
rect 12207 21372 12848 21400
rect 12207 21369 12219 21372
rect 12161 21363 12219 21369
rect 12894 21360 12900 21412
rect 12952 21400 12958 21412
rect 14292 21400 14320 21508
rect 15102 21496 15108 21508
rect 15160 21496 15166 21548
rect 15212 21536 15240 21576
rect 16117 21573 16129 21607
rect 16163 21604 16175 21607
rect 18248 21604 18276 21644
rect 19150 21632 19156 21644
rect 19208 21632 19214 21684
rect 19978 21672 19984 21684
rect 19939 21644 19984 21672
rect 19978 21632 19984 21644
rect 20036 21632 20042 21684
rect 21174 21632 21180 21684
rect 21232 21672 21238 21684
rect 21232 21644 22094 21672
rect 21232 21632 21238 21644
rect 16163 21576 18276 21604
rect 18325 21607 18383 21613
rect 16163 21573 16175 21576
rect 16117 21567 16175 21573
rect 18325 21573 18337 21607
rect 18371 21604 18383 21607
rect 22066 21604 22094 21644
rect 22189 21607 22247 21613
rect 22189 21604 22201 21607
rect 18371 21576 21312 21604
rect 22066 21576 22201 21604
rect 18371 21573 18383 21576
rect 18325 21567 18383 21573
rect 21284 21548 21312 21576
rect 22189 21573 22201 21576
rect 22235 21573 22247 21607
rect 22189 21567 22247 21573
rect 17034 21536 17040 21548
rect 15212 21508 17040 21536
rect 17034 21496 17040 21508
rect 17092 21496 17098 21548
rect 17678 21496 17684 21548
rect 17736 21536 17742 21548
rect 17957 21539 18015 21545
rect 17957 21536 17969 21539
rect 17736 21508 17969 21536
rect 17736 21496 17742 21508
rect 17957 21505 17969 21508
rect 18003 21536 18015 21539
rect 20271 21539 20329 21545
rect 20271 21536 20283 21539
rect 18003 21508 20283 21536
rect 18003 21505 18015 21508
rect 17957 21499 18015 21505
rect 20271 21505 20283 21508
rect 20317 21505 20329 21539
rect 21085 21539 21143 21545
rect 21085 21536 21097 21539
rect 20271 21499 20329 21505
rect 20364 21508 21097 21536
rect 14918 21468 14924 21480
rect 14879 21440 14924 21468
rect 14918 21428 14924 21440
rect 14976 21428 14982 21480
rect 15010 21428 15016 21480
rect 15068 21468 15074 21480
rect 15197 21471 15255 21477
rect 15068 21440 15113 21468
rect 15068 21428 15074 21440
rect 15197 21437 15209 21471
rect 15243 21468 15255 21471
rect 17865 21471 17923 21477
rect 15243 21440 16344 21468
rect 15243 21437 15255 21440
rect 15197 21431 15255 21437
rect 12952 21372 14320 21400
rect 12952 21360 12958 21372
rect 14366 21360 14372 21412
rect 14424 21400 14430 21412
rect 14737 21403 14795 21409
rect 14737 21400 14749 21403
rect 14424 21372 14749 21400
rect 14424 21360 14430 21372
rect 14737 21369 14749 21372
rect 14783 21369 14795 21403
rect 15746 21400 15752 21412
rect 15707 21372 15752 21400
rect 14737 21363 14795 21369
rect 15746 21360 15752 21372
rect 15804 21360 15810 21412
rect 16316 21409 16344 21440
rect 17865 21437 17877 21471
rect 17911 21468 17923 21471
rect 20364 21468 20392 21508
rect 21085 21505 21097 21508
rect 21131 21505 21143 21539
rect 21085 21499 21143 21505
rect 21266 21496 21272 21548
rect 21324 21536 21330 21548
rect 22370 21536 22376 21548
rect 21324 21508 21417 21536
rect 22331 21508 22376 21536
rect 21324 21496 21330 21508
rect 22370 21496 22376 21508
rect 22428 21496 22434 21548
rect 17911 21440 20392 21468
rect 17911 21437 17923 21440
rect 17865 21431 17923 21437
rect 16301 21403 16359 21409
rect 16301 21369 16313 21403
rect 16347 21369 16359 21403
rect 20364 21400 20392 21440
rect 20441 21471 20499 21477
rect 20441 21437 20453 21471
rect 20487 21468 20499 21471
rect 21177 21471 21235 21477
rect 21177 21468 21189 21471
rect 20487 21440 21189 21468
rect 20487 21437 20499 21440
rect 20441 21431 20499 21437
rect 21177 21437 21189 21440
rect 21223 21437 21235 21471
rect 21177 21431 21235 21437
rect 22005 21403 22063 21409
rect 22005 21400 22017 21403
rect 20364 21372 22017 21400
rect 16301 21363 16359 21369
rect 22005 21369 22017 21372
rect 22051 21369 22063 21403
rect 22005 21363 22063 21369
rect 12989 21335 13047 21341
rect 12989 21332 13001 21335
rect 11848 21304 13001 21332
rect 11848 21292 11854 21304
rect 12989 21301 13001 21304
rect 13035 21332 13047 21335
rect 14642 21332 14648 21344
rect 13035 21304 14648 21332
rect 13035 21301 13047 21304
rect 12989 21295 13047 21301
rect 14642 21292 14648 21304
rect 14700 21292 14706 21344
rect 16117 21335 16175 21341
rect 16117 21301 16129 21335
rect 16163 21332 16175 21335
rect 16482 21332 16488 21344
rect 16163 21304 16488 21332
rect 16163 21301 16175 21304
rect 16117 21295 16175 21301
rect 16482 21292 16488 21304
rect 16540 21292 16546 21344
rect 1104 21242 23828 21264
rect 1104 21190 3790 21242
rect 3842 21190 3854 21242
rect 3906 21190 3918 21242
rect 3970 21190 3982 21242
rect 4034 21190 4046 21242
rect 4098 21190 9471 21242
rect 9523 21190 9535 21242
rect 9587 21190 9599 21242
rect 9651 21190 9663 21242
rect 9715 21190 9727 21242
rect 9779 21190 15152 21242
rect 15204 21190 15216 21242
rect 15268 21190 15280 21242
rect 15332 21190 15344 21242
rect 15396 21190 15408 21242
rect 15460 21190 20833 21242
rect 20885 21190 20897 21242
rect 20949 21190 20961 21242
rect 21013 21190 21025 21242
rect 21077 21190 21089 21242
rect 21141 21190 23828 21242
rect 1104 21168 23828 21190
rect 9398 21088 9404 21140
rect 9456 21128 9462 21140
rect 11330 21128 11336 21140
rect 9456 21100 11336 21128
rect 9456 21088 9462 21100
rect 11330 21088 11336 21100
rect 11388 21088 11394 21140
rect 11701 21131 11759 21137
rect 11701 21097 11713 21131
rect 11747 21128 11759 21131
rect 14277 21131 14335 21137
rect 14277 21128 14289 21131
rect 11747 21100 14289 21128
rect 11747 21097 11759 21100
rect 11701 21091 11759 21097
rect 14277 21097 14289 21100
rect 14323 21097 14335 21131
rect 16482 21128 16488 21140
rect 14277 21091 14335 21097
rect 14384 21100 16488 21128
rect 12253 21063 12311 21069
rect 12253 21060 12265 21063
rect 10152 21032 12265 21060
rect 5350 20992 5356 21004
rect 5311 20964 5356 20992
rect 5350 20952 5356 20964
rect 5408 20992 5414 21004
rect 5813 20995 5871 21001
rect 5813 20992 5825 20995
rect 5408 20964 5825 20992
rect 5408 20952 5414 20964
rect 5813 20961 5825 20964
rect 5859 20961 5871 20995
rect 9122 20992 9128 21004
rect 9083 20964 9128 20992
rect 5813 20955 5871 20961
rect 9122 20952 9128 20964
rect 9180 20952 9186 21004
rect 2038 20924 2044 20936
rect 1999 20896 2044 20924
rect 2038 20884 2044 20896
rect 2096 20884 2102 20936
rect 6080 20927 6138 20933
rect 6080 20893 6092 20927
rect 6126 20924 6138 20927
rect 10152 20924 10180 21032
rect 12253 21029 12265 21032
rect 12299 21029 12311 21063
rect 13446 21060 13452 21072
rect 13407 21032 13452 21060
rect 12253 21023 12311 21029
rect 13446 21020 13452 21032
rect 13504 21020 13510 21072
rect 13630 21020 13636 21072
rect 13688 21060 13694 21072
rect 14384 21060 14412 21100
rect 16482 21088 16488 21100
rect 16540 21088 16546 21140
rect 21266 21128 21272 21140
rect 21227 21100 21272 21128
rect 21266 21088 21272 21100
rect 21324 21088 21330 21140
rect 13688 21032 14412 21060
rect 13688 21020 13694 21032
rect 14458 21020 14464 21072
rect 14516 21020 14522 21072
rect 14550 21020 14556 21072
rect 14608 21060 14614 21072
rect 15562 21060 15568 21072
rect 14608 21032 14653 21060
rect 14752 21032 15568 21060
rect 14608 21020 14614 21032
rect 11333 20995 11391 21001
rect 11333 20961 11345 20995
rect 11379 20992 11391 20995
rect 14476 20992 14504 21020
rect 14752 21001 14780 21032
rect 15562 21020 15568 21032
rect 15620 21020 15626 21072
rect 16206 21060 16212 21072
rect 16167 21032 16212 21060
rect 16206 21020 16212 21032
rect 16264 21020 16270 21072
rect 14644 20995 14702 21001
rect 14644 20992 14656 20995
rect 11379 20964 12848 20992
rect 14476 20964 14656 20992
rect 11379 20961 11391 20964
rect 11333 20955 11391 20961
rect 6126 20896 10180 20924
rect 11517 20927 11575 20933
rect 6126 20893 6138 20896
rect 6080 20887 6138 20893
rect 11517 20893 11529 20927
rect 11563 20893 11575 20927
rect 11790 20924 11796 20936
rect 11751 20896 11796 20924
rect 11517 20887 11575 20893
rect 1670 20816 1676 20868
rect 1728 20856 1734 20868
rect 2286 20859 2344 20865
rect 2286 20856 2298 20859
rect 1728 20828 2298 20856
rect 1728 20816 1734 20828
rect 2286 20825 2298 20828
rect 2332 20825 2344 20859
rect 2286 20819 2344 20825
rect 4706 20816 4712 20868
rect 4764 20856 4770 20868
rect 9398 20865 9404 20868
rect 5086 20859 5144 20865
rect 5086 20856 5098 20859
rect 4764 20828 5098 20856
rect 4764 20816 4770 20828
rect 5086 20825 5098 20828
rect 5132 20825 5144 20859
rect 9392 20856 9404 20865
rect 9359 20828 9404 20856
rect 5086 20819 5144 20825
rect 9392 20819 9404 20828
rect 9398 20816 9404 20819
rect 9456 20816 9462 20868
rect 11238 20856 11244 20868
rect 9968 20828 11244 20856
rect 3142 20748 3148 20800
rect 3200 20788 3206 20800
rect 3421 20791 3479 20797
rect 3421 20788 3433 20791
rect 3200 20760 3433 20788
rect 3200 20748 3206 20760
rect 3421 20757 3433 20760
rect 3467 20757 3479 20791
rect 3421 20751 3479 20757
rect 3510 20748 3516 20800
rect 3568 20788 3574 20800
rect 3973 20791 4031 20797
rect 3973 20788 3985 20791
rect 3568 20760 3985 20788
rect 3568 20748 3574 20760
rect 3973 20757 3985 20760
rect 4019 20757 4031 20791
rect 3973 20751 4031 20757
rect 7193 20791 7251 20797
rect 7193 20757 7205 20791
rect 7239 20788 7251 20791
rect 9968 20788 9996 20828
rect 11238 20816 11244 20828
rect 11296 20816 11302 20868
rect 11330 20816 11336 20868
rect 11388 20856 11394 20868
rect 11532 20856 11560 20887
rect 11790 20884 11796 20896
rect 11848 20884 11854 20936
rect 12437 20927 12495 20933
rect 12437 20893 12449 20927
rect 12483 20924 12495 20927
rect 12710 20924 12716 20936
rect 12483 20896 12716 20924
rect 12483 20893 12495 20896
rect 12437 20887 12495 20893
rect 12710 20884 12716 20896
rect 12768 20884 12774 20936
rect 12820 20933 12848 20964
rect 14644 20961 14656 20964
rect 14690 20961 14702 20995
rect 14644 20955 14702 20961
rect 14737 20995 14795 21001
rect 14737 20961 14749 20995
rect 14783 20961 14795 20995
rect 22094 20992 22100 21004
rect 14737 20955 14795 20961
rect 14844 20964 15424 20992
rect 12805 20927 12863 20933
rect 12805 20893 12817 20927
rect 12851 20893 12863 20927
rect 12805 20887 12863 20893
rect 13725 20927 13783 20933
rect 13725 20893 13737 20927
rect 13771 20924 13783 20927
rect 14274 20924 14280 20936
rect 13771 20896 14280 20924
rect 13771 20893 13783 20896
rect 13725 20887 13783 20893
rect 14274 20884 14280 20896
rect 14332 20884 14338 20936
rect 14461 20927 14519 20933
rect 14461 20893 14473 20927
rect 14507 20924 14519 20927
rect 14844 20924 14872 20964
rect 15396 20933 15424 20964
rect 16408 20964 22100 20992
rect 14507 20896 14872 20924
rect 15381 20927 15439 20933
rect 14507 20893 14519 20896
rect 14461 20887 14519 20893
rect 14921 20893 14979 20899
rect 11388 20828 11560 20856
rect 12529 20859 12587 20865
rect 11388 20816 11394 20828
rect 12529 20825 12541 20859
rect 12575 20825 12587 20859
rect 12529 20819 12587 20825
rect 12621 20859 12679 20865
rect 12621 20825 12633 20859
rect 12667 20856 12679 20859
rect 13354 20856 13360 20868
rect 12667 20828 13360 20856
rect 12667 20825 12679 20828
rect 12621 20819 12679 20825
rect 7239 20760 9996 20788
rect 7239 20757 7251 20760
rect 7193 20751 7251 20757
rect 10042 20748 10048 20800
rect 10100 20788 10106 20800
rect 10505 20791 10563 20797
rect 10505 20788 10517 20791
rect 10100 20760 10517 20788
rect 10100 20748 10106 20760
rect 10505 20757 10517 20760
rect 10551 20757 10563 20791
rect 12544 20788 12572 20819
rect 13354 20816 13360 20828
rect 13412 20816 13418 20868
rect 13449 20859 13507 20865
rect 13449 20825 13461 20859
rect 13495 20856 13507 20859
rect 14826 20856 14832 20868
rect 13495 20828 14832 20856
rect 13495 20825 13507 20828
rect 13449 20819 13507 20825
rect 14826 20816 14832 20828
rect 14884 20816 14890 20868
rect 14921 20859 14933 20893
rect 14967 20890 14979 20893
rect 15381 20893 15393 20927
rect 15427 20924 15439 20927
rect 15470 20924 15476 20936
rect 15427 20896 15476 20924
rect 15427 20893 15439 20896
rect 14967 20862 15056 20890
rect 15381 20887 15439 20893
rect 15470 20884 15476 20896
rect 15528 20884 15534 20936
rect 15565 20927 15623 20933
rect 15565 20893 15577 20927
rect 15611 20924 15623 20927
rect 15654 20924 15660 20936
rect 15611 20896 15660 20924
rect 15611 20893 15623 20896
rect 15565 20887 15623 20893
rect 15654 20884 15660 20896
rect 15712 20924 15718 20936
rect 16114 20924 16120 20936
rect 15712 20896 16120 20924
rect 15712 20884 15718 20896
rect 16114 20884 16120 20896
rect 16172 20884 16178 20936
rect 16408 20933 16436 20964
rect 22094 20952 22100 20964
rect 22152 20952 22158 21004
rect 16393 20927 16451 20933
rect 16393 20893 16405 20927
rect 16439 20893 16451 20927
rect 16666 20924 16672 20936
rect 16627 20896 16672 20924
rect 16393 20887 16451 20893
rect 16666 20884 16672 20896
rect 16724 20884 16730 20936
rect 16942 20924 16948 20936
rect 16903 20896 16948 20924
rect 16942 20884 16948 20896
rect 17000 20884 17006 20936
rect 17589 20927 17647 20933
rect 17589 20893 17601 20927
rect 17635 20924 17647 20927
rect 18322 20924 18328 20936
rect 17635 20896 18328 20924
rect 17635 20893 17647 20896
rect 17589 20887 17647 20893
rect 18322 20884 18328 20896
rect 18380 20884 18386 20936
rect 21174 20924 21180 20936
rect 21135 20896 21180 20924
rect 21174 20884 21180 20896
rect 21232 20884 21238 20936
rect 21361 20927 21419 20933
rect 21361 20893 21373 20927
rect 21407 20924 21419 20927
rect 22370 20924 22376 20936
rect 21407 20896 22376 20924
rect 21407 20893 21419 20896
rect 21361 20887 21419 20893
rect 22370 20884 22376 20896
rect 22428 20884 22434 20936
rect 14967 20859 14979 20862
rect 14921 20853 14979 20859
rect 15028 20856 15056 20862
rect 15286 20856 15292 20868
rect 15028 20828 15292 20856
rect 15286 20816 15292 20828
rect 15344 20816 15350 20868
rect 12710 20788 12716 20800
rect 12544 20760 12716 20788
rect 10505 20751 10563 20757
rect 12710 20748 12716 20760
rect 12768 20748 12774 20800
rect 13262 20748 13268 20800
rect 13320 20788 13326 20800
rect 13633 20791 13691 20797
rect 13633 20788 13645 20791
rect 13320 20760 13645 20788
rect 13320 20748 13326 20760
rect 13633 20757 13645 20760
rect 13679 20757 13691 20791
rect 15378 20788 15384 20800
rect 15339 20760 15384 20788
rect 13633 20751 13691 20757
rect 15378 20748 15384 20760
rect 15436 20748 15442 20800
rect 15470 20748 15476 20800
rect 15528 20788 15534 20800
rect 15654 20788 15660 20800
rect 15528 20760 15660 20788
rect 15528 20748 15534 20760
rect 15654 20748 15660 20760
rect 15712 20748 15718 20800
rect 1104 20698 23987 20720
rect 1104 20646 6630 20698
rect 6682 20646 6694 20698
rect 6746 20646 6758 20698
rect 6810 20646 6822 20698
rect 6874 20646 6886 20698
rect 6938 20646 12311 20698
rect 12363 20646 12375 20698
rect 12427 20646 12439 20698
rect 12491 20646 12503 20698
rect 12555 20646 12567 20698
rect 12619 20646 17992 20698
rect 18044 20646 18056 20698
rect 18108 20646 18120 20698
rect 18172 20646 18184 20698
rect 18236 20646 18248 20698
rect 18300 20646 23673 20698
rect 23725 20646 23737 20698
rect 23789 20646 23801 20698
rect 23853 20646 23865 20698
rect 23917 20646 23929 20698
rect 23981 20646 23987 20698
rect 1104 20624 23987 20646
rect 10321 20587 10379 20593
rect 10321 20553 10333 20587
rect 10367 20584 10379 20587
rect 11054 20584 11060 20596
rect 10367 20556 11060 20584
rect 10367 20553 10379 20556
rect 10321 20547 10379 20553
rect 11054 20544 11060 20556
rect 11112 20544 11118 20596
rect 12253 20587 12311 20593
rect 12253 20553 12265 20587
rect 12299 20584 12311 20587
rect 14829 20587 14887 20593
rect 12299 20556 12434 20584
rect 12299 20553 12311 20556
rect 12253 20547 12311 20553
rect 4338 20448 4344 20460
rect 4299 20420 4344 20448
rect 4338 20408 4344 20420
rect 4396 20408 4402 20460
rect 8941 20451 8999 20457
rect 8941 20417 8953 20451
rect 8987 20448 8999 20451
rect 9030 20448 9036 20460
rect 8987 20420 9036 20448
rect 8987 20417 8999 20420
rect 8941 20411 8999 20417
rect 9030 20408 9036 20420
rect 9088 20408 9094 20460
rect 9208 20451 9266 20457
rect 9208 20417 9220 20451
rect 9254 20448 9266 20451
rect 12066 20448 12072 20460
rect 9254 20420 12072 20448
rect 9254 20417 9266 20420
rect 9208 20411 9266 20417
rect 12066 20408 12072 20420
rect 12124 20408 12130 20460
rect 12158 20408 12164 20460
rect 12216 20448 12222 20460
rect 12406 20448 12434 20556
rect 14829 20553 14841 20587
rect 14875 20584 14887 20587
rect 14918 20584 14924 20596
rect 14875 20556 14924 20584
rect 14875 20553 14887 20556
rect 14829 20547 14887 20553
rect 14918 20544 14924 20556
rect 14976 20544 14982 20596
rect 15657 20587 15715 20593
rect 15657 20553 15669 20587
rect 15703 20584 15715 20587
rect 15746 20584 15752 20596
rect 15703 20556 15752 20584
rect 15703 20553 15715 20556
rect 15657 20547 15715 20553
rect 15746 20544 15752 20556
rect 15804 20544 15810 20596
rect 17310 20584 17316 20596
rect 16132 20556 17316 20584
rect 13630 20516 13636 20528
rect 13188 20488 13636 20516
rect 13188 20460 13216 20488
rect 13630 20476 13636 20488
rect 13688 20476 13694 20528
rect 15378 20516 15384 20528
rect 13924 20488 15384 20516
rect 12710 20448 12716 20460
rect 12216 20420 12261 20448
rect 12406 20420 12716 20448
rect 12216 20408 12222 20420
rect 12710 20408 12716 20420
rect 12768 20448 12774 20460
rect 13170 20448 13176 20460
rect 12768 20420 13176 20448
rect 12768 20408 12774 20420
rect 13170 20408 13176 20420
rect 13228 20408 13234 20460
rect 13538 20448 13544 20460
rect 13499 20420 13544 20448
rect 13538 20408 13544 20420
rect 13596 20408 13602 20460
rect 13924 20457 13952 20488
rect 15378 20476 15384 20488
rect 15436 20476 15442 20528
rect 13909 20451 13967 20457
rect 13909 20417 13921 20451
rect 13955 20417 13967 20451
rect 13909 20411 13967 20417
rect 14185 20451 14243 20457
rect 14185 20417 14197 20451
rect 14231 20448 14243 20451
rect 14734 20448 14740 20460
rect 14231 20420 14740 20448
rect 14231 20417 14243 20420
rect 14185 20411 14243 20417
rect 14734 20408 14740 20420
rect 14792 20408 14798 20460
rect 14918 20408 14924 20460
rect 14976 20448 14982 20460
rect 15013 20451 15071 20457
rect 15013 20448 15025 20451
rect 14976 20420 15025 20448
rect 14976 20408 14982 20420
rect 15013 20417 15025 20420
rect 15059 20417 15071 20451
rect 15013 20411 15071 20417
rect 15197 20451 15255 20457
rect 15197 20417 15209 20451
rect 15243 20448 15255 20451
rect 15562 20448 15568 20460
rect 15243 20420 15568 20448
rect 15243 20417 15255 20420
rect 15197 20411 15255 20417
rect 15562 20408 15568 20420
rect 15620 20408 15626 20460
rect 15746 20408 15752 20460
rect 15804 20448 15810 20460
rect 15841 20451 15899 20457
rect 15841 20448 15853 20451
rect 15804 20420 15853 20448
rect 15804 20408 15810 20420
rect 15841 20417 15853 20420
rect 15887 20417 15899 20451
rect 15841 20411 15899 20417
rect 15930 20408 15936 20460
rect 15988 20448 15994 20460
rect 16132 20457 16160 20556
rect 17310 20544 17316 20556
rect 17368 20584 17374 20596
rect 17368 20556 17448 20584
rect 17368 20544 17374 20556
rect 16025 20451 16083 20457
rect 16025 20448 16037 20451
rect 15988 20420 16037 20448
rect 15988 20408 15994 20420
rect 16025 20417 16037 20420
rect 16071 20417 16083 20451
rect 16025 20411 16083 20417
rect 16117 20451 16175 20457
rect 16117 20417 16129 20451
rect 16163 20417 16175 20451
rect 16117 20411 16175 20417
rect 16298 20408 16304 20460
rect 16356 20448 16362 20460
rect 16942 20448 16948 20460
rect 16356 20420 16948 20448
rect 16356 20408 16362 20420
rect 16942 20408 16948 20420
rect 17000 20408 17006 20460
rect 17420 20457 17448 20556
rect 17862 20544 17868 20596
rect 17920 20584 17926 20596
rect 18417 20587 18475 20593
rect 18417 20584 18429 20587
rect 17920 20556 18429 20584
rect 17920 20544 17926 20556
rect 18417 20553 18429 20556
rect 18463 20553 18475 20587
rect 19426 20584 19432 20596
rect 18417 20547 18475 20553
rect 18708 20556 19432 20584
rect 17267 20451 17325 20457
rect 17267 20448 17279 20451
rect 17144 20420 17279 20448
rect 2038 20340 2044 20392
rect 2096 20380 2102 20392
rect 2593 20383 2651 20389
rect 2593 20380 2605 20383
rect 2096 20352 2605 20380
rect 2096 20340 2102 20352
rect 2593 20349 2605 20352
rect 2639 20349 2651 20383
rect 2593 20343 2651 20349
rect 14826 20340 14832 20392
rect 14884 20380 14890 20392
rect 17037 20383 17095 20389
rect 17037 20380 17049 20383
rect 14884 20352 17049 20380
rect 14884 20340 14890 20352
rect 17037 20349 17049 20352
rect 17083 20349 17095 20383
rect 17037 20343 17095 20349
rect 13541 20315 13599 20321
rect 13541 20281 13553 20315
rect 13587 20312 13599 20315
rect 13630 20312 13636 20324
rect 13587 20284 13636 20312
rect 13587 20281 13599 20284
rect 13541 20275 13599 20281
rect 13630 20272 13636 20284
rect 13688 20272 13694 20324
rect 15470 20272 15476 20324
rect 15528 20312 15534 20324
rect 15933 20315 15991 20321
rect 15933 20312 15945 20315
rect 15528 20284 15945 20312
rect 15528 20272 15534 20284
rect 15933 20281 15945 20284
rect 15979 20312 15991 20315
rect 17144 20312 17172 20420
rect 17267 20417 17279 20420
rect 17313 20417 17325 20451
rect 17267 20411 17325 20417
rect 17405 20451 17463 20457
rect 17405 20417 17417 20451
rect 17451 20417 17463 20451
rect 17405 20411 17463 20417
rect 17497 20451 17555 20457
rect 17497 20417 17509 20451
rect 17543 20417 17555 20451
rect 17678 20448 17684 20460
rect 17639 20420 17684 20448
rect 17497 20411 17555 20417
rect 17512 20380 17540 20411
rect 17678 20408 17684 20420
rect 17736 20408 17742 20460
rect 18598 20448 18604 20460
rect 18559 20420 18604 20448
rect 18598 20408 18604 20420
rect 18656 20408 18662 20460
rect 18708 20457 18736 20556
rect 19426 20544 19432 20556
rect 19484 20544 19490 20596
rect 22094 20544 22100 20596
rect 22152 20584 22158 20596
rect 22152 20556 22197 20584
rect 22152 20544 22158 20556
rect 19521 20519 19579 20525
rect 19521 20516 19533 20519
rect 18892 20488 19533 20516
rect 18892 20457 18920 20488
rect 19521 20485 19533 20488
rect 19567 20485 19579 20519
rect 19521 20479 19579 20485
rect 18693 20451 18751 20457
rect 18693 20417 18705 20451
rect 18739 20417 18751 20451
rect 18693 20411 18751 20417
rect 18877 20451 18935 20457
rect 18877 20417 18889 20451
rect 18923 20417 18935 20451
rect 18877 20411 18935 20417
rect 18966 20408 18972 20460
rect 19024 20448 19030 20460
rect 19426 20448 19432 20460
rect 19024 20420 19069 20448
rect 19387 20420 19432 20448
rect 19024 20408 19030 20420
rect 19426 20408 19432 20420
rect 19484 20408 19490 20460
rect 19613 20451 19671 20457
rect 19613 20417 19625 20451
rect 19659 20448 19671 20451
rect 20162 20448 20168 20460
rect 19659 20420 20168 20448
rect 19659 20417 19671 20420
rect 19613 20411 19671 20417
rect 20162 20408 20168 20420
rect 20220 20408 20226 20460
rect 22005 20451 22063 20457
rect 22005 20417 22017 20451
rect 22051 20417 22063 20451
rect 22186 20448 22192 20460
rect 22147 20420 22192 20448
rect 22005 20411 22063 20417
rect 20070 20380 20076 20392
rect 17512 20352 20076 20380
rect 20070 20340 20076 20352
rect 20128 20340 20134 20392
rect 15979 20284 17172 20312
rect 15979 20281 15991 20284
rect 15933 20275 15991 20281
rect 17678 20272 17684 20324
rect 17736 20312 17742 20324
rect 19334 20312 19340 20324
rect 17736 20284 19340 20312
rect 17736 20272 17742 20284
rect 19334 20272 19340 20284
rect 19392 20312 19398 20324
rect 22020 20312 22048 20411
rect 22186 20408 22192 20420
rect 22244 20408 22250 20460
rect 19392 20284 22048 20312
rect 19392 20272 19398 20284
rect 11149 20247 11207 20253
rect 11149 20213 11161 20247
rect 11195 20244 11207 20247
rect 11330 20244 11336 20256
rect 11195 20216 11336 20244
rect 11195 20213 11207 20216
rect 11149 20207 11207 20213
rect 11330 20204 11336 20216
rect 11388 20204 11394 20256
rect 14642 20204 14648 20256
rect 14700 20244 14706 20256
rect 15197 20247 15255 20253
rect 15197 20244 15209 20247
rect 14700 20216 15209 20244
rect 14700 20204 14706 20216
rect 15197 20213 15209 20216
rect 15243 20244 15255 20247
rect 16298 20244 16304 20256
rect 15243 20216 16304 20244
rect 15243 20213 15255 20216
rect 15197 20207 15255 20213
rect 16298 20204 16304 20216
rect 16356 20204 16362 20256
rect 1104 20154 23828 20176
rect 1104 20102 3790 20154
rect 3842 20102 3854 20154
rect 3906 20102 3918 20154
rect 3970 20102 3982 20154
rect 4034 20102 4046 20154
rect 4098 20102 9471 20154
rect 9523 20102 9535 20154
rect 9587 20102 9599 20154
rect 9651 20102 9663 20154
rect 9715 20102 9727 20154
rect 9779 20102 15152 20154
rect 15204 20102 15216 20154
rect 15268 20102 15280 20154
rect 15332 20102 15344 20154
rect 15396 20102 15408 20154
rect 15460 20102 20833 20154
rect 20885 20102 20897 20154
rect 20949 20102 20961 20154
rect 21013 20102 21025 20154
rect 21077 20102 21089 20154
rect 21141 20102 23828 20154
rect 1104 20080 23828 20102
rect 12066 20000 12072 20052
rect 12124 20040 12130 20052
rect 12161 20043 12219 20049
rect 12161 20040 12173 20043
rect 12124 20012 12173 20040
rect 12124 20000 12130 20012
rect 12161 20009 12173 20012
rect 12207 20009 12219 20043
rect 12161 20003 12219 20009
rect 14737 20043 14795 20049
rect 14737 20009 14749 20043
rect 14783 20040 14795 20043
rect 15010 20040 15016 20052
rect 14783 20012 15016 20040
rect 14783 20009 14795 20012
rect 14737 20003 14795 20009
rect 15010 20000 15016 20012
rect 15068 20000 15074 20052
rect 18233 20043 18291 20049
rect 18233 20040 18245 20043
rect 16316 20012 18245 20040
rect 16316 19984 16344 20012
rect 18233 20009 18245 20012
rect 18279 20040 18291 20043
rect 18966 20040 18972 20052
rect 18279 20012 18972 20040
rect 18279 20009 18291 20012
rect 18233 20003 18291 20009
rect 18966 20000 18972 20012
rect 19024 20000 19030 20052
rect 13262 19972 13268 19984
rect 10980 19944 13268 19972
rect 2038 19904 2044 19916
rect 1999 19876 2044 19904
rect 2038 19864 2044 19876
rect 2096 19864 2102 19916
rect 6641 19907 6699 19913
rect 6641 19873 6653 19907
rect 6687 19904 6699 19907
rect 9122 19904 9128 19916
rect 6687 19876 9128 19904
rect 6687 19873 6699 19876
rect 6641 19867 6699 19873
rect 9122 19864 9128 19876
rect 9180 19864 9186 19916
rect 10980 19845 11008 19944
rect 13262 19932 13268 19944
rect 13320 19932 13326 19984
rect 15286 19932 15292 19984
rect 15344 19972 15350 19984
rect 15933 19975 15991 19981
rect 15933 19972 15945 19975
rect 15344 19944 15945 19972
rect 15344 19932 15350 19944
rect 15933 19941 15945 19944
rect 15979 19972 15991 19975
rect 16298 19972 16304 19984
rect 15979 19944 16304 19972
rect 15979 19941 15991 19944
rect 15933 19935 15991 19941
rect 16298 19932 16304 19944
rect 16356 19932 16362 19984
rect 16482 19972 16488 19984
rect 16443 19944 16488 19972
rect 16482 19932 16488 19944
rect 16540 19932 16546 19984
rect 16758 19932 16764 19984
rect 16816 19972 16822 19984
rect 16816 19944 20576 19972
rect 16816 19932 16822 19944
rect 12158 19904 12164 19916
rect 11624 19876 12164 19904
rect 9392 19839 9450 19845
rect 9392 19805 9404 19839
rect 9438 19836 9450 19839
rect 10965 19839 11023 19845
rect 10965 19836 10977 19839
rect 9438 19808 10977 19836
rect 9438 19805 9450 19808
rect 9392 19799 9450 19805
rect 10965 19805 10977 19808
rect 11011 19805 11023 19839
rect 10965 19799 11023 19805
rect 1578 19728 1584 19780
rect 1636 19768 1642 19780
rect 2286 19771 2344 19777
rect 2286 19768 2298 19771
rect 1636 19740 2298 19768
rect 1636 19728 1642 19740
rect 2286 19737 2298 19740
rect 2332 19737 2344 19771
rect 2286 19731 2344 19737
rect 5718 19728 5724 19780
rect 5776 19768 5782 19780
rect 6374 19771 6432 19777
rect 6374 19768 6386 19771
rect 5776 19740 6386 19768
rect 5776 19728 5782 19740
rect 6374 19737 6386 19740
rect 6420 19737 6432 19771
rect 6374 19731 6432 19737
rect 3421 19703 3479 19709
rect 3421 19669 3433 19703
rect 3467 19700 3479 19703
rect 3602 19700 3608 19712
rect 3467 19672 3608 19700
rect 3467 19669 3479 19672
rect 3421 19663 3479 19669
rect 3602 19660 3608 19672
rect 3660 19660 3666 19712
rect 4430 19660 4436 19712
rect 4488 19700 4494 19712
rect 5261 19703 5319 19709
rect 5261 19700 5273 19703
rect 4488 19672 5273 19700
rect 4488 19660 4494 19672
rect 5261 19669 5273 19672
rect 5307 19669 5319 19703
rect 5261 19663 5319 19669
rect 10505 19703 10563 19709
rect 10505 19669 10517 19703
rect 10551 19700 10563 19703
rect 10778 19700 10784 19712
rect 10551 19672 10784 19700
rect 10551 19669 10563 19672
rect 10505 19663 10563 19669
rect 10778 19660 10784 19672
rect 10836 19660 10842 19712
rect 11330 19660 11336 19712
rect 11388 19700 11394 19712
rect 11624 19709 11652 19876
rect 12158 19864 12164 19876
rect 12216 19904 12222 19916
rect 12805 19907 12863 19913
rect 12805 19904 12817 19907
rect 12216 19876 12817 19904
rect 12216 19864 12222 19876
rect 12805 19873 12817 19876
rect 12851 19904 12863 19907
rect 12894 19904 12900 19916
rect 12851 19876 12900 19904
rect 12851 19873 12863 19876
rect 12805 19867 12863 19873
rect 12894 19864 12900 19876
rect 12952 19864 12958 19916
rect 15010 19864 15016 19916
rect 15068 19904 15074 19916
rect 15378 19904 15384 19916
rect 15068 19876 15384 19904
rect 15068 19864 15074 19876
rect 15378 19864 15384 19876
rect 15436 19864 15442 19916
rect 16669 19907 16727 19913
rect 16669 19873 16681 19907
rect 16715 19904 16727 19907
rect 17678 19904 17684 19916
rect 16715 19876 17684 19904
rect 16715 19873 16727 19876
rect 16669 19867 16727 19873
rect 17678 19864 17684 19876
rect 17736 19864 17742 19916
rect 19426 19864 19432 19916
rect 19484 19904 19490 19916
rect 20257 19907 20315 19913
rect 20257 19904 20269 19907
rect 19484 19876 20269 19904
rect 19484 19864 19490 19876
rect 20257 19873 20269 19876
rect 20303 19904 20315 19907
rect 20438 19904 20444 19916
rect 20303 19876 20444 19904
rect 20303 19873 20315 19876
rect 20257 19867 20315 19873
rect 20438 19864 20444 19876
rect 20496 19864 20502 19916
rect 12621 19839 12679 19845
rect 12621 19805 12633 19839
rect 12667 19836 12679 19839
rect 13446 19836 13452 19848
rect 12667 19808 13452 19836
rect 12667 19805 12679 19808
rect 12621 19799 12679 19805
rect 13446 19796 13452 19808
rect 13504 19796 13510 19848
rect 14642 19836 14648 19848
rect 14603 19808 14648 19836
rect 14642 19796 14648 19808
rect 14700 19796 14706 19848
rect 14829 19839 14887 19845
rect 14829 19805 14841 19839
rect 14875 19836 14887 19839
rect 16022 19836 16028 19848
rect 14875 19808 16028 19836
rect 14875 19805 14887 19808
rect 14829 19799 14887 19805
rect 16022 19796 16028 19808
rect 16080 19796 16086 19848
rect 16390 19836 16396 19848
rect 16351 19808 16396 19836
rect 16390 19796 16396 19808
rect 16448 19796 16454 19848
rect 17034 19796 17040 19848
rect 17092 19836 17098 19848
rect 17405 19839 17463 19845
rect 17405 19836 17417 19839
rect 17092 19808 17417 19836
rect 17092 19796 17098 19808
rect 17405 19805 17417 19808
rect 17451 19805 17463 19839
rect 17405 19799 17463 19805
rect 17589 19839 17647 19845
rect 17589 19805 17601 19839
rect 17635 19836 17647 19839
rect 18690 19836 18696 19848
rect 17635 19808 18696 19836
rect 17635 19805 17647 19808
rect 17589 19799 17647 19805
rect 18690 19796 18696 19808
rect 18748 19796 18754 19848
rect 20548 19845 20576 19944
rect 20533 19839 20591 19845
rect 20533 19805 20545 19839
rect 20579 19836 20591 19839
rect 20990 19836 20996 19848
rect 20579 19808 20996 19836
rect 20579 19805 20591 19808
rect 20533 19799 20591 19805
rect 20990 19796 20996 19808
rect 21048 19796 21054 19848
rect 13078 19728 13084 19780
rect 13136 19768 13142 19780
rect 16669 19771 16727 19777
rect 16669 19768 16681 19771
rect 13136 19740 16681 19768
rect 13136 19728 13142 19740
rect 16669 19737 16681 19740
rect 16715 19737 16727 19771
rect 16669 19731 16727 19737
rect 16850 19728 16856 19780
rect 16908 19768 16914 19780
rect 16908 19740 19380 19768
rect 16908 19728 16914 19740
rect 11609 19703 11667 19709
rect 11609 19700 11621 19703
rect 11388 19672 11621 19700
rect 11388 19660 11394 19672
rect 11609 19669 11621 19672
rect 11655 19669 11667 19703
rect 11609 19663 11667 19669
rect 12529 19703 12587 19709
rect 12529 19669 12541 19703
rect 12575 19700 12587 19703
rect 14918 19700 14924 19712
rect 12575 19672 14924 19700
rect 12575 19669 12587 19672
rect 12529 19663 12587 19669
rect 14918 19660 14924 19672
rect 14976 19660 14982 19712
rect 15930 19660 15936 19712
rect 15988 19700 15994 19712
rect 17221 19703 17279 19709
rect 17221 19700 17233 19703
rect 15988 19672 17233 19700
rect 15988 19660 15994 19672
rect 17221 19669 17233 19672
rect 17267 19700 17279 19703
rect 17862 19700 17868 19712
rect 17267 19672 17868 19700
rect 17267 19669 17279 19672
rect 17221 19663 17279 19669
rect 17862 19660 17868 19672
rect 17920 19660 17926 19712
rect 19352 19700 19380 19740
rect 19886 19700 19892 19712
rect 19352 19672 19892 19700
rect 19886 19660 19892 19672
rect 19944 19660 19950 19712
rect 1104 19610 23987 19632
rect 1104 19558 6630 19610
rect 6682 19558 6694 19610
rect 6746 19558 6758 19610
rect 6810 19558 6822 19610
rect 6874 19558 6886 19610
rect 6938 19558 12311 19610
rect 12363 19558 12375 19610
rect 12427 19558 12439 19610
rect 12491 19558 12503 19610
rect 12555 19558 12567 19610
rect 12619 19558 17992 19610
rect 18044 19558 18056 19610
rect 18108 19558 18120 19610
rect 18172 19558 18184 19610
rect 18236 19558 18248 19610
rect 18300 19558 23673 19610
rect 23725 19558 23737 19610
rect 23789 19558 23801 19610
rect 23853 19558 23865 19610
rect 23917 19558 23929 19610
rect 23981 19558 23987 19610
rect 1104 19536 23987 19558
rect 4249 19499 4307 19505
rect 4249 19465 4261 19499
rect 4295 19496 4307 19499
rect 5166 19496 5172 19508
rect 4295 19468 5172 19496
rect 4295 19465 4307 19468
rect 4249 19459 4307 19465
rect 5166 19456 5172 19468
rect 5224 19456 5230 19508
rect 5902 19456 5908 19508
rect 5960 19496 5966 19508
rect 6641 19499 6699 19505
rect 6641 19496 6653 19499
rect 5960 19468 6653 19496
rect 5960 19456 5966 19468
rect 6641 19465 6653 19468
rect 6687 19465 6699 19499
rect 6641 19459 6699 19465
rect 10321 19499 10379 19505
rect 10321 19465 10333 19499
rect 10367 19496 10379 19499
rect 11974 19496 11980 19508
rect 10367 19468 11980 19496
rect 10367 19465 10379 19468
rect 10321 19459 10379 19465
rect 11974 19456 11980 19468
rect 12032 19456 12038 19508
rect 16482 19456 16488 19508
rect 16540 19496 16546 19508
rect 17497 19499 17555 19505
rect 17497 19496 17509 19499
rect 16540 19468 17509 19496
rect 16540 19456 16546 19468
rect 17497 19465 17509 19468
rect 17543 19465 17555 19499
rect 17497 19459 17555 19465
rect 7558 19388 7564 19440
rect 7616 19428 7622 19440
rect 7754 19431 7812 19437
rect 7754 19428 7766 19431
rect 7616 19400 7766 19428
rect 7616 19388 7622 19400
rect 7754 19397 7766 19400
rect 7800 19397 7812 19431
rect 15746 19428 15752 19440
rect 7754 19391 7812 19397
rect 14660 19400 15752 19428
rect 3136 19363 3194 19369
rect 3136 19329 3148 19363
rect 3182 19360 3194 19363
rect 3418 19360 3424 19372
rect 3182 19332 3424 19360
rect 3182 19329 3194 19332
rect 3136 19323 3194 19329
rect 3418 19320 3424 19332
rect 3476 19320 3482 19372
rect 4338 19320 4344 19372
rect 4396 19360 4402 19372
rect 7466 19360 7472 19372
rect 4396 19332 7472 19360
rect 4396 19320 4402 19332
rect 7466 19320 7472 19332
rect 7524 19320 7530 19372
rect 8018 19360 8024 19372
rect 7979 19332 8024 19360
rect 8018 19320 8024 19332
rect 8076 19320 8082 19372
rect 8941 19363 8999 19369
rect 8941 19329 8953 19363
rect 8987 19360 8999 19363
rect 9030 19360 9036 19372
rect 8987 19332 9036 19360
rect 8987 19329 8999 19332
rect 8941 19323 8999 19329
rect 9030 19320 9036 19332
rect 9088 19320 9094 19372
rect 9208 19363 9266 19369
rect 9208 19329 9220 19363
rect 9254 19360 9266 19363
rect 14550 19360 14556 19372
rect 9254 19332 14556 19360
rect 9254 19329 9266 19332
rect 9208 19323 9266 19329
rect 14550 19320 14556 19332
rect 14608 19320 14614 19372
rect 14660 19369 14688 19400
rect 15746 19388 15752 19400
rect 15804 19388 15810 19440
rect 16666 19388 16672 19440
rect 16724 19428 16730 19440
rect 17405 19431 17463 19437
rect 17405 19428 17417 19431
rect 16724 19400 17417 19428
rect 16724 19388 16730 19400
rect 17405 19397 17417 19400
rect 17451 19397 17463 19431
rect 17405 19391 17463 19397
rect 18690 19388 18696 19440
rect 18748 19428 18754 19440
rect 20441 19431 20499 19437
rect 20441 19428 20453 19431
rect 18748 19400 20453 19428
rect 18748 19388 18754 19400
rect 20441 19397 20453 19400
rect 20487 19397 20499 19431
rect 20441 19391 20499 19397
rect 14645 19363 14703 19369
rect 14645 19329 14657 19363
rect 14691 19329 14703 19363
rect 14645 19323 14703 19329
rect 14734 19320 14740 19372
rect 14792 19360 14798 19372
rect 14829 19363 14887 19369
rect 14829 19360 14841 19363
rect 14792 19332 14841 19360
rect 14792 19320 14798 19332
rect 14829 19329 14841 19332
rect 14875 19329 14887 19363
rect 14829 19323 14887 19329
rect 15194 19320 15200 19372
rect 15252 19360 15258 19372
rect 15289 19363 15347 19369
rect 15289 19360 15301 19363
rect 15252 19332 15301 19360
rect 15252 19320 15258 19332
rect 15289 19329 15301 19332
rect 15335 19329 15347 19363
rect 15930 19360 15936 19372
rect 15289 19323 15347 19329
rect 15396 19332 15936 19360
rect 2774 19252 2780 19304
rect 2832 19292 2838 19304
rect 2869 19295 2927 19301
rect 2869 19292 2881 19295
rect 2832 19264 2881 19292
rect 2832 19252 2838 19264
rect 2869 19261 2881 19264
rect 2915 19261 2927 19295
rect 2869 19255 2927 19261
rect 12986 19252 12992 19304
rect 13044 19292 13050 19304
rect 15396 19292 15424 19332
rect 15930 19320 15936 19332
rect 15988 19320 15994 19372
rect 17126 19320 17132 19372
rect 17184 19320 17190 19372
rect 17310 19360 17316 19372
rect 17271 19332 17316 19360
rect 17310 19320 17316 19332
rect 17368 19320 17374 19372
rect 17773 19363 17831 19369
rect 17773 19329 17785 19363
rect 17819 19360 17831 19363
rect 18506 19360 18512 19372
rect 17819 19332 18512 19360
rect 17819 19329 17831 19332
rect 17773 19323 17831 19329
rect 18506 19320 18512 19332
rect 18564 19320 18570 19372
rect 19334 19360 19340 19372
rect 19295 19332 19340 19360
rect 19334 19320 19340 19332
rect 19392 19320 19398 19372
rect 19518 19360 19524 19372
rect 19479 19332 19524 19360
rect 19518 19320 19524 19332
rect 19576 19320 19582 19372
rect 19610 19320 19616 19372
rect 19668 19360 19674 19372
rect 20254 19360 20260 19372
rect 19668 19332 19713 19360
rect 20215 19332 20260 19360
rect 19668 19320 19674 19332
rect 20254 19320 20260 19332
rect 20312 19320 20318 19372
rect 20533 19363 20591 19369
rect 20533 19329 20545 19363
rect 20579 19360 20591 19363
rect 21174 19360 21180 19372
rect 20579 19332 21180 19360
rect 20579 19329 20591 19332
rect 20533 19323 20591 19329
rect 21174 19320 21180 19332
rect 21232 19320 21238 19372
rect 21269 19363 21327 19369
rect 21269 19329 21281 19363
rect 21315 19360 21327 19363
rect 22094 19360 22100 19372
rect 21315 19332 22100 19360
rect 21315 19329 21327 19332
rect 21269 19323 21327 19329
rect 22094 19320 22100 19332
rect 22152 19320 22158 19372
rect 13044 19264 15424 19292
rect 15473 19295 15531 19301
rect 13044 19252 13050 19264
rect 15473 19261 15485 19295
rect 15519 19292 15531 19295
rect 15654 19292 15660 19304
rect 15519 19264 15660 19292
rect 15519 19261 15531 19264
rect 15473 19255 15531 19261
rect 15654 19252 15660 19264
rect 15712 19252 15718 19304
rect 17144 19292 17172 19320
rect 18966 19292 18972 19304
rect 17144 19264 18972 19292
rect 18966 19252 18972 19264
rect 19024 19252 19030 19304
rect 19150 19292 19156 19304
rect 19111 19264 19156 19292
rect 19150 19252 19156 19264
rect 19208 19252 19214 19304
rect 20070 19292 20076 19304
rect 20031 19264 20076 19292
rect 20070 19252 20076 19264
rect 20128 19252 20134 19304
rect 20990 19292 20996 19304
rect 20951 19264 20996 19292
rect 20990 19252 20996 19264
rect 21048 19292 21054 19304
rect 21358 19292 21364 19304
rect 21048 19264 21364 19292
rect 21048 19252 21054 19264
rect 21358 19252 21364 19264
rect 21416 19252 21422 19304
rect 14182 19184 14188 19236
rect 14240 19224 14246 19236
rect 15194 19224 15200 19236
rect 14240 19196 15200 19224
rect 14240 19184 14246 19196
rect 15194 19184 15200 19196
rect 15252 19184 15258 19236
rect 15562 19184 15568 19236
rect 15620 19224 15626 19236
rect 22370 19224 22376 19236
rect 15620 19196 22376 19224
rect 15620 19184 15626 19196
rect 22370 19184 22376 19196
rect 22428 19184 22434 19236
rect 14458 19116 14464 19168
rect 14516 19156 14522 19168
rect 14737 19159 14795 19165
rect 14737 19156 14749 19159
rect 14516 19128 14749 19156
rect 14516 19116 14522 19128
rect 14737 19125 14749 19128
rect 14783 19125 14795 19159
rect 14737 19119 14795 19125
rect 14826 19116 14832 19168
rect 14884 19156 14890 19168
rect 19702 19156 19708 19168
rect 14884 19128 19708 19156
rect 14884 19116 14890 19128
rect 19702 19116 19708 19128
rect 19760 19156 19766 19168
rect 21726 19156 21732 19168
rect 19760 19128 21732 19156
rect 19760 19116 19766 19128
rect 21726 19116 21732 19128
rect 21784 19116 21790 19168
rect 1104 19066 23828 19088
rect 1104 19014 3790 19066
rect 3842 19014 3854 19066
rect 3906 19014 3918 19066
rect 3970 19014 3982 19066
rect 4034 19014 4046 19066
rect 4098 19014 9471 19066
rect 9523 19014 9535 19066
rect 9587 19014 9599 19066
rect 9651 19014 9663 19066
rect 9715 19014 9727 19066
rect 9779 19014 15152 19066
rect 15204 19014 15216 19066
rect 15268 19014 15280 19066
rect 15332 19014 15344 19066
rect 15396 19014 15408 19066
rect 15460 19014 20833 19066
rect 20885 19014 20897 19066
rect 20949 19014 20961 19066
rect 21013 19014 21025 19066
rect 21077 19014 21089 19066
rect 21141 19014 23828 19066
rect 1104 18992 23828 19014
rect 5810 18952 5816 18964
rect 5771 18924 5816 18952
rect 5810 18912 5816 18924
rect 5868 18912 5874 18964
rect 7466 18912 7472 18964
rect 7524 18952 7530 18964
rect 7653 18955 7711 18961
rect 7653 18952 7665 18955
rect 7524 18924 7665 18952
rect 7524 18912 7530 18924
rect 7653 18921 7665 18924
rect 7699 18921 7711 18955
rect 14274 18952 14280 18964
rect 14235 18924 14280 18952
rect 7653 18915 7711 18921
rect 14274 18912 14280 18924
rect 14332 18912 14338 18964
rect 14550 18912 14556 18964
rect 14608 18952 14614 18964
rect 15286 18952 15292 18964
rect 14608 18924 15292 18952
rect 14608 18912 14614 18924
rect 15286 18912 15292 18924
rect 15344 18952 15350 18964
rect 15654 18952 15660 18964
rect 15344 18924 15660 18952
rect 15344 18912 15350 18924
rect 15654 18912 15660 18924
rect 15712 18912 15718 18964
rect 16022 18952 16028 18964
rect 15983 18924 16028 18952
rect 16022 18912 16028 18924
rect 16080 18912 16086 18964
rect 18322 18952 18328 18964
rect 18283 18924 18328 18952
rect 18322 18912 18328 18924
rect 18380 18912 18386 18964
rect 18874 18952 18880 18964
rect 18524 18924 18880 18952
rect 14826 18884 14832 18896
rect 13280 18856 14832 18884
rect 13280 18828 13308 18856
rect 14826 18844 14832 18856
rect 14884 18844 14890 18896
rect 16853 18887 16911 18893
rect 16853 18853 16865 18887
rect 16899 18884 16911 18887
rect 18524 18884 18552 18924
rect 18874 18912 18880 18924
rect 18932 18912 18938 18964
rect 19429 18955 19487 18961
rect 19429 18921 19441 18955
rect 19475 18952 19487 18955
rect 19610 18952 19616 18964
rect 19475 18924 19616 18952
rect 19475 18921 19487 18924
rect 19429 18915 19487 18921
rect 19610 18912 19616 18924
rect 19668 18912 19674 18964
rect 22370 18952 22376 18964
rect 22331 18924 22376 18952
rect 22370 18912 22376 18924
rect 22428 18912 22434 18964
rect 20714 18884 20720 18896
rect 16899 18856 18552 18884
rect 18616 18856 20720 18884
rect 16899 18853 16911 18856
rect 16853 18847 16911 18853
rect 9122 18816 9128 18828
rect 9083 18788 9128 18816
rect 9122 18776 9128 18788
rect 9180 18776 9186 18828
rect 12894 18776 12900 18828
rect 12952 18816 12958 18828
rect 13173 18819 13231 18825
rect 13173 18816 13185 18819
rect 12952 18788 13185 18816
rect 12952 18776 12958 18788
rect 13173 18785 13185 18788
rect 13219 18785 13231 18819
rect 13173 18779 13231 18785
rect 13262 18776 13268 18828
rect 13320 18816 13326 18828
rect 13541 18819 13599 18825
rect 13320 18788 13413 18816
rect 13320 18776 13326 18788
rect 13541 18785 13553 18819
rect 13587 18816 13599 18819
rect 15381 18819 15439 18825
rect 15381 18816 15393 18819
rect 13587 18788 15393 18816
rect 13587 18785 13599 18788
rect 13541 18779 13599 18785
rect 15381 18785 15393 18788
rect 15427 18785 15439 18819
rect 15381 18779 15439 18785
rect 16574 18776 16580 18828
rect 16632 18816 16638 18828
rect 18616 18825 18644 18856
rect 20714 18844 20720 18856
rect 20772 18844 20778 18896
rect 18601 18819 18659 18825
rect 16632 18788 17816 18816
rect 16632 18776 16638 18788
rect 2774 18708 2780 18760
rect 2832 18748 2838 18760
rect 3421 18751 3479 18757
rect 3421 18748 3433 18751
rect 2832 18720 3433 18748
rect 2832 18708 2838 18720
rect 3421 18717 3433 18720
rect 3467 18717 3479 18751
rect 3421 18711 3479 18717
rect 5810 18708 5816 18760
rect 5868 18748 5874 18760
rect 6365 18751 6423 18757
rect 6365 18748 6377 18751
rect 5868 18720 6377 18748
rect 5868 18708 5874 18720
rect 6365 18717 6377 18720
rect 6411 18717 6423 18751
rect 6365 18711 6423 18717
rect 12986 18708 12992 18760
rect 13044 18748 13050 18760
rect 13081 18751 13139 18757
rect 13081 18748 13093 18751
rect 13044 18720 13093 18748
rect 13044 18708 13050 18720
rect 13081 18717 13093 18720
rect 13127 18717 13139 18751
rect 13354 18748 13360 18760
rect 13315 18720 13360 18748
rect 13081 18711 13139 18717
rect 13354 18708 13360 18720
rect 13412 18708 13418 18760
rect 14458 18748 14464 18760
rect 14419 18720 14464 18748
rect 14458 18708 14464 18720
rect 14516 18708 14522 18760
rect 14921 18751 14979 18757
rect 14921 18717 14933 18751
rect 14967 18748 14979 18751
rect 15746 18748 15752 18760
rect 14967 18720 15608 18748
rect 15707 18720 15752 18748
rect 14967 18717 14979 18720
rect 14921 18711 14979 18717
rect 3176 18683 3234 18689
rect 3176 18649 3188 18683
rect 3222 18680 3234 18683
rect 8294 18680 8300 18692
rect 3222 18652 8300 18680
rect 3222 18649 3234 18652
rect 3176 18643 3234 18649
rect 8294 18640 8300 18652
rect 8352 18640 8358 18692
rect 9392 18683 9450 18689
rect 9392 18649 9404 18683
rect 9438 18680 9450 18683
rect 10870 18680 10876 18692
rect 9438 18652 10876 18680
rect 9438 18649 9450 18652
rect 9392 18643 9450 18649
rect 10870 18640 10876 18652
rect 10928 18640 10934 18692
rect 12066 18640 12072 18692
rect 12124 18680 12130 18692
rect 14366 18680 14372 18692
rect 12124 18652 14372 18680
rect 12124 18640 12130 18652
rect 14366 18640 14372 18652
rect 14424 18640 14430 18692
rect 14550 18680 14556 18692
rect 14511 18652 14556 18680
rect 14550 18640 14556 18652
rect 14608 18640 14614 18692
rect 14645 18683 14703 18689
rect 14645 18649 14657 18683
rect 14691 18649 14703 18683
rect 14645 18643 14703 18649
rect 2041 18615 2099 18621
rect 2041 18581 2053 18615
rect 2087 18612 2099 18615
rect 2590 18612 2596 18624
rect 2087 18584 2596 18612
rect 2087 18581 2099 18584
rect 2041 18575 2099 18581
rect 2590 18572 2596 18584
rect 2648 18572 2654 18624
rect 10505 18615 10563 18621
rect 10505 18581 10517 18615
rect 10551 18612 10563 18615
rect 10594 18612 10600 18624
rect 10551 18584 10600 18612
rect 10551 18581 10563 18584
rect 10505 18575 10563 18581
rect 10594 18572 10600 18584
rect 10652 18572 10658 18624
rect 14458 18572 14464 18624
rect 14516 18612 14522 18624
rect 14660 18612 14688 18643
rect 14734 18640 14740 18692
rect 14792 18689 14798 18692
rect 14792 18683 14821 18689
rect 14809 18649 14821 18683
rect 14792 18643 14821 18649
rect 14792 18640 14798 18643
rect 15286 18640 15292 18692
rect 15344 18680 15350 18692
rect 15473 18683 15531 18689
rect 15473 18680 15485 18683
rect 15344 18652 15485 18680
rect 15344 18640 15350 18652
rect 15473 18649 15485 18652
rect 15519 18649 15531 18683
rect 15580 18680 15608 18720
rect 15746 18708 15752 18720
rect 15804 18708 15810 18760
rect 15841 18751 15899 18757
rect 15841 18717 15853 18751
rect 15887 18748 15899 18751
rect 16482 18748 16488 18760
rect 15887 18720 16488 18748
rect 15887 18717 15899 18720
rect 15841 18711 15899 18717
rect 16482 18708 16488 18720
rect 16540 18708 16546 18760
rect 16666 18748 16672 18760
rect 16627 18720 16672 18748
rect 16666 18708 16672 18720
rect 16724 18708 16730 18760
rect 16942 18708 16948 18760
rect 17000 18748 17006 18760
rect 17000 18720 17045 18748
rect 17000 18708 17006 18720
rect 17788 18692 17816 18788
rect 18601 18785 18613 18819
rect 18647 18785 18659 18819
rect 18601 18779 18659 18785
rect 18874 18776 18880 18828
rect 18932 18816 18938 18828
rect 18932 18788 19840 18816
rect 18932 18776 18938 18788
rect 18506 18748 18512 18760
rect 18467 18720 18512 18748
rect 18506 18708 18512 18720
rect 18564 18708 18570 18760
rect 18693 18751 18751 18757
rect 18693 18717 18705 18751
rect 18739 18717 18751 18751
rect 18693 18711 18751 18717
rect 17126 18680 17132 18692
rect 15580 18652 17132 18680
rect 15473 18643 15531 18649
rect 17126 18640 17132 18652
rect 17184 18640 17190 18692
rect 17770 18640 17776 18692
rect 17828 18680 17834 18692
rect 18708 18680 18736 18711
rect 18782 18708 18788 18760
rect 18840 18748 18846 18760
rect 18840 18720 18885 18748
rect 18840 18708 18846 18720
rect 18966 18708 18972 18760
rect 19024 18748 19030 18760
rect 19567 18751 19625 18757
rect 19567 18748 19579 18751
rect 19024 18720 19579 18748
rect 19024 18708 19030 18720
rect 19567 18717 19579 18720
rect 19613 18717 19625 18751
rect 19702 18748 19708 18760
rect 19663 18720 19708 18748
rect 19567 18711 19625 18717
rect 19702 18708 19708 18720
rect 19760 18708 19766 18760
rect 19812 18689 19840 18788
rect 19886 18708 19892 18760
rect 19944 18757 19950 18760
rect 19944 18751 19983 18757
rect 19971 18717 19983 18751
rect 19944 18711 19983 18717
rect 19944 18708 19950 18711
rect 20070 18708 20076 18760
rect 20128 18748 20134 18760
rect 20254 18748 20260 18760
rect 20128 18720 20260 18748
rect 20128 18708 20134 18720
rect 20254 18708 20260 18720
rect 20312 18708 20318 18760
rect 20438 18708 20444 18760
rect 20496 18748 20502 18760
rect 20717 18751 20775 18757
rect 20717 18748 20729 18751
rect 20496 18720 20729 18748
rect 20496 18708 20502 18720
rect 20717 18717 20729 18720
rect 20763 18717 20775 18751
rect 20717 18711 20775 18717
rect 20993 18751 21051 18757
rect 20993 18717 21005 18751
rect 21039 18748 21051 18751
rect 21174 18748 21180 18760
rect 21039 18720 21180 18748
rect 21039 18717 21051 18720
rect 20993 18711 21051 18717
rect 21174 18708 21180 18720
rect 21232 18748 21238 18760
rect 22097 18751 22155 18757
rect 22097 18748 22109 18751
rect 21232 18720 22109 18748
rect 21232 18708 21238 18720
rect 22097 18717 22109 18720
rect 22143 18717 22155 18751
rect 22097 18711 22155 18717
rect 17828 18652 18736 18680
rect 19797 18683 19855 18689
rect 17828 18640 17834 18652
rect 19797 18649 19809 18683
rect 19843 18680 19855 18683
rect 20622 18680 20628 18692
rect 19843 18652 20628 18680
rect 19843 18649 19855 18652
rect 19797 18643 19855 18649
rect 20622 18640 20628 18652
rect 20680 18640 20686 18692
rect 22281 18683 22339 18689
rect 22281 18649 22293 18683
rect 22327 18649 22339 18683
rect 22281 18643 22339 18649
rect 14516 18584 14688 18612
rect 14516 18572 14522 18584
rect 15654 18572 15660 18624
rect 15712 18612 15718 18624
rect 16485 18615 16543 18621
rect 16485 18612 16497 18615
rect 15712 18584 16497 18612
rect 15712 18572 15718 18584
rect 16485 18581 16497 18584
rect 16531 18581 16543 18615
rect 16485 18575 16543 18581
rect 17402 18572 17408 18624
rect 17460 18612 17466 18624
rect 20533 18615 20591 18621
rect 20533 18612 20545 18615
rect 17460 18584 20545 18612
rect 17460 18572 17466 18584
rect 20533 18581 20545 18584
rect 20579 18581 20591 18615
rect 20898 18612 20904 18624
rect 20859 18584 20904 18612
rect 20533 18575 20591 18581
rect 20898 18572 20904 18584
rect 20956 18572 20962 18624
rect 22094 18572 22100 18624
rect 22152 18612 22158 18624
rect 22296 18612 22324 18643
rect 22152 18584 22324 18612
rect 22152 18572 22158 18584
rect 1104 18522 23987 18544
rect 1104 18470 6630 18522
rect 6682 18470 6694 18522
rect 6746 18470 6758 18522
rect 6810 18470 6822 18522
rect 6874 18470 6886 18522
rect 6938 18470 12311 18522
rect 12363 18470 12375 18522
rect 12427 18470 12439 18522
rect 12491 18470 12503 18522
rect 12555 18470 12567 18522
rect 12619 18470 17992 18522
rect 18044 18470 18056 18522
rect 18108 18470 18120 18522
rect 18172 18470 18184 18522
rect 18236 18470 18248 18522
rect 18300 18470 23673 18522
rect 23725 18470 23737 18522
rect 23789 18470 23801 18522
rect 23853 18470 23865 18522
rect 23917 18470 23929 18522
rect 23981 18470 23987 18522
rect 1104 18448 23987 18470
rect 9122 18408 9128 18420
rect 9083 18380 9128 18408
rect 9122 18368 9128 18380
rect 9180 18368 9186 18420
rect 13538 18408 13544 18420
rect 13499 18380 13544 18408
rect 13538 18368 13544 18380
rect 13596 18368 13602 18420
rect 14645 18411 14703 18417
rect 14645 18377 14657 18411
rect 14691 18408 14703 18411
rect 14734 18408 14740 18420
rect 14691 18380 14740 18408
rect 14691 18377 14703 18380
rect 14645 18371 14703 18377
rect 14734 18368 14740 18380
rect 14792 18368 14798 18420
rect 16482 18368 16488 18420
rect 16540 18408 16546 18420
rect 17218 18408 17224 18420
rect 16540 18380 17224 18408
rect 16540 18368 16546 18380
rect 17218 18368 17224 18380
rect 17276 18408 17282 18420
rect 17276 18380 18736 18408
rect 17276 18368 17282 18380
rect 7466 18300 7472 18352
rect 7524 18340 7530 18352
rect 7837 18343 7895 18349
rect 7837 18340 7849 18343
rect 7524 18312 7849 18340
rect 7524 18300 7530 18312
rect 7837 18309 7849 18312
rect 7883 18309 7895 18343
rect 13998 18340 14004 18352
rect 7837 18303 7895 18309
rect 13096 18312 14004 18340
rect 2314 18232 2320 18284
rect 2372 18272 2378 18284
rect 13096 18281 13124 18312
rect 13998 18300 14004 18312
rect 14056 18300 14062 18352
rect 14277 18343 14335 18349
rect 14277 18309 14289 18343
rect 14323 18340 14335 18343
rect 16114 18340 16120 18352
rect 14323 18312 16120 18340
rect 14323 18309 14335 18312
rect 14277 18303 14335 18309
rect 16114 18300 16120 18312
rect 16172 18300 16178 18352
rect 18708 18340 18736 18380
rect 18782 18368 18788 18420
rect 18840 18408 18846 18420
rect 19797 18411 19855 18417
rect 19797 18408 19809 18411
rect 18840 18380 19809 18408
rect 18840 18368 18846 18380
rect 19797 18377 19809 18380
rect 19843 18377 19855 18411
rect 19797 18371 19855 18377
rect 19886 18368 19892 18420
rect 19944 18408 19950 18420
rect 20901 18411 20959 18417
rect 20901 18408 20913 18411
rect 19944 18380 20913 18408
rect 19944 18368 19950 18380
rect 20901 18377 20913 18380
rect 20947 18408 20959 18411
rect 21450 18408 21456 18420
rect 20947 18380 21456 18408
rect 20947 18377 20959 18380
rect 20901 18371 20959 18377
rect 21450 18368 21456 18380
rect 21508 18368 21514 18420
rect 22005 18411 22063 18417
rect 22005 18377 22017 18411
rect 22051 18408 22063 18411
rect 22186 18408 22192 18420
rect 22051 18380 22192 18408
rect 22051 18377 22063 18380
rect 22005 18371 22063 18377
rect 22186 18368 22192 18380
rect 22244 18368 22250 18420
rect 22370 18408 22376 18420
rect 22296 18380 22376 18408
rect 19242 18340 19248 18352
rect 18708 18312 19248 18340
rect 19242 18300 19248 18312
rect 19300 18300 19306 18352
rect 20346 18340 20352 18352
rect 20088 18312 20352 18340
rect 2869 18275 2927 18281
rect 2869 18272 2881 18275
rect 2372 18244 2881 18272
rect 2372 18232 2378 18244
rect 2869 18241 2881 18244
rect 2915 18241 2927 18275
rect 2869 18235 2927 18241
rect 13081 18275 13139 18281
rect 13081 18241 13093 18275
rect 13127 18241 13139 18275
rect 13081 18235 13139 18241
rect 13365 18278 13423 18281
rect 13365 18275 13492 18278
rect 13365 18241 13377 18275
rect 13411 18272 13492 18275
rect 14185 18275 14243 18281
rect 13411 18250 14136 18272
rect 13411 18241 13423 18250
rect 13464 18244 14136 18250
rect 13365 18235 13423 18241
rect 2593 18207 2651 18213
rect 2593 18173 2605 18207
rect 2639 18204 2651 18207
rect 2774 18204 2780 18216
rect 2639 18176 2780 18204
rect 2639 18173 2651 18176
rect 2593 18167 2651 18173
rect 2774 18164 2780 18176
rect 2832 18164 2838 18216
rect 12894 18164 12900 18216
rect 12952 18204 12958 18216
rect 13173 18207 13231 18213
rect 13173 18204 13185 18207
rect 12952 18176 13185 18204
rect 12952 18164 12958 18176
rect 13173 18173 13185 18176
rect 13219 18173 13231 18207
rect 13173 18167 13231 18173
rect 13287 18207 13345 18213
rect 13287 18173 13299 18207
rect 13333 18173 13345 18207
rect 13287 18167 13345 18173
rect 13290 18080 13318 18167
rect 3326 18028 3332 18080
rect 3384 18068 3390 18080
rect 4157 18071 4215 18077
rect 4157 18068 4169 18071
rect 3384 18040 4169 18068
rect 3384 18028 3390 18040
rect 4157 18037 4169 18040
rect 4203 18037 4215 18071
rect 4157 18031 4215 18037
rect 13262 18028 13268 18080
rect 13320 18028 13326 18080
rect 14108 18068 14136 18244
rect 14185 18241 14197 18275
rect 14231 18241 14243 18275
rect 14185 18235 14243 18241
rect 14461 18275 14519 18281
rect 14461 18241 14473 18275
rect 14507 18272 14519 18275
rect 14826 18272 14832 18284
rect 14507 18244 14832 18272
rect 14507 18241 14519 18244
rect 14461 18235 14519 18241
rect 14200 18204 14228 18235
rect 14826 18232 14832 18244
rect 14884 18232 14890 18284
rect 16945 18275 17003 18281
rect 16945 18241 16957 18275
rect 16991 18241 17003 18275
rect 16945 18235 17003 18241
rect 17129 18275 17187 18281
rect 17129 18241 17141 18275
rect 17175 18272 17187 18275
rect 18690 18272 18696 18284
rect 17175 18244 18696 18272
rect 17175 18241 17187 18244
rect 17129 18235 17187 18241
rect 15470 18204 15476 18216
rect 14200 18176 15476 18204
rect 15470 18164 15476 18176
rect 15528 18164 15534 18216
rect 16960 18204 16988 18235
rect 18690 18232 18696 18244
rect 18748 18232 18754 18284
rect 19702 18232 19708 18284
rect 19760 18272 19766 18284
rect 20088 18281 20116 18312
rect 20346 18300 20352 18312
rect 20404 18300 20410 18352
rect 22296 18340 22324 18380
rect 22370 18368 22376 18380
rect 22428 18368 22434 18420
rect 22296 18312 22416 18340
rect 22388 18284 22416 18312
rect 20159 18281 20165 18284
rect 20053 18275 20116 18281
rect 20053 18272 20065 18275
rect 19760 18244 20065 18272
rect 19760 18232 19766 18244
rect 20053 18241 20065 18244
rect 20099 18244 20116 18275
rect 20146 18275 20165 18281
rect 20099 18241 20111 18244
rect 20053 18235 20111 18241
rect 20146 18241 20158 18275
rect 20146 18235 20165 18241
rect 20159 18232 20165 18235
rect 20217 18232 20223 18284
rect 20254 18232 20260 18284
rect 20312 18281 20318 18284
rect 20312 18272 20320 18281
rect 20441 18275 20499 18281
rect 20312 18244 20357 18272
rect 20312 18235 20320 18244
rect 20441 18241 20453 18275
rect 20487 18241 20499 18275
rect 22278 18272 22284 18284
rect 22239 18244 22284 18272
rect 20441 18235 20499 18241
rect 20312 18232 20318 18235
rect 18414 18204 18420 18216
rect 16960 18176 18420 18204
rect 18414 18164 18420 18176
rect 18472 18164 18478 18216
rect 20456 18204 20484 18235
rect 22278 18232 22284 18244
rect 22336 18232 22342 18284
rect 22370 18278 22428 18284
rect 22370 18244 22382 18278
rect 22416 18244 22428 18278
rect 22370 18238 22428 18244
rect 22462 18232 22468 18284
rect 22520 18272 22526 18284
rect 22646 18272 22652 18284
rect 22520 18244 22565 18272
rect 22607 18244 22652 18272
rect 22520 18232 22526 18244
rect 22646 18232 22652 18244
rect 22704 18232 22710 18284
rect 22664 18204 22692 18232
rect 19904 18176 22692 18204
rect 14458 18096 14464 18148
rect 14516 18136 14522 18148
rect 15657 18139 15715 18145
rect 15657 18136 15669 18139
rect 14516 18108 15669 18136
rect 14516 18096 14522 18108
rect 15657 18105 15669 18108
rect 15703 18136 15715 18139
rect 16850 18136 16856 18148
rect 15703 18108 16856 18136
rect 15703 18105 15715 18108
rect 15657 18099 15715 18105
rect 16850 18096 16856 18108
rect 16908 18096 16914 18148
rect 19904 18080 19932 18176
rect 15197 18071 15255 18077
rect 15197 18068 15209 18071
rect 14108 18040 15209 18068
rect 15197 18037 15209 18040
rect 15243 18068 15255 18071
rect 16022 18068 16028 18080
rect 15243 18040 16028 18068
rect 15243 18037 15255 18040
rect 15197 18031 15255 18037
rect 16022 18028 16028 18040
rect 16080 18028 16086 18080
rect 16114 18028 16120 18080
rect 16172 18068 16178 18080
rect 16209 18071 16267 18077
rect 16209 18068 16221 18071
rect 16172 18040 16221 18068
rect 16172 18028 16178 18040
rect 16209 18037 16221 18040
rect 16255 18037 16267 18071
rect 16942 18068 16948 18080
rect 16903 18040 16948 18068
rect 16209 18031 16267 18037
rect 16942 18028 16948 18040
rect 17000 18028 17006 18080
rect 17310 18028 17316 18080
rect 17368 18068 17374 18080
rect 17589 18071 17647 18077
rect 17589 18068 17601 18071
rect 17368 18040 17601 18068
rect 17368 18028 17374 18040
rect 17589 18037 17601 18040
rect 17635 18037 17647 18071
rect 17589 18031 17647 18037
rect 19337 18071 19395 18077
rect 19337 18037 19349 18071
rect 19383 18068 19395 18071
rect 19886 18068 19892 18080
rect 19383 18040 19892 18068
rect 19383 18037 19395 18040
rect 19337 18031 19395 18037
rect 19886 18028 19892 18040
rect 19944 18028 19950 18080
rect 1104 17978 23828 18000
rect 1104 17926 3790 17978
rect 3842 17926 3854 17978
rect 3906 17926 3918 17978
rect 3970 17926 3982 17978
rect 4034 17926 4046 17978
rect 4098 17926 9471 17978
rect 9523 17926 9535 17978
rect 9587 17926 9599 17978
rect 9651 17926 9663 17978
rect 9715 17926 9727 17978
rect 9779 17926 15152 17978
rect 15204 17926 15216 17978
rect 15268 17926 15280 17978
rect 15332 17926 15344 17978
rect 15396 17926 15408 17978
rect 15460 17926 20833 17978
rect 20885 17926 20897 17978
rect 20949 17926 20961 17978
rect 21013 17926 21025 17978
rect 21077 17926 21089 17978
rect 21141 17926 23828 17978
rect 1104 17904 23828 17926
rect 13265 17867 13323 17873
rect 13265 17833 13277 17867
rect 13311 17864 13323 17867
rect 14550 17864 14556 17876
rect 13311 17836 14556 17864
rect 13311 17833 13323 17836
rect 13265 17827 13323 17833
rect 14550 17824 14556 17836
rect 14608 17824 14614 17876
rect 18506 17824 18512 17876
rect 18564 17864 18570 17876
rect 19429 17867 19487 17873
rect 19429 17864 19441 17867
rect 18564 17836 19441 17864
rect 18564 17824 18570 17836
rect 19429 17833 19441 17836
rect 19475 17833 19487 17867
rect 19794 17864 19800 17876
rect 19755 17836 19800 17864
rect 19429 17827 19487 17833
rect 19794 17824 19800 17836
rect 19852 17824 19858 17876
rect 22646 17864 22652 17876
rect 22607 17836 22652 17864
rect 22646 17824 22652 17836
rect 22704 17824 22710 17876
rect 12158 17756 12164 17808
rect 12216 17796 12222 17808
rect 12216 17768 18920 17796
rect 12216 17756 12222 17768
rect 7098 17688 7104 17740
rect 7156 17728 7162 17740
rect 8018 17728 8024 17740
rect 7156 17700 8024 17728
rect 7156 17688 7162 17700
rect 8018 17688 8024 17700
rect 8076 17688 8082 17740
rect 9122 17728 9128 17740
rect 9083 17700 9128 17728
rect 9122 17688 9128 17700
rect 9180 17688 9186 17740
rect 17681 17731 17739 17737
rect 17681 17697 17693 17731
rect 17727 17728 17739 17731
rect 17770 17728 17776 17740
rect 17727 17700 17776 17728
rect 17727 17697 17739 17700
rect 17681 17691 17739 17697
rect 17770 17688 17776 17700
rect 17828 17688 17834 17740
rect 2041 17663 2099 17669
rect 2041 17629 2053 17663
rect 2087 17660 2099 17663
rect 2682 17660 2688 17672
rect 2087 17632 2688 17660
rect 2087 17629 2099 17632
rect 2041 17623 2099 17629
rect 2682 17620 2688 17632
rect 2740 17620 2746 17672
rect 9392 17663 9450 17669
rect 9392 17629 9404 17663
rect 9438 17660 9450 17663
rect 12066 17660 12072 17672
rect 9438 17632 12072 17660
rect 9438 17629 9450 17632
rect 9392 17623 9450 17629
rect 12066 17620 12072 17632
rect 12124 17620 12130 17672
rect 12805 17663 12863 17669
rect 12805 17629 12817 17663
rect 12851 17629 12863 17663
rect 12805 17623 12863 17629
rect 13081 17663 13139 17669
rect 13081 17629 13093 17663
rect 13127 17660 13139 17663
rect 13127 17632 13768 17660
rect 13127 17629 13139 17632
rect 13081 17623 13139 17629
rect 2308 17595 2366 17601
rect 2308 17561 2320 17595
rect 2354 17592 2366 17595
rect 2406 17592 2412 17604
rect 2354 17564 2412 17592
rect 2354 17561 2366 17564
rect 2308 17555 2366 17561
rect 2406 17552 2412 17564
rect 2464 17552 2470 17604
rect 6362 17552 6368 17604
rect 6420 17592 6426 17604
rect 6834 17595 6892 17601
rect 6834 17592 6846 17595
rect 6420 17564 6846 17592
rect 6420 17552 6426 17564
rect 6834 17561 6846 17564
rect 6880 17561 6892 17595
rect 12820 17592 12848 17623
rect 13262 17592 13268 17604
rect 12820 17564 13268 17592
rect 6834 17555 6892 17561
rect 13262 17552 13268 17564
rect 13320 17552 13326 17604
rect 13740 17592 13768 17632
rect 13814 17620 13820 17672
rect 13872 17660 13878 17672
rect 14458 17660 14464 17672
rect 13872 17632 14464 17660
rect 13872 17620 13878 17632
rect 14458 17620 14464 17632
rect 14516 17620 14522 17672
rect 16209 17663 16267 17669
rect 16209 17629 16221 17663
rect 16255 17660 16267 17663
rect 16298 17660 16304 17672
rect 16255 17632 16304 17660
rect 16255 17629 16267 17632
rect 16209 17623 16267 17629
rect 16298 17620 16304 17632
rect 16356 17620 16362 17672
rect 16482 17660 16488 17672
rect 16443 17632 16488 17660
rect 16482 17620 16488 17632
rect 16540 17620 16546 17672
rect 17405 17663 17463 17669
rect 17405 17629 17417 17663
rect 17451 17629 17463 17663
rect 17405 17623 17463 17629
rect 14826 17592 14832 17604
rect 13740 17564 14832 17592
rect 14826 17552 14832 17564
rect 14884 17592 14890 17604
rect 14921 17595 14979 17601
rect 14921 17592 14933 17595
rect 14884 17564 14933 17592
rect 14884 17552 14890 17564
rect 14921 17561 14933 17564
rect 14967 17592 14979 17595
rect 15473 17595 15531 17601
rect 15473 17592 15485 17595
rect 14967 17564 15485 17592
rect 14967 17561 14979 17564
rect 14921 17555 14979 17561
rect 15473 17561 15485 17564
rect 15519 17592 15531 17595
rect 17310 17592 17316 17604
rect 15519 17564 17316 17592
rect 15519 17561 15531 17564
rect 15473 17555 15531 17561
rect 17310 17552 17316 17564
rect 17368 17552 17374 17604
rect 17420 17592 17448 17623
rect 17494 17620 17500 17672
rect 17552 17660 17558 17672
rect 17589 17663 17647 17669
rect 17589 17660 17601 17663
rect 17552 17632 17601 17660
rect 17552 17620 17558 17632
rect 17589 17629 17601 17632
rect 17635 17629 17647 17663
rect 17589 17623 17647 17629
rect 17862 17620 17868 17672
rect 17920 17660 17926 17672
rect 18141 17663 18199 17669
rect 18141 17660 18153 17663
rect 17920 17632 18153 17660
rect 17920 17620 17926 17632
rect 18141 17629 18153 17632
rect 18187 17629 18199 17663
rect 18141 17623 18199 17629
rect 18233 17663 18291 17669
rect 18233 17629 18245 17663
rect 18279 17660 18291 17663
rect 18322 17660 18328 17672
rect 18279 17632 18328 17660
rect 18279 17629 18291 17632
rect 18233 17623 18291 17629
rect 18322 17620 18328 17632
rect 18380 17620 18386 17672
rect 18892 17669 18920 17768
rect 19702 17728 19708 17740
rect 19663 17700 19708 17728
rect 19702 17688 19708 17700
rect 19760 17688 19766 17740
rect 18877 17663 18935 17669
rect 18877 17629 18889 17663
rect 18923 17660 18935 17663
rect 19797 17663 19855 17669
rect 19797 17660 19809 17663
rect 18923 17632 19809 17660
rect 18923 17629 18935 17632
rect 18877 17623 18935 17629
rect 19797 17629 19809 17632
rect 19843 17660 19855 17663
rect 19978 17660 19984 17672
rect 19843 17632 19984 17660
rect 19843 17629 19855 17632
rect 19797 17623 19855 17629
rect 19978 17620 19984 17632
rect 20036 17620 20042 17672
rect 20070 17620 20076 17672
rect 20128 17660 20134 17672
rect 21818 17660 21824 17672
rect 20128 17632 21824 17660
rect 20128 17620 20134 17632
rect 21818 17620 21824 17632
rect 21876 17620 21882 17672
rect 22097 17663 22155 17669
rect 22097 17629 22109 17663
rect 22143 17629 22155 17663
rect 22097 17623 22155 17629
rect 19334 17592 19340 17604
rect 17420 17564 19340 17592
rect 19334 17552 19340 17564
rect 19392 17552 19398 17604
rect 19426 17552 19432 17604
rect 19484 17592 19490 17604
rect 22112 17592 22140 17623
rect 19484 17564 22140 17592
rect 19484 17552 19490 17564
rect 2958 17484 2964 17536
rect 3016 17524 3022 17536
rect 3421 17527 3479 17533
rect 3421 17524 3433 17527
rect 3016 17496 3433 17524
rect 3016 17484 3022 17496
rect 3421 17493 3433 17496
rect 3467 17493 3479 17527
rect 3421 17487 3479 17493
rect 5534 17484 5540 17536
rect 5592 17524 5598 17536
rect 5721 17527 5779 17533
rect 5721 17524 5733 17527
rect 5592 17496 5733 17524
rect 5592 17484 5598 17496
rect 5721 17493 5733 17496
rect 5767 17493 5779 17527
rect 5721 17487 5779 17493
rect 10410 17484 10416 17536
rect 10468 17524 10474 17536
rect 10505 17527 10563 17533
rect 10505 17524 10517 17527
rect 10468 17496 10517 17524
rect 10468 17484 10474 17496
rect 10505 17493 10517 17496
rect 10551 17493 10563 17527
rect 10505 17487 10563 17493
rect 11790 17484 11796 17536
rect 11848 17524 11854 17536
rect 12894 17524 12900 17536
rect 11848 17496 12900 17524
rect 11848 17484 11854 17496
rect 12894 17484 12900 17496
rect 12952 17524 12958 17536
rect 14369 17527 14427 17533
rect 14369 17524 14381 17527
rect 12952 17496 14381 17524
rect 12952 17484 12958 17496
rect 14369 17493 14381 17496
rect 14415 17493 14427 17527
rect 14369 17487 14427 17493
rect 15838 17484 15844 17536
rect 15896 17524 15902 17536
rect 16025 17527 16083 17533
rect 16025 17524 16037 17527
rect 15896 17496 16037 17524
rect 15896 17484 15902 17496
rect 16025 17493 16037 17496
rect 16071 17493 16083 17527
rect 16390 17524 16396 17536
rect 16351 17496 16396 17524
rect 16025 17487 16083 17493
rect 16390 17484 16396 17496
rect 16448 17484 16454 17536
rect 16574 17484 16580 17536
rect 16632 17524 16638 17536
rect 17221 17527 17279 17533
rect 17221 17524 17233 17527
rect 16632 17496 17233 17524
rect 16632 17484 16638 17496
rect 17221 17493 17233 17496
rect 17267 17493 17279 17527
rect 17221 17487 17279 17493
rect 17586 17484 17592 17536
rect 17644 17524 17650 17536
rect 20806 17524 20812 17536
rect 17644 17496 20812 17524
rect 17644 17484 17650 17496
rect 20806 17484 20812 17496
rect 20864 17484 20870 17536
rect 20898 17484 20904 17536
rect 20956 17524 20962 17536
rect 21637 17527 21695 17533
rect 21637 17524 21649 17527
rect 20956 17496 21649 17524
rect 20956 17484 20962 17496
rect 21637 17493 21649 17496
rect 21683 17493 21695 17527
rect 22002 17524 22008 17536
rect 21963 17496 22008 17524
rect 21637 17487 21695 17493
rect 22002 17484 22008 17496
rect 22060 17484 22066 17536
rect 1104 17434 23987 17456
rect 1104 17382 6630 17434
rect 6682 17382 6694 17434
rect 6746 17382 6758 17434
rect 6810 17382 6822 17434
rect 6874 17382 6886 17434
rect 6938 17382 12311 17434
rect 12363 17382 12375 17434
rect 12427 17382 12439 17434
rect 12491 17382 12503 17434
rect 12555 17382 12567 17434
rect 12619 17382 17992 17434
rect 18044 17382 18056 17434
rect 18108 17382 18120 17434
rect 18172 17382 18184 17434
rect 18236 17382 18248 17434
rect 18300 17382 23673 17434
rect 23725 17382 23737 17434
rect 23789 17382 23801 17434
rect 23853 17382 23865 17434
rect 23917 17382 23929 17434
rect 23981 17382 23987 17434
rect 1104 17360 23987 17382
rect 12158 17320 12164 17332
rect 12119 17292 12164 17320
rect 12158 17280 12164 17292
rect 12216 17280 12222 17332
rect 12621 17323 12679 17329
rect 12621 17320 12633 17323
rect 12406 17292 12633 17320
rect 10870 17212 10876 17264
rect 10928 17252 10934 17264
rect 12406 17252 12434 17292
rect 12621 17289 12633 17292
rect 12667 17289 12679 17323
rect 13998 17320 14004 17332
rect 13959 17292 14004 17320
rect 12621 17283 12679 17289
rect 13998 17280 14004 17292
rect 14056 17280 14062 17332
rect 14090 17280 14096 17332
rect 14148 17320 14154 17332
rect 14148 17292 16804 17320
rect 14148 17280 14154 17292
rect 15010 17252 15016 17264
rect 10928 17224 12434 17252
rect 12912 17224 15016 17252
rect 10928 17212 10934 17224
rect 8018 17144 8024 17196
rect 8076 17184 8082 17196
rect 8202 17184 8208 17196
rect 8076 17156 8208 17184
rect 8076 17144 8082 17156
rect 8202 17144 8208 17156
rect 8260 17184 8266 17196
rect 12912 17193 12940 17224
rect 15010 17212 15016 17224
rect 15068 17212 15074 17264
rect 16776 17252 16804 17292
rect 18874 17280 18880 17332
rect 18932 17320 18938 17332
rect 19061 17323 19119 17329
rect 19061 17320 19073 17323
rect 18932 17292 19073 17320
rect 18932 17280 18938 17292
rect 19061 17289 19073 17292
rect 19107 17289 19119 17323
rect 19061 17283 19119 17289
rect 19518 17280 19524 17332
rect 19576 17320 19582 17332
rect 19705 17323 19763 17329
rect 19705 17320 19717 17323
rect 19576 17292 19717 17320
rect 19576 17280 19582 17292
rect 19705 17289 19717 17292
rect 19751 17289 19763 17323
rect 20714 17320 20720 17332
rect 20675 17292 20720 17320
rect 19705 17283 19763 17289
rect 20714 17280 20720 17292
rect 20772 17280 20778 17332
rect 16945 17255 17003 17261
rect 16776 17224 16896 17252
rect 8849 17187 8907 17193
rect 8849 17184 8861 17187
rect 8260 17156 8861 17184
rect 8260 17144 8266 17156
rect 8849 17153 8861 17156
rect 8895 17153 8907 17187
rect 8849 17147 8907 17153
rect 12805 17187 12863 17193
rect 12805 17153 12817 17187
rect 12851 17153 12863 17187
rect 12805 17147 12863 17153
rect 12897 17187 12955 17193
rect 12897 17153 12909 17187
rect 12943 17153 12955 17187
rect 13170 17184 13176 17196
rect 13131 17156 13176 17184
rect 12897 17147 12955 17153
rect 2682 17116 2688 17128
rect 2643 17088 2688 17116
rect 2682 17076 2688 17088
rect 2740 17076 2746 17128
rect 2961 17119 3019 17125
rect 2961 17085 2973 17119
rect 3007 17116 3019 17119
rect 5074 17116 5080 17128
rect 3007 17088 5080 17116
rect 3007 17085 3019 17088
rect 2961 17079 3019 17085
rect 5074 17076 5080 17088
rect 5132 17076 5138 17128
rect 9125 17119 9183 17125
rect 9125 17085 9137 17119
rect 9171 17116 9183 17119
rect 12820 17116 12848 17147
rect 13170 17144 13176 17156
rect 13228 17144 13234 17196
rect 14277 17187 14335 17193
rect 14277 17153 14289 17187
rect 14323 17184 14335 17187
rect 14550 17184 14556 17196
rect 14323 17156 14556 17184
rect 14323 17153 14335 17156
rect 14277 17147 14335 17153
rect 14550 17144 14556 17156
rect 14608 17144 14614 17196
rect 15473 17187 15531 17193
rect 15473 17153 15485 17187
rect 15519 17184 15531 17187
rect 15930 17184 15936 17196
rect 15519 17156 15936 17184
rect 15519 17153 15531 17156
rect 15473 17147 15531 17153
rect 15930 17144 15936 17156
rect 15988 17144 15994 17196
rect 16868 17193 16896 17224
rect 16945 17221 16957 17255
rect 16991 17252 17003 17255
rect 17310 17252 17316 17264
rect 16991 17224 17316 17252
rect 16991 17221 17003 17224
rect 16945 17215 17003 17221
rect 17310 17212 17316 17224
rect 17368 17212 17374 17264
rect 20070 17252 20076 17264
rect 17880 17224 20076 17252
rect 16853 17187 16911 17193
rect 16853 17153 16865 17187
rect 16899 17184 16911 17187
rect 17034 17184 17040 17196
rect 16899 17156 17040 17184
rect 16899 17153 16911 17156
rect 16853 17147 16911 17153
rect 17034 17144 17040 17156
rect 17092 17144 17098 17196
rect 17880 17193 17908 17224
rect 20070 17212 20076 17224
rect 20128 17212 20134 17264
rect 17129 17187 17187 17193
rect 17129 17153 17141 17187
rect 17175 17184 17187 17187
rect 17865 17187 17923 17193
rect 17865 17184 17877 17187
rect 17175 17156 17877 17184
rect 17175 17153 17187 17156
rect 17129 17147 17187 17153
rect 17865 17153 17877 17156
rect 17911 17153 17923 17187
rect 17865 17147 17923 17153
rect 13630 17116 13636 17128
rect 9171 17088 11100 17116
rect 12820 17088 13636 17116
rect 9171 17085 9183 17088
rect 9125 17079 9183 17085
rect 11072 17057 11100 17088
rect 13630 17076 13636 17088
rect 13688 17076 13694 17128
rect 14090 17076 14096 17128
rect 14148 17116 14154 17128
rect 14185 17119 14243 17125
rect 14185 17116 14197 17119
rect 14148 17088 14197 17116
rect 14148 17076 14154 17088
rect 14185 17085 14197 17088
rect 14231 17085 14243 17119
rect 14185 17079 14243 17085
rect 14369 17119 14427 17125
rect 14369 17085 14381 17119
rect 14415 17085 14427 17119
rect 14369 17079 14427 17085
rect 11057 17051 11115 17057
rect 11057 17017 11069 17051
rect 11103 17048 11115 17051
rect 11882 17048 11888 17060
rect 11103 17020 11888 17048
rect 11103 17017 11115 17020
rect 11057 17011 11115 17017
rect 11882 17008 11888 17020
rect 11940 17008 11946 17060
rect 13078 17048 13084 17060
rect 13039 17020 13084 17048
rect 13078 17008 13084 17020
rect 13136 17008 13142 17060
rect 14274 17008 14280 17060
rect 14332 17048 14338 17060
rect 14384 17048 14412 17079
rect 14458 17076 14464 17128
rect 14516 17116 14522 17128
rect 15102 17116 15108 17128
rect 14516 17088 15108 17116
rect 14516 17076 14522 17088
rect 15102 17076 15108 17088
rect 15160 17076 15166 17128
rect 15286 17076 15292 17128
rect 15344 17116 15350 17128
rect 15746 17116 15752 17128
rect 15344 17088 15752 17116
rect 15344 17076 15350 17088
rect 15746 17076 15752 17088
rect 15804 17116 15810 17128
rect 16390 17116 16396 17128
rect 15804 17088 16396 17116
rect 15804 17076 15810 17088
rect 16390 17076 16396 17088
rect 16448 17116 16454 17128
rect 17144 17116 17172 17147
rect 18414 17144 18420 17196
rect 18472 17184 18478 17196
rect 18969 17187 19027 17193
rect 18969 17184 18981 17187
rect 18472 17156 18981 17184
rect 18472 17144 18478 17156
rect 18969 17153 18981 17156
rect 19015 17153 19027 17187
rect 18969 17147 19027 17153
rect 19242 17144 19248 17196
rect 19300 17184 19306 17196
rect 19337 17187 19395 17193
rect 19337 17184 19349 17187
rect 19300 17156 19349 17184
rect 19300 17144 19306 17156
rect 19337 17153 19349 17156
rect 19383 17153 19395 17187
rect 20898 17184 20904 17196
rect 20859 17156 20904 17184
rect 19337 17147 19395 17153
rect 20898 17144 20904 17156
rect 20956 17144 20962 17196
rect 20993 17187 21051 17193
rect 20993 17153 21005 17187
rect 21039 17184 21051 17187
rect 22278 17184 22284 17196
rect 21039 17156 22284 17184
rect 21039 17153 21051 17156
rect 20993 17147 21051 17153
rect 22278 17144 22284 17156
rect 22336 17144 22342 17196
rect 16448 17088 17172 17116
rect 18141 17119 18199 17125
rect 16448 17076 16454 17088
rect 18141 17085 18153 17119
rect 18187 17116 18199 17119
rect 18782 17116 18788 17128
rect 18187 17088 18788 17116
rect 18187 17085 18199 17088
rect 18141 17079 18199 17085
rect 18782 17076 18788 17088
rect 18840 17076 18846 17128
rect 20714 17116 20720 17128
rect 20675 17088 20720 17116
rect 20714 17076 20720 17088
rect 20772 17076 20778 17128
rect 20806 17076 20812 17128
rect 20864 17116 20870 17128
rect 22370 17116 22376 17128
rect 20864 17088 22376 17116
rect 20864 17076 20870 17088
rect 22370 17076 22376 17088
rect 22428 17076 22434 17128
rect 14332 17020 14412 17048
rect 14332 17008 14338 17020
rect 14734 17008 14740 17060
rect 14792 17048 14798 17060
rect 17126 17048 17132 17060
rect 14792 17020 16528 17048
rect 17087 17020 17132 17048
rect 14792 17008 14798 17020
rect 4249 16983 4307 16989
rect 4249 16949 4261 16983
rect 4295 16980 4307 16983
rect 5350 16980 5356 16992
rect 4295 16952 5356 16980
rect 4295 16949 4307 16952
rect 4249 16943 4307 16949
rect 5350 16940 5356 16952
rect 5408 16940 5414 16992
rect 8386 16980 8392 16992
rect 8299 16952 8392 16980
rect 8386 16940 8392 16952
rect 8444 16980 8450 16992
rect 9214 16980 9220 16992
rect 8444 16952 9220 16980
rect 8444 16940 8450 16952
rect 9214 16940 9220 16952
rect 9272 16940 9278 16992
rect 10413 16983 10471 16989
rect 10413 16949 10425 16983
rect 10459 16980 10471 16983
rect 11698 16980 11704 16992
rect 10459 16952 11704 16980
rect 10459 16949 10471 16952
rect 10413 16943 10471 16949
rect 11698 16940 11704 16952
rect 11756 16940 11762 16992
rect 14366 16940 14372 16992
rect 14424 16980 14430 16992
rect 15286 16980 15292 16992
rect 14424 16952 15292 16980
rect 14424 16940 14430 16952
rect 15286 16940 15292 16952
rect 15344 16940 15350 16992
rect 16022 16980 16028 16992
rect 15983 16952 16028 16980
rect 16022 16940 16028 16952
rect 16080 16940 16086 16992
rect 16500 16980 16528 17020
rect 17126 17008 17132 17020
rect 17184 17008 17190 17060
rect 17862 17008 17868 17060
rect 17920 17048 17926 17060
rect 19429 17051 19487 17057
rect 19429 17048 19441 17051
rect 17920 17020 19441 17048
rect 17920 17008 17926 17020
rect 19429 17017 19441 17020
rect 19475 17048 19487 17051
rect 19702 17048 19708 17060
rect 19475 17020 19708 17048
rect 19475 17017 19487 17020
rect 19429 17011 19487 17017
rect 19702 17008 19708 17020
rect 19760 17008 19766 17060
rect 20257 17051 20315 17057
rect 20257 17017 20269 17051
rect 20303 17048 20315 17051
rect 20346 17048 20352 17060
rect 20303 17020 20352 17048
rect 20303 17017 20315 17020
rect 20257 17011 20315 17017
rect 20346 17008 20352 17020
rect 20404 17048 20410 17060
rect 20404 17020 20944 17048
rect 20404 17008 20410 17020
rect 17586 16980 17592 16992
rect 16500 16952 17592 16980
rect 17586 16940 17592 16952
rect 17644 16940 17650 16992
rect 17681 16983 17739 16989
rect 17681 16949 17693 16983
rect 17727 16980 17739 16983
rect 17770 16980 17776 16992
rect 17727 16952 17776 16980
rect 17727 16949 17739 16952
rect 17681 16943 17739 16949
rect 17770 16940 17776 16952
rect 17828 16940 17834 16992
rect 18046 16980 18052 16992
rect 18007 16952 18052 16980
rect 18046 16940 18052 16952
rect 18104 16980 18110 16992
rect 18966 16980 18972 16992
rect 18104 16952 18972 16980
rect 18104 16940 18110 16952
rect 18966 16940 18972 16952
rect 19024 16940 19030 16992
rect 19242 16980 19248 16992
rect 19203 16952 19248 16980
rect 19242 16940 19248 16952
rect 19300 16940 19306 16992
rect 20916 16980 20944 17020
rect 22738 16980 22744 16992
rect 20916 16952 22744 16980
rect 22738 16940 22744 16952
rect 22796 16940 22802 16992
rect 1104 16890 23828 16912
rect 1104 16838 3790 16890
rect 3842 16838 3854 16890
rect 3906 16838 3918 16890
rect 3970 16838 3982 16890
rect 4034 16838 4046 16890
rect 4098 16838 9471 16890
rect 9523 16838 9535 16890
rect 9587 16838 9599 16890
rect 9651 16838 9663 16890
rect 9715 16838 9727 16890
rect 9779 16838 15152 16890
rect 15204 16838 15216 16890
rect 15268 16838 15280 16890
rect 15332 16838 15344 16890
rect 15396 16838 15408 16890
rect 15460 16838 20833 16890
rect 20885 16838 20897 16890
rect 20949 16838 20961 16890
rect 21013 16838 21025 16890
rect 21077 16838 21089 16890
rect 21141 16838 23828 16890
rect 1104 16816 23828 16838
rect 13262 16776 13268 16788
rect 12912 16748 13268 16776
rect 12912 16708 12940 16748
rect 13262 16736 13268 16748
rect 13320 16736 13326 16788
rect 14274 16736 14280 16788
rect 14332 16776 14338 16788
rect 14826 16776 14832 16788
rect 14332 16748 14832 16776
rect 14332 16736 14338 16748
rect 14826 16736 14832 16748
rect 14884 16736 14890 16788
rect 14918 16736 14924 16788
rect 14976 16776 14982 16788
rect 15473 16779 15531 16785
rect 15473 16776 15485 16779
rect 14976 16748 15485 16776
rect 14976 16736 14982 16748
rect 15473 16745 15485 16748
rect 15519 16745 15531 16779
rect 15473 16739 15531 16745
rect 17310 16736 17316 16788
rect 17368 16776 17374 16788
rect 18506 16776 18512 16788
rect 17368 16748 18512 16776
rect 17368 16736 17374 16748
rect 18506 16736 18512 16748
rect 18564 16736 18570 16788
rect 22005 16779 22063 16785
rect 22005 16745 22017 16779
rect 22051 16776 22063 16779
rect 22189 16779 22247 16785
rect 22051 16748 22141 16776
rect 22051 16745 22063 16748
rect 22005 16739 22063 16745
rect 12834 16680 12940 16708
rect 6641 16643 6699 16649
rect 6641 16609 6653 16643
rect 6687 16640 6699 16643
rect 7098 16640 7104 16652
rect 6687 16612 7104 16640
rect 6687 16609 6699 16612
rect 6641 16603 6699 16609
rect 7098 16600 7104 16612
rect 7156 16600 7162 16652
rect 8202 16600 8208 16652
rect 8260 16640 8266 16652
rect 9125 16643 9183 16649
rect 9125 16640 9137 16643
rect 8260 16612 9137 16640
rect 8260 16600 8266 16612
rect 9125 16609 9137 16612
rect 9171 16609 9183 16643
rect 9125 16603 9183 16609
rect 9401 16643 9459 16649
rect 9401 16609 9413 16643
rect 9447 16640 9459 16643
rect 11790 16640 11796 16652
rect 9447 16612 11796 16640
rect 9447 16609 9459 16612
rect 9401 16603 9459 16609
rect 11790 16600 11796 16612
rect 11848 16600 11854 16652
rect 12621 16643 12679 16649
rect 12621 16609 12633 16643
rect 12667 16640 12679 16643
rect 12710 16640 12716 16652
rect 12667 16612 12716 16640
rect 12667 16609 12679 16612
rect 12621 16603 12679 16609
rect 12710 16600 12716 16612
rect 12768 16600 12774 16652
rect 12834 16591 12862 16680
rect 14090 16668 14096 16720
rect 14148 16708 14154 16720
rect 14734 16708 14740 16720
rect 14148 16680 14740 16708
rect 14148 16668 14154 16680
rect 12819 16585 12877 16591
rect 2041 16575 2099 16581
rect 2041 16541 2053 16575
rect 2087 16572 2099 16575
rect 2682 16572 2688 16584
rect 2087 16544 2688 16572
rect 2087 16541 2099 16544
rect 2041 16535 2099 16541
rect 2682 16532 2688 16544
rect 2740 16572 2746 16584
rect 3050 16572 3056 16584
rect 2740 16544 3056 16572
rect 2740 16532 2746 16544
rect 3050 16532 3056 16544
rect 3108 16532 3114 16584
rect 7368 16575 7426 16581
rect 7368 16541 7380 16575
rect 7414 16572 7426 16575
rect 8386 16572 8392 16584
rect 7414 16544 8392 16572
rect 7414 16541 7426 16544
rect 7368 16535 7426 16541
rect 8386 16532 8392 16544
rect 8444 16532 8450 16584
rect 11882 16572 11888 16584
rect 11795 16544 11888 16572
rect 11882 16532 11888 16544
rect 11940 16532 11946 16584
rect 12069 16575 12127 16581
rect 12069 16541 12081 16575
rect 12115 16572 12127 16575
rect 12158 16572 12164 16584
rect 12115 16544 12164 16572
rect 12115 16541 12127 16544
rect 12069 16535 12127 16541
rect 12158 16532 12164 16544
rect 12216 16532 12222 16584
rect 12819 16551 12831 16585
rect 12865 16551 12877 16585
rect 12986 16581 12992 16584
rect 12819 16545 12877 16551
rect 12970 16575 12992 16581
rect 12970 16541 12982 16575
rect 12970 16535 12992 16541
rect 12986 16532 12992 16535
rect 13044 16532 13050 16584
rect 13078 16532 13084 16584
rect 13136 16581 13142 16584
rect 13136 16575 13151 16581
rect 13139 16541 13151 16575
rect 13136 16535 13151 16541
rect 13183 16575 13241 16581
rect 13183 16541 13195 16575
rect 13229 16572 13241 16575
rect 14182 16572 14188 16584
rect 13229 16544 14188 16572
rect 13229 16541 13241 16544
rect 13183 16535 13241 16541
rect 13136 16532 13142 16535
rect 14182 16532 14188 16544
rect 14240 16532 14246 16584
rect 14366 16572 14372 16584
rect 14327 16544 14372 16572
rect 14366 16532 14372 16544
rect 14424 16532 14430 16584
rect 14568 16581 14596 16680
rect 14734 16668 14740 16680
rect 14792 16668 14798 16720
rect 15013 16711 15071 16717
rect 15013 16677 15025 16711
rect 15059 16708 15071 16711
rect 15746 16708 15752 16720
rect 15059 16680 15752 16708
rect 15059 16677 15071 16680
rect 15013 16671 15071 16677
rect 15746 16668 15752 16680
rect 15804 16668 15810 16720
rect 16022 16708 16028 16720
rect 15856 16680 16028 16708
rect 14642 16600 14648 16652
rect 14700 16600 14706 16652
rect 15856 16640 15884 16680
rect 16022 16668 16028 16680
rect 16080 16668 16086 16720
rect 16298 16668 16304 16720
rect 16356 16708 16362 16720
rect 16485 16711 16543 16717
rect 16485 16708 16497 16711
rect 16356 16680 16497 16708
rect 16356 16668 16362 16680
rect 16485 16677 16497 16680
rect 16531 16677 16543 16711
rect 16485 16671 16543 16677
rect 17034 16668 17040 16720
rect 17092 16708 17098 16720
rect 19242 16708 19248 16720
rect 17092 16680 19248 16708
rect 17092 16668 17098 16680
rect 19242 16668 19248 16680
rect 19300 16668 19306 16720
rect 20165 16711 20223 16717
rect 20165 16677 20177 16711
rect 20211 16708 20223 16711
rect 20530 16708 20536 16720
rect 20211 16680 20536 16708
rect 20211 16677 20223 16680
rect 20165 16671 20223 16677
rect 20530 16668 20536 16680
rect 20588 16668 20594 16720
rect 22113 16708 22141 16748
rect 22189 16745 22201 16779
rect 22235 16776 22247 16779
rect 22370 16776 22376 16788
rect 22235 16748 22376 16776
rect 22235 16745 22247 16748
rect 22189 16739 22247 16745
rect 22370 16736 22376 16748
rect 22428 16736 22434 16788
rect 22278 16708 22284 16720
rect 22113 16680 22284 16708
rect 22278 16668 22284 16680
rect 22336 16668 22342 16720
rect 15488 16612 15884 16640
rect 15933 16643 15991 16649
rect 14517 16575 14596 16581
rect 14517 16541 14529 16575
rect 14563 16544 14596 16575
rect 14660 16572 14688 16600
rect 14834 16575 14892 16581
rect 14834 16572 14846 16575
rect 14660 16544 14846 16572
rect 14563 16541 14575 16544
rect 14517 16535 14575 16541
rect 14834 16541 14846 16544
rect 14880 16541 14892 16575
rect 15488 16572 15516 16612
rect 15933 16609 15945 16643
rect 15979 16640 15991 16643
rect 17129 16643 17187 16649
rect 17129 16640 17141 16643
rect 15979 16612 17141 16640
rect 15979 16609 15991 16612
rect 15933 16603 15991 16609
rect 17129 16609 17141 16612
rect 17175 16609 17187 16643
rect 17402 16640 17408 16652
rect 17129 16603 17187 16609
rect 17236 16612 17408 16640
rect 15654 16572 15660 16584
rect 14834 16535 14892 16541
rect 15304 16544 15516 16572
rect 15615 16544 15660 16572
rect 2308 16507 2366 16513
rect 2308 16473 2320 16507
rect 2354 16504 2366 16507
rect 2774 16504 2780 16516
rect 2354 16476 2780 16504
rect 2354 16473 2366 16476
rect 2308 16467 2366 16473
rect 2774 16464 2780 16476
rect 2832 16464 2838 16516
rect 6374 16507 6432 16513
rect 6374 16473 6386 16507
rect 6420 16473 6432 16507
rect 11900 16504 11928 16532
rect 14645 16507 14703 16513
rect 11900 16476 12572 16504
rect 6374 16467 6432 16473
rect 3421 16439 3479 16445
rect 3421 16405 3433 16439
rect 3467 16436 3479 16439
rect 4890 16436 4896 16448
rect 3467 16408 4896 16436
rect 3467 16405 3479 16408
rect 3421 16399 3479 16405
rect 4890 16396 4896 16408
rect 4948 16396 4954 16448
rect 5258 16436 5264 16448
rect 5219 16408 5264 16436
rect 5258 16396 5264 16408
rect 5316 16396 5322 16448
rect 6380 16436 6408 16467
rect 6454 16436 6460 16448
rect 6380 16408 6460 16436
rect 6454 16396 6460 16408
rect 6512 16396 6518 16448
rect 8478 16436 8484 16448
rect 8439 16408 8484 16436
rect 8478 16396 8484 16408
rect 8536 16396 8542 16448
rect 10686 16436 10692 16448
rect 10647 16408 10692 16436
rect 10686 16396 10692 16408
rect 10744 16396 10750 16448
rect 12066 16436 12072 16448
rect 12027 16408 12072 16436
rect 12066 16396 12072 16408
rect 12124 16396 12130 16448
rect 12544 16436 12572 16476
rect 14645 16473 14657 16507
rect 14691 16473 14703 16507
rect 14645 16467 14703 16473
rect 14737 16507 14795 16513
rect 14737 16473 14749 16507
rect 14783 16504 14795 16507
rect 15304 16504 15332 16544
rect 15654 16532 15660 16544
rect 15712 16532 15718 16584
rect 15749 16575 15807 16581
rect 15749 16541 15761 16575
rect 15795 16572 15807 16575
rect 15838 16572 15844 16584
rect 15795 16544 15844 16572
rect 15795 16541 15807 16544
rect 15749 16535 15807 16541
rect 15838 16532 15844 16544
rect 15896 16532 15902 16584
rect 16025 16575 16083 16581
rect 16025 16541 16037 16575
rect 16071 16572 16083 16575
rect 17034 16572 17040 16584
rect 16071 16544 17040 16572
rect 16071 16541 16083 16544
rect 16025 16535 16083 16541
rect 17034 16532 17040 16544
rect 17092 16572 17098 16584
rect 17236 16572 17264 16612
rect 17402 16600 17408 16612
rect 17460 16600 17466 16652
rect 17770 16640 17776 16652
rect 17731 16612 17776 16640
rect 17770 16600 17776 16612
rect 17828 16600 17834 16652
rect 18322 16600 18328 16652
rect 18380 16600 18386 16652
rect 18506 16600 18512 16652
rect 18564 16640 18570 16652
rect 20346 16640 20352 16652
rect 18564 16612 20116 16640
rect 20307 16612 20352 16640
rect 18564 16600 18570 16612
rect 17092 16544 17264 16572
rect 17313 16575 17371 16581
rect 17092 16532 17098 16544
rect 17313 16541 17325 16575
rect 17359 16572 17371 16575
rect 18340 16572 18368 16600
rect 20088 16581 20116 16612
rect 20346 16600 20352 16612
rect 20404 16600 20410 16652
rect 17359 16544 18368 16572
rect 20073 16575 20131 16581
rect 17359 16541 17371 16544
rect 17313 16535 17371 16541
rect 20073 16541 20085 16575
rect 20119 16541 20131 16575
rect 20073 16535 20131 16541
rect 20257 16575 20315 16581
rect 20257 16541 20269 16575
rect 20303 16541 20315 16575
rect 20257 16535 20315 16541
rect 16942 16504 16948 16516
rect 14783 16476 15332 16504
rect 15396 16476 16948 16504
rect 14783 16473 14795 16476
rect 14737 16467 14795 16473
rect 13725 16439 13783 16445
rect 13725 16436 13737 16439
rect 12544 16408 13737 16436
rect 13725 16405 13737 16408
rect 13771 16436 13783 16439
rect 14366 16436 14372 16448
rect 13771 16408 14372 16436
rect 13771 16405 13783 16408
rect 13725 16399 13783 16405
rect 14366 16396 14372 16408
rect 14424 16396 14430 16448
rect 14660 16436 14688 16467
rect 15396 16436 15424 16476
rect 16942 16464 16948 16476
rect 17000 16464 17006 16516
rect 17402 16504 17408 16516
rect 17363 16476 17408 16504
rect 17402 16464 17408 16476
rect 17460 16464 17466 16516
rect 17497 16507 17555 16513
rect 17497 16473 17509 16507
rect 17543 16473 17555 16507
rect 17497 16467 17555 16473
rect 17635 16507 17693 16513
rect 17635 16473 17647 16507
rect 17681 16504 17693 16507
rect 18322 16504 18328 16516
rect 17681 16476 18328 16504
rect 17681 16473 17693 16476
rect 17635 16467 17693 16473
rect 14660 16408 15424 16436
rect 16666 16396 16672 16448
rect 16724 16436 16730 16448
rect 17512 16436 17540 16467
rect 18322 16464 18328 16476
rect 18380 16464 18386 16516
rect 18782 16464 18788 16516
rect 18840 16504 18846 16516
rect 20272 16504 20300 16535
rect 20438 16532 20444 16584
rect 20496 16572 20502 16584
rect 20533 16575 20591 16581
rect 20533 16572 20545 16575
rect 20496 16544 20545 16572
rect 20496 16532 20502 16544
rect 20533 16541 20545 16544
rect 20579 16541 20591 16575
rect 20533 16535 20591 16541
rect 22373 16507 22431 16513
rect 22373 16504 22385 16507
rect 18840 16476 22385 16504
rect 18840 16464 18846 16476
rect 22373 16473 22385 16476
rect 22419 16504 22431 16507
rect 23290 16504 23296 16516
rect 22419 16476 23296 16504
rect 22419 16473 22431 16476
rect 22373 16467 22431 16473
rect 23290 16464 23296 16476
rect 23348 16464 23354 16516
rect 17862 16436 17868 16448
rect 16724 16408 17868 16436
rect 16724 16396 16730 16408
rect 17862 16396 17868 16408
rect 17920 16396 17926 16448
rect 18874 16436 18880 16448
rect 18835 16408 18880 16436
rect 18874 16396 18880 16408
rect 18932 16396 18938 16448
rect 19889 16439 19947 16445
rect 19889 16405 19901 16439
rect 19935 16436 19947 16439
rect 20162 16436 20168 16448
rect 19935 16408 20168 16436
rect 19935 16405 19947 16408
rect 19889 16399 19947 16405
rect 20162 16396 20168 16408
rect 20220 16396 20226 16448
rect 20990 16436 20996 16448
rect 20951 16408 20996 16436
rect 20990 16396 20996 16408
rect 21048 16396 21054 16448
rect 22173 16439 22231 16445
rect 22173 16405 22185 16439
rect 22219 16436 22231 16439
rect 22278 16436 22284 16448
rect 22219 16408 22284 16436
rect 22219 16405 22231 16408
rect 22173 16399 22231 16405
rect 22278 16396 22284 16408
rect 22336 16396 22342 16448
rect 1104 16346 23987 16368
rect 1104 16294 6630 16346
rect 6682 16294 6694 16346
rect 6746 16294 6758 16346
rect 6810 16294 6822 16346
rect 6874 16294 6886 16346
rect 6938 16294 12311 16346
rect 12363 16294 12375 16346
rect 12427 16294 12439 16346
rect 12491 16294 12503 16346
rect 12555 16294 12567 16346
rect 12619 16294 17992 16346
rect 18044 16294 18056 16346
rect 18108 16294 18120 16346
rect 18172 16294 18184 16346
rect 18236 16294 18248 16346
rect 18300 16294 23673 16346
rect 23725 16294 23737 16346
rect 23789 16294 23801 16346
rect 23853 16294 23865 16346
rect 23917 16294 23929 16346
rect 23981 16294 23987 16346
rect 1104 16272 23987 16294
rect 8202 16192 8208 16244
rect 8260 16232 8266 16244
rect 9125 16235 9183 16241
rect 9125 16232 9137 16235
rect 8260 16204 9137 16232
rect 8260 16192 8266 16204
rect 9125 16201 9137 16204
rect 9171 16201 9183 16235
rect 9125 16195 9183 16201
rect 9214 16192 9220 16244
rect 9272 16232 9278 16244
rect 14734 16232 14740 16244
rect 9272 16204 14740 16232
rect 9272 16192 9278 16204
rect 14734 16192 14740 16204
rect 14792 16192 14798 16244
rect 18322 16232 18328 16244
rect 18283 16204 18328 16232
rect 18322 16192 18328 16204
rect 18380 16192 18386 16244
rect 20254 16192 20260 16244
rect 20312 16232 20318 16244
rect 20441 16235 20499 16241
rect 20441 16232 20453 16235
rect 20312 16204 20453 16232
rect 20312 16192 20318 16204
rect 20441 16201 20453 16204
rect 20487 16201 20499 16235
rect 20990 16232 20996 16244
rect 20441 16195 20499 16201
rect 20729 16204 20996 16232
rect 4338 16164 4344 16176
rect 4299 16136 4344 16164
rect 4338 16124 4344 16136
rect 4396 16164 4402 16176
rect 7837 16167 7895 16173
rect 7837 16164 7849 16167
rect 4396 16136 7849 16164
rect 4396 16124 4402 16136
rect 7837 16133 7849 16136
rect 7883 16133 7895 16167
rect 17126 16164 17132 16176
rect 7837 16127 7895 16133
rect 11716 16136 13124 16164
rect 11716 16108 11744 16136
rect 11698 16096 11704 16108
rect 11659 16068 11704 16096
rect 11698 16056 11704 16068
rect 11756 16056 11762 16108
rect 11974 16096 11980 16108
rect 11935 16068 11980 16096
rect 11974 16056 11980 16068
rect 12032 16056 12038 16108
rect 13096 16105 13124 16136
rect 16868 16136 17132 16164
rect 12713 16099 12771 16105
rect 12713 16065 12725 16099
rect 12759 16065 12771 16099
rect 12713 16059 12771 16065
rect 13081 16099 13139 16105
rect 13081 16065 13093 16099
rect 13127 16065 13139 16099
rect 13081 16059 13139 16065
rect 11793 16031 11851 16037
rect 11793 15997 11805 16031
rect 11839 16028 11851 16031
rect 12158 16028 12164 16040
rect 11839 16000 12164 16028
rect 11839 15997 11851 16000
rect 11793 15991 11851 15997
rect 12158 15988 12164 16000
rect 12216 16028 12222 16040
rect 12728 16028 12756 16059
rect 12216 16000 12756 16028
rect 12216 15988 12222 16000
rect 14090 15988 14096 16040
rect 14148 16028 14154 16040
rect 14185 16031 14243 16037
rect 14185 16028 14197 16031
rect 14148 16000 14197 16028
rect 14148 15988 14154 16000
rect 14185 15997 14197 16000
rect 14231 16028 14243 16031
rect 16117 16031 16175 16037
rect 16117 16028 16129 16031
rect 14231 16000 16129 16028
rect 14231 15997 14243 16000
rect 14185 15991 14243 15997
rect 16117 15997 16129 16000
rect 16163 16028 16175 16031
rect 16482 16028 16488 16040
rect 16163 16000 16488 16028
rect 16163 15997 16175 16000
rect 16117 15991 16175 15997
rect 16482 15988 16488 16000
rect 16540 15988 16546 16040
rect 16868 16028 16896 16136
rect 17126 16124 17132 16136
rect 17184 16124 17190 16176
rect 20162 16124 20168 16176
rect 20220 16164 20226 16176
rect 20729 16164 20757 16204
rect 20990 16192 20996 16204
rect 21048 16192 21054 16244
rect 20220 16136 20757 16164
rect 20220 16124 20226 16136
rect 17037 16099 17095 16105
rect 17037 16065 17049 16099
rect 17083 16065 17095 16099
rect 17037 16059 17095 16065
rect 17313 16099 17371 16105
rect 17313 16065 17325 16099
rect 17359 16096 17371 16099
rect 18414 16096 18420 16108
rect 17359 16068 18420 16096
rect 17359 16065 17371 16068
rect 17313 16059 17371 16065
rect 16945 16031 17003 16037
rect 16945 16028 16957 16031
rect 16868 16000 16957 16028
rect 16945 15997 16957 16000
rect 16991 15997 17003 16031
rect 16945 15991 17003 15997
rect 17052 15972 17080 16059
rect 18414 16056 18420 16068
rect 18472 16056 18478 16108
rect 18693 16099 18751 16105
rect 18693 16065 18705 16099
rect 18739 16096 18751 16099
rect 19426 16096 19432 16108
rect 18739 16068 19432 16096
rect 18739 16065 18751 16068
rect 18693 16059 18751 16065
rect 19426 16056 19432 16068
rect 19484 16056 19490 16108
rect 19610 16096 19616 16108
rect 19571 16068 19616 16096
rect 19610 16056 19616 16068
rect 19668 16056 19674 16108
rect 19794 16096 19800 16108
rect 19755 16068 19800 16096
rect 19794 16056 19800 16068
rect 19852 16056 19858 16108
rect 20729 16105 20757 16136
rect 20806 16124 20812 16176
rect 20864 16164 20870 16176
rect 20864 16136 20909 16164
rect 20864 16124 20870 16136
rect 20625 16099 20683 16105
rect 20625 16065 20637 16099
rect 20671 16065 20683 16099
rect 20625 16059 20683 16065
rect 20717 16099 20775 16105
rect 20717 16065 20729 16099
rect 20763 16065 20775 16099
rect 20990 16096 20996 16108
rect 20951 16068 20996 16096
rect 20717 16059 20775 16065
rect 17221 16031 17279 16037
rect 17221 15997 17233 16031
rect 17267 16028 17279 16031
rect 17586 16028 17592 16040
rect 17267 16000 17592 16028
rect 17267 15997 17279 16000
rect 17221 15991 17279 15997
rect 17586 15988 17592 16000
rect 17644 15988 17650 16040
rect 18601 16031 18659 16037
rect 18601 15997 18613 16031
rect 18647 16028 18659 16031
rect 19150 16028 19156 16040
rect 18647 16000 19156 16028
rect 18647 15997 18659 16000
rect 18601 15991 18659 15997
rect 19150 15988 19156 16000
rect 19208 15988 19214 16040
rect 20640 16028 20668 16059
rect 20990 16056 20996 16068
rect 21048 16056 21054 16108
rect 21085 16099 21143 16105
rect 21085 16065 21097 16099
rect 21131 16096 21143 16099
rect 21818 16096 21824 16108
rect 21131 16068 21824 16096
rect 21131 16065 21143 16068
rect 21085 16059 21143 16065
rect 21818 16056 21824 16068
rect 21876 16056 21882 16108
rect 21910 16028 21916 16040
rect 20640 16000 21916 16028
rect 21910 15988 21916 16000
rect 21968 15988 21974 16040
rect 22097 16031 22155 16037
rect 22097 15997 22109 16031
rect 22143 16028 22155 16031
rect 22554 16028 22560 16040
rect 22143 16000 22560 16028
rect 22143 15997 22155 16000
rect 22097 15991 22155 15997
rect 22554 15988 22560 16000
rect 22612 15988 22618 16040
rect 2682 15920 2688 15972
rect 2740 15960 2746 15972
rect 3142 15960 3148 15972
rect 2740 15932 3148 15960
rect 2740 15920 2746 15932
rect 3142 15920 3148 15932
rect 3200 15920 3206 15972
rect 12066 15920 12072 15972
rect 12124 15960 12130 15972
rect 15562 15960 15568 15972
rect 12124 15932 15568 15960
rect 12124 15920 12130 15932
rect 15562 15920 15568 15932
rect 15620 15920 15626 15972
rect 17034 15920 17040 15972
rect 17092 15960 17098 15972
rect 17770 15960 17776 15972
rect 17092 15932 17776 15960
rect 17092 15920 17098 15932
rect 17770 15920 17776 15932
rect 17828 15920 17834 15972
rect 19889 15963 19947 15969
rect 19889 15929 19901 15963
rect 19935 15960 19947 15963
rect 21174 15960 21180 15972
rect 19935 15932 21180 15960
rect 19935 15929 19947 15932
rect 19889 15923 19947 15929
rect 21174 15920 21180 15932
rect 21232 15920 21238 15972
rect 3050 15892 3056 15904
rect 3011 15864 3056 15892
rect 3050 15852 3056 15864
rect 3108 15852 3114 15904
rect 12161 15895 12219 15901
rect 12161 15861 12173 15895
rect 12207 15892 12219 15895
rect 13078 15892 13084 15904
rect 12207 15864 13084 15892
rect 12207 15861 12219 15864
rect 12161 15855 12219 15861
rect 13078 15852 13084 15864
rect 13136 15852 13142 15904
rect 13906 15852 13912 15904
rect 13964 15892 13970 15904
rect 15013 15895 15071 15901
rect 15013 15892 15025 15895
rect 13964 15864 15025 15892
rect 13964 15852 13970 15864
rect 15013 15861 15025 15864
rect 15059 15861 15071 15895
rect 15654 15892 15660 15904
rect 15615 15864 15660 15892
rect 15013 15855 15071 15861
rect 15654 15852 15660 15864
rect 15712 15852 15718 15904
rect 17126 15892 17132 15904
rect 17087 15864 17132 15892
rect 17126 15852 17132 15864
rect 17184 15852 17190 15904
rect 18693 15895 18751 15901
rect 18693 15861 18705 15895
rect 18739 15892 18751 15895
rect 19702 15892 19708 15904
rect 18739 15864 19708 15892
rect 18739 15861 18751 15864
rect 18693 15855 18751 15861
rect 19702 15852 19708 15864
rect 19760 15852 19766 15904
rect 20990 15852 20996 15904
rect 21048 15892 21054 15904
rect 21266 15892 21272 15904
rect 21048 15864 21272 15892
rect 21048 15852 21054 15864
rect 21266 15852 21272 15864
rect 21324 15852 21330 15904
rect 22646 15892 22652 15904
rect 22607 15864 22652 15892
rect 22646 15852 22652 15864
rect 22704 15852 22710 15904
rect 1104 15802 23828 15824
rect 1104 15750 3790 15802
rect 3842 15750 3854 15802
rect 3906 15750 3918 15802
rect 3970 15750 3982 15802
rect 4034 15750 4046 15802
rect 4098 15750 9471 15802
rect 9523 15750 9535 15802
rect 9587 15750 9599 15802
rect 9651 15750 9663 15802
rect 9715 15750 9727 15802
rect 9779 15750 15152 15802
rect 15204 15750 15216 15802
rect 15268 15750 15280 15802
rect 15332 15750 15344 15802
rect 15396 15750 15408 15802
rect 15460 15750 20833 15802
rect 20885 15750 20897 15802
rect 20949 15750 20961 15802
rect 21013 15750 21025 15802
rect 21077 15750 21089 15802
rect 21141 15750 23828 15802
rect 1104 15728 23828 15750
rect 13262 15648 13268 15700
rect 13320 15688 13326 15700
rect 14277 15691 14335 15697
rect 14277 15688 14289 15691
rect 13320 15660 14289 15688
rect 13320 15648 13326 15660
rect 14277 15657 14289 15660
rect 14323 15657 14335 15691
rect 14277 15651 14335 15657
rect 15010 15648 15016 15700
rect 15068 15688 15074 15700
rect 15105 15691 15163 15697
rect 15105 15688 15117 15691
rect 15068 15660 15117 15688
rect 15068 15648 15074 15660
rect 15105 15657 15117 15660
rect 15151 15657 15163 15691
rect 19242 15688 19248 15700
rect 15105 15651 15163 15657
rect 15304 15660 19248 15688
rect 10686 15580 10692 15632
rect 10744 15620 10750 15632
rect 10744 15592 12434 15620
rect 10744 15580 10750 15592
rect 3050 15512 3056 15564
rect 3108 15552 3114 15564
rect 4985 15555 5043 15561
rect 4985 15552 4997 15555
rect 3108 15524 4997 15552
rect 3108 15512 3114 15524
rect 4985 15521 4997 15524
rect 5031 15521 5043 15555
rect 4985 15515 5043 15521
rect 8202 15512 8208 15564
rect 8260 15552 8266 15564
rect 9125 15555 9183 15561
rect 9125 15552 9137 15555
rect 8260 15524 9137 15552
rect 8260 15512 8266 15524
rect 9125 15521 9137 15524
rect 9171 15521 9183 15555
rect 9125 15515 9183 15521
rect 10134 15512 10140 15564
rect 10192 15552 10198 15564
rect 10192 15524 11376 15552
rect 10192 15512 10198 15524
rect 2225 15487 2283 15493
rect 2225 15453 2237 15487
rect 2271 15453 2283 15487
rect 2498 15484 2504 15496
rect 2459 15456 2504 15484
rect 2225 15447 2283 15453
rect 2240 15416 2268 15447
rect 2498 15444 2504 15456
rect 2556 15444 2562 15496
rect 3694 15444 3700 15496
rect 3752 15484 3758 15496
rect 3973 15487 4031 15493
rect 3973 15484 3985 15487
rect 3752 15456 3985 15484
rect 3752 15444 3758 15456
rect 3973 15453 3985 15456
rect 4019 15453 4031 15487
rect 11238 15484 11244 15496
rect 11199 15456 11244 15484
rect 3973 15447 4031 15453
rect 11238 15444 11244 15456
rect 11296 15444 11302 15496
rect 11348 15493 11376 15524
rect 11422 15512 11428 15564
rect 11480 15552 11486 15564
rect 11977 15555 12035 15561
rect 11977 15552 11989 15555
rect 11480 15524 11989 15552
rect 11480 15512 11486 15524
rect 11977 15521 11989 15524
rect 12023 15521 12035 15555
rect 12406 15552 12434 15592
rect 15010 15552 15016 15564
rect 12406 15524 15016 15552
rect 11977 15515 12035 15521
rect 15010 15512 15016 15524
rect 15068 15512 15074 15564
rect 15304 15561 15332 15660
rect 19242 15648 19248 15660
rect 19300 15648 19306 15700
rect 19610 15648 19616 15700
rect 19668 15688 19674 15700
rect 19981 15691 20039 15697
rect 19981 15688 19993 15691
rect 19668 15660 19993 15688
rect 19668 15648 19674 15660
rect 19981 15657 19993 15660
rect 20027 15688 20039 15691
rect 20346 15688 20352 15700
rect 20027 15660 20352 15688
rect 20027 15657 20039 15660
rect 19981 15651 20039 15657
rect 20346 15648 20352 15660
rect 20404 15648 20410 15700
rect 22002 15648 22008 15700
rect 22060 15688 22066 15700
rect 22097 15691 22155 15697
rect 22097 15688 22109 15691
rect 22060 15660 22109 15688
rect 22060 15648 22066 15660
rect 22097 15657 22109 15660
rect 22143 15657 22155 15691
rect 22738 15688 22744 15700
rect 22699 15660 22744 15688
rect 22097 15651 22155 15657
rect 22738 15648 22744 15660
rect 22796 15648 22802 15700
rect 16669 15623 16727 15629
rect 16669 15589 16681 15623
rect 16715 15589 16727 15623
rect 16669 15583 16727 15589
rect 15289 15555 15347 15561
rect 15289 15521 15301 15555
rect 15335 15521 15347 15555
rect 15289 15515 15347 15521
rect 15381 15555 15439 15561
rect 15381 15521 15393 15555
rect 15427 15552 15439 15555
rect 16684 15552 16712 15583
rect 16850 15580 16856 15632
rect 16908 15620 16914 15632
rect 18141 15623 18199 15629
rect 18141 15620 18153 15623
rect 16908 15592 18153 15620
rect 16908 15580 16914 15592
rect 18141 15589 18153 15592
rect 18187 15589 18199 15623
rect 18141 15583 18199 15589
rect 15427 15524 16712 15552
rect 15427 15521 15439 15524
rect 15381 15515 15439 15521
rect 11333 15487 11391 15493
rect 11333 15453 11345 15487
rect 11379 15453 11391 15487
rect 11333 15447 11391 15453
rect 11517 15487 11575 15493
rect 11517 15453 11529 15487
rect 11563 15484 11575 15487
rect 11790 15484 11796 15496
rect 11563 15456 11796 15484
rect 11563 15453 11575 15456
rect 11517 15447 11575 15453
rect 11790 15444 11796 15456
rect 11848 15444 11854 15496
rect 11882 15444 11888 15496
rect 11940 15484 11946 15496
rect 12529 15487 12587 15493
rect 12529 15484 12541 15487
rect 11940 15456 12541 15484
rect 11940 15444 11946 15456
rect 12529 15453 12541 15456
rect 12575 15453 12587 15487
rect 12529 15447 12587 15453
rect 13538 15444 13544 15496
rect 13596 15484 13602 15496
rect 13633 15487 13691 15493
rect 13633 15484 13645 15487
rect 13596 15456 13645 15484
rect 13596 15444 13602 15456
rect 13633 15453 13645 15456
rect 13679 15453 13691 15487
rect 13633 15447 13691 15453
rect 13906 15444 13912 15496
rect 13964 15484 13970 15496
rect 14277 15487 14335 15493
rect 14277 15484 14289 15487
rect 13964 15456 14289 15484
rect 13964 15444 13970 15456
rect 14277 15453 14289 15456
rect 14323 15453 14335 15487
rect 14277 15447 14335 15453
rect 14461 15487 14519 15493
rect 14461 15453 14473 15487
rect 14507 15484 14519 15487
rect 14734 15484 14740 15496
rect 14507 15456 14740 15484
rect 14507 15453 14519 15456
rect 14461 15447 14519 15453
rect 14734 15444 14740 15456
rect 14792 15444 14798 15496
rect 15194 15444 15200 15496
rect 15252 15484 15258 15496
rect 15473 15487 15531 15493
rect 15473 15484 15485 15487
rect 15252 15456 15485 15484
rect 15252 15444 15258 15456
rect 15473 15453 15485 15456
rect 15519 15453 15531 15487
rect 15473 15447 15531 15453
rect 15565 15487 15623 15493
rect 15565 15453 15577 15487
rect 15611 15484 15623 15487
rect 15654 15484 15660 15496
rect 15611 15456 15660 15484
rect 15611 15453 15623 15456
rect 15565 15447 15623 15453
rect 15654 15444 15660 15456
rect 15712 15484 15718 15496
rect 16206 15484 16212 15496
rect 15712 15456 16212 15484
rect 15712 15444 15718 15456
rect 16206 15444 16212 15456
rect 16264 15444 16270 15496
rect 16666 15484 16672 15496
rect 16627 15456 16672 15484
rect 16666 15444 16672 15456
rect 16724 15444 16730 15496
rect 18156 15484 18184 15583
rect 18966 15580 18972 15632
rect 19024 15620 19030 15632
rect 22554 15620 22560 15632
rect 19024 15592 22560 15620
rect 19024 15580 19030 15592
rect 22554 15580 22560 15592
rect 22612 15580 22618 15632
rect 18782 15512 18788 15564
rect 18840 15552 18846 15564
rect 19429 15555 19487 15561
rect 19429 15552 19441 15555
rect 18840 15524 19441 15552
rect 18840 15512 18846 15524
rect 19429 15521 19441 15524
rect 19475 15552 19487 15555
rect 19886 15552 19892 15564
rect 19475 15524 19892 15552
rect 19475 15521 19487 15524
rect 19429 15515 19487 15521
rect 19886 15512 19892 15524
rect 19944 15512 19950 15564
rect 18693 15487 18751 15493
rect 18693 15484 18705 15487
rect 18156 15456 18705 15484
rect 18693 15453 18705 15456
rect 18739 15453 18751 15487
rect 18693 15447 18751 15453
rect 18877 15487 18935 15493
rect 18877 15453 18889 15487
rect 18923 15484 18935 15487
rect 19518 15484 19524 15496
rect 18923 15456 19524 15484
rect 18923 15453 18935 15456
rect 18877 15447 18935 15453
rect 19518 15444 19524 15456
rect 19576 15444 19582 15496
rect 21085 15487 21143 15493
rect 21085 15453 21097 15487
rect 21131 15484 21143 15487
rect 21358 15484 21364 15496
rect 21131 15456 21364 15484
rect 21131 15453 21143 15456
rect 21085 15447 21143 15453
rect 21358 15444 21364 15456
rect 21416 15444 21422 15496
rect 22281 15487 22339 15493
rect 22281 15453 22293 15487
rect 22327 15484 22339 15487
rect 22646 15484 22652 15496
rect 22327 15456 22652 15484
rect 22327 15453 22339 15456
rect 22281 15447 22339 15453
rect 22646 15444 22652 15456
rect 22704 15484 22710 15496
rect 23014 15484 23020 15496
rect 22704 15456 23020 15484
rect 22704 15444 22710 15456
rect 23014 15444 23020 15456
rect 23072 15444 23078 15496
rect 2682 15416 2688 15428
rect 2240 15388 2688 15416
rect 2682 15376 2688 15388
rect 2740 15416 2746 15428
rect 2740 15388 3280 15416
rect 2740 15376 2746 15388
rect 2041 15351 2099 15357
rect 2041 15317 2053 15351
rect 2087 15348 2099 15351
rect 2222 15348 2228 15360
rect 2087 15320 2228 15348
rect 2087 15317 2099 15320
rect 2041 15311 2099 15317
rect 2222 15308 2228 15320
rect 2280 15308 2286 15360
rect 2409 15351 2467 15357
rect 2409 15317 2421 15351
rect 2455 15348 2467 15351
rect 3053 15351 3111 15357
rect 3053 15348 3065 15351
rect 2455 15320 3065 15348
rect 2455 15317 2467 15320
rect 2409 15311 2467 15317
rect 3053 15317 3065 15320
rect 3099 15348 3111 15351
rect 3142 15348 3148 15360
rect 3099 15320 3148 15348
rect 3099 15317 3111 15320
rect 3053 15311 3111 15317
rect 3142 15308 3148 15320
rect 3200 15308 3206 15360
rect 3252 15348 3280 15388
rect 3326 15376 3332 15428
rect 3384 15416 3390 15428
rect 4246 15416 4252 15428
rect 3384 15388 3429 15416
rect 4207 15388 4252 15416
rect 3384 15376 3390 15388
rect 4246 15376 4252 15388
rect 4304 15376 4310 15428
rect 5252 15419 5310 15425
rect 5252 15385 5264 15419
rect 5298 15416 5310 15419
rect 6546 15416 6552 15428
rect 5298 15388 6552 15416
rect 5298 15385 5310 15388
rect 5252 15379 5310 15385
rect 6546 15376 6552 15388
rect 6604 15376 6610 15428
rect 9392 15419 9450 15425
rect 9392 15385 9404 15419
rect 9438 15416 9450 15419
rect 12894 15416 12900 15428
rect 9438 15388 11468 15416
rect 12855 15388 12900 15416
rect 9438 15385 9450 15388
rect 9392 15379 9450 15385
rect 4522 15348 4528 15360
rect 3252 15320 4528 15348
rect 4522 15308 4528 15320
rect 4580 15308 4586 15360
rect 6365 15351 6423 15357
rect 6365 15317 6377 15351
rect 6411 15348 6423 15351
rect 7926 15348 7932 15360
rect 6411 15320 7932 15348
rect 6411 15317 6423 15320
rect 6365 15311 6423 15317
rect 7926 15308 7932 15320
rect 7984 15308 7990 15360
rect 10505 15351 10563 15357
rect 10505 15317 10517 15351
rect 10551 15348 10563 15351
rect 11146 15348 11152 15360
rect 10551 15320 11152 15348
rect 10551 15317 10563 15320
rect 10505 15311 10563 15317
rect 11146 15308 11152 15320
rect 11204 15308 11210 15360
rect 11440 15348 11468 15388
rect 12894 15376 12900 15388
rect 12952 15376 12958 15428
rect 16574 15416 16580 15428
rect 13556 15388 16580 15416
rect 13556 15348 13584 15388
rect 16574 15376 16580 15388
rect 16632 15376 16638 15428
rect 16761 15419 16819 15425
rect 16761 15385 16773 15419
rect 16807 15385 16819 15419
rect 16761 15379 16819 15385
rect 16945 15419 17003 15425
rect 16945 15385 16957 15419
rect 16991 15416 17003 15419
rect 17402 15416 17408 15428
rect 16991 15388 17408 15416
rect 16991 15385 17003 15388
rect 16945 15379 17003 15385
rect 11440 15320 13584 15348
rect 14734 15308 14740 15360
rect 14792 15348 14798 15360
rect 16114 15348 16120 15360
rect 14792 15320 16120 15348
rect 14792 15308 14798 15320
rect 16114 15308 16120 15320
rect 16172 15348 16178 15360
rect 16209 15351 16267 15357
rect 16209 15348 16221 15351
rect 16172 15320 16221 15348
rect 16172 15308 16178 15320
rect 16209 15317 16221 15320
rect 16255 15348 16267 15351
rect 16390 15348 16396 15360
rect 16255 15320 16396 15348
rect 16255 15317 16267 15320
rect 16209 15311 16267 15317
rect 16390 15308 16396 15320
rect 16448 15308 16454 15360
rect 16482 15308 16488 15360
rect 16540 15348 16546 15360
rect 16776 15348 16804 15379
rect 17402 15376 17408 15388
rect 17460 15416 17466 15428
rect 18785 15419 18843 15425
rect 18785 15416 18797 15419
rect 17460 15388 18797 15416
rect 17460 15376 17466 15388
rect 18785 15385 18797 15388
rect 18831 15385 18843 15419
rect 18785 15379 18843 15385
rect 19058 15376 19064 15428
rect 19116 15416 19122 15428
rect 19794 15416 19800 15428
rect 19116 15388 19800 15416
rect 19116 15376 19122 15388
rect 19794 15376 19800 15388
rect 19852 15376 19858 15428
rect 20806 15416 20812 15428
rect 20767 15388 20812 15416
rect 20806 15376 20812 15388
rect 20864 15376 20870 15428
rect 16540 15320 16804 15348
rect 16540 15308 16546 15320
rect 1104 15258 23987 15280
rect 1104 15206 6630 15258
rect 6682 15206 6694 15258
rect 6746 15206 6758 15258
rect 6810 15206 6822 15258
rect 6874 15206 6886 15258
rect 6938 15206 12311 15258
rect 12363 15206 12375 15258
rect 12427 15206 12439 15258
rect 12491 15206 12503 15258
rect 12555 15206 12567 15258
rect 12619 15206 17992 15258
rect 18044 15206 18056 15258
rect 18108 15206 18120 15258
rect 18172 15206 18184 15258
rect 18236 15206 18248 15258
rect 18300 15206 23673 15258
rect 23725 15206 23737 15258
rect 23789 15206 23801 15258
rect 23853 15206 23865 15258
rect 23917 15206 23929 15258
rect 23981 15206 23987 15258
rect 1104 15184 23987 15206
rect 3234 15144 3240 15156
rect 1596 15116 3240 15144
rect 1596 15017 1624 15116
rect 3234 15104 3240 15116
rect 3292 15104 3298 15156
rect 3418 15104 3424 15156
rect 3476 15144 3482 15156
rect 4801 15147 4859 15153
rect 4801 15144 4813 15147
rect 3476 15116 4813 15144
rect 3476 15104 3482 15116
rect 4801 15113 4813 15116
rect 4847 15113 4859 15147
rect 4801 15107 4859 15113
rect 6270 15104 6276 15156
rect 6328 15144 6334 15156
rect 11701 15147 11759 15153
rect 6328 15116 6868 15144
rect 6328 15104 6334 15116
rect 1854 15076 1860 15088
rect 1767 15048 1860 15076
rect 1854 15036 1860 15048
rect 1912 15076 1918 15088
rect 2130 15076 2136 15088
rect 1912 15048 2136 15076
rect 1912 15036 1918 15048
rect 2130 15036 2136 15048
rect 2188 15036 2194 15088
rect 4154 15036 4160 15088
rect 4212 15076 4218 15088
rect 5169 15079 5227 15085
rect 5169 15076 5181 15079
rect 4212 15048 5181 15076
rect 4212 15036 4218 15048
rect 5169 15045 5181 15048
rect 5215 15045 5227 15079
rect 5169 15039 5227 15045
rect 5258 15036 5264 15088
rect 5316 15076 5322 15088
rect 6549 15079 6607 15085
rect 6549 15076 6561 15079
rect 5316 15048 6561 15076
rect 5316 15036 5322 15048
rect 6549 15045 6561 15048
rect 6595 15045 6607 15079
rect 6549 15039 6607 15045
rect 1581 15011 1639 15017
rect 1581 14977 1593 15011
rect 1627 14977 1639 15011
rect 1762 15008 1768 15020
rect 1723 14980 1768 15008
rect 1581 14971 1639 14977
rect 1762 14968 1768 14980
rect 1820 14968 1826 15020
rect 1949 15011 2007 15017
rect 1949 14977 1961 15011
rect 1995 15008 2007 15011
rect 2314 15008 2320 15020
rect 1995 14980 2320 15008
rect 1995 14977 2007 14980
rect 1949 14971 2007 14977
rect 2314 14968 2320 14980
rect 2372 14968 2378 15020
rect 3050 15008 3056 15020
rect 2884 14980 3056 15008
rect 2685 14943 2743 14949
rect 2685 14909 2697 14943
rect 2731 14940 2743 14943
rect 2884 14940 2912 14980
rect 3050 14968 3056 14980
rect 3108 14968 3114 15020
rect 4982 15008 4988 15020
rect 4943 14980 4988 15008
rect 4982 14968 4988 14980
rect 5040 14968 5046 15020
rect 5077 15011 5135 15017
rect 5077 14977 5089 15011
rect 5123 14977 5135 15011
rect 5077 14971 5135 14977
rect 5353 15011 5411 15017
rect 5353 14977 5365 15011
rect 5399 14977 5411 15011
rect 5353 14971 5411 14977
rect 2731 14912 2912 14940
rect 2961 14943 3019 14949
rect 2731 14909 2743 14912
rect 2685 14903 2743 14909
rect 2961 14909 2973 14943
rect 3007 14940 3019 14943
rect 4614 14940 4620 14952
rect 3007 14912 4620 14940
rect 3007 14909 3019 14912
rect 2961 14903 3019 14909
rect 4614 14900 4620 14912
rect 4672 14900 4678 14952
rect 4982 14832 4988 14884
rect 5040 14872 5046 14884
rect 5092 14872 5120 14971
rect 5368 14940 5396 14971
rect 5626 14968 5632 15020
rect 5684 15008 5690 15020
rect 6840 15017 6868 15116
rect 11701 15113 11713 15147
rect 11747 15144 11759 15147
rect 11882 15144 11888 15156
rect 11747 15116 11888 15144
rect 11747 15113 11759 15116
rect 11701 15107 11759 15113
rect 11882 15104 11888 15116
rect 11940 15104 11946 15156
rect 15470 15104 15476 15156
rect 15528 15144 15534 15156
rect 16482 15144 16488 15156
rect 15528 15116 16488 15144
rect 15528 15104 15534 15116
rect 16482 15104 16488 15116
rect 16540 15104 16546 15156
rect 19242 15104 19248 15156
rect 19300 15144 19306 15156
rect 20349 15147 20407 15153
rect 20349 15144 20361 15147
rect 19300 15116 20361 15144
rect 19300 15104 19306 15116
rect 20349 15113 20361 15116
rect 20395 15113 20407 15147
rect 20349 15107 20407 15113
rect 22462 15104 22468 15156
rect 22520 15144 22526 15156
rect 22649 15147 22707 15153
rect 22649 15144 22661 15147
rect 22520 15116 22661 15144
rect 22520 15104 22526 15116
rect 22649 15113 22661 15116
rect 22695 15113 22707 15147
rect 22649 15107 22707 15113
rect 11790 15036 11796 15088
rect 11848 15076 11854 15088
rect 12894 15076 12900 15088
rect 11848 15048 12900 15076
rect 11848 15036 11854 15048
rect 12894 15036 12900 15048
rect 12952 15036 12958 15088
rect 18506 15076 18512 15088
rect 13832 15048 18512 15076
rect 5997 15011 6055 15017
rect 5997 15008 6009 15011
rect 5684 14980 6009 15008
rect 5684 14968 5690 14980
rect 5997 14977 6009 14980
rect 6043 15008 6055 15011
rect 6733 15011 6791 15017
rect 6733 15008 6745 15011
rect 6043 14980 6745 15008
rect 6043 14977 6055 14980
rect 5997 14971 6055 14977
rect 6733 14977 6745 14980
rect 6779 14977 6791 15011
rect 6733 14971 6791 14977
rect 6825 15011 6883 15017
rect 6825 14977 6837 15011
rect 6871 14977 6883 15011
rect 6825 14971 6883 14977
rect 8202 14968 8208 15020
rect 8260 15008 8266 15020
rect 9677 15011 9735 15017
rect 9677 15008 9689 15011
rect 8260 14980 9689 15008
rect 8260 14968 8266 14980
rect 9677 14977 9689 14980
rect 9723 14977 9735 15011
rect 9677 14971 9735 14977
rect 12529 15011 12587 15017
rect 12529 14977 12541 15011
rect 12575 15008 12587 15011
rect 12618 15008 12624 15020
rect 12575 14980 12624 15008
rect 12575 14977 12587 14980
rect 12529 14971 12587 14977
rect 12618 14968 12624 14980
rect 12676 14968 12682 15020
rect 13078 15008 13084 15020
rect 13039 14980 13084 15008
rect 13078 14968 13084 14980
rect 13136 14968 13142 15020
rect 13262 15008 13268 15020
rect 13223 14980 13268 15008
rect 13262 14968 13268 14980
rect 13320 14968 13326 15020
rect 13832 15017 13860 15048
rect 18506 15036 18512 15048
rect 18564 15036 18570 15088
rect 19334 15076 19340 15088
rect 19295 15048 19340 15076
rect 19334 15036 19340 15048
rect 19392 15036 19398 15088
rect 13357 15011 13415 15017
rect 13357 14977 13369 15011
rect 13403 15008 13415 15011
rect 13817 15011 13875 15017
rect 13817 15008 13829 15011
rect 13403 14980 13829 15008
rect 13403 14977 13415 14980
rect 13357 14971 13415 14977
rect 13817 14977 13829 14980
rect 13863 14977 13875 15011
rect 13817 14971 13875 14977
rect 14737 15011 14795 15017
rect 14737 14977 14749 15011
rect 14783 15008 14795 15011
rect 14918 15008 14924 15020
rect 14783 14980 14924 15008
rect 14783 14977 14795 14980
rect 14737 14971 14795 14977
rect 14918 14968 14924 14980
rect 14976 14968 14982 15020
rect 15562 15008 15568 15020
rect 15523 14980 15568 15008
rect 15562 14968 15568 14980
rect 15620 14968 15626 15020
rect 15841 15011 15899 15017
rect 15841 14977 15853 15011
rect 15887 15008 15899 15011
rect 16942 15008 16948 15020
rect 15887 14980 16948 15008
rect 15887 14977 15899 14980
rect 15841 14971 15899 14977
rect 7834 14940 7840 14952
rect 5368 14912 7840 14940
rect 7834 14900 7840 14912
rect 7892 14900 7898 14952
rect 9401 14943 9459 14949
rect 9401 14909 9413 14943
rect 9447 14940 9459 14943
rect 10229 14943 10287 14949
rect 10229 14940 10241 14943
rect 9447 14912 10241 14940
rect 9447 14909 9459 14912
rect 9401 14903 9459 14909
rect 10229 14909 10241 14912
rect 10275 14940 10287 14943
rect 12894 14940 12900 14952
rect 10275 14912 12900 14940
rect 10275 14909 10287 14912
rect 10229 14903 10287 14909
rect 12894 14900 12900 14912
rect 12952 14900 12958 14952
rect 14093 14943 14151 14949
rect 14093 14909 14105 14943
rect 14139 14940 14151 14943
rect 14182 14940 14188 14952
rect 14139 14912 14188 14940
rect 14139 14909 14151 14912
rect 14093 14903 14151 14909
rect 14182 14900 14188 14912
rect 14240 14900 14246 14952
rect 15013 14943 15071 14949
rect 15013 14940 15025 14943
rect 14292 14912 15025 14940
rect 5040 14844 5120 14872
rect 5040 14832 5046 14844
rect 6178 14832 6184 14884
rect 6236 14872 6242 14884
rect 6638 14872 6644 14884
rect 6236 14844 6644 14872
rect 6236 14832 6242 14844
rect 6638 14832 6644 14844
rect 6696 14832 6702 14884
rect 11149 14875 11207 14881
rect 11149 14841 11161 14875
rect 11195 14872 11207 14875
rect 11790 14872 11796 14884
rect 11195 14844 11796 14872
rect 11195 14841 11207 14844
rect 11149 14835 11207 14841
rect 11790 14832 11796 14844
rect 11848 14832 11854 14884
rect 13538 14832 13544 14884
rect 13596 14872 13602 14884
rect 14292 14872 14320 14912
rect 15013 14909 15025 14912
rect 15059 14909 15071 14943
rect 15013 14903 15071 14909
rect 14826 14872 14832 14884
rect 13596 14844 14320 14872
rect 14787 14844 14832 14872
rect 13596 14832 13602 14844
rect 14826 14832 14832 14844
rect 14884 14832 14890 14884
rect 15028 14872 15056 14903
rect 15194 14900 15200 14952
rect 15252 14940 15258 14952
rect 15856 14940 15884 14971
rect 16942 14968 16948 14980
rect 17000 14968 17006 15020
rect 19242 14968 19248 15020
rect 19300 15008 19306 15020
rect 19513 15011 19571 15017
rect 19513 15008 19525 15011
rect 19300 14980 19525 15008
rect 19300 14968 19306 14980
rect 19513 14977 19525 14980
rect 19559 14977 19571 15011
rect 19513 14971 19571 14977
rect 19613 15011 19671 15017
rect 19613 14977 19625 15011
rect 19659 14977 19671 15011
rect 19794 15008 19800 15020
rect 19755 14980 19800 15008
rect 19613 14971 19671 14977
rect 15252 14912 15884 14940
rect 15252 14900 15258 14912
rect 16574 14900 16580 14952
rect 16632 14940 16638 14952
rect 17310 14940 17316 14952
rect 16632 14912 17316 14940
rect 16632 14900 16638 14912
rect 17310 14900 17316 14912
rect 17368 14940 17374 14952
rect 18322 14940 18328 14952
rect 17368 14912 18328 14940
rect 17368 14900 17374 14912
rect 18322 14900 18328 14912
rect 18380 14900 18386 14952
rect 18877 14943 18935 14949
rect 18877 14909 18889 14943
rect 18923 14940 18935 14943
rect 18923 14912 19334 14940
rect 18923 14909 18935 14912
rect 18877 14903 18935 14909
rect 16298 14872 16304 14884
rect 15028 14844 16304 14872
rect 16298 14832 16304 14844
rect 16356 14872 16362 14884
rect 18892 14872 18920 14903
rect 16356 14844 18920 14872
rect 16356 14832 16362 14844
rect 2133 14807 2191 14813
rect 2133 14773 2145 14807
rect 2179 14804 2191 14807
rect 2866 14804 2872 14816
rect 2179 14776 2872 14804
rect 2179 14773 2191 14776
rect 2133 14767 2191 14773
rect 2866 14764 2872 14776
rect 2924 14764 2930 14816
rect 3142 14764 3148 14816
rect 3200 14804 3206 14816
rect 3418 14804 3424 14816
rect 3200 14776 3424 14804
rect 3200 14764 3206 14776
rect 3418 14764 3424 14776
rect 3476 14764 3482 14816
rect 4249 14807 4307 14813
rect 4249 14773 4261 14807
rect 4295 14804 4307 14807
rect 5994 14804 6000 14816
rect 4295 14776 6000 14804
rect 4295 14773 4307 14776
rect 4249 14767 4307 14773
rect 5994 14764 6000 14776
rect 6052 14764 6058 14816
rect 6086 14764 6092 14816
rect 6144 14804 6150 14816
rect 6549 14807 6607 14813
rect 6549 14804 6561 14807
rect 6144 14776 6561 14804
rect 6144 14764 6150 14776
rect 6549 14773 6561 14776
rect 6595 14773 6607 14807
rect 6549 14767 6607 14773
rect 7650 14764 7656 14816
rect 7708 14804 7714 14816
rect 8113 14807 8171 14813
rect 8113 14804 8125 14807
rect 7708 14776 8125 14804
rect 7708 14764 7714 14776
rect 8113 14773 8125 14776
rect 8159 14773 8171 14807
rect 8113 14767 8171 14773
rect 13354 14764 13360 14816
rect 13412 14804 13418 14816
rect 14737 14807 14795 14813
rect 14737 14804 14749 14807
rect 13412 14776 14749 14804
rect 13412 14764 13418 14776
rect 14737 14773 14749 14776
rect 14783 14773 14795 14807
rect 14737 14767 14795 14773
rect 16206 14764 16212 14816
rect 16264 14804 16270 14816
rect 16853 14807 16911 14813
rect 16853 14804 16865 14807
rect 16264 14776 16865 14804
rect 16264 14764 16270 14776
rect 16853 14773 16865 14776
rect 16899 14804 16911 14807
rect 18782 14804 18788 14816
rect 16899 14776 18788 14804
rect 16899 14773 16911 14776
rect 16853 14767 16911 14773
rect 18782 14764 18788 14776
rect 18840 14764 18846 14816
rect 19306 14804 19334 14912
rect 19628 14804 19656 14971
rect 19794 14968 19800 14980
rect 19852 14968 19858 15020
rect 19886 14968 19892 15020
rect 19944 15008 19950 15020
rect 19944 14980 19989 15008
rect 19944 14968 19950 14980
rect 20254 14968 20260 15020
rect 20312 15008 20318 15020
rect 20901 15011 20959 15017
rect 20901 15008 20913 15011
rect 20312 14980 20913 15008
rect 20312 14968 20318 14980
rect 20901 14977 20913 14980
rect 20947 14977 20959 15011
rect 20901 14971 20959 14977
rect 21085 15011 21143 15017
rect 21085 14977 21097 15011
rect 21131 15008 21143 15011
rect 21174 15008 21180 15020
rect 21131 14980 21180 15008
rect 21131 14977 21143 14980
rect 21085 14971 21143 14977
rect 21174 14968 21180 14980
rect 21232 14968 21238 15020
rect 22002 15008 22008 15020
rect 21963 14980 22008 15008
rect 22002 14968 22008 14980
rect 22060 14968 22066 15020
rect 22094 14968 22100 15020
rect 22152 15008 22158 15020
rect 22278 15008 22284 15020
rect 22152 14980 22197 15008
rect 22239 14980 22284 15008
rect 22152 14968 22158 14980
rect 22278 14968 22284 14980
rect 22336 14968 22342 15020
rect 22373 15011 22431 15017
rect 22373 14977 22385 15011
rect 22419 14977 22431 15011
rect 22373 14971 22431 14977
rect 22511 15011 22569 15017
rect 22511 14977 22523 15011
rect 22557 15008 22569 15011
rect 22830 15008 22836 15020
rect 22557 14980 22836 15008
rect 22557 14977 22569 14980
rect 22511 14971 22569 14977
rect 20625 14943 20683 14949
rect 20625 14909 20637 14943
rect 20671 14940 20683 14943
rect 20806 14940 20812 14952
rect 20671 14912 20812 14940
rect 20671 14909 20683 14912
rect 20625 14903 20683 14909
rect 20806 14900 20812 14912
rect 20864 14940 20870 14952
rect 22020 14940 22048 14968
rect 20864 14912 22048 14940
rect 20864 14900 20870 14912
rect 20717 14875 20775 14881
rect 20717 14841 20729 14875
rect 20763 14872 20775 14875
rect 21358 14872 21364 14884
rect 20763 14844 21364 14872
rect 20763 14841 20775 14844
rect 20717 14835 20775 14841
rect 21358 14832 21364 14844
rect 21416 14832 21422 14884
rect 22278 14832 22284 14884
rect 22336 14872 22342 14884
rect 22388 14872 22416 14971
rect 22830 14968 22836 14980
rect 22888 14968 22894 15020
rect 22336 14844 22416 14872
rect 22336 14832 22342 14844
rect 19306 14776 19656 14804
rect 20809 14807 20867 14813
rect 20809 14773 20821 14807
rect 20855 14804 20867 14807
rect 21818 14804 21824 14816
rect 20855 14776 21824 14804
rect 20855 14773 20867 14776
rect 20809 14767 20867 14773
rect 21818 14764 21824 14776
rect 21876 14764 21882 14816
rect 23106 14804 23112 14816
rect 23067 14776 23112 14804
rect 23106 14764 23112 14776
rect 23164 14764 23170 14816
rect 1104 14714 23828 14736
rect 1104 14662 3790 14714
rect 3842 14662 3854 14714
rect 3906 14662 3918 14714
rect 3970 14662 3982 14714
rect 4034 14662 4046 14714
rect 4098 14662 9471 14714
rect 9523 14662 9535 14714
rect 9587 14662 9599 14714
rect 9651 14662 9663 14714
rect 9715 14662 9727 14714
rect 9779 14662 15152 14714
rect 15204 14662 15216 14714
rect 15268 14662 15280 14714
rect 15332 14662 15344 14714
rect 15396 14662 15408 14714
rect 15460 14662 20833 14714
rect 20885 14662 20897 14714
rect 20949 14662 20961 14714
rect 21013 14662 21025 14714
rect 21077 14662 21089 14714
rect 21141 14662 23828 14714
rect 1104 14640 23828 14662
rect 1670 14560 1676 14612
rect 1728 14600 1734 14612
rect 2041 14603 2099 14609
rect 2041 14600 2053 14603
rect 1728 14572 2053 14600
rect 1728 14560 1734 14572
rect 2041 14569 2053 14572
rect 2087 14569 2099 14603
rect 4706 14600 4712 14612
rect 2041 14563 2099 14569
rect 3068 14572 4384 14600
rect 4667 14572 4712 14600
rect 3068 14532 3096 14572
rect 4246 14532 4252 14544
rect 2424 14504 3096 14532
rect 3160 14504 4252 14532
rect 2424 14473 2452 14504
rect 2409 14467 2467 14473
rect 2409 14433 2421 14467
rect 2455 14433 2467 14467
rect 2409 14427 2467 14433
rect 2222 14396 2228 14408
rect 2183 14368 2228 14396
rect 2222 14356 2228 14368
rect 2280 14356 2286 14408
rect 2314 14356 2320 14408
rect 2372 14396 2378 14408
rect 2682 14396 2688 14408
rect 2372 14368 2688 14396
rect 2372 14356 2378 14368
rect 2682 14356 2688 14368
rect 2740 14396 2746 14408
rect 3160 14405 3188 14504
rect 4246 14492 4252 14504
rect 4304 14492 4310 14544
rect 3234 14424 3240 14476
rect 3292 14464 3298 14476
rect 3510 14464 3516 14476
rect 3292 14436 3516 14464
rect 3292 14424 3298 14436
rect 3510 14424 3516 14436
rect 3568 14464 3574 14476
rect 4157 14467 4215 14473
rect 4157 14464 4169 14467
rect 3568 14436 4169 14464
rect 3568 14424 3574 14436
rect 4157 14433 4169 14436
rect 4203 14433 4215 14467
rect 4356 14464 4384 14572
rect 4706 14560 4712 14572
rect 4764 14560 4770 14612
rect 5813 14603 5871 14609
rect 5813 14569 5825 14603
rect 5859 14569 5871 14603
rect 5813 14563 5871 14569
rect 4614 14492 4620 14544
rect 4672 14532 4678 14544
rect 5828 14532 5856 14563
rect 6546 14560 6552 14612
rect 6604 14600 6610 14612
rect 6825 14603 6883 14609
rect 6825 14600 6837 14603
rect 6604 14572 6837 14600
rect 6604 14560 6610 14572
rect 6825 14569 6837 14572
rect 6871 14569 6883 14603
rect 6825 14563 6883 14569
rect 8294 14560 8300 14612
rect 8352 14600 8358 14612
rect 9125 14603 9183 14609
rect 9125 14600 9137 14603
rect 8352 14572 9137 14600
rect 8352 14560 8358 14572
rect 9125 14569 9137 14572
rect 9171 14569 9183 14603
rect 9125 14563 9183 14569
rect 12621 14603 12679 14609
rect 12621 14569 12633 14603
rect 12667 14600 12679 14603
rect 12802 14600 12808 14612
rect 12667 14572 12808 14600
rect 12667 14569 12679 14572
rect 12621 14563 12679 14569
rect 12802 14560 12808 14572
rect 12860 14560 12866 14612
rect 13814 14560 13820 14612
rect 13872 14600 13878 14612
rect 13872 14572 14872 14600
rect 13872 14560 13878 14572
rect 4672 14504 5856 14532
rect 4672 14492 4678 14504
rect 5994 14492 6000 14544
rect 6052 14532 6058 14544
rect 6052 14504 6408 14532
rect 6052 14492 6058 14504
rect 6086 14464 6092 14476
rect 4157 14427 4215 14433
rect 4264 14436 6092 14464
rect 4264 14405 4292 14436
rect 6086 14424 6092 14436
rect 6144 14424 6150 14476
rect 6380 14464 6408 14504
rect 7190 14492 7196 14544
rect 7248 14532 7254 14544
rect 9306 14532 9312 14544
rect 7248 14504 9312 14532
rect 7248 14492 7254 14504
rect 9306 14492 9312 14504
rect 9364 14492 9370 14544
rect 10502 14492 10508 14544
rect 10560 14532 10566 14544
rect 10689 14535 10747 14541
rect 10689 14532 10701 14535
rect 10560 14504 10701 14532
rect 10560 14492 10566 14504
rect 10689 14501 10701 14504
rect 10735 14501 10747 14535
rect 11882 14532 11888 14544
rect 10689 14495 10747 14501
rect 10796 14504 11888 14532
rect 7282 14464 7288 14476
rect 6380 14436 7288 14464
rect 3053 14399 3111 14405
rect 3053 14396 3065 14399
rect 2740 14368 3065 14396
rect 2740 14356 2746 14368
rect 3053 14365 3065 14368
rect 3099 14365 3111 14399
rect 3053 14359 3111 14365
rect 3145 14399 3203 14405
rect 3145 14365 3157 14399
rect 3191 14365 3203 14399
rect 3145 14359 3203 14365
rect 3421 14399 3479 14405
rect 3421 14365 3433 14399
rect 3467 14365 3479 14399
rect 3421 14359 3479 14365
rect 4249 14399 4307 14405
rect 4249 14365 4261 14399
rect 4295 14365 4307 14399
rect 4249 14359 4307 14365
rect 4341 14399 4399 14405
rect 4341 14365 4353 14399
rect 4387 14396 4399 14399
rect 4614 14396 4620 14408
rect 4387 14368 4620 14396
rect 4387 14365 4399 14368
rect 4341 14359 4399 14365
rect 1946 14288 1952 14340
rect 2004 14328 2010 14340
rect 3160 14328 3188 14359
rect 2004 14300 3188 14328
rect 2004 14288 2010 14300
rect 3234 14288 3240 14340
rect 3292 14328 3298 14340
rect 3436 14328 3464 14359
rect 4614 14356 4620 14368
rect 4672 14396 4678 14408
rect 5258 14396 5264 14408
rect 4672 14368 5264 14396
rect 4672 14356 4678 14368
rect 5258 14356 5264 14368
rect 5316 14356 5322 14408
rect 5442 14356 5448 14408
rect 5500 14396 5506 14408
rect 6380 14405 6408 14436
rect 7282 14424 7288 14436
rect 7340 14424 7346 14476
rect 10796 14464 10824 14504
rect 11882 14492 11888 14504
rect 11940 14492 11946 14544
rect 13354 14532 13360 14544
rect 12176 14504 13360 14532
rect 11054 14464 11060 14476
rect 8404 14436 10824 14464
rect 11015 14436 11060 14464
rect 5997 14399 6055 14405
rect 5997 14396 6009 14399
rect 5500 14368 6009 14396
rect 5500 14356 5506 14368
rect 5997 14365 6009 14368
rect 6043 14365 6055 14399
rect 5997 14359 6055 14365
rect 6365 14399 6423 14405
rect 6365 14365 6377 14399
rect 6411 14365 6423 14399
rect 7006 14396 7012 14408
rect 6967 14368 7012 14396
rect 6365 14359 6423 14365
rect 7006 14356 7012 14368
rect 7064 14356 7070 14408
rect 7374 14396 7380 14408
rect 7335 14368 7380 14396
rect 7374 14356 7380 14368
rect 7432 14356 7438 14408
rect 7926 14396 7932 14408
rect 7887 14368 7932 14396
rect 7926 14356 7932 14368
rect 7984 14356 7990 14408
rect 3510 14328 3516 14340
rect 3292 14300 3337 14328
rect 3436 14300 3516 14328
rect 3292 14288 3298 14300
rect 3510 14288 3516 14300
rect 3568 14288 3574 14340
rect 6086 14328 6092 14340
rect 6047 14300 6092 14328
rect 6086 14288 6092 14300
rect 6144 14288 6150 14340
rect 6178 14288 6184 14340
rect 6236 14328 6242 14340
rect 7101 14331 7159 14337
rect 7101 14328 7113 14331
rect 6236 14300 6281 14328
rect 7024 14300 7113 14328
rect 6236 14288 6242 14300
rect 7024 14272 7052 14300
rect 7101 14297 7113 14300
rect 7147 14297 7159 14331
rect 7101 14291 7159 14297
rect 7193 14331 7251 14337
rect 7193 14297 7205 14331
rect 7239 14328 7251 14331
rect 8294 14328 8300 14340
rect 7239 14300 8300 14328
rect 7239 14297 7251 14300
rect 7193 14291 7251 14297
rect 8294 14288 8300 14300
rect 8352 14288 8358 14340
rect 8404 14337 8432 14436
rect 11054 14424 11060 14436
rect 11112 14424 11118 14476
rect 12176 14473 12204 14504
rect 13354 14492 13360 14504
rect 13412 14492 13418 14544
rect 14844 14532 14872 14572
rect 14918 14560 14924 14612
rect 14976 14600 14982 14612
rect 15013 14603 15071 14609
rect 15013 14600 15025 14603
rect 14976 14572 15025 14600
rect 14976 14560 14982 14572
rect 15013 14569 15025 14572
rect 15059 14569 15071 14603
rect 17402 14600 17408 14612
rect 15013 14563 15071 14569
rect 15120 14572 17408 14600
rect 15120 14532 15148 14572
rect 17402 14560 17408 14572
rect 17460 14560 17466 14612
rect 19334 14560 19340 14612
rect 19392 14600 19398 14612
rect 19429 14603 19487 14609
rect 19429 14600 19441 14603
rect 19392 14572 19441 14600
rect 19392 14560 19398 14572
rect 19429 14569 19441 14572
rect 19475 14569 19487 14603
rect 19429 14563 19487 14569
rect 19536 14572 19840 14600
rect 14844 14504 15148 14532
rect 15194 14492 15200 14544
rect 15252 14532 15258 14544
rect 16390 14532 16396 14544
rect 15252 14504 16396 14532
rect 15252 14492 15258 14504
rect 16390 14492 16396 14504
rect 16448 14532 16454 14544
rect 19536 14532 19564 14572
rect 16448 14504 19564 14532
rect 16448 14492 16454 14504
rect 19702 14492 19708 14544
rect 19760 14492 19766 14544
rect 19812 14532 19840 14572
rect 20346 14560 20352 14612
rect 20404 14600 20410 14612
rect 20441 14603 20499 14609
rect 20441 14600 20453 14603
rect 20404 14572 20453 14600
rect 20404 14560 20410 14572
rect 20441 14569 20453 14572
rect 20487 14569 20499 14603
rect 20441 14563 20499 14569
rect 20714 14560 20720 14612
rect 20772 14600 20778 14612
rect 22373 14603 22431 14609
rect 22373 14600 22385 14603
rect 20772 14572 22385 14600
rect 20772 14560 20778 14572
rect 22373 14569 22385 14572
rect 22419 14569 22431 14603
rect 22373 14563 22431 14569
rect 21266 14532 21272 14544
rect 19812 14504 21272 14532
rect 21266 14492 21272 14504
rect 21324 14492 21330 14544
rect 12161 14467 12219 14473
rect 12161 14433 12173 14467
rect 12207 14433 12219 14467
rect 12342 14464 12348 14476
rect 12303 14436 12348 14464
rect 12161 14427 12219 14433
rect 12342 14424 12348 14436
rect 12400 14424 12406 14476
rect 12437 14467 12495 14473
rect 12437 14433 12449 14467
rect 12483 14464 12495 14467
rect 12710 14464 12716 14476
rect 12483 14436 12716 14464
rect 12483 14433 12495 14436
rect 12437 14427 12495 14433
rect 12710 14424 12716 14436
rect 12768 14424 12774 14476
rect 14182 14424 14188 14476
rect 14240 14464 14246 14476
rect 14240 14436 14780 14464
rect 14240 14424 14246 14436
rect 9306 14396 9312 14408
rect 9267 14368 9312 14396
rect 9306 14356 9312 14368
rect 9364 14356 9370 14408
rect 9674 14396 9680 14408
rect 9635 14368 9680 14396
rect 9674 14356 9680 14368
rect 9732 14356 9738 14408
rect 12253 14399 12311 14405
rect 12253 14365 12265 14399
rect 12299 14365 12311 14399
rect 12802 14396 12808 14408
rect 12253 14359 12311 14365
rect 12406 14368 12808 14396
rect 8389 14331 8447 14337
rect 8389 14297 8401 14331
rect 8435 14297 8447 14331
rect 9398 14328 9404 14340
rect 9359 14300 9404 14328
rect 8389 14291 8447 14297
rect 2866 14260 2872 14272
rect 2827 14232 2872 14260
rect 2866 14220 2872 14232
rect 2924 14220 2930 14272
rect 7006 14220 7012 14272
rect 7064 14260 7070 14272
rect 8404 14260 8432 14291
rect 9398 14288 9404 14300
rect 9456 14288 9462 14340
rect 9493 14331 9551 14337
rect 9493 14297 9505 14331
rect 9539 14297 9551 14331
rect 11146 14328 11152 14340
rect 11107 14300 11152 14328
rect 9493 14291 9551 14297
rect 7064 14232 8432 14260
rect 7064 14220 7070 14232
rect 9214 14220 9220 14272
rect 9272 14260 9278 14272
rect 9508 14260 9536 14291
rect 11146 14288 11152 14300
rect 11204 14288 11210 14340
rect 11241 14331 11299 14337
rect 11241 14297 11253 14331
rect 11287 14328 11299 14331
rect 11790 14328 11796 14340
rect 11287 14300 11796 14328
rect 11287 14297 11299 14300
rect 11241 14291 11299 14297
rect 11790 14288 11796 14300
rect 11848 14288 11854 14340
rect 12268 14328 12296 14359
rect 12406 14328 12434 14368
rect 12802 14356 12808 14368
rect 12860 14396 12866 14408
rect 13538 14396 13544 14408
rect 12860 14368 13544 14396
rect 12860 14356 12866 14368
rect 13538 14356 13544 14368
rect 13596 14356 13602 14408
rect 14274 14396 14280 14408
rect 14235 14368 14280 14396
rect 14274 14356 14280 14368
rect 14332 14356 14338 14408
rect 14369 14399 14427 14405
rect 14369 14365 14381 14399
rect 14415 14365 14427 14399
rect 14550 14396 14556 14408
rect 14511 14368 14556 14396
rect 14369 14359 14427 14365
rect 12268 14300 12434 14328
rect 13354 14288 13360 14340
rect 13412 14328 13418 14340
rect 13449 14331 13507 14337
rect 13449 14328 13461 14331
rect 13412 14300 13461 14328
rect 13412 14288 13418 14300
rect 13449 14297 13461 14300
rect 13495 14297 13507 14331
rect 13449 14291 13507 14297
rect 13998 14288 14004 14340
rect 14056 14328 14062 14340
rect 14182 14328 14188 14340
rect 14056 14300 14188 14328
rect 14056 14288 14062 14300
rect 14182 14288 14188 14300
rect 14240 14328 14246 14340
rect 14384 14328 14412 14359
rect 14550 14356 14556 14368
rect 14608 14356 14614 14408
rect 14752 14405 14780 14436
rect 15378 14424 15384 14476
rect 15436 14464 15442 14476
rect 16206 14464 16212 14476
rect 15436 14436 16212 14464
rect 15436 14424 15442 14436
rect 16206 14424 16212 14436
rect 16264 14424 16270 14476
rect 17126 14424 17132 14476
rect 17184 14464 17190 14476
rect 17497 14467 17555 14473
rect 17497 14464 17509 14467
rect 17184 14436 17509 14464
rect 17184 14424 17190 14436
rect 17497 14433 17509 14436
rect 17543 14433 17555 14467
rect 19720 14464 19748 14492
rect 19720 14436 19932 14464
rect 17497 14427 17555 14433
rect 14737 14399 14795 14405
rect 14737 14365 14749 14399
rect 14783 14396 14795 14399
rect 15930 14396 15936 14408
rect 14783 14368 15936 14396
rect 14783 14365 14795 14368
rect 14737 14359 14795 14365
rect 15930 14356 15936 14368
rect 15988 14396 15994 14408
rect 16758 14396 16764 14408
rect 15988 14368 16764 14396
rect 15988 14356 15994 14368
rect 16758 14356 16764 14368
rect 16816 14356 16822 14408
rect 17310 14396 17316 14408
rect 17271 14368 17316 14396
rect 17310 14356 17316 14368
rect 17368 14356 17374 14408
rect 17402 14356 17408 14408
rect 17460 14396 17466 14408
rect 17589 14399 17647 14405
rect 17460 14368 17553 14396
rect 17460 14356 17466 14368
rect 17589 14365 17601 14399
rect 17635 14396 17647 14399
rect 19334 14396 19340 14408
rect 17635 14368 19340 14396
rect 17635 14365 17647 14368
rect 17589 14359 17647 14365
rect 19334 14356 19340 14368
rect 19392 14356 19398 14408
rect 19610 14396 19616 14408
rect 19571 14368 19616 14396
rect 19610 14356 19616 14368
rect 19668 14356 19674 14408
rect 19904 14405 19932 14436
rect 19996 14436 22140 14464
rect 19996 14405 20024 14436
rect 22112 14408 22140 14436
rect 19705 14399 19763 14405
rect 19705 14365 19717 14399
rect 19751 14365 19763 14399
rect 19705 14359 19763 14365
rect 19889 14399 19947 14405
rect 19889 14365 19901 14399
rect 19935 14365 19947 14399
rect 19889 14359 19947 14365
rect 19981 14399 20039 14405
rect 19981 14365 19993 14399
rect 20027 14365 20039 14399
rect 19981 14359 20039 14365
rect 21085 14399 21143 14405
rect 21085 14365 21097 14399
rect 21131 14396 21143 14399
rect 21450 14396 21456 14408
rect 21131 14368 21456 14396
rect 21131 14365 21143 14368
rect 21085 14359 21143 14365
rect 14642 14328 14648 14340
rect 14240 14300 14412 14328
rect 14555 14300 14648 14328
rect 14240 14288 14246 14300
rect 14642 14288 14648 14300
rect 14700 14328 14706 14340
rect 15470 14328 15476 14340
rect 14700 14300 15476 14328
rect 14700 14288 14706 14300
rect 15470 14288 15476 14300
rect 15528 14288 15534 14340
rect 16025 14331 16083 14337
rect 16025 14297 16037 14331
rect 16071 14328 16083 14331
rect 17420 14328 17448 14356
rect 16071 14300 17172 14328
rect 16071 14297 16083 14300
rect 16025 14291 16083 14297
rect 9272 14232 9536 14260
rect 9272 14220 9278 14232
rect 11330 14220 11336 14272
rect 11388 14260 11394 14272
rect 15378 14260 15384 14272
rect 11388 14232 15384 14260
rect 11388 14220 11394 14232
rect 15378 14220 15384 14232
rect 15436 14220 15442 14272
rect 15654 14260 15660 14272
rect 15615 14232 15660 14260
rect 15654 14220 15660 14232
rect 15712 14220 15718 14272
rect 16114 14260 16120 14272
rect 16075 14232 16120 14260
rect 16114 14220 16120 14232
rect 16172 14220 16178 14272
rect 17144 14269 17172 14300
rect 17236 14300 17448 14328
rect 17236 14272 17264 14300
rect 19150 14288 19156 14340
rect 19208 14328 19214 14340
rect 19720 14328 19748 14359
rect 19208 14300 19748 14328
rect 19904 14328 19932 14359
rect 21450 14356 21456 14368
rect 21508 14356 21514 14408
rect 21726 14396 21732 14408
rect 21687 14368 21732 14396
rect 21726 14356 21732 14368
rect 21784 14356 21790 14408
rect 22094 14356 22100 14408
rect 22152 14396 22158 14408
rect 22557 14399 22615 14405
rect 22557 14396 22569 14399
rect 22152 14368 22569 14396
rect 22152 14356 22158 14368
rect 22557 14365 22569 14368
rect 22603 14365 22615 14399
rect 22830 14396 22836 14408
rect 22791 14368 22836 14396
rect 22557 14359 22615 14365
rect 22830 14356 22836 14368
rect 22888 14356 22894 14408
rect 20070 14328 20076 14340
rect 19904 14300 20076 14328
rect 19208 14288 19214 14300
rect 20070 14288 20076 14300
rect 20128 14288 20134 14340
rect 17129 14263 17187 14269
rect 17129 14229 17141 14263
rect 17175 14229 17187 14263
rect 17129 14223 17187 14229
rect 17218 14220 17224 14272
rect 17276 14220 17282 14272
rect 18690 14220 18696 14272
rect 18748 14260 18754 14272
rect 20254 14260 20260 14272
rect 18748 14232 20260 14260
rect 18748 14220 18754 14232
rect 20254 14220 20260 14232
rect 20312 14220 20318 14272
rect 21821 14263 21879 14269
rect 21821 14229 21833 14263
rect 21867 14260 21879 14263
rect 22462 14260 22468 14272
rect 21867 14232 22468 14260
rect 21867 14229 21879 14232
rect 21821 14223 21879 14229
rect 22462 14220 22468 14232
rect 22520 14220 22526 14272
rect 22741 14263 22799 14269
rect 22741 14229 22753 14263
rect 22787 14260 22799 14263
rect 22922 14260 22928 14272
rect 22787 14232 22928 14260
rect 22787 14229 22799 14232
rect 22741 14223 22799 14229
rect 22922 14220 22928 14232
rect 22980 14220 22986 14272
rect 1104 14170 23987 14192
rect 1104 14118 6630 14170
rect 6682 14118 6694 14170
rect 6746 14118 6758 14170
rect 6810 14118 6822 14170
rect 6874 14118 6886 14170
rect 6938 14118 12311 14170
rect 12363 14118 12375 14170
rect 12427 14118 12439 14170
rect 12491 14118 12503 14170
rect 12555 14118 12567 14170
rect 12619 14118 17992 14170
rect 18044 14118 18056 14170
rect 18108 14118 18120 14170
rect 18172 14118 18184 14170
rect 18236 14118 18248 14170
rect 18300 14118 23673 14170
rect 23725 14118 23737 14170
rect 23789 14118 23801 14170
rect 23853 14118 23865 14170
rect 23917 14118 23929 14170
rect 23981 14118 23987 14170
rect 1104 14096 23987 14118
rect 3050 14016 3056 14068
rect 3108 14016 3114 14068
rect 3694 14016 3700 14068
rect 3752 14056 3758 14068
rect 3973 14059 4031 14065
rect 3973 14056 3985 14059
rect 3752 14028 3985 14056
rect 3752 14016 3758 14028
rect 3973 14025 3985 14028
rect 4019 14025 4031 14059
rect 5074 14056 5080 14068
rect 5035 14028 5080 14056
rect 3973 14019 4031 14025
rect 5074 14016 5080 14028
rect 5132 14016 5138 14068
rect 9585 14059 9643 14065
rect 9585 14025 9597 14059
rect 9631 14056 9643 14059
rect 10134 14056 10140 14068
rect 9631 14028 10140 14056
rect 9631 14025 9643 14028
rect 9585 14019 9643 14025
rect 10134 14016 10140 14028
rect 10192 14016 10198 14068
rect 12802 14056 12808 14068
rect 12763 14028 12808 14056
rect 12802 14016 12808 14028
rect 12860 14016 12866 14068
rect 15565 14059 15623 14065
rect 15565 14025 15577 14059
rect 15611 14056 15623 14059
rect 16114 14056 16120 14068
rect 15611 14028 16120 14056
rect 15611 14025 15623 14028
rect 15565 14019 15623 14025
rect 16114 14016 16120 14028
rect 16172 14016 16178 14068
rect 16942 14016 16948 14068
rect 17000 14056 17006 14068
rect 17402 14056 17408 14068
rect 17000 14028 17408 14056
rect 17000 14016 17006 14028
rect 17402 14016 17408 14028
rect 17460 14056 17466 14068
rect 17460 14028 18276 14056
rect 17460 14016 17466 14028
rect 2866 13997 2872 14000
rect 2860 13988 2872 13997
rect 2827 13960 2872 13988
rect 2860 13951 2872 13960
rect 2866 13948 2872 13951
rect 2924 13948 2930 14000
rect 2133 13923 2191 13929
rect 2133 13889 2145 13923
rect 2179 13920 2191 13923
rect 2498 13920 2504 13932
rect 2179 13892 2504 13920
rect 2179 13889 2191 13892
rect 2133 13883 2191 13889
rect 2498 13880 2504 13892
rect 2556 13880 2562 13932
rect 2593 13923 2651 13929
rect 2593 13889 2605 13923
rect 2639 13920 2651 13923
rect 3068 13920 3096 14016
rect 8472 13991 8530 13997
rect 8472 13957 8484 13991
rect 8518 13988 8530 13991
rect 13078 13988 13084 14000
rect 8518 13960 13084 13988
rect 8518 13957 8530 13960
rect 8472 13951 8530 13957
rect 13078 13948 13084 13960
rect 13136 13948 13142 14000
rect 15194 13988 15200 14000
rect 14757 13960 15200 13988
rect 5442 13920 5448 13932
rect 2639 13892 3096 13920
rect 5403 13892 5448 13920
rect 2639 13889 2651 13892
rect 2593 13883 2651 13889
rect 5442 13880 5448 13892
rect 5500 13880 5506 13932
rect 5537 13923 5595 13929
rect 5537 13889 5549 13923
rect 5583 13920 5595 13923
rect 6178 13920 6184 13932
rect 5583 13892 6184 13920
rect 5583 13889 5595 13892
rect 5537 13883 5595 13889
rect 6178 13880 6184 13892
rect 6236 13880 6242 13932
rect 8202 13920 8208 13932
rect 8163 13892 8208 13920
rect 8202 13880 8208 13892
rect 8260 13880 8266 13932
rect 9674 13920 9680 13932
rect 8312 13892 9680 13920
rect 1854 13852 1860 13864
rect 1815 13824 1860 13852
rect 1854 13812 1860 13824
rect 1912 13812 1918 13864
rect 5350 13812 5356 13864
rect 5408 13852 5414 13864
rect 5629 13855 5687 13861
rect 5629 13852 5641 13855
rect 5408 13824 5641 13852
rect 5408 13812 5414 13824
rect 5629 13821 5641 13824
rect 5675 13852 5687 13855
rect 5902 13852 5908 13864
rect 5675 13824 5908 13852
rect 5675 13821 5687 13824
rect 5629 13815 5687 13821
rect 5902 13812 5908 13824
rect 5960 13812 5966 13864
rect 7834 13812 7840 13864
rect 7892 13852 7898 13864
rect 8312 13852 8340 13892
rect 9674 13880 9680 13892
rect 9732 13880 9738 13932
rect 10042 13920 10048 13932
rect 10003 13892 10048 13920
rect 10042 13880 10048 13892
rect 10100 13880 10106 13932
rect 10229 13923 10287 13929
rect 10229 13889 10241 13923
rect 10275 13920 10287 13923
rect 10686 13920 10692 13932
rect 10275 13892 10692 13920
rect 10275 13889 10287 13892
rect 10229 13883 10287 13889
rect 10686 13880 10692 13892
rect 10744 13880 10750 13932
rect 10778 13880 10784 13932
rect 10836 13920 10842 13932
rect 10903 13923 10961 13929
rect 10903 13920 10915 13923
rect 10836 13892 10915 13920
rect 10836 13880 10842 13892
rect 10903 13889 10915 13892
rect 10949 13889 10961 13923
rect 10903 13883 10961 13889
rect 11057 13923 11115 13929
rect 11057 13889 11069 13923
rect 11103 13920 11115 13923
rect 12710 13920 12716 13932
rect 11103 13892 12716 13920
rect 11103 13889 11115 13892
rect 11057 13883 11115 13889
rect 12710 13880 12716 13892
rect 12768 13880 12774 13932
rect 14458 13880 14464 13932
rect 14516 13920 14522 13932
rect 14553 13923 14611 13929
rect 14553 13920 14565 13923
rect 14516 13892 14565 13920
rect 14516 13880 14522 13892
rect 14553 13889 14565 13892
rect 14599 13889 14611 13923
rect 14553 13883 14611 13889
rect 14645 13923 14703 13929
rect 14645 13889 14657 13923
rect 14691 13920 14703 13923
rect 14757 13920 14785 13960
rect 15194 13948 15200 13960
rect 15252 13948 15258 14000
rect 15838 13988 15844 14000
rect 15799 13960 15844 13988
rect 15838 13948 15844 13960
rect 15896 13948 15902 14000
rect 16022 13948 16028 14000
rect 16080 13988 16086 14000
rect 16080 13960 18184 13988
rect 16080 13948 16086 13960
rect 14691 13892 14785 13920
rect 14829 13923 14887 13929
rect 14691 13889 14703 13892
rect 14645 13883 14703 13889
rect 14829 13889 14841 13923
rect 14875 13889 14887 13923
rect 14829 13883 14887 13889
rect 11790 13852 11796 13864
rect 7892 13824 8340 13852
rect 11751 13824 11796 13852
rect 7892 13812 7898 13824
rect 11790 13812 11796 13824
rect 11848 13812 11854 13864
rect 14274 13812 14280 13864
rect 14332 13852 14338 13864
rect 14844 13852 14872 13883
rect 14918 13880 14924 13932
rect 14976 13920 14982 13932
rect 15746 13920 15752 13932
rect 14976 13892 15021 13920
rect 15707 13892 15752 13920
rect 14976 13880 14982 13892
rect 15746 13880 15752 13892
rect 15804 13880 15810 13932
rect 15930 13880 15936 13932
rect 15988 13920 15994 13932
rect 16117 13923 16175 13929
rect 15988 13892 16033 13920
rect 15988 13880 15994 13892
rect 16117 13889 16129 13923
rect 16163 13920 16175 13923
rect 16942 13920 16948 13932
rect 16163 13892 16948 13920
rect 16163 13889 16175 13892
rect 16117 13883 16175 13889
rect 16942 13880 16948 13892
rect 17000 13880 17006 13932
rect 17865 13923 17923 13929
rect 17865 13889 17877 13923
rect 17911 13889 17923 13923
rect 17865 13883 17923 13889
rect 15654 13852 15660 13864
rect 14332 13824 15660 13852
rect 14332 13812 14338 13824
rect 15654 13812 15660 13824
rect 15712 13812 15718 13864
rect 17880 13852 17908 13883
rect 17954 13880 17960 13932
rect 18012 13920 18018 13932
rect 18156 13929 18184 13960
rect 18248 13932 18276 14028
rect 19794 14016 19800 14068
rect 19852 14056 19858 14068
rect 20349 14059 20407 14065
rect 20349 14056 20361 14059
rect 19852 14028 20361 14056
rect 19852 14016 19858 14028
rect 20349 14025 20361 14028
rect 20395 14025 20407 14059
rect 21450 14056 21456 14068
rect 20349 14019 20407 14025
rect 20732 14028 21456 14056
rect 18141 13923 18199 13929
rect 18012 13892 18057 13920
rect 18012 13880 18018 13892
rect 18141 13889 18153 13923
rect 18187 13889 18199 13923
rect 18141 13883 18199 13889
rect 18230 13880 18236 13932
rect 18288 13920 18294 13932
rect 19245 13923 19303 13929
rect 18288 13892 18333 13920
rect 18288 13880 18294 13892
rect 19245 13889 19257 13923
rect 19291 13920 19303 13923
rect 20254 13920 20260 13932
rect 19291 13892 20260 13920
rect 19291 13889 19303 13892
rect 19245 13883 19303 13889
rect 20254 13880 20260 13892
rect 20312 13880 20318 13932
rect 20732 13929 20760 14028
rect 21450 14016 21456 14028
rect 21508 14016 21514 14068
rect 22649 13991 22707 13997
rect 22649 13988 22661 13991
rect 21928 13960 22661 13988
rect 20990 13929 20996 13932
rect 20625 13923 20683 13929
rect 20625 13889 20637 13923
rect 20671 13889 20683 13923
rect 20625 13883 20683 13889
rect 20717 13923 20775 13929
rect 20717 13889 20729 13923
rect 20763 13889 20775 13923
rect 20809 13923 20867 13929
rect 20809 13898 20821 13923
rect 20855 13898 20867 13923
rect 20717 13883 20775 13889
rect 19061 13855 19119 13861
rect 19061 13852 19073 13855
rect 17880 13824 19073 13852
rect 19061 13821 19073 13824
rect 19107 13821 19119 13855
rect 19061 13815 19119 13821
rect 19150 13812 19156 13864
rect 19208 13852 19214 13864
rect 19337 13855 19395 13861
rect 19337 13852 19349 13855
rect 19208 13824 19349 13852
rect 19208 13812 19214 13824
rect 19337 13821 19349 13824
rect 19383 13821 19395 13855
rect 19337 13815 19395 13821
rect 19429 13855 19487 13861
rect 19429 13821 19441 13855
rect 19475 13821 19487 13855
rect 19429 13815 19487 13821
rect 1949 13787 2007 13793
rect 1949 13753 1961 13787
rect 1995 13784 2007 13787
rect 2314 13784 2320 13796
rect 1995 13756 2320 13784
rect 1995 13753 2007 13756
rect 1949 13747 2007 13753
rect 2314 13744 2320 13756
rect 2372 13744 2378 13796
rect 17678 13784 17684 13796
rect 17639 13756 17684 13784
rect 17678 13744 17684 13756
rect 17736 13744 17742 13796
rect 2038 13716 2044 13728
rect 1999 13688 2044 13716
rect 2038 13676 2044 13688
rect 2096 13676 2102 13728
rect 3694 13676 3700 13728
rect 3752 13716 3758 13728
rect 5718 13716 5724 13728
rect 3752 13688 5724 13716
rect 3752 13676 3758 13688
rect 5718 13676 5724 13688
rect 5776 13676 5782 13728
rect 7006 13676 7012 13728
rect 7064 13716 7070 13728
rect 7469 13719 7527 13725
rect 7469 13716 7481 13719
rect 7064 13688 7481 13716
rect 7064 13676 7070 13688
rect 7469 13685 7481 13688
rect 7515 13685 7527 13719
rect 7469 13679 7527 13685
rect 10229 13719 10287 13725
rect 10229 13685 10241 13719
rect 10275 13716 10287 13719
rect 10318 13716 10324 13728
rect 10275 13688 10324 13716
rect 10275 13685 10287 13688
rect 10229 13679 10287 13685
rect 10318 13676 10324 13688
rect 10376 13676 10382 13728
rect 10873 13719 10931 13725
rect 10873 13685 10885 13719
rect 10919 13716 10931 13719
rect 11606 13716 11612 13728
rect 10919 13688 11612 13716
rect 10919 13685 10931 13688
rect 10873 13679 10931 13685
rect 11606 13676 11612 13688
rect 11664 13676 11670 13728
rect 14090 13716 14096 13728
rect 14051 13688 14096 13716
rect 14090 13676 14096 13688
rect 14148 13676 14154 13728
rect 15105 13719 15163 13725
rect 15105 13685 15117 13719
rect 15151 13716 15163 13719
rect 15470 13716 15476 13728
rect 15151 13688 15476 13716
rect 15151 13685 15163 13688
rect 15105 13679 15163 13685
rect 15470 13676 15476 13688
rect 15528 13676 15534 13728
rect 15654 13676 15660 13728
rect 15712 13716 15718 13728
rect 16945 13719 17003 13725
rect 16945 13716 16957 13719
rect 15712 13688 16957 13716
rect 15712 13676 15718 13688
rect 16945 13685 16957 13688
rect 16991 13716 17003 13719
rect 18874 13716 18880 13728
rect 16991 13688 18880 13716
rect 16991 13685 17003 13688
rect 16945 13679 17003 13685
rect 18874 13676 18880 13688
rect 18932 13716 18938 13728
rect 19444 13716 19472 13815
rect 19518 13812 19524 13864
rect 19576 13852 19582 13864
rect 19576 13824 19621 13852
rect 19576 13812 19582 13824
rect 20640 13784 20668 13883
rect 20806 13846 20812 13898
rect 20864 13846 20870 13898
rect 20987 13883 20996 13929
rect 21048 13920 21054 13932
rect 21048 13892 21087 13920
rect 20990 13880 20996 13883
rect 21048 13880 21054 13892
rect 21634 13880 21640 13932
rect 21692 13920 21698 13932
rect 21928 13920 21956 13960
rect 22649 13957 22661 13960
rect 22695 13957 22707 13991
rect 22649 13951 22707 13957
rect 22738 13948 22744 14000
rect 22796 13988 22802 14000
rect 22796 13960 23244 13988
rect 22796 13948 22802 13960
rect 22278 13920 22284 13932
rect 21692 13892 21956 13920
rect 22239 13892 22284 13920
rect 21692 13880 21698 13892
rect 22278 13880 22284 13892
rect 22336 13880 22342 13932
rect 22554 13920 22560 13932
rect 22515 13892 22560 13920
rect 22554 13880 22560 13892
rect 22612 13880 22618 13932
rect 22833 13923 22891 13929
rect 22833 13889 22845 13923
rect 22879 13920 22891 13923
rect 23106 13920 23112 13932
rect 22879 13892 23112 13920
rect 22879 13889 22891 13892
rect 22833 13883 22891 13889
rect 21818 13784 21824 13796
rect 20640 13756 21824 13784
rect 21818 13744 21824 13756
rect 21876 13744 21882 13796
rect 22940 13784 22968 13892
rect 23106 13880 23112 13892
rect 23164 13880 23170 13932
rect 23017 13855 23075 13861
rect 23017 13821 23029 13855
rect 23063 13852 23075 13855
rect 23216 13852 23244 13960
rect 23063 13824 23244 13852
rect 23063 13821 23075 13824
rect 23017 13815 23075 13821
rect 23382 13784 23388 13796
rect 22940 13756 23388 13784
rect 23382 13744 23388 13756
rect 23440 13744 23446 13796
rect 18932 13688 19472 13716
rect 18932 13676 18938 13688
rect 19978 13676 19984 13728
rect 20036 13716 20042 13728
rect 22278 13716 22284 13728
rect 20036 13688 22284 13716
rect 20036 13676 20042 13688
rect 22278 13676 22284 13688
rect 22336 13676 22342 13728
rect 1104 13626 23828 13648
rect 1104 13574 3790 13626
rect 3842 13574 3854 13626
rect 3906 13574 3918 13626
rect 3970 13574 3982 13626
rect 4034 13574 4046 13626
rect 4098 13574 9471 13626
rect 9523 13574 9535 13626
rect 9587 13574 9599 13626
rect 9651 13574 9663 13626
rect 9715 13574 9727 13626
rect 9779 13574 15152 13626
rect 15204 13574 15216 13626
rect 15268 13574 15280 13626
rect 15332 13574 15344 13626
rect 15396 13574 15408 13626
rect 15460 13574 20833 13626
rect 20885 13574 20897 13626
rect 20949 13574 20961 13626
rect 21013 13574 21025 13626
rect 21077 13574 21089 13626
rect 21141 13574 23828 13626
rect 1104 13552 23828 13574
rect 2498 13472 2504 13524
rect 2556 13512 2562 13524
rect 4433 13515 4491 13521
rect 2556 13484 4384 13512
rect 2556 13472 2562 13484
rect 2685 13447 2743 13453
rect 2685 13413 2697 13447
rect 2731 13444 2743 13447
rect 3694 13444 3700 13456
rect 2731 13416 3700 13444
rect 2731 13413 2743 13416
rect 2685 13407 2743 13413
rect 3694 13404 3700 13416
rect 3752 13404 3758 13456
rect 3510 13376 3516 13388
rect 2148 13348 3516 13376
rect 2148 13317 2176 13348
rect 3510 13336 3516 13348
rect 3568 13336 3574 13388
rect 4246 13336 4252 13388
rect 4304 13336 4310 13388
rect 2133 13311 2191 13317
rect 2133 13277 2145 13311
rect 2179 13277 2191 13311
rect 2314 13308 2320 13320
rect 2275 13280 2320 13308
rect 2133 13271 2191 13277
rect 2314 13268 2320 13280
rect 2372 13268 2378 13320
rect 2501 13311 2559 13317
rect 2501 13277 2513 13311
rect 2547 13308 2559 13311
rect 2682 13308 2688 13320
rect 2547 13280 2688 13308
rect 2547 13277 2559 13280
rect 2501 13271 2559 13277
rect 2682 13268 2688 13280
rect 2740 13268 2746 13320
rect 3421 13311 3479 13317
rect 3421 13277 3433 13311
rect 3467 13308 3479 13311
rect 4264 13308 4292 13336
rect 3467 13280 4292 13308
rect 3467 13277 3479 13280
rect 3421 13271 3479 13277
rect 4356 13252 4384 13484
rect 4433 13481 4445 13515
rect 4479 13481 4491 13515
rect 4614 13512 4620 13524
rect 4575 13484 4620 13512
rect 4433 13475 4491 13481
rect 4448 13444 4476 13475
rect 4614 13472 4620 13484
rect 4672 13472 4678 13524
rect 4982 13472 4988 13524
rect 5040 13512 5046 13524
rect 5261 13515 5319 13521
rect 5261 13512 5273 13515
rect 5040 13484 5273 13512
rect 5040 13472 5046 13484
rect 5261 13481 5273 13484
rect 5307 13481 5319 13515
rect 5261 13475 5319 13481
rect 6178 13472 6184 13524
rect 6236 13512 6242 13524
rect 6641 13515 6699 13521
rect 6641 13512 6653 13515
rect 6236 13484 6653 13512
rect 6236 13472 6242 13484
rect 6641 13481 6653 13484
rect 6687 13481 6699 13515
rect 6641 13475 6699 13481
rect 9677 13515 9735 13521
rect 9677 13481 9689 13515
rect 9723 13512 9735 13515
rect 11330 13512 11336 13524
rect 9723 13484 11336 13512
rect 9723 13481 9735 13484
rect 9677 13475 9735 13481
rect 11330 13472 11336 13484
rect 11388 13472 11394 13524
rect 15657 13515 15715 13521
rect 15657 13481 15669 13515
rect 15703 13512 15715 13515
rect 15746 13512 15752 13524
rect 15703 13484 15752 13512
rect 15703 13481 15715 13484
rect 15657 13475 15715 13481
rect 15746 13472 15752 13484
rect 15804 13472 15810 13524
rect 16577 13515 16635 13521
rect 16577 13481 16589 13515
rect 16623 13512 16635 13515
rect 17310 13512 17316 13524
rect 16623 13484 17316 13512
rect 16623 13481 16635 13484
rect 16577 13475 16635 13481
rect 17310 13472 17316 13484
rect 17368 13472 17374 13524
rect 19429 13515 19487 13521
rect 19429 13481 19441 13515
rect 19475 13512 19487 13515
rect 19610 13512 19616 13524
rect 19475 13484 19616 13512
rect 19475 13481 19487 13484
rect 19429 13475 19487 13481
rect 19610 13472 19616 13484
rect 19668 13472 19674 13524
rect 19702 13472 19708 13524
rect 19760 13472 19766 13524
rect 19794 13472 19800 13524
rect 19852 13512 19858 13524
rect 20625 13515 20683 13521
rect 20625 13512 20637 13515
rect 19852 13484 20637 13512
rect 19852 13472 19858 13484
rect 20625 13481 20637 13484
rect 20671 13481 20683 13515
rect 21450 13512 21456 13524
rect 21411 13484 21456 13512
rect 20625 13475 20683 13481
rect 21450 13472 21456 13484
rect 21508 13472 21514 13524
rect 4522 13444 4528 13456
rect 4448 13416 4528 13444
rect 4522 13404 4528 13416
rect 4580 13404 4586 13456
rect 6549 13447 6607 13453
rect 6549 13413 6561 13447
rect 6595 13444 6607 13447
rect 7098 13444 7104 13456
rect 6595 13416 7104 13444
rect 6595 13413 6607 13416
rect 6549 13407 6607 13413
rect 7098 13404 7104 13416
rect 7156 13404 7162 13456
rect 10042 13404 10048 13456
rect 10100 13444 10106 13456
rect 11241 13447 11299 13453
rect 10100 13416 10640 13444
rect 10100 13404 10106 13416
rect 5442 13336 5448 13388
rect 5500 13376 5506 13388
rect 6181 13379 6239 13385
rect 6181 13376 6193 13379
rect 5500 13348 6193 13376
rect 5500 13336 5506 13348
rect 6181 13345 6193 13348
rect 6227 13345 6239 13379
rect 6181 13339 6239 13345
rect 6270 13336 6276 13388
rect 6328 13376 6334 13388
rect 10318 13376 10324 13388
rect 6328 13348 7880 13376
rect 10279 13348 10324 13376
rect 6328 13336 6334 13348
rect 5166 13308 5172 13320
rect 5127 13280 5172 13308
rect 5166 13268 5172 13280
rect 5224 13268 5230 13320
rect 5258 13268 5264 13320
rect 5316 13308 5322 13320
rect 7852 13317 7880 13348
rect 10318 13336 10324 13348
rect 10376 13336 10382 13388
rect 10612 13317 10640 13416
rect 11241 13413 11253 13447
rect 11287 13444 11299 13447
rect 13354 13444 13360 13456
rect 11287 13416 13360 13444
rect 11287 13413 11299 13416
rect 11241 13407 11299 13413
rect 7193 13311 7251 13317
rect 7193 13308 7205 13311
rect 5316 13280 7205 13308
rect 5316 13268 5322 13280
rect 7193 13277 7205 13280
rect 7239 13277 7251 13311
rect 7193 13271 7251 13277
rect 7837 13311 7895 13317
rect 7837 13277 7849 13311
rect 7883 13277 7895 13311
rect 7837 13271 7895 13277
rect 10229 13311 10287 13317
rect 10229 13277 10241 13311
rect 10275 13277 10287 13311
rect 10229 13271 10287 13277
rect 10597 13311 10655 13317
rect 10597 13277 10609 13311
rect 10643 13277 10655 13311
rect 10597 13271 10655 13277
rect 2409 13243 2467 13249
rect 2409 13209 2421 13243
rect 2455 13240 2467 13243
rect 2774 13240 2780 13252
rect 2455 13212 2780 13240
rect 2455 13209 2467 13212
rect 2409 13203 2467 13209
rect 2774 13200 2780 13212
rect 2832 13240 2838 13252
rect 2832 13212 3280 13240
rect 2832 13200 2838 13212
rect 3252 13181 3280 13212
rect 3510 13200 3516 13252
rect 3568 13240 3574 13252
rect 3970 13240 3976 13252
rect 3568 13212 3976 13240
rect 3568 13200 3574 13212
rect 3970 13200 3976 13212
rect 4028 13240 4034 13252
rect 4246 13240 4252 13252
rect 4028 13212 4252 13240
rect 4028 13200 4034 13212
rect 4246 13200 4252 13212
rect 4304 13200 4310 13252
rect 4338 13200 4344 13252
rect 4396 13240 4402 13252
rect 4449 13243 4507 13249
rect 4449 13240 4461 13243
rect 4396 13212 4461 13240
rect 4396 13200 4402 13212
rect 4449 13209 4461 13212
rect 4495 13209 4507 13243
rect 4449 13203 4507 13209
rect 6546 13200 6552 13252
rect 6604 13240 6610 13252
rect 10134 13240 10140 13252
rect 6604 13212 10140 13240
rect 6604 13200 6610 13212
rect 10134 13200 10140 13212
rect 10192 13200 10198 13252
rect 10244 13240 10272 13271
rect 10686 13268 10692 13320
rect 10744 13308 10750 13320
rect 10744 13280 10789 13308
rect 10744 13268 10750 13280
rect 11256 13240 11284 13407
rect 13354 13404 13360 13416
rect 13412 13404 13418 13456
rect 14829 13447 14887 13453
rect 14829 13413 14841 13447
rect 14875 13444 14887 13447
rect 16022 13444 16028 13456
rect 14875 13416 16028 13444
rect 14875 13413 14887 13416
rect 14829 13407 14887 13413
rect 16022 13404 16028 13416
rect 16080 13404 16086 13456
rect 18414 13444 18420 13456
rect 17144 13416 18420 13444
rect 14734 13336 14740 13388
rect 14792 13376 14798 13388
rect 16942 13376 16948 13388
rect 14792 13348 16948 13376
rect 14792 13336 14798 13348
rect 11698 13268 11704 13320
rect 11756 13308 11762 13320
rect 11885 13311 11943 13317
rect 11885 13308 11897 13311
rect 11756 13280 11897 13308
rect 11756 13268 11762 13280
rect 11885 13277 11897 13280
rect 11931 13277 11943 13311
rect 11885 13271 11943 13277
rect 12066 13268 12072 13320
rect 12124 13308 12130 13320
rect 12437 13311 12495 13317
rect 12437 13308 12449 13311
rect 12124 13280 12449 13308
rect 12124 13268 12130 13280
rect 12437 13277 12449 13280
rect 12483 13277 12495 13311
rect 14274 13308 14280 13320
rect 14235 13280 14280 13308
rect 12437 13271 12495 13277
rect 14274 13268 14280 13280
rect 14332 13308 14338 13320
rect 14458 13308 14464 13320
rect 14332 13280 14464 13308
rect 14332 13268 14338 13280
rect 14458 13268 14464 13280
rect 14516 13268 14522 13320
rect 14553 13311 14611 13317
rect 14553 13277 14565 13311
rect 14599 13308 14611 13311
rect 14642 13308 14648 13320
rect 14599 13280 14648 13308
rect 14599 13277 14611 13280
rect 14553 13271 14611 13277
rect 14642 13268 14648 13280
rect 14700 13268 14706 13320
rect 15286 13308 15292 13320
rect 15247 13280 15292 13308
rect 15286 13268 15292 13280
rect 15344 13268 15350 13320
rect 15470 13308 15476 13320
rect 15431 13280 15476 13308
rect 15470 13268 15476 13280
rect 15528 13268 15534 13320
rect 16132 13317 16160 13348
rect 16942 13336 16948 13348
rect 17000 13336 17006 13388
rect 16117 13311 16175 13317
rect 16117 13277 16129 13311
rect 16163 13277 16175 13311
rect 16117 13271 16175 13277
rect 16393 13311 16451 13317
rect 16393 13277 16405 13311
rect 16439 13308 16451 13311
rect 16850 13308 16856 13320
rect 16439 13280 16856 13308
rect 16439 13277 16451 13280
rect 16393 13271 16451 13277
rect 16850 13268 16856 13280
rect 16908 13268 16914 13320
rect 17144 13317 17172 13416
rect 18414 13404 18420 13416
rect 18472 13404 18478 13456
rect 17954 13376 17960 13388
rect 17236 13348 17960 13376
rect 17037 13311 17095 13317
rect 17037 13277 17049 13311
rect 17083 13277 17095 13311
rect 17037 13271 17095 13277
rect 17129 13311 17187 13317
rect 17129 13277 17141 13311
rect 17175 13277 17187 13311
rect 17129 13271 17187 13277
rect 10244 13212 11284 13240
rect 3237 13175 3295 13181
rect 3237 13141 3249 13175
rect 3283 13141 3295 13175
rect 3237 13135 3295 13141
rect 3326 13132 3332 13184
rect 3384 13172 3390 13184
rect 5258 13172 5264 13184
rect 3384 13144 5264 13172
rect 3384 13132 3390 13144
rect 5258 13132 5264 13144
rect 5316 13132 5322 13184
rect 7190 13172 7196 13184
rect 7151 13144 7196 13172
rect 7190 13132 7196 13144
rect 7248 13172 7254 13184
rect 7742 13172 7748 13184
rect 7248 13144 7748 13172
rect 7248 13132 7254 13144
rect 7742 13132 7748 13144
rect 7800 13132 7806 13184
rect 11882 13132 11888 13184
rect 11940 13172 11946 13184
rect 12084 13172 12112 13268
rect 12986 13200 12992 13252
rect 13044 13200 13050 13252
rect 14660 13240 14688 13268
rect 15838 13240 15844 13252
rect 14660 13212 15844 13240
rect 15838 13200 15844 13212
rect 15896 13200 15902 13252
rect 16209 13243 16267 13249
rect 16209 13209 16221 13243
rect 16255 13240 16267 13243
rect 16574 13240 16580 13252
rect 16255 13212 16580 13240
rect 16255 13209 16267 13212
rect 16209 13203 16267 13209
rect 16574 13200 16580 13212
rect 16632 13200 16638 13252
rect 16758 13200 16764 13252
rect 16816 13240 16822 13252
rect 17052 13240 17080 13271
rect 17236 13240 17264 13348
rect 17954 13336 17960 13348
rect 18012 13336 18018 13388
rect 18782 13336 18788 13388
rect 18840 13376 18846 13388
rect 19518 13376 19524 13388
rect 18840 13348 19524 13376
rect 18840 13336 18846 13348
rect 19518 13336 19524 13348
rect 19576 13336 19582 13388
rect 19613 13379 19671 13385
rect 19613 13345 19625 13379
rect 19659 13345 19671 13379
rect 19720 13376 19748 13472
rect 19889 13379 19947 13385
rect 19889 13376 19901 13379
rect 19720 13348 19901 13376
rect 19613 13339 19671 13345
rect 19889 13345 19901 13348
rect 19935 13345 19947 13379
rect 20898 13376 20904 13388
rect 19889 13339 19947 13345
rect 20732 13348 20904 13376
rect 17313 13311 17371 13317
rect 17313 13277 17325 13311
rect 17359 13277 17371 13311
rect 17313 13271 17371 13277
rect 17405 13311 17463 13317
rect 17405 13277 17417 13311
rect 17451 13308 17463 13311
rect 17586 13308 17592 13320
rect 17451 13280 17592 13308
rect 17451 13277 17463 13280
rect 17405 13271 17463 13277
rect 16816 13212 17264 13240
rect 17328 13240 17356 13271
rect 17586 13268 17592 13280
rect 17644 13308 17650 13320
rect 19242 13308 19248 13320
rect 17644 13280 19248 13308
rect 17644 13268 17650 13280
rect 19242 13268 19248 13280
rect 19300 13268 19306 13320
rect 19628 13252 19656 13339
rect 19706 13311 19764 13317
rect 19706 13277 19718 13311
rect 19752 13277 19764 13311
rect 19706 13271 19764 13277
rect 19797 13311 19855 13317
rect 19797 13277 19809 13311
rect 19843 13308 19855 13311
rect 20732 13308 20760 13348
rect 20898 13336 20904 13348
rect 20956 13376 20962 13388
rect 20993 13379 21051 13385
rect 20993 13376 21005 13379
rect 20956 13348 21005 13376
rect 20956 13336 20962 13348
rect 20993 13345 21005 13348
rect 21039 13376 21051 13379
rect 21542 13376 21548 13388
rect 21039 13348 21548 13376
rect 21039 13345 21051 13348
rect 20993 13339 21051 13345
rect 21542 13336 21548 13348
rect 21600 13336 21606 13388
rect 22094 13376 22100 13388
rect 21652 13348 22100 13376
rect 21652 13317 21680 13348
rect 22094 13336 22100 13348
rect 22152 13336 22158 13388
rect 19843 13280 20760 13308
rect 20809 13311 20867 13317
rect 19843 13277 19855 13280
rect 19797 13271 19855 13277
rect 20809 13277 20821 13311
rect 20855 13277 20867 13311
rect 20809 13271 20867 13277
rect 21637 13311 21695 13317
rect 21637 13277 21649 13311
rect 21683 13277 21695 13311
rect 21637 13271 21695 13277
rect 21913 13311 21971 13317
rect 21913 13277 21925 13311
rect 21959 13308 21971 13311
rect 21959 13280 22094 13308
rect 21959 13277 21971 13280
rect 21913 13271 21971 13277
rect 19150 13240 19156 13252
rect 17328 13212 19156 13240
rect 16816 13200 16822 13212
rect 11940 13144 12112 13172
rect 11940 13132 11946 13144
rect 13998 13132 14004 13184
rect 14056 13172 14062 13184
rect 14461 13175 14519 13181
rect 14461 13172 14473 13175
rect 14056 13144 14473 13172
rect 14056 13132 14062 13144
rect 14461 13141 14473 13144
rect 14507 13172 14519 13175
rect 14550 13172 14556 13184
rect 14507 13144 14556 13172
rect 14507 13141 14519 13144
rect 14461 13135 14519 13141
rect 14550 13132 14556 13144
rect 14608 13132 14614 13184
rect 14642 13132 14648 13184
rect 14700 13172 14706 13184
rect 14700 13144 14745 13172
rect 14700 13132 14706 13144
rect 15286 13132 15292 13184
rect 15344 13172 15350 13184
rect 15470 13172 15476 13184
rect 15344 13144 15476 13172
rect 15344 13132 15350 13144
rect 15470 13132 15476 13144
rect 15528 13172 15534 13184
rect 16114 13172 16120 13184
rect 15528 13144 16120 13172
rect 15528 13132 15534 13144
rect 16114 13132 16120 13144
rect 16172 13132 16178 13184
rect 16298 13132 16304 13184
rect 16356 13172 16362 13184
rect 17328 13172 17356 13212
rect 19150 13200 19156 13212
rect 19208 13240 19214 13252
rect 19208 13212 19334 13240
rect 19208 13200 19214 13212
rect 16356 13144 17356 13172
rect 17589 13175 17647 13181
rect 16356 13132 16362 13144
rect 17589 13141 17601 13175
rect 17635 13172 17647 13175
rect 17770 13172 17776 13184
rect 17635 13144 17776 13172
rect 17635 13141 17647 13144
rect 17589 13135 17647 13141
rect 17770 13132 17776 13144
rect 17828 13132 17834 13184
rect 18874 13172 18880 13184
rect 18835 13144 18880 13172
rect 18874 13132 18880 13144
rect 18932 13132 18938 13184
rect 19306 13172 19334 13212
rect 19610 13200 19616 13252
rect 19668 13200 19674 13252
rect 19721 13240 19749 13271
rect 19978 13240 19984 13252
rect 19721 13212 19984 13240
rect 19978 13200 19984 13212
rect 20036 13200 20042 13252
rect 20346 13200 20352 13252
rect 20404 13240 20410 13252
rect 20824 13240 20852 13271
rect 20404 13212 20852 13240
rect 22066 13240 22094 13280
rect 22462 13268 22468 13320
rect 22520 13308 22526 13320
rect 22741 13311 22799 13317
rect 22741 13308 22753 13311
rect 22520 13280 22753 13308
rect 22520 13268 22526 13280
rect 22741 13277 22753 13280
rect 22787 13277 22799 13311
rect 22741 13271 22799 13277
rect 22922 13240 22928 13252
rect 22066 13212 22928 13240
rect 20404 13200 20410 13212
rect 22922 13200 22928 13212
rect 22980 13200 22986 13252
rect 23017 13243 23075 13249
rect 23017 13209 23029 13243
rect 23063 13240 23075 13243
rect 23106 13240 23112 13252
rect 23063 13212 23112 13240
rect 23063 13209 23075 13212
rect 23017 13203 23075 13209
rect 23106 13200 23112 13212
rect 23164 13200 23170 13252
rect 21821 13175 21879 13181
rect 21821 13172 21833 13175
rect 19306 13144 21833 13172
rect 21821 13141 21833 13144
rect 21867 13172 21879 13175
rect 22646 13172 22652 13184
rect 21867 13144 22652 13172
rect 21867 13141 21879 13144
rect 21821 13135 21879 13141
rect 22646 13132 22652 13144
rect 22704 13132 22710 13184
rect 1104 13082 23987 13104
rect 1104 13030 6630 13082
rect 6682 13030 6694 13082
rect 6746 13030 6758 13082
rect 6810 13030 6822 13082
rect 6874 13030 6886 13082
rect 6938 13030 12311 13082
rect 12363 13030 12375 13082
rect 12427 13030 12439 13082
rect 12491 13030 12503 13082
rect 12555 13030 12567 13082
rect 12619 13030 17992 13082
rect 18044 13030 18056 13082
rect 18108 13030 18120 13082
rect 18172 13030 18184 13082
rect 18236 13030 18248 13082
rect 18300 13030 23673 13082
rect 23725 13030 23737 13082
rect 23789 13030 23801 13082
rect 23853 13030 23865 13082
rect 23917 13030 23929 13082
rect 23981 13030 23987 13082
rect 1104 13008 23987 13030
rect 2038 12928 2044 12980
rect 2096 12968 2102 12980
rect 3322 12971 3380 12977
rect 3322 12968 3334 12971
rect 2096 12940 3334 12968
rect 2096 12928 2102 12940
rect 3322 12937 3334 12940
rect 3368 12937 3380 12971
rect 3322 12931 3380 12937
rect 4183 12971 4241 12977
rect 4183 12937 4195 12971
rect 4229 12968 4241 12971
rect 4338 12968 4344 12980
rect 4229 12940 4344 12968
rect 4229 12937 4241 12940
rect 4183 12931 4241 12937
rect 4338 12928 4344 12940
rect 4396 12928 4402 12980
rect 6546 12928 6552 12980
rect 6604 12968 6610 12980
rect 7834 12968 7840 12980
rect 6604 12940 7840 12968
rect 6604 12928 6610 12940
rect 7834 12928 7840 12940
rect 7892 12928 7898 12980
rect 8205 12971 8263 12977
rect 8205 12937 8217 12971
rect 8251 12968 8263 12971
rect 9214 12968 9220 12980
rect 8251 12940 9220 12968
rect 8251 12937 8263 12940
rect 8205 12931 8263 12937
rect 9214 12928 9220 12940
rect 9272 12928 9278 12980
rect 11882 12928 11888 12980
rect 11940 12968 11946 12980
rect 17678 12968 17684 12980
rect 11940 12940 12296 12968
rect 11940 12928 11946 12940
rect 2590 12900 2596 12912
rect 2551 12872 2596 12900
rect 2590 12860 2596 12872
rect 2648 12860 2654 12912
rect 2774 12860 2780 12912
rect 2832 12900 2838 12912
rect 3421 12903 3479 12909
rect 3421 12900 3433 12903
rect 2832 12872 3433 12900
rect 2832 12860 2838 12872
rect 3421 12869 3433 12872
rect 3467 12869 3479 12903
rect 3970 12900 3976 12912
rect 3931 12872 3976 12900
rect 3421 12863 3479 12869
rect 3970 12860 3976 12872
rect 4028 12860 4034 12912
rect 4982 12900 4988 12912
rect 4080 12872 4988 12900
rect 2608 12696 2636 12860
rect 2682 12792 2688 12844
rect 2740 12832 2746 12844
rect 3145 12835 3203 12841
rect 3145 12832 3157 12835
rect 2740 12804 3157 12832
rect 2740 12792 2746 12804
rect 3145 12801 3157 12804
rect 3191 12801 3203 12835
rect 3145 12795 3203 12801
rect 3237 12835 3295 12841
rect 3237 12801 3249 12835
rect 3283 12832 3295 12835
rect 3326 12832 3332 12844
rect 3283 12804 3332 12832
rect 3283 12801 3295 12804
rect 3237 12795 3295 12801
rect 3326 12792 3332 12804
rect 3384 12832 3390 12844
rect 4080 12832 4108 12872
rect 4982 12860 4988 12872
rect 5040 12860 5046 12912
rect 6564 12900 6592 12928
rect 5088 12872 6592 12900
rect 3384 12804 4108 12832
rect 3384 12792 3390 12804
rect 4246 12792 4252 12844
rect 4304 12832 4310 12844
rect 5088 12832 5116 12872
rect 7742 12860 7748 12912
rect 7800 12900 7806 12912
rect 8662 12900 8668 12912
rect 7800 12872 8668 12900
rect 7800 12860 7806 12872
rect 8662 12860 8668 12872
rect 8720 12860 8726 12912
rect 10134 12860 10140 12912
rect 10192 12900 10198 12912
rect 10192 12872 10548 12900
rect 10192 12860 10198 12872
rect 5258 12832 5264 12844
rect 4304 12804 5116 12832
rect 5219 12804 5264 12832
rect 4304 12792 4310 12804
rect 5258 12792 5264 12804
rect 5316 12792 5322 12844
rect 5353 12835 5411 12841
rect 5353 12801 5365 12835
rect 5399 12832 5411 12835
rect 5626 12832 5632 12844
rect 5399 12804 5632 12832
rect 5399 12801 5411 12804
rect 5353 12795 5411 12801
rect 5626 12792 5632 12804
rect 5684 12792 5690 12844
rect 5994 12792 6000 12844
rect 6052 12832 6058 12844
rect 7285 12835 7343 12841
rect 7285 12832 7297 12835
rect 6052 12804 7297 12832
rect 6052 12792 6058 12804
rect 7285 12801 7297 12804
rect 7331 12801 7343 12835
rect 7285 12795 7343 12801
rect 7377 12835 7435 12841
rect 7377 12801 7389 12835
rect 7423 12801 7435 12835
rect 7558 12832 7564 12844
rect 7519 12804 7564 12832
rect 7377 12795 7435 12801
rect 7392 12764 7420 12795
rect 7558 12792 7564 12804
rect 7616 12792 7622 12844
rect 7653 12835 7711 12841
rect 7653 12801 7665 12835
rect 7699 12832 7711 12835
rect 7760 12832 7788 12860
rect 8110 12832 8116 12844
rect 7699 12804 7788 12832
rect 8071 12804 8116 12832
rect 7699 12801 7711 12804
rect 7653 12795 7711 12801
rect 8110 12792 8116 12804
rect 8168 12792 8174 12844
rect 8294 12832 8300 12844
rect 8255 12804 8300 12832
rect 8294 12792 8300 12804
rect 8352 12792 8358 12844
rect 8938 12832 8944 12844
rect 8899 12804 8944 12832
rect 8938 12792 8944 12804
rect 8996 12792 9002 12844
rect 9030 12792 9036 12844
rect 9088 12832 9094 12844
rect 9306 12832 9312 12844
rect 9088 12804 9133 12832
rect 9219 12804 9312 12832
rect 9088 12792 9094 12804
rect 9306 12792 9312 12804
rect 9364 12792 9370 12844
rect 10410 12832 10416 12844
rect 10371 12804 10416 12832
rect 10410 12792 10416 12804
rect 10468 12792 10474 12844
rect 10520 12841 10548 12872
rect 11698 12860 11704 12912
rect 11756 12900 11762 12912
rect 12066 12900 12072 12912
rect 11756 12872 12072 12900
rect 11756 12860 11762 12872
rect 10505 12835 10563 12841
rect 10505 12801 10517 12835
rect 10551 12801 10563 12835
rect 10505 12795 10563 12801
rect 10689 12835 10747 12841
rect 10689 12801 10701 12835
rect 10735 12832 10747 12835
rect 11790 12832 11796 12844
rect 10735 12804 11796 12832
rect 10735 12801 10747 12804
rect 10689 12795 10747 12801
rect 11790 12792 11796 12804
rect 11848 12792 11854 12844
rect 11900 12841 11928 12872
rect 12066 12860 12072 12872
rect 12124 12860 12130 12912
rect 11885 12835 11943 12841
rect 11885 12801 11897 12835
rect 11931 12801 11943 12835
rect 11885 12795 11943 12801
rect 11974 12792 11980 12844
rect 12032 12832 12038 12844
rect 12161 12835 12219 12841
rect 12161 12832 12173 12835
rect 12032 12804 12173 12832
rect 12032 12792 12038 12804
rect 12161 12801 12173 12804
rect 12207 12801 12219 12835
rect 12268 12832 12296 12940
rect 17352 12940 17684 12968
rect 12529 12903 12587 12909
rect 12529 12869 12541 12903
rect 12575 12900 12587 12903
rect 12710 12900 12716 12912
rect 12575 12872 12716 12900
rect 12575 12869 12587 12872
rect 12529 12863 12587 12869
rect 12710 12860 12716 12872
rect 12768 12860 12774 12912
rect 13354 12860 13360 12912
rect 13412 12900 13418 12912
rect 14645 12903 14703 12909
rect 13412 12872 14044 12900
rect 13412 12860 13418 12872
rect 12345 12835 12403 12841
rect 12345 12832 12357 12835
rect 12268 12804 12357 12832
rect 12161 12795 12219 12801
rect 12345 12801 12357 12804
rect 12391 12801 12403 12835
rect 12345 12795 12403 12801
rect 12894 12792 12900 12844
rect 12952 12832 12958 12844
rect 13170 12832 13176 12844
rect 12952 12804 13176 12832
rect 12952 12792 12958 12804
rect 13170 12792 13176 12804
rect 13228 12832 13234 12844
rect 14016 12841 14044 12872
rect 14645 12869 14657 12903
rect 14691 12900 14703 12903
rect 14734 12900 14740 12912
rect 14691 12872 14740 12900
rect 14691 12869 14703 12872
rect 14645 12863 14703 12869
rect 14734 12860 14740 12872
rect 14792 12860 14798 12912
rect 15289 12903 15347 12909
rect 15289 12869 15301 12903
rect 15335 12900 15347 12903
rect 15654 12900 15660 12912
rect 15335 12872 15660 12900
rect 15335 12869 15347 12872
rect 15289 12863 15347 12869
rect 15654 12860 15660 12872
rect 15712 12860 15718 12912
rect 17218 12900 17224 12912
rect 17179 12872 17224 12900
rect 17218 12860 17224 12872
rect 17276 12860 17282 12912
rect 13633 12835 13691 12841
rect 13633 12832 13645 12835
rect 13228 12804 13645 12832
rect 13228 12792 13234 12804
rect 13633 12801 13645 12804
rect 13679 12801 13691 12835
rect 13633 12795 13691 12801
rect 14001 12835 14059 12841
rect 14001 12801 14013 12835
rect 14047 12801 14059 12835
rect 14001 12795 14059 12801
rect 15841 12835 15899 12841
rect 15841 12801 15853 12835
rect 15887 12832 15899 12835
rect 16853 12835 16911 12841
rect 16853 12832 16865 12835
rect 15887 12804 16865 12832
rect 15887 12801 15899 12804
rect 15841 12795 15899 12801
rect 16853 12801 16865 12804
rect 16899 12801 16911 12835
rect 16853 12795 16911 12801
rect 4080 12736 7328 12764
rect 7392 12736 7604 12764
rect 3418 12696 3424 12708
rect 2608 12668 3424 12696
rect 3418 12656 3424 12668
rect 3476 12656 3482 12708
rect 1765 12631 1823 12637
rect 1765 12597 1777 12631
rect 1811 12628 1823 12631
rect 1946 12628 1952 12640
rect 1811 12600 1952 12628
rect 1811 12597 1823 12600
rect 1765 12591 1823 12597
rect 1946 12588 1952 12600
rect 2004 12588 2010 12640
rect 2501 12631 2559 12637
rect 2501 12597 2513 12631
rect 2547 12628 2559 12631
rect 2590 12628 2596 12640
rect 2547 12600 2596 12628
rect 2547 12597 2559 12600
rect 2501 12591 2559 12597
rect 2590 12588 2596 12600
rect 2648 12628 2654 12640
rect 4080 12628 4108 12736
rect 4341 12699 4399 12705
rect 4341 12665 4353 12699
rect 4387 12696 4399 12699
rect 5442 12696 5448 12708
rect 4387 12668 5448 12696
rect 4387 12665 4399 12668
rect 4341 12659 4399 12665
rect 5442 12656 5448 12668
rect 5500 12656 5506 12708
rect 7098 12656 7104 12708
rect 7156 12696 7162 12708
rect 7300 12696 7328 12736
rect 7576 12696 7604 12736
rect 8846 12724 8852 12776
rect 8904 12764 8910 12776
rect 9217 12767 9275 12773
rect 9217 12764 9229 12767
rect 8904 12736 9229 12764
rect 8904 12724 8910 12736
rect 9217 12733 9229 12736
rect 9263 12733 9275 12767
rect 9217 12727 9275 12733
rect 7834 12696 7840 12708
rect 7156 12668 7201 12696
rect 7300 12668 7512 12696
rect 7576 12668 7840 12696
rect 7156 12656 7162 12668
rect 2648 12600 4108 12628
rect 4157 12631 4215 12637
rect 2648 12588 2654 12600
rect 4157 12597 4169 12631
rect 4203 12628 4215 12631
rect 4246 12628 4252 12640
rect 4203 12600 4252 12628
rect 4203 12597 4215 12600
rect 4157 12591 4215 12597
rect 4246 12588 4252 12600
rect 4304 12588 4310 12640
rect 5718 12588 5724 12640
rect 5776 12628 5782 12640
rect 6549 12631 6607 12637
rect 6549 12628 6561 12631
rect 5776 12600 6561 12628
rect 5776 12588 5782 12600
rect 6549 12597 6561 12600
rect 6595 12628 6607 12631
rect 7006 12628 7012 12640
rect 6595 12600 7012 12628
rect 6595 12597 6607 12600
rect 6549 12591 6607 12597
rect 7006 12588 7012 12600
rect 7064 12588 7070 12640
rect 7484 12628 7512 12668
rect 7834 12656 7840 12668
rect 7892 12656 7898 12708
rect 9324 12696 9352 12792
rect 11146 12764 11152 12776
rect 11107 12736 11152 12764
rect 11146 12724 11152 12736
rect 11204 12724 11210 12776
rect 13722 12764 13728 12776
rect 13683 12736 13728 12764
rect 13722 12724 13728 12736
rect 13780 12724 13786 12776
rect 14090 12724 14096 12776
rect 14148 12764 14154 12776
rect 14185 12767 14243 12773
rect 14185 12764 14197 12767
rect 14148 12736 14197 12764
rect 14148 12724 14154 12736
rect 14185 12733 14197 12736
rect 14231 12764 14243 12767
rect 15654 12764 15660 12776
rect 14231 12736 15660 12764
rect 14231 12733 14243 12736
rect 14185 12727 14243 12733
rect 15654 12724 15660 12736
rect 15712 12724 15718 12776
rect 15930 12764 15936 12776
rect 15891 12736 15936 12764
rect 15930 12724 15936 12736
rect 15988 12724 15994 12776
rect 16025 12767 16083 12773
rect 16025 12733 16037 12767
rect 16071 12733 16083 12767
rect 16025 12727 16083 12733
rect 8036 12668 9352 12696
rect 16040 12696 16068 12727
rect 16114 12724 16120 12776
rect 16172 12764 16178 12776
rect 16868 12764 16896 12795
rect 16942 12792 16948 12844
rect 17000 12832 17006 12844
rect 17126 12832 17132 12844
rect 17000 12804 17045 12832
rect 17087 12804 17132 12832
rect 17000 12792 17006 12804
rect 17126 12792 17132 12804
rect 17184 12792 17190 12844
rect 17352 12841 17380 12940
rect 17678 12928 17684 12940
rect 17736 12928 17742 12980
rect 19334 12928 19340 12980
rect 19392 12968 19398 12980
rect 19429 12971 19487 12977
rect 19429 12968 19441 12971
rect 19392 12940 19441 12968
rect 19392 12928 19398 12940
rect 19429 12937 19441 12940
rect 19475 12937 19487 12971
rect 19978 12968 19984 12980
rect 19429 12931 19487 12937
rect 19628 12940 19984 12968
rect 17586 12860 17592 12912
rect 17644 12900 17650 12912
rect 19628 12900 19656 12940
rect 19978 12928 19984 12940
rect 20036 12928 20042 12980
rect 20254 12928 20260 12980
rect 20312 12968 20318 12980
rect 22278 12968 22284 12980
rect 20312 12940 21864 12968
rect 22239 12940 22284 12968
rect 20312 12928 20318 12940
rect 21358 12900 21364 12912
rect 17644 12872 19656 12900
rect 19720 12872 21364 12900
rect 17644 12860 17650 12872
rect 17337 12835 17395 12841
rect 17337 12801 17349 12835
rect 17383 12801 17395 12835
rect 17337 12795 17395 12801
rect 17862 12792 17868 12844
rect 17920 12832 17926 12844
rect 19334 12832 19340 12844
rect 17920 12804 19340 12832
rect 17920 12792 17926 12804
rect 19334 12792 19340 12804
rect 19392 12832 19398 12844
rect 19720 12841 19748 12872
rect 21358 12860 21364 12872
rect 21416 12860 21422 12912
rect 21453 12903 21511 12909
rect 21453 12869 21465 12903
rect 21499 12900 21511 12903
rect 21726 12900 21732 12912
rect 21499 12872 21732 12900
rect 21499 12869 21511 12872
rect 21453 12863 21511 12869
rect 19613 12835 19671 12841
rect 19613 12832 19625 12835
rect 19392 12804 19625 12832
rect 19392 12792 19398 12804
rect 19613 12801 19625 12804
rect 19659 12801 19671 12835
rect 19613 12795 19671 12801
rect 19705 12835 19763 12841
rect 19705 12801 19717 12835
rect 19751 12801 19763 12835
rect 19886 12832 19892 12844
rect 19847 12804 19892 12832
rect 19705 12795 19763 12801
rect 19886 12792 19892 12804
rect 19944 12792 19950 12844
rect 20073 12835 20131 12841
rect 20073 12801 20085 12835
rect 20119 12832 20131 12835
rect 20254 12832 20260 12844
rect 20119 12804 20260 12832
rect 20119 12801 20131 12804
rect 20073 12795 20131 12801
rect 20254 12792 20260 12804
rect 20312 12792 20318 12844
rect 20346 12792 20352 12844
rect 20404 12832 20410 12844
rect 20622 12832 20628 12844
rect 20404 12804 20628 12832
rect 20404 12792 20410 12804
rect 20622 12792 20628 12804
rect 20680 12792 20686 12844
rect 20714 12792 20720 12844
rect 20772 12832 20778 12844
rect 21085 12835 21143 12841
rect 21085 12832 21097 12835
rect 20772 12804 21097 12832
rect 20772 12792 20778 12804
rect 21085 12801 21097 12804
rect 21131 12801 21143 12835
rect 21085 12795 21143 12801
rect 21266 12792 21272 12844
rect 21324 12832 21330 12844
rect 21468 12832 21496 12863
rect 21726 12860 21732 12872
rect 21784 12860 21790 12912
rect 21324 12804 21496 12832
rect 21836 12832 21864 12940
rect 22278 12928 22284 12940
rect 22336 12928 22342 12980
rect 22738 12860 22744 12912
rect 22796 12909 22802 12912
rect 22796 12903 22825 12909
rect 22813 12869 22825 12903
rect 22796 12863 22825 12869
rect 22796 12860 22802 12863
rect 22465 12835 22523 12841
rect 22465 12832 22477 12835
rect 21836 12804 22477 12832
rect 21324 12792 21330 12804
rect 22465 12801 22477 12804
rect 22511 12801 22523 12835
rect 22465 12795 22523 12801
rect 22557 12835 22615 12841
rect 22557 12801 22569 12835
rect 22603 12801 22615 12835
rect 22557 12795 22615 12801
rect 22094 12764 22100 12776
rect 16172 12736 16217 12764
rect 16868 12736 22100 12764
rect 16172 12724 16178 12736
rect 22094 12724 22100 12736
rect 22152 12724 22158 12776
rect 16666 12696 16672 12708
rect 16040 12668 16672 12696
rect 8036 12640 8064 12668
rect 16666 12656 16672 12668
rect 16724 12696 16730 12708
rect 18049 12699 18107 12705
rect 16724 12668 17080 12696
rect 16724 12656 16730 12668
rect 8018 12628 8024 12640
rect 7484 12600 8024 12628
rect 8018 12588 8024 12600
rect 8076 12588 8082 12640
rect 8754 12628 8760 12640
rect 8715 12600 8760 12628
rect 8754 12588 8760 12600
rect 8812 12588 8818 12640
rect 11790 12588 11796 12640
rect 11848 12628 11854 12640
rect 12526 12628 12532 12640
rect 11848 12600 12532 12628
rect 11848 12588 11854 12600
rect 12526 12588 12532 12600
rect 12584 12588 12590 12640
rect 16301 12631 16359 12637
rect 16301 12597 16313 12631
rect 16347 12628 16359 12631
rect 16850 12628 16856 12640
rect 16347 12600 16856 12628
rect 16347 12597 16359 12600
rect 16301 12591 16359 12597
rect 16850 12588 16856 12600
rect 16908 12588 16914 12640
rect 17052 12628 17080 12668
rect 17420 12668 17724 12696
rect 17420 12628 17448 12668
rect 17052 12600 17448 12628
rect 17497 12631 17555 12637
rect 17497 12597 17509 12631
rect 17543 12628 17555 12631
rect 17586 12628 17592 12640
rect 17543 12600 17592 12628
rect 17543 12597 17555 12600
rect 17497 12591 17555 12597
rect 17586 12588 17592 12600
rect 17644 12588 17650 12640
rect 17696 12628 17724 12668
rect 18049 12665 18061 12699
rect 18095 12696 18107 12699
rect 18506 12696 18512 12708
rect 18095 12668 18512 12696
rect 18095 12665 18107 12668
rect 18049 12659 18107 12665
rect 18506 12656 18512 12668
rect 18564 12656 18570 12708
rect 19794 12656 19800 12708
rect 19852 12696 19858 12708
rect 19852 12668 19897 12696
rect 19852 12656 19858 12668
rect 18598 12628 18604 12640
rect 17696 12600 18604 12628
rect 18598 12588 18604 12600
rect 18656 12588 18662 12640
rect 19334 12588 19340 12640
rect 19392 12628 19398 12640
rect 20622 12628 20628 12640
rect 19392 12600 20628 12628
rect 19392 12588 19398 12600
rect 20622 12588 20628 12600
rect 20680 12588 20686 12640
rect 22480 12628 22508 12795
rect 22572 12696 22600 12795
rect 22646 12792 22652 12844
rect 22704 12832 22710 12844
rect 22922 12832 22928 12844
rect 22704 12804 22749 12832
rect 22883 12804 22928 12832
rect 22704 12792 22710 12804
rect 22922 12792 22928 12804
rect 22980 12792 22986 12844
rect 23014 12696 23020 12708
rect 22572 12668 23020 12696
rect 23014 12656 23020 12668
rect 23072 12656 23078 12708
rect 22738 12628 22744 12640
rect 22480 12600 22744 12628
rect 22738 12588 22744 12600
rect 22796 12588 22802 12640
rect 1104 12538 23828 12560
rect 1104 12486 3790 12538
rect 3842 12486 3854 12538
rect 3906 12486 3918 12538
rect 3970 12486 3982 12538
rect 4034 12486 4046 12538
rect 4098 12486 9471 12538
rect 9523 12486 9535 12538
rect 9587 12486 9599 12538
rect 9651 12486 9663 12538
rect 9715 12486 9727 12538
rect 9779 12486 15152 12538
rect 15204 12486 15216 12538
rect 15268 12486 15280 12538
rect 15332 12486 15344 12538
rect 15396 12486 15408 12538
rect 15460 12486 20833 12538
rect 20885 12486 20897 12538
rect 20949 12486 20961 12538
rect 21013 12486 21025 12538
rect 21077 12486 21089 12538
rect 21141 12486 23828 12538
rect 1104 12464 23828 12486
rect 1578 12384 1584 12436
rect 1636 12424 1642 12436
rect 4065 12427 4123 12433
rect 1636 12396 4016 12424
rect 1636 12384 1642 12396
rect 2038 12316 2044 12368
rect 2096 12316 2102 12368
rect 3988 12356 4016 12396
rect 4065 12393 4077 12427
rect 4111 12424 4123 12427
rect 4154 12424 4160 12436
rect 4111 12396 4160 12424
rect 4111 12393 4123 12396
rect 4065 12387 4123 12393
rect 4154 12384 4160 12396
rect 4212 12384 4218 12436
rect 5626 12384 5632 12436
rect 5684 12424 5690 12436
rect 5997 12427 6055 12433
rect 5997 12424 6009 12427
rect 5684 12396 6009 12424
rect 5684 12384 5690 12396
rect 5997 12393 6009 12396
rect 6043 12424 6055 12427
rect 7190 12424 7196 12436
rect 6043 12396 7196 12424
rect 6043 12393 6055 12396
rect 5997 12387 6055 12393
rect 7190 12384 7196 12396
rect 7248 12384 7254 12436
rect 7374 12424 7380 12436
rect 7335 12396 7380 12424
rect 7374 12384 7380 12396
rect 7432 12384 7438 12436
rect 7558 12384 7564 12436
rect 7616 12424 7622 12436
rect 8113 12427 8171 12433
rect 8113 12424 8125 12427
rect 7616 12396 8125 12424
rect 7616 12384 7622 12396
rect 8113 12393 8125 12396
rect 8159 12393 8171 12427
rect 8113 12387 8171 12393
rect 10686 12384 10692 12436
rect 10744 12424 10750 12436
rect 10962 12424 10968 12436
rect 10744 12396 10968 12424
rect 10744 12384 10750 12396
rect 10962 12384 10968 12396
rect 11020 12424 11026 12436
rect 11517 12427 11575 12433
rect 11517 12424 11529 12427
rect 11020 12396 11529 12424
rect 11020 12384 11026 12396
rect 11517 12393 11529 12396
rect 11563 12393 11575 12427
rect 11974 12424 11980 12436
rect 11935 12396 11980 12424
rect 11517 12387 11575 12393
rect 11974 12384 11980 12396
rect 12032 12384 12038 12436
rect 12158 12384 12164 12436
rect 12216 12424 12222 12436
rect 13633 12427 13691 12433
rect 13633 12424 13645 12427
rect 12216 12396 13645 12424
rect 12216 12384 12222 12396
rect 13633 12393 13645 12396
rect 13679 12393 13691 12427
rect 13633 12387 13691 12393
rect 15381 12427 15439 12433
rect 15381 12393 15393 12427
rect 15427 12424 15439 12427
rect 15470 12424 15476 12436
rect 15427 12396 15476 12424
rect 15427 12393 15439 12396
rect 15381 12387 15439 12393
rect 15470 12384 15476 12396
rect 15528 12384 15534 12436
rect 16298 12424 16304 12436
rect 16259 12396 16304 12424
rect 16298 12384 16304 12396
rect 16356 12384 16362 12436
rect 18966 12384 18972 12436
rect 19024 12424 19030 12436
rect 19150 12424 19156 12436
rect 19024 12396 19156 12424
rect 19024 12384 19030 12396
rect 19150 12384 19156 12396
rect 19208 12424 19214 12436
rect 19429 12427 19487 12433
rect 19429 12424 19441 12427
rect 19208 12396 19441 12424
rect 19208 12384 19214 12396
rect 19429 12393 19441 12396
rect 19475 12393 19487 12427
rect 19429 12387 19487 12393
rect 20346 12384 20352 12436
rect 20404 12424 20410 12436
rect 20717 12427 20775 12433
rect 20717 12424 20729 12427
rect 20404 12396 20729 12424
rect 20404 12384 20410 12396
rect 20717 12393 20729 12396
rect 20763 12393 20775 12427
rect 20717 12387 20775 12393
rect 6733 12359 6791 12365
rect 6733 12356 6745 12359
rect 2424 12328 3188 12356
rect 3988 12328 6745 12356
rect 2056 12288 2084 12316
rect 2225 12291 2283 12297
rect 2225 12288 2237 12291
rect 2056 12260 2237 12288
rect 2225 12257 2237 12260
rect 2271 12257 2283 12291
rect 2225 12251 2283 12257
rect 2041 12223 2099 12229
rect 2041 12189 2053 12223
rect 2087 12220 2099 12223
rect 2130 12220 2136 12232
rect 2087 12192 2136 12220
rect 2087 12189 2099 12192
rect 2041 12183 2099 12189
rect 2130 12180 2136 12192
rect 2188 12220 2194 12232
rect 2314 12220 2320 12232
rect 2188 12192 2320 12220
rect 2188 12180 2194 12192
rect 2314 12180 2320 12192
rect 2372 12180 2378 12232
rect 2424 12229 2452 12328
rect 2590 12248 2596 12300
rect 2648 12288 2654 12300
rect 2648 12260 2774 12288
rect 2648 12248 2654 12260
rect 2409 12223 2467 12229
rect 2409 12189 2421 12223
rect 2455 12189 2467 12223
rect 2608 12220 2636 12248
rect 2409 12183 2467 12189
rect 2516 12192 2636 12220
rect 2746 12220 2774 12260
rect 3160 12229 3188 12328
rect 6733 12325 6745 12328
rect 6779 12325 6791 12359
rect 6733 12319 6791 12325
rect 7282 12316 7288 12368
rect 7340 12356 7346 12368
rect 8202 12356 8208 12368
rect 7340 12328 8208 12356
rect 7340 12316 7346 12328
rect 8202 12316 8208 12328
rect 8260 12316 8266 12368
rect 12526 12356 12532 12368
rect 12487 12328 12532 12356
rect 12526 12316 12532 12328
rect 12584 12316 12590 12368
rect 13170 12316 13176 12368
rect 13228 12356 13234 12368
rect 15562 12356 15568 12368
rect 13228 12328 15568 12356
rect 13228 12316 13234 12328
rect 15562 12316 15568 12328
rect 15620 12316 15626 12368
rect 16485 12359 16543 12365
rect 16485 12325 16497 12359
rect 16531 12325 16543 12359
rect 16485 12319 16543 12325
rect 21085 12359 21143 12365
rect 21085 12325 21097 12359
rect 21131 12356 21143 12359
rect 21266 12356 21272 12368
rect 21131 12328 21272 12356
rect 21131 12325 21143 12328
rect 21085 12319 21143 12325
rect 6270 12248 6276 12300
rect 6328 12288 6334 12300
rect 8294 12288 8300 12300
rect 6328 12260 6776 12288
rect 6328 12248 6334 12260
rect 2961 12223 3019 12229
rect 2961 12220 2973 12223
rect 2746 12192 2973 12220
rect 1946 12112 1952 12164
rect 2004 12152 2010 12164
rect 2424 12152 2452 12183
rect 2004 12124 2452 12152
rect 2004 12112 2010 12124
rect 1670 12044 1676 12096
rect 1728 12084 1734 12096
rect 2133 12087 2191 12093
rect 2133 12084 2145 12087
rect 1728 12056 2145 12084
rect 1728 12044 1734 12056
rect 2133 12053 2145 12056
rect 2179 12053 2191 12087
rect 2133 12047 2191 12053
rect 2222 12044 2228 12096
rect 2280 12084 2286 12096
rect 2317 12087 2375 12093
rect 2317 12084 2329 12087
rect 2280 12056 2329 12084
rect 2280 12044 2286 12056
rect 2317 12053 2329 12056
rect 2363 12084 2375 12087
rect 2516 12084 2544 12192
rect 2961 12189 2973 12192
rect 3007 12189 3019 12223
rect 2961 12183 3019 12189
rect 3145 12223 3203 12229
rect 3145 12189 3157 12223
rect 3191 12189 3203 12223
rect 3145 12183 3203 12189
rect 3694 12180 3700 12232
rect 3752 12220 3758 12232
rect 3973 12223 4031 12229
rect 3973 12220 3985 12223
rect 3752 12192 3985 12220
rect 3752 12180 3758 12192
rect 3973 12189 3985 12192
rect 4019 12189 4031 12223
rect 3973 12183 4031 12189
rect 4154 12180 4160 12232
rect 4212 12222 4218 12232
rect 4212 12220 4226 12222
rect 6546 12220 6552 12232
rect 4212 12192 5028 12220
rect 6507 12192 6552 12220
rect 4212 12180 4218 12192
rect 2869 12155 2927 12161
rect 2869 12121 2881 12155
rect 2915 12152 2927 12155
rect 3326 12152 3332 12164
rect 2915 12124 3332 12152
rect 2915 12121 2927 12124
rect 2869 12115 2927 12121
rect 3326 12112 3332 12124
rect 3384 12112 3390 12164
rect 5000 12152 5028 12192
rect 6546 12180 6552 12192
rect 6604 12180 6610 12232
rect 6748 12229 6776 12260
rect 6840 12260 8300 12288
rect 6733 12223 6791 12229
rect 6733 12189 6745 12223
rect 6779 12189 6791 12223
rect 6733 12183 6791 12189
rect 6840 12152 6868 12260
rect 8294 12248 8300 12260
rect 8352 12288 8358 12300
rect 8352 12260 10088 12288
rect 8352 12248 8358 12260
rect 7190 12220 7196 12232
rect 7151 12192 7196 12220
rect 7190 12180 7196 12192
rect 7248 12180 7254 12232
rect 7377 12223 7435 12229
rect 7377 12222 7389 12223
rect 7300 12194 7389 12222
rect 5000 12124 6868 12152
rect 7006 12112 7012 12164
rect 7064 12152 7070 12164
rect 7300 12152 7328 12194
rect 7377 12189 7389 12194
rect 7423 12189 7435 12223
rect 7377 12183 7435 12189
rect 8202 12180 8208 12232
rect 8260 12220 8266 12232
rect 10060 12229 10088 12260
rect 10778 12248 10784 12300
rect 10836 12288 10842 12300
rect 11793 12291 11851 12297
rect 11793 12288 11805 12291
rect 10836 12260 11805 12288
rect 10836 12248 10842 12260
rect 11793 12257 11805 12260
rect 11839 12257 11851 12291
rect 12066 12288 12072 12300
rect 11793 12251 11851 12257
rect 11900 12260 12072 12288
rect 8389 12223 8447 12229
rect 8389 12220 8401 12223
rect 8260 12192 8401 12220
rect 8260 12180 8266 12192
rect 8389 12189 8401 12192
rect 8435 12189 8447 12223
rect 8389 12183 8447 12189
rect 10045 12223 10103 12229
rect 10045 12189 10057 12223
rect 10091 12189 10103 12223
rect 10045 12183 10103 12189
rect 10413 12223 10471 12229
rect 10413 12189 10425 12223
rect 10459 12220 10471 12223
rect 10502 12220 10508 12232
rect 10459 12192 10508 12220
rect 10459 12189 10471 12192
rect 10413 12183 10471 12189
rect 10502 12180 10508 12192
rect 10560 12180 10566 12232
rect 10686 12220 10692 12232
rect 10647 12192 10692 12220
rect 10686 12180 10692 12192
rect 10744 12180 10750 12232
rect 11701 12223 11759 12229
rect 11701 12189 11713 12223
rect 11747 12220 11759 12223
rect 11900 12220 11928 12260
rect 12066 12248 12072 12260
rect 12124 12248 12130 12300
rect 12544 12288 12572 12316
rect 13262 12288 13268 12300
rect 12544 12260 13268 12288
rect 13262 12248 13268 12260
rect 13320 12248 13326 12300
rect 14366 12288 14372 12300
rect 13556 12260 14372 12288
rect 13556 12229 13584 12260
rect 14366 12248 14372 12260
rect 14424 12248 14430 12300
rect 15010 12288 15016 12300
rect 14752 12260 15016 12288
rect 14752 12232 14780 12260
rect 15010 12248 15016 12260
rect 15068 12248 15074 12300
rect 16500 12288 16528 12319
rect 21266 12316 21272 12328
rect 21324 12316 21330 12368
rect 21634 12316 21640 12368
rect 21692 12316 21698 12368
rect 22830 12356 22836 12368
rect 21744 12328 22836 12356
rect 16500 12260 17632 12288
rect 11747 12192 11928 12220
rect 13541 12223 13599 12229
rect 11747 12189 11759 12192
rect 11701 12183 11759 12189
rect 13541 12189 13553 12223
rect 13587 12189 13599 12223
rect 13541 12183 13599 12189
rect 13725 12223 13783 12229
rect 13725 12189 13737 12223
rect 13771 12189 13783 12223
rect 13725 12183 13783 12189
rect 7064 12124 7328 12152
rect 7064 12112 7070 12124
rect 7834 12112 7840 12164
rect 7892 12152 7898 12164
rect 8113 12155 8171 12161
rect 8113 12152 8125 12155
rect 7892 12124 8125 12152
rect 7892 12112 7898 12124
rect 8113 12121 8125 12124
rect 8159 12152 8171 12155
rect 9217 12155 9275 12161
rect 9217 12152 9229 12155
rect 8159 12124 9229 12152
rect 8159 12121 8171 12124
rect 8113 12115 8171 12121
rect 9217 12121 9229 12124
rect 9263 12152 9275 12155
rect 10704 12152 10732 12180
rect 9263 12124 10732 12152
rect 9263 12121 9275 12124
rect 9217 12115 9275 12121
rect 11882 12112 11888 12164
rect 11940 12152 11946 12164
rect 11977 12155 12035 12161
rect 11977 12152 11989 12155
rect 11940 12124 11989 12152
rect 11940 12112 11946 12124
rect 11977 12121 11989 12124
rect 12023 12121 12035 12155
rect 13740 12152 13768 12183
rect 13998 12180 14004 12232
rect 14056 12220 14062 12232
rect 14274 12220 14280 12232
rect 14056 12192 14280 12220
rect 14056 12180 14062 12192
rect 14274 12180 14280 12192
rect 14332 12180 14338 12232
rect 14461 12223 14519 12229
rect 14461 12189 14473 12223
rect 14507 12220 14519 12223
rect 14734 12220 14740 12232
rect 14507 12192 14740 12220
rect 14507 12189 14519 12192
rect 14461 12183 14519 12189
rect 14734 12180 14740 12192
rect 14792 12180 14798 12232
rect 14829 12223 14887 12229
rect 14829 12189 14841 12223
rect 14875 12220 14887 12223
rect 14875 12192 16804 12220
rect 14875 12189 14887 12192
rect 14829 12183 14887 12189
rect 16022 12152 16028 12164
rect 13740 12124 16028 12152
rect 11977 12115 12035 12121
rect 16022 12112 16028 12124
rect 16080 12112 16086 12164
rect 16114 12112 16120 12164
rect 16172 12152 16178 12164
rect 16776 12152 16804 12192
rect 16850 12180 16856 12232
rect 16908 12220 16914 12232
rect 17604 12229 17632 12260
rect 17954 12248 17960 12300
rect 18012 12288 18018 12300
rect 19702 12288 19708 12300
rect 18012 12260 19708 12288
rect 18012 12248 18018 12260
rect 19702 12248 19708 12260
rect 19760 12248 19766 12300
rect 21652 12288 21680 12316
rect 20732 12260 21680 12288
rect 17497 12223 17555 12229
rect 17497 12220 17509 12223
rect 16908 12192 17509 12220
rect 16908 12180 16914 12192
rect 17497 12189 17509 12192
rect 17543 12189 17555 12223
rect 17497 12183 17555 12189
rect 17589 12223 17647 12229
rect 17589 12189 17601 12223
rect 17635 12189 17647 12223
rect 17589 12183 17647 12189
rect 17678 12180 17684 12232
rect 17736 12220 17742 12232
rect 17862 12220 17868 12232
rect 17736 12192 17781 12220
rect 17823 12192 17868 12220
rect 17736 12180 17742 12192
rect 17862 12180 17868 12192
rect 17920 12180 17926 12232
rect 18414 12180 18420 12232
rect 18472 12220 18478 12232
rect 20732 12229 20760 12260
rect 20717 12223 20775 12229
rect 20717 12220 20729 12223
rect 18472 12192 20729 12220
rect 18472 12180 18478 12192
rect 20717 12189 20729 12192
rect 20763 12189 20775 12223
rect 20717 12183 20775 12189
rect 20806 12180 20812 12232
rect 20864 12220 20870 12232
rect 20864 12192 20909 12220
rect 20864 12180 20870 12192
rect 21634 12180 21640 12232
rect 21692 12220 21698 12232
rect 21744 12229 21772 12328
rect 22830 12316 22836 12328
rect 22888 12316 22894 12368
rect 22278 12288 22284 12300
rect 21836 12260 22284 12288
rect 21836 12229 21864 12260
rect 22278 12248 22284 12260
rect 22336 12288 22342 12300
rect 22922 12288 22928 12300
rect 22336 12260 22928 12288
rect 22336 12248 22342 12260
rect 22922 12248 22928 12260
rect 22980 12248 22986 12300
rect 21729 12223 21787 12229
rect 21729 12220 21741 12223
rect 21692 12192 21741 12220
rect 21692 12180 21698 12192
rect 21729 12189 21741 12192
rect 21775 12189 21787 12223
rect 21729 12183 21787 12189
rect 21821 12223 21879 12229
rect 21821 12189 21833 12223
rect 21867 12189 21879 12223
rect 22002 12220 22008 12232
rect 21963 12192 22008 12220
rect 21821 12183 21879 12189
rect 22002 12180 22008 12192
rect 22060 12180 22066 12232
rect 22097 12223 22155 12229
rect 22097 12189 22109 12223
rect 22143 12220 22155 12223
rect 22186 12220 22192 12232
rect 22143 12192 22192 12220
rect 22143 12189 22155 12192
rect 22097 12183 22155 12189
rect 22186 12180 22192 12192
rect 22244 12180 22250 12232
rect 23109 12223 23167 12229
rect 23109 12189 23121 12223
rect 23155 12220 23167 12223
rect 23198 12220 23204 12232
rect 23155 12192 23204 12220
rect 23155 12189 23167 12192
rect 23109 12183 23167 12189
rect 23198 12180 23204 12192
rect 23256 12180 23262 12232
rect 16942 12152 16948 12164
rect 16172 12124 16712 12152
rect 16776 12124 16948 12152
rect 16172 12112 16178 12124
rect 2363 12056 2544 12084
rect 2363 12053 2375 12056
rect 2317 12047 2375 12053
rect 4338 12044 4344 12096
rect 4396 12084 4402 12096
rect 4617 12087 4675 12093
rect 4617 12084 4629 12087
rect 4396 12056 4629 12084
rect 4396 12044 4402 12056
rect 4617 12053 4629 12056
rect 4663 12053 4675 12087
rect 4617 12047 4675 12053
rect 5902 12044 5908 12096
rect 5960 12084 5966 12096
rect 8297 12087 8355 12093
rect 8297 12084 8309 12087
rect 5960 12056 8309 12084
rect 5960 12044 5966 12056
rect 8297 12053 8309 12056
rect 8343 12053 8355 12087
rect 8297 12047 8355 12053
rect 9306 12044 9312 12096
rect 9364 12084 9370 12096
rect 9769 12087 9827 12093
rect 9769 12084 9781 12087
rect 9364 12056 9781 12084
rect 9364 12044 9370 12056
rect 9769 12053 9781 12056
rect 9815 12053 9827 12087
rect 9769 12047 9827 12053
rect 13081 12087 13139 12093
rect 13081 12053 13093 12087
rect 13127 12084 13139 12087
rect 13354 12084 13360 12096
rect 13127 12056 13360 12084
rect 13127 12053 13139 12056
rect 13081 12047 13139 12053
rect 13354 12044 13360 12056
rect 13412 12044 13418 12096
rect 15746 12044 15752 12096
rect 15804 12084 15810 12096
rect 16317 12087 16375 12093
rect 16317 12084 16329 12087
rect 15804 12056 16329 12084
rect 15804 12044 15810 12056
rect 16317 12053 16329 12056
rect 16363 12053 16375 12087
rect 16684 12084 16712 12124
rect 16942 12112 16948 12124
rect 17000 12112 17006 12164
rect 17144 12124 17954 12152
rect 17144 12084 17172 12124
rect 16684 12056 17172 12084
rect 17221 12087 17279 12093
rect 16317 12047 16375 12053
rect 17221 12053 17233 12087
rect 17267 12084 17279 12087
rect 17402 12084 17408 12096
rect 17267 12056 17408 12084
rect 17267 12053 17279 12056
rect 17221 12047 17279 12053
rect 17402 12044 17408 12056
rect 17460 12044 17466 12096
rect 17926 12084 17954 12124
rect 18598 12112 18604 12164
rect 18656 12152 18662 12164
rect 20162 12152 20168 12164
rect 18656 12124 20168 12152
rect 18656 12112 18662 12124
rect 20162 12112 20168 12124
rect 20220 12152 20226 12164
rect 21266 12152 21272 12164
rect 20220 12124 21272 12152
rect 20220 12112 20226 12124
rect 21266 12112 21272 12124
rect 21324 12112 21330 12164
rect 21542 12112 21548 12164
rect 21600 12152 21606 12164
rect 21600 12124 21645 12152
rect 21600 12112 21606 12124
rect 22370 12112 22376 12164
rect 22428 12152 22434 12164
rect 22646 12152 22652 12164
rect 22428 12124 22652 12152
rect 22428 12112 22434 12124
rect 22646 12112 22652 12124
rect 22704 12152 22710 12164
rect 22833 12155 22891 12161
rect 22833 12152 22845 12155
rect 22704 12124 22845 12152
rect 22704 12112 22710 12124
rect 22833 12121 22845 12124
rect 22879 12121 22891 12155
rect 22833 12115 22891 12121
rect 18417 12087 18475 12093
rect 18417 12084 18429 12087
rect 17926 12056 18429 12084
rect 18417 12053 18429 12056
rect 18463 12084 18475 12087
rect 20073 12087 20131 12093
rect 20073 12084 20085 12087
rect 18463 12056 20085 12084
rect 18463 12053 18475 12056
rect 18417 12047 18475 12053
rect 20073 12053 20085 12056
rect 20119 12084 20131 12087
rect 21174 12084 21180 12096
rect 20119 12056 21180 12084
rect 20119 12053 20131 12056
rect 20073 12047 20131 12053
rect 21174 12044 21180 12056
rect 21232 12084 21238 12096
rect 21450 12084 21456 12096
rect 21232 12056 21456 12084
rect 21232 12044 21238 12056
rect 21450 12044 21456 12056
rect 21508 12044 21514 12096
rect 1104 11994 23987 12016
rect 1104 11942 6630 11994
rect 6682 11942 6694 11994
rect 6746 11942 6758 11994
rect 6810 11942 6822 11994
rect 6874 11942 6886 11994
rect 6938 11942 12311 11994
rect 12363 11942 12375 11994
rect 12427 11942 12439 11994
rect 12491 11942 12503 11994
rect 12555 11942 12567 11994
rect 12619 11942 17992 11994
rect 18044 11942 18056 11994
rect 18108 11942 18120 11994
rect 18172 11942 18184 11994
rect 18236 11942 18248 11994
rect 18300 11942 23673 11994
rect 23725 11942 23737 11994
rect 23789 11942 23801 11994
rect 23853 11942 23865 11994
rect 23917 11942 23929 11994
rect 23981 11942 23987 11994
rect 1104 11920 23987 11942
rect 1762 11840 1768 11892
rect 1820 11880 1826 11892
rect 1857 11883 1915 11889
rect 1857 11880 1869 11883
rect 1820 11852 1869 11880
rect 1820 11840 1826 11852
rect 1857 11849 1869 11852
rect 1903 11849 1915 11883
rect 2498 11880 2504 11892
rect 2459 11852 2504 11880
rect 1857 11843 1915 11849
rect 2498 11840 2504 11852
rect 2556 11840 2562 11892
rect 2682 11880 2688 11892
rect 2643 11852 2688 11880
rect 2682 11840 2688 11852
rect 2740 11840 2746 11892
rect 2958 11840 2964 11892
rect 3016 11880 3022 11892
rect 4801 11883 4859 11889
rect 4801 11880 4813 11883
rect 3016 11852 4813 11880
rect 3016 11840 3022 11852
rect 4801 11849 4813 11852
rect 4847 11849 4859 11883
rect 4801 11843 4859 11849
rect 4890 11840 4896 11892
rect 4948 11880 4954 11892
rect 4948 11852 5488 11880
rect 4948 11840 4954 11852
rect 2700 11812 2728 11840
rect 1596 11784 2728 11812
rect 2869 11815 2927 11821
rect 1596 11753 1624 11784
rect 2869 11781 2881 11815
rect 2915 11812 2927 11815
rect 2915 11784 3004 11812
rect 2915 11781 2927 11784
rect 2869 11775 2927 11781
rect 2976 11756 3004 11784
rect 3326 11772 3332 11824
rect 3384 11812 3390 11824
rect 5166 11812 5172 11824
rect 3384 11784 4108 11812
rect 5127 11784 5172 11812
rect 3384 11772 3390 11784
rect 1581 11747 1639 11753
rect 1581 11713 1593 11747
rect 1627 11713 1639 11747
rect 1581 11707 1639 11713
rect 1670 11704 1676 11756
rect 1728 11744 1734 11756
rect 1728 11716 1773 11744
rect 1728 11704 1734 11716
rect 2958 11704 2964 11756
rect 3016 11704 3022 11756
rect 3510 11704 3516 11756
rect 3568 11744 3574 11756
rect 4080 11753 4108 11784
rect 5166 11772 5172 11784
rect 5224 11772 5230 11824
rect 5460 11756 5488 11852
rect 5626 11840 5632 11892
rect 5684 11880 5690 11892
rect 5905 11883 5963 11889
rect 5905 11880 5917 11883
rect 5684 11852 5917 11880
rect 5684 11840 5690 11852
rect 5905 11849 5917 11852
rect 5951 11849 5963 11883
rect 5905 11843 5963 11849
rect 7006 11840 7012 11892
rect 7064 11880 7070 11892
rect 7929 11883 7987 11889
rect 7929 11880 7941 11883
rect 7064 11852 7941 11880
rect 7064 11840 7070 11852
rect 7929 11849 7941 11852
rect 7975 11880 7987 11883
rect 9214 11880 9220 11892
rect 7975 11852 9220 11880
rect 7975 11849 7987 11852
rect 7929 11843 7987 11849
rect 9214 11840 9220 11852
rect 9272 11840 9278 11892
rect 11606 11840 11612 11892
rect 11664 11880 11670 11892
rect 11885 11883 11943 11889
rect 11885 11880 11897 11883
rect 11664 11852 11897 11880
rect 11664 11840 11670 11852
rect 11885 11849 11897 11852
rect 11931 11849 11943 11883
rect 11885 11843 11943 11849
rect 12069 11883 12127 11889
rect 12069 11849 12081 11883
rect 12115 11880 12127 11883
rect 13170 11880 13176 11892
rect 12115 11852 13176 11880
rect 12115 11849 12127 11852
rect 12069 11843 12127 11849
rect 13170 11840 13176 11852
rect 13228 11840 13234 11892
rect 17494 11840 17500 11892
rect 17552 11880 17558 11892
rect 17865 11883 17923 11889
rect 17865 11880 17877 11883
rect 17552 11852 17877 11880
rect 17552 11840 17558 11852
rect 17865 11849 17877 11852
rect 17911 11849 17923 11883
rect 17865 11843 17923 11849
rect 19150 11840 19156 11892
rect 19208 11880 19214 11892
rect 19705 11883 19763 11889
rect 19705 11880 19717 11883
rect 19208 11852 19717 11880
rect 19208 11840 19214 11852
rect 19705 11849 19717 11852
rect 19751 11849 19763 11883
rect 19705 11843 19763 11849
rect 19794 11840 19800 11892
rect 19852 11880 19858 11892
rect 19981 11883 20039 11889
rect 19981 11880 19993 11883
rect 19852 11852 19993 11880
rect 19852 11840 19858 11852
rect 19981 11849 19993 11852
rect 20027 11849 20039 11883
rect 21358 11880 21364 11892
rect 21319 11852 21364 11880
rect 19981 11843 20039 11849
rect 21358 11840 21364 11852
rect 21416 11840 21422 11892
rect 23014 11880 23020 11892
rect 22975 11852 23020 11880
rect 23014 11840 23020 11852
rect 23072 11840 23078 11892
rect 7190 11772 7196 11824
rect 7248 11812 7254 11824
rect 9401 11815 9459 11821
rect 7248 11784 7411 11812
rect 7248 11772 7254 11784
rect 3973 11747 4031 11753
rect 3973 11744 3985 11747
rect 3568 11716 3985 11744
rect 3568 11704 3574 11716
rect 3973 11713 3985 11716
rect 4019 11713 4031 11747
rect 3973 11707 4031 11713
rect 4066 11747 4124 11753
rect 4066 11713 4078 11747
rect 4112 11713 4124 11747
rect 4982 11744 4988 11756
rect 4943 11716 4988 11744
rect 4066 11707 4124 11713
rect 4982 11704 4988 11716
rect 5040 11704 5046 11756
rect 5077 11747 5135 11753
rect 5077 11713 5089 11747
rect 5123 11713 5135 11747
rect 5077 11707 5135 11713
rect 5287 11747 5345 11753
rect 5287 11713 5299 11747
rect 5333 11713 5345 11747
rect 5287 11707 5345 11713
rect 1854 11676 1860 11688
rect 1815 11648 1860 11676
rect 1854 11636 1860 11648
rect 1912 11636 1918 11688
rect 1946 11636 1952 11688
rect 2004 11676 2010 11688
rect 3329 11679 3387 11685
rect 3329 11676 3341 11679
rect 2004 11648 3341 11676
rect 2004 11636 2010 11648
rect 3329 11645 3341 11648
rect 3375 11676 3387 11679
rect 4614 11676 4620 11688
rect 3375 11648 4620 11676
rect 3375 11645 3387 11648
rect 3329 11639 3387 11645
rect 4614 11636 4620 11648
rect 4672 11636 4678 11688
rect 4890 11636 4896 11688
rect 4948 11676 4954 11688
rect 5088 11676 5116 11707
rect 4948 11648 5116 11676
rect 5292 11668 5320 11707
rect 5442 11704 5448 11756
rect 5500 11744 5506 11756
rect 5500 11716 5593 11744
rect 5500 11704 5506 11716
rect 6270 11704 6276 11756
rect 6328 11744 6334 11756
rect 7285 11747 7343 11753
rect 7285 11744 7297 11747
rect 6328 11716 7297 11744
rect 6328 11704 6334 11716
rect 7285 11713 7297 11716
rect 7331 11713 7343 11747
rect 7383 11744 7411 11784
rect 8128 11784 9260 11812
rect 7834 11744 7840 11756
rect 7383 11716 7840 11744
rect 7285 11707 7343 11713
rect 7834 11704 7840 11716
rect 7892 11704 7898 11756
rect 8128 11753 8156 11784
rect 8113 11747 8171 11753
rect 8113 11713 8125 11747
rect 8159 11713 8171 11747
rect 8662 11744 8668 11756
rect 8623 11716 8668 11744
rect 8113 11707 8171 11713
rect 8662 11704 8668 11716
rect 8720 11744 8726 11756
rect 9122 11744 9128 11756
rect 8720 11716 9128 11744
rect 8720 11704 8726 11716
rect 9122 11704 9128 11716
rect 9180 11704 9186 11756
rect 9232 11753 9260 11784
rect 9401 11781 9413 11815
rect 9447 11812 9459 11815
rect 11054 11812 11060 11824
rect 9447 11784 11060 11812
rect 9447 11781 9459 11784
rect 9401 11775 9459 11781
rect 11054 11772 11060 11784
rect 11112 11772 11118 11824
rect 11698 11812 11704 11824
rect 11659 11784 11704 11812
rect 11698 11772 11704 11784
rect 11756 11772 11762 11824
rect 11974 11772 11980 11824
rect 12032 11812 12038 11824
rect 12710 11812 12716 11824
rect 12032 11784 12716 11812
rect 12032 11772 12038 11784
rect 12710 11772 12716 11784
rect 12768 11812 12774 11824
rect 13449 11815 13507 11821
rect 13449 11812 13461 11815
rect 12768 11784 13461 11812
rect 12768 11772 12774 11784
rect 13449 11781 13461 11784
rect 13495 11781 13507 11815
rect 13449 11775 13507 11781
rect 14182 11772 14188 11824
rect 14240 11812 14246 11824
rect 14277 11815 14335 11821
rect 14277 11812 14289 11815
rect 14240 11784 14289 11812
rect 14240 11772 14246 11784
rect 14277 11781 14289 11784
rect 14323 11781 14335 11815
rect 14277 11775 14335 11781
rect 15102 11772 15108 11824
rect 15160 11812 15166 11824
rect 18782 11812 18788 11824
rect 15160 11784 18788 11812
rect 15160 11772 15166 11784
rect 18782 11772 18788 11784
rect 18840 11772 18846 11824
rect 19518 11772 19524 11824
rect 19576 11812 19582 11824
rect 19613 11815 19671 11821
rect 19613 11812 19625 11815
rect 19576 11784 19625 11812
rect 19576 11772 19582 11784
rect 19613 11781 19625 11784
rect 19659 11812 19671 11815
rect 22922 11812 22928 11824
rect 19659 11784 22928 11812
rect 19659 11781 19671 11784
rect 19613 11775 19671 11781
rect 22922 11772 22928 11784
rect 22980 11812 22986 11824
rect 23290 11812 23296 11824
rect 22980 11784 23296 11812
rect 22980 11772 22986 11784
rect 23290 11772 23296 11784
rect 23348 11772 23354 11824
rect 9217 11747 9275 11753
rect 9217 11713 9229 11747
rect 9263 11744 9275 11747
rect 9306 11744 9312 11756
rect 9263 11716 9312 11744
rect 9263 11713 9275 11716
rect 9217 11707 9275 11713
rect 9306 11704 9312 11716
rect 9364 11704 9370 11756
rect 10226 11704 10232 11756
rect 10284 11744 10290 11756
rect 10321 11747 10379 11753
rect 10321 11744 10333 11747
rect 10284 11716 10333 11744
rect 10284 11704 10290 11716
rect 10321 11713 10333 11716
rect 10367 11713 10379 11747
rect 10321 11707 10379 11713
rect 10502 11704 10508 11756
rect 10560 11744 10566 11756
rect 10778 11744 10784 11756
rect 10560 11716 10784 11744
rect 10560 11704 10566 11716
rect 10778 11704 10784 11716
rect 10836 11744 10842 11756
rect 10965 11747 11023 11753
rect 10965 11744 10977 11747
rect 10836 11716 10977 11744
rect 10836 11704 10842 11716
rect 10965 11713 10977 11716
rect 11011 11713 11023 11747
rect 10965 11707 11023 11713
rect 11149 11747 11207 11753
rect 11149 11713 11161 11747
rect 11195 11744 11207 11747
rect 11238 11744 11244 11756
rect 11195 11716 11244 11744
rect 11195 11713 11207 11716
rect 11149 11707 11207 11713
rect 11238 11704 11244 11716
rect 11296 11704 11302 11756
rect 12066 11704 12072 11756
rect 12124 11744 12130 11756
rect 13357 11747 13415 11753
rect 13357 11744 13369 11747
rect 12124 11716 13369 11744
rect 12124 11704 12130 11716
rect 13357 11713 13369 11716
rect 13403 11713 13415 11747
rect 13817 11747 13875 11753
rect 13817 11744 13829 11747
rect 13357 11707 13415 11713
rect 13464 11716 13829 11744
rect 13464 11688 13492 11716
rect 13817 11713 13829 11716
rect 13863 11713 13875 11747
rect 17402 11744 17408 11756
rect 17363 11716 17408 11744
rect 13817 11707 13875 11713
rect 17402 11704 17408 11716
rect 17460 11704 17466 11756
rect 17586 11744 17592 11756
rect 17547 11716 17592 11744
rect 17586 11704 17592 11716
rect 17644 11704 17650 11756
rect 17681 11747 17739 11753
rect 17681 11713 17693 11747
rect 17727 11744 17739 11747
rect 17770 11744 17776 11756
rect 17727 11716 17776 11744
rect 17727 11713 17739 11716
rect 17681 11707 17739 11713
rect 17770 11704 17776 11716
rect 17828 11704 17834 11756
rect 18966 11704 18972 11756
rect 19024 11744 19030 11756
rect 19429 11747 19487 11753
rect 19429 11744 19441 11747
rect 19024 11716 19441 11744
rect 19024 11704 19030 11716
rect 5626 11676 5632 11688
rect 4948 11636 4954 11648
rect 5292 11640 5396 11668
rect 5368 11608 5396 11640
rect 5552 11648 5632 11676
rect 5552 11608 5580 11648
rect 5626 11636 5632 11648
rect 5684 11636 5690 11688
rect 7009 11679 7067 11685
rect 7009 11676 7021 11679
rect 6472 11648 7021 11676
rect 5368 11580 5580 11608
rect 2130 11500 2136 11552
rect 2188 11540 2194 11552
rect 2685 11543 2743 11549
rect 2685 11540 2697 11543
rect 2188 11512 2697 11540
rect 2188 11500 2194 11512
rect 2685 11509 2697 11512
rect 2731 11540 2743 11543
rect 2774 11540 2780 11552
rect 2731 11512 2780 11540
rect 2731 11509 2743 11512
rect 2685 11503 2743 11509
rect 2774 11500 2780 11512
rect 2832 11500 2838 11552
rect 4157 11543 4215 11549
rect 4157 11509 4169 11543
rect 4203 11540 4215 11543
rect 6472 11540 6500 11648
rect 7009 11645 7021 11648
rect 7055 11645 7067 11679
rect 7009 11639 7067 11645
rect 7101 11679 7159 11685
rect 7101 11645 7113 11679
rect 7147 11645 7159 11679
rect 7101 11639 7159 11645
rect 4203 11512 6500 11540
rect 4203 11509 4215 11512
rect 4157 11503 4215 11509
rect 6546 11500 6552 11552
rect 6604 11540 6610 11552
rect 6825 11543 6883 11549
rect 6825 11540 6837 11543
rect 6604 11512 6837 11540
rect 6604 11500 6610 11512
rect 6825 11509 6837 11512
rect 6871 11509 6883 11543
rect 7024 11540 7052 11639
rect 7116 11608 7144 11639
rect 7190 11636 7196 11688
rect 7248 11676 7254 11688
rect 10042 11676 10048 11688
rect 7248 11648 7293 11676
rect 10003 11648 10048 11676
rect 7248 11636 7254 11648
rect 10042 11636 10048 11648
rect 10100 11636 10106 11688
rect 13446 11636 13452 11688
rect 13504 11636 13510 11688
rect 13541 11679 13599 11685
rect 13541 11645 13553 11679
rect 13587 11676 13599 11679
rect 13722 11676 13728 11688
rect 13587 11648 13728 11676
rect 13587 11645 13599 11648
rect 13541 11639 13599 11645
rect 13722 11636 13728 11648
rect 13780 11636 13786 11688
rect 15654 11636 15660 11688
rect 15712 11676 15718 11688
rect 15712 11648 16068 11676
rect 15712 11636 15718 11648
rect 7650 11608 7656 11620
rect 7116 11580 7656 11608
rect 7650 11568 7656 11580
rect 7708 11568 7714 11620
rect 16040 11608 16068 11648
rect 17310 11636 17316 11688
rect 17368 11676 17374 11688
rect 17497 11679 17555 11685
rect 17497 11676 17509 11679
rect 17368 11648 17509 11676
rect 17368 11636 17374 11648
rect 17497 11645 17509 11648
rect 17543 11645 17555 11679
rect 17497 11639 17555 11645
rect 19260 11608 19288 11716
rect 19429 11713 19441 11716
rect 19475 11713 19487 11747
rect 19429 11707 19487 11713
rect 19797 11747 19855 11753
rect 19797 11713 19809 11747
rect 19843 11744 19855 11747
rect 19978 11744 19984 11756
rect 19843 11716 19984 11744
rect 19843 11713 19855 11716
rect 19797 11707 19855 11713
rect 19334 11636 19340 11688
rect 19392 11676 19398 11688
rect 19812 11676 19840 11707
rect 19978 11704 19984 11716
rect 20036 11704 20042 11756
rect 21269 11747 21327 11753
rect 21269 11713 21281 11747
rect 21315 11744 21327 11747
rect 21358 11744 21364 11756
rect 21315 11716 21364 11744
rect 21315 11713 21327 11716
rect 21269 11707 21327 11713
rect 21358 11704 21364 11716
rect 21416 11704 21422 11756
rect 21453 11747 21511 11753
rect 21453 11713 21465 11747
rect 21499 11744 21511 11747
rect 21726 11744 21732 11756
rect 21499 11716 21732 11744
rect 21499 11713 21511 11716
rect 21453 11707 21511 11713
rect 21726 11704 21732 11716
rect 21784 11704 21790 11756
rect 22094 11704 22100 11756
rect 22152 11744 22158 11756
rect 23014 11744 23020 11756
rect 22152 11716 22197 11744
rect 22975 11716 23020 11744
rect 22152 11704 22158 11716
rect 23014 11704 23020 11716
rect 23072 11704 23078 11756
rect 23106 11704 23112 11756
rect 23164 11744 23170 11756
rect 23201 11747 23259 11753
rect 23201 11744 23213 11747
rect 23164 11716 23213 11744
rect 23164 11704 23170 11716
rect 23201 11713 23213 11716
rect 23247 11713 23259 11747
rect 23201 11707 23259 11713
rect 19392 11648 19840 11676
rect 22373 11679 22431 11685
rect 19392 11636 19398 11648
rect 22373 11645 22385 11679
rect 22419 11676 22431 11679
rect 22646 11676 22652 11688
rect 22419 11648 22652 11676
rect 22419 11645 22431 11648
rect 22373 11639 22431 11645
rect 22646 11636 22652 11648
rect 22704 11636 22710 11688
rect 20441 11611 20499 11617
rect 20441 11608 20453 11611
rect 13648 11580 15976 11608
rect 16040 11580 18828 11608
rect 19260 11580 20453 11608
rect 8110 11540 8116 11552
rect 7024 11512 8116 11540
rect 6825 11503 6883 11509
rect 8110 11500 8116 11512
rect 8168 11500 8174 11552
rect 9858 11500 9864 11552
rect 9916 11540 9922 11552
rect 10781 11543 10839 11549
rect 10781 11540 10793 11543
rect 9916 11512 10793 11540
rect 9916 11500 9922 11512
rect 10781 11509 10793 11512
rect 10827 11509 10839 11543
rect 10781 11503 10839 11509
rect 10962 11500 10968 11552
rect 11020 11540 11026 11552
rect 11885 11543 11943 11549
rect 11885 11540 11897 11543
rect 11020 11512 11897 11540
rect 11020 11500 11026 11512
rect 11885 11509 11897 11512
rect 11931 11509 11943 11543
rect 11885 11503 11943 11509
rect 13538 11500 13544 11552
rect 13596 11540 13602 11552
rect 13648 11540 13676 11580
rect 15948 11552 15976 11580
rect 18800 11552 18828 11580
rect 20441 11577 20453 11580
rect 20487 11577 20499 11611
rect 20441 11571 20499 11577
rect 13596 11512 13676 11540
rect 13596 11500 13602 11512
rect 14366 11500 14372 11552
rect 14424 11540 14430 11552
rect 14734 11540 14740 11552
rect 14424 11512 14740 11540
rect 14424 11500 14430 11512
rect 14734 11500 14740 11512
rect 14792 11500 14798 11552
rect 15381 11543 15439 11549
rect 15381 11509 15393 11543
rect 15427 11540 15439 11543
rect 15562 11540 15568 11552
rect 15427 11512 15568 11540
rect 15427 11509 15439 11512
rect 15381 11503 15439 11509
rect 15562 11500 15568 11512
rect 15620 11500 15626 11552
rect 15930 11540 15936 11552
rect 15891 11512 15936 11540
rect 15930 11500 15936 11512
rect 15988 11500 15994 11552
rect 18414 11540 18420 11552
rect 18375 11512 18420 11540
rect 18414 11500 18420 11512
rect 18472 11500 18478 11552
rect 18782 11500 18788 11552
rect 18840 11540 18846 11552
rect 18969 11543 19027 11549
rect 18969 11540 18981 11543
rect 18840 11512 18981 11540
rect 18840 11500 18846 11512
rect 18969 11509 18981 11512
rect 19015 11540 19027 11543
rect 19978 11540 19984 11552
rect 19015 11512 19984 11540
rect 19015 11509 19027 11512
rect 18969 11503 19027 11509
rect 19978 11500 19984 11512
rect 20036 11500 20042 11552
rect 1104 11450 23828 11472
rect 1104 11398 3790 11450
rect 3842 11398 3854 11450
rect 3906 11398 3918 11450
rect 3970 11398 3982 11450
rect 4034 11398 4046 11450
rect 4098 11398 9471 11450
rect 9523 11398 9535 11450
rect 9587 11398 9599 11450
rect 9651 11398 9663 11450
rect 9715 11398 9727 11450
rect 9779 11398 15152 11450
rect 15204 11398 15216 11450
rect 15268 11398 15280 11450
rect 15332 11398 15344 11450
rect 15396 11398 15408 11450
rect 15460 11398 20833 11450
rect 20885 11398 20897 11450
rect 20949 11398 20961 11450
rect 21013 11398 21025 11450
rect 21077 11398 21089 11450
rect 21141 11398 23828 11450
rect 1104 11376 23828 11398
rect 3234 11296 3240 11348
rect 3292 11336 3298 11348
rect 4617 11339 4675 11345
rect 4617 11336 4629 11339
rect 3292 11308 4629 11336
rect 3292 11296 3298 11308
rect 4617 11305 4629 11308
rect 4663 11305 4675 11339
rect 4617 11299 4675 11305
rect 7466 11296 7472 11348
rect 7524 11336 7530 11348
rect 9125 11339 9183 11345
rect 9125 11336 9137 11339
rect 7524 11308 9137 11336
rect 7524 11296 7530 11308
rect 9125 11305 9137 11308
rect 9171 11305 9183 11339
rect 13078 11336 13084 11348
rect 9125 11299 9183 11305
rect 12176 11308 13084 11336
rect 1854 11228 1860 11280
rect 1912 11268 1918 11280
rect 3145 11271 3203 11277
rect 3145 11268 3157 11271
rect 1912 11240 3157 11268
rect 1912 11228 1918 11240
rect 3145 11237 3157 11240
rect 3191 11268 3203 11271
rect 3878 11268 3884 11280
rect 3191 11240 3884 11268
rect 3191 11237 3203 11240
rect 3145 11231 3203 11237
rect 3878 11228 3884 11240
rect 3936 11228 3942 11280
rect 4338 11268 4344 11280
rect 4080 11240 4344 11268
rect 4080 11212 4108 11240
rect 4338 11228 4344 11240
rect 4396 11228 4402 11280
rect 7926 11228 7932 11280
rect 7984 11268 7990 11280
rect 7984 11240 10824 11268
rect 7984 11228 7990 11240
rect 4062 11200 4068 11212
rect 2792 11172 4068 11200
rect 1578 11132 1584 11144
rect 1539 11104 1584 11132
rect 1578 11092 1584 11104
rect 1636 11092 1642 11144
rect 2406 11132 2412 11144
rect 2367 11104 2412 11132
rect 2406 11092 2412 11104
rect 2464 11092 2470 11144
rect 2792 11141 2820 11172
rect 4062 11160 4068 11172
rect 4120 11160 4126 11212
rect 4154 11160 4160 11212
rect 4212 11200 4218 11212
rect 4433 11203 4491 11209
rect 4433 11200 4445 11203
rect 4212 11172 4445 11200
rect 4212 11160 4218 11172
rect 4433 11169 4445 11172
rect 4479 11169 4491 11203
rect 4433 11163 4491 11169
rect 4614 11160 4620 11212
rect 4672 11200 4678 11212
rect 5537 11203 5595 11209
rect 5537 11200 5549 11203
rect 4672 11172 5549 11200
rect 4672 11160 4678 11172
rect 5537 11169 5549 11172
rect 5583 11200 5595 11203
rect 5718 11200 5724 11212
rect 5583 11172 5724 11200
rect 5583 11169 5595 11172
rect 5537 11163 5595 11169
rect 5718 11160 5724 11172
rect 5776 11160 5782 11212
rect 7834 11160 7840 11212
rect 7892 11200 7898 11212
rect 8481 11203 8539 11209
rect 8481 11200 8493 11203
rect 7892 11172 8493 11200
rect 7892 11160 7898 11172
rect 8481 11169 8493 11172
rect 8527 11169 8539 11203
rect 9858 11200 9864 11212
rect 8481 11163 8539 11169
rect 9508 11172 9864 11200
rect 2777 11135 2835 11141
rect 2777 11101 2789 11135
rect 2823 11101 2835 11135
rect 2777 11095 2835 11101
rect 2866 11092 2872 11144
rect 2924 11132 2930 11144
rect 2961 11135 3019 11141
rect 2961 11132 2973 11135
rect 2924 11104 2973 11132
rect 2924 11092 2930 11104
rect 2961 11101 2973 11104
rect 3007 11132 3019 11135
rect 3510 11132 3516 11144
rect 3007 11104 3516 11132
rect 3007 11101 3019 11104
rect 2961 11095 3019 11101
rect 3510 11092 3516 11104
rect 3568 11132 3574 11144
rect 3973 11135 4031 11141
rect 3973 11132 3985 11135
rect 3568 11104 3985 11132
rect 3568 11092 3574 11104
rect 3973 11101 3985 11104
rect 4019 11101 4031 11135
rect 4338 11132 4344 11144
rect 4299 11104 4344 11132
rect 3973 11095 4031 11101
rect 4338 11092 4344 11104
rect 4396 11092 4402 11144
rect 5902 11092 5908 11144
rect 5960 11132 5966 11144
rect 6641 11135 6699 11141
rect 6641 11132 6653 11135
rect 5960 11104 6653 11132
rect 5960 11092 5966 11104
rect 6641 11101 6653 11104
rect 6687 11101 6699 11135
rect 6641 11095 6699 11101
rect 7282 11092 7288 11144
rect 7340 11132 7346 11144
rect 7377 11135 7435 11141
rect 7377 11132 7389 11135
rect 7340 11104 7389 11132
rect 7340 11092 7346 11104
rect 7377 11101 7389 11104
rect 7423 11132 7435 11135
rect 7466 11132 7472 11144
rect 7423 11104 7472 11132
rect 7423 11101 7435 11104
rect 7377 11095 7435 11101
rect 7466 11092 7472 11104
rect 7524 11092 7530 11144
rect 9214 11092 9220 11144
rect 9272 11132 9278 11144
rect 9508 11141 9536 11172
rect 9858 11160 9864 11172
rect 9916 11160 9922 11212
rect 9309 11135 9367 11141
rect 9309 11132 9321 11135
rect 9272 11104 9321 11132
rect 9272 11092 9278 11104
rect 9309 11101 9321 11104
rect 9355 11101 9367 11135
rect 9309 11095 9367 11101
rect 9493 11135 9551 11141
rect 9493 11101 9505 11135
rect 9539 11101 9551 11135
rect 9766 11132 9772 11144
rect 9727 11104 9772 11132
rect 9493 11095 9551 11101
rect 9766 11092 9772 11104
rect 9824 11092 9830 11144
rect 10594 11132 10600 11144
rect 10555 11104 10600 11132
rect 10594 11092 10600 11104
rect 10652 11092 10658 11144
rect 10796 11141 10824 11240
rect 12176 11200 12204 11308
rect 13078 11296 13084 11308
rect 13136 11336 13142 11348
rect 13538 11336 13544 11348
rect 13136 11308 13544 11336
rect 13136 11296 13142 11308
rect 13538 11296 13544 11308
rect 13596 11296 13602 11348
rect 13633 11339 13691 11345
rect 13633 11305 13645 11339
rect 13679 11336 13691 11339
rect 14642 11336 14648 11348
rect 13679 11308 14648 11336
rect 13679 11305 13691 11308
rect 13633 11299 13691 11305
rect 14642 11296 14648 11308
rect 14700 11296 14706 11348
rect 16022 11296 16028 11348
rect 16080 11336 16086 11348
rect 19521 11339 19579 11345
rect 19521 11336 19533 11339
rect 16080 11308 19533 11336
rect 16080 11296 16086 11308
rect 19521 11305 19533 11308
rect 19567 11305 19579 11339
rect 19521 11299 19579 11305
rect 19610 11296 19616 11348
rect 19668 11336 19674 11348
rect 22278 11336 22284 11348
rect 19668 11308 19713 11336
rect 22239 11308 22284 11336
rect 19668 11296 19674 11308
rect 22278 11296 22284 11308
rect 22336 11296 22342 11348
rect 14921 11271 14979 11277
rect 14921 11237 14933 11271
rect 14967 11268 14979 11271
rect 15010 11268 15016 11280
rect 14967 11240 15016 11268
rect 14967 11237 14979 11240
rect 14921 11231 14979 11237
rect 15010 11228 15016 11240
rect 15068 11228 15074 11280
rect 15562 11268 15568 11280
rect 15475 11240 15568 11268
rect 15562 11228 15568 11240
rect 15620 11268 15626 11280
rect 16850 11268 16856 11280
rect 15620 11240 16856 11268
rect 15620 11228 15626 11240
rect 16850 11228 16856 11240
rect 16908 11228 16914 11280
rect 16942 11228 16948 11280
rect 17000 11268 17006 11280
rect 20809 11271 20867 11277
rect 17000 11240 19380 11268
rect 17000 11228 17006 11240
rect 15378 11200 15384 11212
rect 12084 11172 12204 11200
rect 14568 11172 15384 11200
rect 10781 11135 10839 11141
rect 10781 11101 10793 11135
rect 10827 11101 10839 11135
rect 11882 11132 11888 11144
rect 11843 11104 11888 11132
rect 10781 11095 10839 11101
rect 11882 11092 11888 11104
rect 11940 11092 11946 11144
rect 12084 11141 12112 11172
rect 12069 11135 12127 11141
rect 12069 11101 12081 11135
rect 12115 11101 12127 11135
rect 12069 11095 12127 11101
rect 12161 11135 12219 11141
rect 12161 11101 12173 11135
rect 12207 11101 12219 11135
rect 12618 11132 12624 11144
rect 12579 11104 12624 11132
rect 12161 11095 12219 11101
rect 2424 11064 2452 11092
rect 4246 11064 4252 11076
rect 2424 11036 4252 11064
rect 4172 11005 4200 11036
rect 4246 11024 4252 11036
rect 4304 11024 4310 11076
rect 6086 11024 6092 11076
rect 6144 11064 6150 11076
rect 6144 11036 6486 11064
rect 6144 11024 6150 11036
rect 8570 11024 8576 11076
rect 8628 11064 8634 11076
rect 9401 11067 9459 11073
rect 9401 11064 9413 11067
rect 8628 11036 9413 11064
rect 8628 11024 8634 11036
rect 9401 11033 9413 11036
rect 9447 11033 9459 11067
rect 9401 11027 9459 11033
rect 9631 11067 9689 11073
rect 9631 11033 9643 11067
rect 9677 11064 9689 11067
rect 10042 11064 10048 11076
rect 9677 11036 10048 11064
rect 9677 11033 9689 11036
rect 9631 11027 9689 11033
rect 10042 11024 10048 11036
rect 10100 11024 10106 11076
rect 10689 11067 10747 11073
rect 10689 11033 10701 11067
rect 10735 11064 10747 11067
rect 10962 11064 10968 11076
rect 10735 11036 10968 11064
rect 10735 11033 10747 11036
rect 10689 11027 10747 11033
rect 10962 11024 10968 11036
rect 11020 11024 11026 11076
rect 12176 11064 12204 11095
rect 12618 11092 12624 11104
rect 12676 11092 12682 11144
rect 13078 11132 13084 11144
rect 13039 11104 13084 11132
rect 13078 11092 13084 11104
rect 13136 11092 13142 11144
rect 13446 11132 13452 11144
rect 13407 11104 13452 11132
rect 13446 11092 13452 11104
rect 13504 11092 13510 11144
rect 13814 11092 13820 11144
rect 13872 11132 13878 11144
rect 14274 11132 14280 11144
rect 13872 11104 14280 11132
rect 13872 11092 13878 11104
rect 14274 11092 14280 11104
rect 14332 11092 14338 11144
rect 14370 11135 14428 11141
rect 14370 11101 14382 11135
rect 14416 11101 14428 11135
rect 14370 11095 14428 11101
rect 12986 11064 12992 11076
rect 12176 11036 12992 11064
rect 12986 11024 12992 11036
rect 13044 11064 13050 11076
rect 13265 11067 13323 11073
rect 13265 11064 13277 11067
rect 13044 11036 13277 11064
rect 13044 11024 13050 11036
rect 13265 11033 13277 11036
rect 13311 11033 13323 11067
rect 13265 11027 13323 11033
rect 4157 10999 4215 11005
rect 4157 10965 4169 10999
rect 4203 10965 4215 10999
rect 4157 10959 4215 10965
rect 5810 10956 5816 11008
rect 5868 10996 5874 11008
rect 7374 10996 7380 11008
rect 5868 10968 7380 10996
rect 5868 10956 5874 10968
rect 7374 10956 7380 10968
rect 7432 10996 7438 11008
rect 9766 10996 9772 11008
rect 7432 10968 9772 10996
rect 7432 10956 7438 10968
rect 9766 10956 9772 10968
rect 9824 10956 9830 11008
rect 11425 10999 11483 11005
rect 11425 10965 11437 10999
rect 11471 10996 11483 10999
rect 12158 10996 12164 11008
rect 11471 10968 12164 10996
rect 11471 10965 11483 10968
rect 11425 10959 11483 10965
rect 12158 10956 12164 10968
rect 12216 10956 12222 11008
rect 13280 10996 13308 11027
rect 13354 11024 13360 11076
rect 13412 11064 13418 11076
rect 13412 11036 13457 11064
rect 13412 11024 13418 11036
rect 14182 11024 14188 11076
rect 14240 11064 14246 11076
rect 14384 11064 14412 11095
rect 14568 11073 14596 11172
rect 15378 11160 15384 11172
rect 15436 11160 15442 11212
rect 14742 11135 14800 11141
rect 14742 11101 14754 11135
rect 14788 11126 14800 11135
rect 14788 11101 14872 11126
rect 14742 11098 14872 11101
rect 14742 11095 14800 11098
rect 14240 11036 14412 11064
rect 14553 11067 14611 11073
rect 14240 11024 14246 11036
rect 14553 11033 14565 11067
rect 14599 11033 14611 11067
rect 14553 11027 14611 11033
rect 14645 11067 14703 11073
rect 14645 11033 14657 11067
rect 14691 11064 14703 11067
rect 14844 11064 14872 11098
rect 14918 11092 14924 11144
rect 14976 11132 14982 11144
rect 15473 11135 15531 11141
rect 15473 11132 15485 11135
rect 14976 11104 15485 11132
rect 14976 11092 14982 11104
rect 15473 11101 15485 11104
rect 15519 11132 15531 11135
rect 15580 11132 15608 11228
rect 15746 11200 15752 11212
rect 15707 11172 15752 11200
rect 15746 11160 15752 11172
rect 15804 11160 15810 11212
rect 15930 11160 15936 11212
rect 15988 11200 15994 11212
rect 18417 11203 18475 11209
rect 18417 11200 18429 11203
rect 15988 11172 18429 11200
rect 15988 11160 15994 11172
rect 18417 11169 18429 11172
rect 18463 11200 18475 11203
rect 19352 11208 19380 11240
rect 20809 11237 20821 11271
rect 20855 11268 20867 11271
rect 21174 11268 21180 11280
rect 20855 11240 21180 11268
rect 20855 11237 20867 11240
rect 20809 11231 20867 11237
rect 21174 11228 21180 11240
rect 21232 11268 21238 11280
rect 23382 11268 23388 11280
rect 21232 11240 23388 11268
rect 21232 11228 21238 11240
rect 23382 11228 23388 11240
rect 23440 11228 23446 11280
rect 19429 11208 19487 11209
rect 19352 11203 19487 11208
rect 18463 11172 18920 11200
rect 19352 11180 19441 11203
rect 18463 11169 18475 11172
rect 18417 11163 18475 11169
rect 15519 11104 15608 11132
rect 15657 11135 15715 11141
rect 15519 11101 15531 11104
rect 15473 11095 15531 11101
rect 15657 11101 15669 11135
rect 15703 11132 15715 11135
rect 16114 11132 16120 11144
rect 15703 11104 16120 11132
rect 15703 11101 15715 11104
rect 15657 11095 15715 11101
rect 16114 11092 16120 11104
rect 16172 11092 16178 11144
rect 16850 11132 16856 11144
rect 16763 11104 16856 11132
rect 16850 11092 16856 11104
rect 16908 11132 16914 11144
rect 17405 11135 17463 11141
rect 17405 11132 17417 11135
rect 16908 11104 17417 11132
rect 16908 11092 16914 11104
rect 17405 11101 17417 11104
rect 17451 11132 17463 11135
rect 17770 11132 17776 11144
rect 17451 11104 17776 11132
rect 17451 11101 17463 11104
rect 17405 11095 17463 11101
rect 17770 11092 17776 11104
rect 17828 11092 17834 11144
rect 18230 11092 18236 11144
rect 18288 11132 18294 11144
rect 18325 11135 18383 11141
rect 18325 11132 18337 11135
rect 18288 11104 18337 11132
rect 18288 11092 18294 11104
rect 18325 11101 18337 11104
rect 18371 11101 18383 11135
rect 18598 11132 18604 11144
rect 18559 11104 18604 11132
rect 18325 11095 18383 11101
rect 18598 11092 18604 11104
rect 18656 11092 18662 11144
rect 18693 11135 18751 11141
rect 18693 11101 18705 11135
rect 18739 11132 18751 11135
rect 18782 11132 18788 11144
rect 18739 11104 18788 11132
rect 18739 11101 18751 11104
rect 18693 11095 18751 11101
rect 18782 11092 18788 11104
rect 18840 11092 18846 11144
rect 18892 11132 18920 11172
rect 19429 11169 19441 11180
rect 19475 11169 19487 11203
rect 22833 11203 22891 11209
rect 22833 11200 22845 11203
rect 19429 11163 19487 11169
rect 19536 11172 20300 11200
rect 19536 11132 19564 11172
rect 18892 11104 19564 11132
rect 19702 11092 19708 11144
rect 19760 11132 19766 11144
rect 19760 11104 19805 11132
rect 19760 11092 19766 11104
rect 15102 11064 15108 11076
rect 14691 11036 14780 11064
rect 14844 11036 15108 11064
rect 14691 11033 14703 11036
rect 14645 11027 14703 11033
rect 14568 10996 14596 11027
rect 13280 10968 14596 10996
rect 14752 10996 14780 11036
rect 15102 11024 15108 11036
rect 15160 11064 15166 11076
rect 16301 11067 16359 11073
rect 16301 11064 16313 11067
rect 15160 11036 16313 11064
rect 15160 11024 15166 11036
rect 16301 11033 16313 11036
rect 16347 11064 16359 11067
rect 17862 11064 17868 11076
rect 16347 11036 17868 11064
rect 16347 11033 16359 11036
rect 16301 11027 16359 11033
rect 17862 11024 17868 11036
rect 17920 11024 17926 11076
rect 18874 11064 18880 11076
rect 18787 11036 18880 11064
rect 18874 11024 18880 11036
rect 18932 11064 18938 11076
rect 19610 11064 19616 11076
rect 18932 11036 19616 11064
rect 18932 11024 18938 11036
rect 19610 11024 19616 11036
rect 19668 11024 19674 11076
rect 20272 11073 20300 11172
rect 22112 11172 22845 11200
rect 21450 11092 21456 11144
rect 21508 11132 21514 11144
rect 22112 11141 22140 11172
rect 22833 11169 22845 11172
rect 22879 11200 22891 11203
rect 23014 11200 23020 11212
rect 22879 11172 23020 11200
rect 22879 11169 22891 11172
rect 22833 11163 22891 11169
rect 23014 11160 23020 11172
rect 23072 11160 23078 11212
rect 22097 11135 22155 11141
rect 22097 11132 22109 11135
rect 21508 11104 22109 11132
rect 21508 11092 21514 11104
rect 22097 11101 22109 11104
rect 22143 11101 22155 11135
rect 22097 11095 22155 11101
rect 22373 11135 22431 11141
rect 22373 11101 22385 11135
rect 22419 11132 22431 11135
rect 22419 11104 22453 11132
rect 22419 11101 22431 11104
rect 22373 11095 22431 11101
rect 20257 11067 20315 11073
rect 20257 11033 20269 11067
rect 20303 11064 20315 11067
rect 22388 11064 22416 11095
rect 22646 11064 22652 11076
rect 20303 11036 22652 11064
rect 20303 11033 20315 11036
rect 20257 11027 20315 11033
rect 22646 11024 22652 11036
rect 22704 11064 22710 11076
rect 23290 11064 23296 11076
rect 22704 11036 23296 11064
rect 22704 11024 22710 11036
rect 23290 11024 23296 11036
rect 23348 11024 23354 11076
rect 15654 10996 15660 11008
rect 14752 10968 15660 10996
rect 15654 10956 15660 10968
rect 15712 10956 15718 11008
rect 15746 10956 15752 11008
rect 15804 10996 15810 11008
rect 16482 10996 16488 11008
rect 15804 10968 16488 10996
rect 15804 10956 15810 10968
rect 16482 10956 16488 10968
rect 16540 10996 16546 11008
rect 18414 10996 18420 11008
rect 16540 10968 18420 10996
rect 16540 10956 16546 10968
rect 18414 10956 18420 10968
rect 18472 10996 18478 11008
rect 18782 10996 18788 11008
rect 18472 10968 18788 10996
rect 18472 10956 18478 10968
rect 18782 10956 18788 10968
rect 18840 10956 18846 11008
rect 21358 10996 21364 11008
rect 21271 10968 21364 10996
rect 21358 10956 21364 10968
rect 21416 10996 21422 11008
rect 21726 10996 21732 11008
rect 21416 10968 21732 10996
rect 21416 10956 21422 10968
rect 21726 10956 21732 10968
rect 21784 10956 21790 11008
rect 1104 10906 23987 10928
rect 1104 10854 6630 10906
rect 6682 10854 6694 10906
rect 6746 10854 6758 10906
rect 6810 10854 6822 10906
rect 6874 10854 6886 10906
rect 6938 10854 12311 10906
rect 12363 10854 12375 10906
rect 12427 10854 12439 10906
rect 12491 10854 12503 10906
rect 12555 10854 12567 10906
rect 12619 10854 17992 10906
rect 18044 10854 18056 10906
rect 18108 10854 18120 10906
rect 18172 10854 18184 10906
rect 18236 10854 18248 10906
rect 18300 10854 23673 10906
rect 23725 10854 23737 10906
rect 23789 10854 23801 10906
rect 23853 10854 23865 10906
rect 23917 10854 23929 10906
rect 23981 10854 23987 10906
rect 1104 10832 23987 10854
rect 1578 10752 1584 10804
rect 1636 10792 1642 10804
rect 1765 10795 1823 10801
rect 1765 10792 1777 10795
rect 1636 10764 1777 10792
rect 1636 10752 1642 10764
rect 1765 10761 1777 10764
rect 1811 10761 1823 10795
rect 2958 10792 2964 10804
rect 1765 10755 1823 10761
rect 1964 10764 2964 10792
rect 1964 10665 1992 10764
rect 2958 10752 2964 10764
rect 3016 10792 3022 10804
rect 4246 10792 4252 10804
rect 3016 10764 4252 10792
rect 3016 10752 3022 10764
rect 4246 10752 4252 10764
rect 4304 10752 4310 10804
rect 4338 10752 4344 10804
rect 4396 10792 4402 10804
rect 4706 10792 4712 10804
rect 4396 10764 4712 10792
rect 4396 10752 4402 10764
rect 4706 10752 4712 10764
rect 4764 10792 4770 10804
rect 5277 10795 5335 10801
rect 5277 10792 5289 10795
rect 4764 10764 5289 10792
rect 4764 10752 4770 10764
rect 5277 10761 5289 10764
rect 5323 10761 5335 10795
rect 5277 10755 5335 10761
rect 6362 10752 6368 10804
rect 6420 10792 6426 10804
rect 6641 10795 6699 10801
rect 6641 10792 6653 10795
rect 6420 10764 6653 10792
rect 6420 10752 6426 10764
rect 6641 10761 6653 10764
rect 6687 10761 6699 10795
rect 10870 10792 10876 10804
rect 6641 10755 6699 10761
rect 6932 10764 10876 10792
rect 2038 10684 2044 10736
rect 2096 10724 2102 10736
rect 2225 10727 2283 10733
rect 2225 10724 2237 10727
rect 2096 10696 2237 10724
rect 2096 10684 2102 10696
rect 2225 10693 2237 10696
rect 2271 10724 2283 10727
rect 2271 10696 3648 10724
rect 2271 10693 2283 10696
rect 2225 10687 2283 10693
rect 1949 10659 2007 10665
rect 1949 10625 1961 10659
rect 1995 10625 2007 10659
rect 1949 10619 2007 10625
rect 2685 10659 2743 10665
rect 2685 10625 2697 10659
rect 2731 10625 2743 10659
rect 2685 10619 2743 10625
rect 2133 10591 2191 10597
rect 2133 10557 2145 10591
rect 2179 10588 2191 10591
rect 2314 10588 2320 10600
rect 2179 10560 2320 10588
rect 2179 10557 2191 10560
rect 2133 10551 2191 10557
rect 2314 10548 2320 10560
rect 2372 10548 2378 10600
rect 2590 10520 2596 10532
rect 2148 10492 2596 10520
rect 2148 10464 2176 10492
rect 2590 10480 2596 10492
rect 2648 10520 2654 10532
rect 2700 10520 2728 10619
rect 2774 10616 2780 10668
rect 2832 10656 2838 10668
rect 3620 10665 3648 10696
rect 4062 10684 4068 10736
rect 4120 10724 4126 10736
rect 4525 10727 4583 10733
rect 4525 10724 4537 10727
rect 4120 10696 4537 10724
rect 4120 10684 4126 10696
rect 4525 10693 4537 10696
rect 4571 10693 4583 10727
rect 4525 10687 4583 10693
rect 2869 10659 2927 10665
rect 2869 10656 2881 10659
rect 2832 10628 2881 10656
rect 2832 10616 2838 10628
rect 2869 10625 2881 10628
rect 2915 10625 2927 10659
rect 2869 10619 2927 10625
rect 3605 10659 3663 10665
rect 3605 10625 3617 10659
rect 3651 10625 3663 10659
rect 4540 10656 4568 10687
rect 4614 10684 4620 10736
rect 4672 10724 4678 10736
rect 5077 10727 5135 10733
rect 5077 10724 5089 10727
rect 4672 10696 5089 10724
rect 4672 10684 4678 10696
rect 5077 10693 5089 10696
rect 5123 10693 5135 10727
rect 5077 10687 5135 10693
rect 5718 10656 5724 10668
rect 4540 10628 5724 10656
rect 3605 10619 3663 10625
rect 3326 10548 3332 10600
rect 3384 10588 3390 10600
rect 3513 10591 3571 10597
rect 3513 10588 3525 10591
rect 3384 10560 3525 10588
rect 3384 10548 3390 10560
rect 3513 10557 3525 10560
rect 3559 10557 3571 10591
rect 3620 10588 3648 10619
rect 5718 10616 5724 10628
rect 5776 10616 5782 10668
rect 6546 10616 6552 10668
rect 6604 10656 6610 10668
rect 6932 10665 6960 10764
rect 10870 10752 10876 10764
rect 10928 10752 10934 10804
rect 11149 10795 11207 10801
rect 11149 10761 11161 10795
rect 11195 10792 11207 10795
rect 11882 10792 11888 10804
rect 11195 10764 11888 10792
rect 11195 10761 11207 10764
rect 11149 10755 11207 10761
rect 11882 10752 11888 10764
rect 11940 10792 11946 10804
rect 13354 10792 13360 10804
rect 11940 10764 13360 10792
rect 11940 10752 11946 10764
rect 13354 10752 13360 10764
rect 13412 10752 13418 10804
rect 13630 10792 13636 10804
rect 13591 10764 13636 10792
rect 13630 10752 13636 10764
rect 13688 10752 13694 10804
rect 14461 10795 14519 10801
rect 14461 10761 14473 10795
rect 14507 10792 14519 10795
rect 14826 10792 14832 10804
rect 14507 10764 14832 10792
rect 14507 10761 14519 10764
rect 14461 10755 14519 10761
rect 14826 10752 14832 10764
rect 14884 10752 14890 10804
rect 15746 10792 15752 10804
rect 15707 10764 15752 10792
rect 15746 10752 15752 10764
rect 15804 10752 15810 10804
rect 15933 10795 15991 10801
rect 15933 10761 15945 10795
rect 15979 10792 15991 10795
rect 16206 10792 16212 10804
rect 15979 10764 16212 10792
rect 15979 10761 15991 10764
rect 15933 10755 15991 10761
rect 16206 10752 16212 10764
rect 16264 10752 16270 10804
rect 17586 10752 17592 10804
rect 17644 10792 17650 10804
rect 19150 10792 19156 10804
rect 17644 10764 19156 10792
rect 17644 10752 17650 10764
rect 7006 10684 7012 10736
rect 7064 10724 7070 10736
rect 7147 10727 7205 10733
rect 7147 10724 7159 10727
rect 7064 10696 7109 10724
rect 7064 10684 7070 10696
rect 7142 10693 7159 10724
rect 7193 10724 7205 10727
rect 7193 10696 8248 10724
rect 7193 10693 7205 10696
rect 7142 10687 7205 10693
rect 6825 10659 6883 10665
rect 6825 10656 6837 10659
rect 6604 10628 6837 10656
rect 6604 10616 6610 10628
rect 6825 10625 6837 10628
rect 6871 10625 6883 10659
rect 6825 10619 6883 10625
rect 6917 10659 6975 10665
rect 6917 10625 6929 10659
rect 6963 10625 6975 10659
rect 6917 10619 6975 10625
rect 4614 10588 4620 10600
rect 3620 10560 4620 10588
rect 3513 10551 3571 10557
rect 4614 10548 4620 10560
rect 4672 10548 4678 10600
rect 5350 10548 5356 10600
rect 5408 10588 5414 10600
rect 5626 10588 5632 10600
rect 5408 10560 5632 10588
rect 5408 10548 5414 10560
rect 5626 10548 5632 10560
rect 5684 10588 5690 10600
rect 7142 10588 7170 10687
rect 7926 10656 7932 10668
rect 7887 10628 7932 10656
rect 7926 10616 7932 10628
rect 7984 10616 7990 10668
rect 8021 10659 8079 10665
rect 8021 10625 8033 10659
rect 8067 10625 8079 10659
rect 8021 10619 8079 10625
rect 8113 10659 8171 10665
rect 8113 10625 8125 10659
rect 8159 10625 8171 10659
rect 8113 10619 8171 10625
rect 7282 10588 7288 10600
rect 5684 10560 7170 10588
rect 7243 10560 7288 10588
rect 5684 10548 5690 10560
rect 7282 10548 7288 10560
rect 7340 10548 7346 10600
rect 7742 10548 7748 10600
rect 7800 10588 7806 10600
rect 8036 10588 8064 10619
rect 7800 10560 8064 10588
rect 7800 10548 7806 10560
rect 2648 10492 2728 10520
rect 3973 10523 4031 10529
rect 2648 10480 2654 10492
rect 3973 10489 3985 10523
rect 4019 10520 4031 10523
rect 4154 10520 4160 10532
rect 4019 10492 4160 10520
rect 4019 10489 4031 10492
rect 3973 10483 4031 10489
rect 4154 10480 4160 10492
rect 4212 10480 4218 10532
rect 5534 10480 5540 10532
rect 5592 10520 5598 10532
rect 5592 10492 6040 10520
rect 5592 10480 5598 10492
rect 2130 10452 2136 10464
rect 2091 10424 2136 10452
rect 2130 10412 2136 10424
rect 2188 10412 2194 10464
rect 2869 10455 2927 10461
rect 2869 10421 2881 10455
rect 2915 10452 2927 10455
rect 3510 10452 3516 10464
rect 2915 10424 3516 10452
rect 2915 10421 2927 10424
rect 2869 10415 2927 10421
rect 3510 10412 3516 10424
rect 3568 10412 3574 10464
rect 4798 10412 4804 10464
rect 4856 10452 4862 10464
rect 5261 10455 5319 10461
rect 5261 10452 5273 10455
rect 4856 10424 5273 10452
rect 4856 10412 4862 10424
rect 5261 10421 5273 10424
rect 5307 10421 5319 10455
rect 5261 10415 5319 10421
rect 5445 10455 5503 10461
rect 5445 10421 5457 10455
rect 5491 10452 5503 10455
rect 5810 10452 5816 10464
rect 5491 10424 5816 10452
rect 5491 10421 5503 10424
rect 5445 10415 5503 10421
rect 5810 10412 5816 10424
rect 5868 10412 5874 10464
rect 6012 10461 6040 10492
rect 6822 10480 6828 10532
rect 6880 10520 6886 10532
rect 8128 10520 8156 10619
rect 8220 10588 8248 10696
rect 9122 10684 9128 10736
rect 9180 10724 9186 10736
rect 9217 10727 9275 10733
rect 9217 10724 9229 10727
rect 9180 10696 9229 10724
rect 9180 10684 9186 10696
rect 9217 10693 9229 10696
rect 9263 10693 9275 10727
rect 9217 10687 9275 10693
rect 11698 10684 11704 10736
rect 11756 10724 11762 10736
rect 11977 10727 12035 10733
rect 11977 10724 11989 10727
rect 11756 10696 11989 10724
rect 11756 10684 11762 10696
rect 11977 10693 11989 10696
rect 12023 10724 12035 10727
rect 12894 10724 12900 10736
rect 12023 10696 12900 10724
rect 12023 10693 12035 10696
rect 11977 10687 12035 10693
rect 12894 10684 12900 10696
rect 12952 10684 12958 10736
rect 13801 10727 13859 10733
rect 13801 10693 13813 10727
rect 13847 10724 13859 10727
rect 13906 10724 13912 10736
rect 13847 10696 13912 10724
rect 13847 10693 13859 10696
rect 13801 10687 13859 10693
rect 13906 10684 13912 10696
rect 13964 10684 13970 10736
rect 14001 10727 14059 10733
rect 14001 10693 14013 10727
rect 14047 10724 14059 10727
rect 15470 10724 15476 10736
rect 14047 10696 15476 10724
rect 14047 10693 14059 10696
rect 14001 10687 14059 10693
rect 15470 10684 15476 10696
rect 15528 10684 15534 10736
rect 15562 10684 15568 10736
rect 15620 10724 15626 10736
rect 16117 10727 16175 10733
rect 15620 10696 15976 10724
rect 15620 10684 15626 10696
rect 9033 10659 9091 10665
rect 9033 10625 9045 10659
rect 9079 10656 9091 10659
rect 9306 10656 9312 10668
rect 9079 10628 9312 10656
rect 9079 10625 9091 10628
rect 9033 10619 9091 10625
rect 9306 10616 9312 10628
rect 9364 10616 9370 10668
rect 12437 10659 12495 10665
rect 12437 10625 12449 10659
rect 12483 10656 12495 10659
rect 12713 10659 12771 10665
rect 12483 10628 12517 10656
rect 12483 10625 12495 10628
rect 12437 10619 12495 10625
rect 12713 10625 12725 10659
rect 12759 10656 12771 10659
rect 13078 10656 13084 10668
rect 12759 10628 13084 10656
rect 12759 10625 12771 10628
rect 12713 10619 12771 10625
rect 10042 10588 10048 10600
rect 8220 10560 10048 10588
rect 10042 10548 10048 10560
rect 10100 10588 10106 10600
rect 12452 10588 12480 10619
rect 13078 10616 13084 10628
rect 13136 10616 13142 10668
rect 14642 10616 14648 10668
rect 14700 10656 14706 10668
rect 14737 10659 14795 10665
rect 14737 10656 14749 10659
rect 14700 10628 14749 10656
rect 14700 10616 14706 10628
rect 14737 10625 14749 10628
rect 14783 10625 14795 10659
rect 14737 10619 14795 10625
rect 14829 10659 14887 10665
rect 14829 10625 14841 10659
rect 14875 10625 14887 10659
rect 14829 10619 14887 10625
rect 12802 10588 12808 10600
rect 10100 10560 12808 10588
rect 10100 10548 10106 10560
rect 12802 10548 12808 10560
rect 12860 10548 12866 10600
rect 6880 10492 8156 10520
rect 9401 10523 9459 10529
rect 6880 10480 6886 10492
rect 9401 10489 9413 10523
rect 9447 10520 9459 10523
rect 10226 10520 10232 10532
rect 9447 10492 10232 10520
rect 9447 10489 9459 10492
rect 9401 10483 9459 10489
rect 10226 10480 10232 10492
rect 10284 10480 10290 10532
rect 12621 10523 12679 10529
rect 12621 10489 12633 10523
rect 12667 10520 12679 10523
rect 12894 10520 12900 10532
rect 12667 10492 12900 10520
rect 12667 10489 12679 10492
rect 12621 10483 12679 10489
rect 12894 10480 12900 10492
rect 12952 10480 12958 10532
rect 14844 10520 14872 10619
rect 14918 10616 14924 10668
rect 14976 10656 14982 10668
rect 15105 10659 15163 10665
rect 14976 10628 15021 10656
rect 14976 10616 14982 10628
rect 15105 10625 15117 10659
rect 15151 10625 15163 10659
rect 15105 10619 15163 10625
rect 15010 10548 15016 10600
rect 15068 10588 15074 10600
rect 15120 10588 15148 10619
rect 15378 10616 15384 10668
rect 15436 10656 15442 10668
rect 15841 10659 15899 10665
rect 15841 10656 15853 10659
rect 15436 10628 15853 10656
rect 15436 10616 15442 10628
rect 15841 10625 15853 10628
rect 15887 10625 15899 10659
rect 15948 10656 15976 10696
rect 16117 10693 16129 10727
rect 16163 10724 16175 10727
rect 16390 10724 16396 10736
rect 16163 10696 16396 10724
rect 16163 10693 16175 10696
rect 16117 10687 16175 10693
rect 16390 10684 16396 10696
rect 16448 10684 16454 10736
rect 17037 10727 17095 10733
rect 17037 10693 17049 10727
rect 17083 10724 17095 10727
rect 17126 10724 17132 10736
rect 17083 10696 17132 10724
rect 17083 10693 17095 10696
rect 17037 10687 17095 10693
rect 17126 10684 17132 10696
rect 17184 10684 17190 10736
rect 17696 10696 18645 10724
rect 17696 10665 17724 10696
rect 17681 10659 17739 10665
rect 17681 10656 17693 10659
rect 15948 10628 17693 10656
rect 15841 10619 15899 10625
rect 17681 10625 17693 10628
rect 17727 10625 17739 10659
rect 18046 10656 18052 10668
rect 18007 10628 18052 10656
rect 17681 10619 17739 10625
rect 15068 10560 15148 10588
rect 15856 10588 15884 10619
rect 18046 10616 18052 10628
rect 18104 10616 18110 10668
rect 18617 10659 18645 10696
rect 18693 10659 18751 10665
rect 18617 10631 18705 10659
rect 18693 10625 18705 10631
rect 18739 10625 18751 10659
rect 18693 10619 18751 10625
rect 18877 10659 18935 10665
rect 18877 10625 18889 10659
rect 18923 10656 18935 10659
rect 18984 10656 19012 10764
rect 19150 10752 19156 10764
rect 19208 10752 19214 10804
rect 19337 10795 19395 10801
rect 19337 10761 19349 10795
rect 19383 10792 19395 10795
rect 21634 10792 21640 10804
rect 19383 10764 21640 10792
rect 19383 10761 19395 10764
rect 19337 10755 19395 10761
rect 21634 10752 21640 10764
rect 21692 10752 21698 10804
rect 22554 10792 22560 10804
rect 21744 10764 22560 10792
rect 19168 10702 19334 10724
rect 19150 10690 19156 10702
rect 19119 10662 19156 10690
rect 18923 10628 19012 10656
rect 19150 10650 19156 10662
rect 19208 10696 19334 10702
rect 19208 10665 19214 10696
rect 19208 10659 19233 10665
rect 19168 10628 19187 10650
rect 18923 10625 18935 10628
rect 18877 10619 18935 10625
rect 19175 10625 19187 10628
rect 19221 10625 19233 10659
rect 19306 10656 19334 10696
rect 19978 10684 19984 10736
rect 20036 10724 20042 10736
rect 21269 10727 21327 10733
rect 21269 10724 21281 10727
rect 20036 10696 21281 10724
rect 20036 10684 20042 10696
rect 21269 10693 21281 10696
rect 21315 10724 21327 10727
rect 21744 10724 21772 10764
rect 22554 10752 22560 10764
rect 22612 10752 22618 10804
rect 23106 10792 23112 10804
rect 23032 10764 23112 10792
rect 22830 10724 22836 10736
rect 21315 10696 21772 10724
rect 21836 10696 22836 10724
rect 21315 10693 21327 10696
rect 21269 10687 21327 10693
rect 19702 10656 19708 10668
rect 19306 10628 19708 10656
rect 19175 10619 19233 10625
rect 19702 10616 19708 10628
rect 19760 10616 19766 10668
rect 19794 10616 19800 10668
rect 19852 10656 19858 10668
rect 19889 10659 19947 10665
rect 19889 10656 19901 10659
rect 19852 10628 19901 10656
rect 19852 10616 19858 10628
rect 19889 10625 19901 10628
rect 19935 10625 19947 10659
rect 20070 10656 20076 10668
rect 20031 10628 20076 10656
rect 19889 10619 19947 10625
rect 20070 10616 20076 10628
rect 20128 10616 20134 10668
rect 21542 10616 21548 10668
rect 21600 10656 21606 10668
rect 21836 10656 21864 10696
rect 22830 10684 22836 10696
rect 22888 10724 22894 10736
rect 23032 10733 23060 10764
rect 23106 10752 23112 10764
rect 23164 10752 23170 10804
rect 23017 10727 23075 10733
rect 23017 10724 23029 10727
rect 22888 10696 23029 10724
rect 22888 10684 22894 10696
rect 23017 10693 23029 10696
rect 23063 10693 23075 10727
rect 23017 10687 23075 10693
rect 21600 10628 21864 10656
rect 22281 10659 22339 10665
rect 21600 10616 21606 10628
rect 22281 10625 22293 10659
rect 22327 10656 22339 10659
rect 22646 10656 22652 10668
rect 22327 10628 22652 10656
rect 22327 10625 22339 10628
rect 22281 10619 22339 10625
rect 22646 10616 22652 10628
rect 22704 10616 22710 10668
rect 17586 10588 17592 10600
rect 15856 10560 17592 10588
rect 15068 10548 15074 10560
rect 17586 10548 17592 10560
rect 17644 10548 17650 10600
rect 18233 10591 18291 10597
rect 18233 10557 18245 10591
rect 18279 10588 18291 10591
rect 18598 10588 18604 10600
rect 18279 10560 18604 10588
rect 18279 10557 18291 10560
rect 18233 10551 18291 10557
rect 18598 10548 18604 10560
rect 18656 10548 18662 10600
rect 18969 10591 19027 10597
rect 18969 10557 18981 10591
rect 19015 10588 19027 10591
rect 19610 10588 19616 10600
rect 19015 10560 19616 10588
rect 19015 10557 19027 10560
rect 18969 10551 19027 10557
rect 16666 10520 16672 10532
rect 14844 10492 16672 10520
rect 16666 10480 16672 10492
rect 16724 10480 16730 10532
rect 18046 10480 18052 10532
rect 18104 10520 18110 10532
rect 18984 10520 19012 10551
rect 19610 10548 19616 10560
rect 19668 10588 19674 10600
rect 20530 10588 20536 10600
rect 19668 10560 20536 10588
rect 19668 10548 19674 10560
rect 20530 10548 20536 10560
rect 20588 10548 20594 10600
rect 20714 10548 20720 10600
rect 20772 10588 20778 10600
rect 22097 10591 22155 10597
rect 22097 10588 22109 10591
rect 20772 10560 22109 10588
rect 20772 10548 20778 10560
rect 22097 10557 22109 10560
rect 22143 10557 22155 10591
rect 22097 10551 22155 10557
rect 22189 10591 22247 10597
rect 22189 10557 22201 10591
rect 22235 10557 22247 10591
rect 22189 10551 22247 10557
rect 22373 10591 22431 10597
rect 22373 10557 22385 10591
rect 22419 10588 22431 10591
rect 22462 10588 22468 10600
rect 22419 10560 22468 10588
rect 22419 10557 22431 10560
rect 22373 10551 22431 10557
rect 18104 10492 19012 10520
rect 18104 10480 18110 10492
rect 19058 10480 19064 10532
rect 19116 10520 19122 10532
rect 19116 10492 19161 10520
rect 19116 10480 19122 10492
rect 19242 10480 19248 10532
rect 19300 10520 19306 10532
rect 19981 10523 20039 10529
rect 19981 10520 19993 10523
rect 19300 10492 19993 10520
rect 19300 10480 19306 10492
rect 19981 10489 19993 10492
rect 20027 10489 20039 10523
rect 22204 10520 22232 10551
rect 22462 10548 22468 10560
rect 22520 10548 22526 10600
rect 22204 10492 22416 10520
rect 19981 10483 20039 10489
rect 22388 10464 22416 10492
rect 5997 10455 6055 10461
rect 5997 10421 6009 10455
rect 6043 10452 6055 10455
rect 7282 10452 7288 10464
rect 6043 10424 7288 10452
rect 6043 10421 6055 10424
rect 5997 10415 6055 10421
rect 7282 10412 7288 10424
rect 7340 10412 7346 10464
rect 7650 10412 7656 10464
rect 7708 10452 7714 10464
rect 7745 10455 7803 10461
rect 7745 10452 7757 10455
rect 7708 10424 7757 10452
rect 7708 10412 7714 10424
rect 7745 10421 7757 10424
rect 7791 10421 7803 10455
rect 7745 10415 7803 10421
rect 10413 10455 10471 10461
rect 10413 10421 10425 10455
rect 10459 10452 10471 10455
rect 10502 10452 10508 10464
rect 10459 10424 10508 10452
rect 10459 10421 10471 10424
rect 10413 10415 10471 10421
rect 10502 10412 10508 10424
rect 10560 10412 10566 10464
rect 12250 10412 12256 10464
rect 12308 10452 12314 10464
rect 13446 10452 13452 10464
rect 12308 10424 13452 10452
rect 12308 10412 12314 10424
rect 13446 10412 13452 10424
rect 13504 10412 13510 10464
rect 13817 10455 13875 10461
rect 13817 10421 13829 10455
rect 13863 10452 13875 10455
rect 16482 10452 16488 10464
rect 13863 10424 16488 10452
rect 13863 10421 13875 10424
rect 13817 10415 13875 10421
rect 16482 10412 16488 10424
rect 16540 10412 16546 10464
rect 17402 10412 17408 10464
rect 17460 10452 17466 10464
rect 19518 10452 19524 10464
rect 17460 10424 19524 10452
rect 17460 10412 17466 10424
rect 19518 10412 19524 10424
rect 19576 10412 19582 10464
rect 19794 10412 19800 10464
rect 19852 10452 19858 10464
rect 20809 10455 20867 10461
rect 20809 10452 20821 10455
rect 19852 10424 20821 10452
rect 19852 10412 19858 10424
rect 20809 10421 20821 10424
rect 20855 10452 20867 10455
rect 21542 10452 21548 10464
rect 20855 10424 21548 10452
rect 20855 10421 20867 10424
rect 20809 10415 20867 10421
rect 21542 10412 21548 10424
rect 21600 10412 21606 10464
rect 22370 10412 22376 10464
rect 22428 10412 22434 10464
rect 22554 10452 22560 10464
rect 22515 10424 22560 10452
rect 22554 10412 22560 10424
rect 22612 10412 22618 10464
rect 1104 10362 23828 10384
rect 1104 10310 3790 10362
rect 3842 10310 3854 10362
rect 3906 10310 3918 10362
rect 3970 10310 3982 10362
rect 4034 10310 4046 10362
rect 4098 10310 9471 10362
rect 9523 10310 9535 10362
rect 9587 10310 9599 10362
rect 9651 10310 9663 10362
rect 9715 10310 9727 10362
rect 9779 10310 15152 10362
rect 15204 10310 15216 10362
rect 15268 10310 15280 10362
rect 15332 10310 15344 10362
rect 15396 10310 15408 10362
rect 15460 10310 20833 10362
rect 20885 10310 20897 10362
rect 20949 10310 20961 10362
rect 21013 10310 21025 10362
rect 21077 10310 21089 10362
rect 21141 10310 23828 10362
rect 1104 10288 23828 10310
rect 2498 10208 2504 10260
rect 2556 10248 2562 10260
rect 4801 10251 4859 10257
rect 4801 10248 4813 10251
rect 2556 10220 4813 10248
rect 2556 10208 2562 10220
rect 4801 10217 4813 10220
rect 4847 10217 4859 10251
rect 4801 10211 4859 10217
rect 4982 10208 4988 10260
rect 5040 10248 5046 10260
rect 6181 10251 6239 10257
rect 6181 10248 6193 10251
rect 5040 10220 6193 10248
rect 5040 10208 5046 10220
rect 6181 10217 6193 10220
rect 6227 10217 6239 10251
rect 6181 10211 6239 10217
rect 6454 10208 6460 10260
rect 6512 10248 6518 10260
rect 8570 10248 8576 10260
rect 6512 10220 8432 10248
rect 8531 10220 8576 10248
rect 6512 10208 6518 10220
rect 2225 10183 2283 10189
rect 2225 10149 2237 10183
rect 2271 10180 2283 10183
rect 2682 10180 2688 10192
rect 2271 10152 2688 10180
rect 2271 10149 2283 10152
rect 2225 10143 2283 10149
rect 2682 10140 2688 10152
rect 2740 10140 2746 10192
rect 3050 10140 3056 10192
rect 3108 10180 3114 10192
rect 4341 10183 4399 10189
rect 4341 10180 4353 10183
rect 3108 10152 4353 10180
rect 3108 10140 3114 10152
rect 4341 10149 4353 10152
rect 4387 10180 4399 10183
rect 5534 10180 5540 10192
rect 4387 10152 5540 10180
rect 4387 10149 4399 10152
rect 4341 10143 4399 10149
rect 5534 10140 5540 10152
rect 5592 10140 5598 10192
rect 6270 10140 6276 10192
rect 6328 10180 6334 10192
rect 6328 10152 6684 10180
rect 6328 10140 6334 10152
rect 3326 10112 3332 10124
rect 2332 10084 3332 10112
rect 2332 10053 2360 10084
rect 3326 10072 3332 10084
rect 3384 10072 3390 10124
rect 4154 10072 4160 10124
rect 4212 10112 4218 10124
rect 6656 10121 6684 10152
rect 7098 10140 7104 10192
rect 7156 10180 7162 10192
rect 7558 10180 7564 10192
rect 7156 10152 7564 10180
rect 7156 10140 7162 10152
rect 7558 10140 7564 10152
rect 7616 10140 7622 10192
rect 8404 10180 8432 10220
rect 8570 10208 8576 10220
rect 8628 10208 8634 10260
rect 13538 10248 13544 10260
rect 13499 10220 13544 10248
rect 13538 10208 13544 10220
rect 13596 10208 13602 10260
rect 13906 10208 13912 10260
rect 13964 10248 13970 10260
rect 14921 10251 14979 10257
rect 14921 10248 14933 10251
rect 13964 10220 14933 10248
rect 13964 10208 13970 10220
rect 14921 10217 14933 10220
rect 14967 10217 14979 10251
rect 15746 10248 15752 10260
rect 14921 10211 14979 10217
rect 15028 10220 15752 10248
rect 10505 10183 10563 10189
rect 10505 10180 10517 10183
rect 8404 10152 10517 10180
rect 10505 10149 10517 10152
rect 10551 10149 10563 10183
rect 12250 10180 12256 10192
rect 12211 10152 12256 10180
rect 10505 10143 10563 10149
rect 12250 10140 12256 10152
rect 12308 10140 12314 10192
rect 13354 10140 13360 10192
rect 13412 10180 13418 10192
rect 14369 10183 14427 10189
rect 14369 10180 14381 10183
rect 13412 10152 14381 10180
rect 13412 10140 13418 10152
rect 14369 10149 14381 10152
rect 14415 10180 14427 10183
rect 15028 10180 15056 10220
rect 15746 10208 15752 10220
rect 15804 10208 15810 10260
rect 17678 10248 17684 10260
rect 17639 10220 17684 10248
rect 17678 10208 17684 10220
rect 17736 10208 17742 10260
rect 18506 10248 18512 10260
rect 17788 10220 18512 10248
rect 15654 10180 15660 10192
rect 14415 10152 15056 10180
rect 15212 10152 15660 10180
rect 14415 10149 14427 10152
rect 14369 10143 14427 10149
rect 6365 10115 6423 10121
rect 6365 10112 6377 10115
rect 4212 10084 6377 10112
rect 4212 10072 4218 10084
rect 6365 10081 6377 10084
rect 6411 10081 6423 10115
rect 6365 10075 6423 10081
rect 6641 10115 6699 10121
rect 6641 10081 6653 10115
rect 6687 10081 6699 10115
rect 6641 10075 6699 10081
rect 6822 10072 6828 10124
rect 6880 10112 6886 10124
rect 7929 10115 7987 10121
rect 7929 10112 7941 10115
rect 6880 10084 7941 10112
rect 6880 10072 6886 10084
rect 7929 10081 7941 10084
rect 7975 10081 7987 10115
rect 7929 10075 7987 10081
rect 8018 10072 8024 10124
rect 8076 10112 8082 10124
rect 8113 10115 8171 10121
rect 8113 10112 8125 10115
rect 8076 10084 8125 10112
rect 8076 10072 8082 10084
rect 8113 10081 8125 10084
rect 8159 10081 8171 10115
rect 8113 10075 8171 10081
rect 9674 10072 9680 10124
rect 9732 10112 9738 10124
rect 12897 10115 12955 10121
rect 9732 10084 11100 10112
rect 9732 10072 9738 10084
rect 2317 10047 2375 10053
rect 2317 10013 2329 10047
rect 2363 10013 2375 10047
rect 2317 10007 2375 10013
rect 2501 10047 2559 10053
rect 2501 10013 2513 10047
rect 2547 10044 2559 10047
rect 3050 10044 3056 10056
rect 2547 10016 3056 10044
rect 2547 10013 2559 10016
rect 2501 10007 2559 10013
rect 3050 10004 3056 10016
rect 3108 10004 3114 10056
rect 3418 10044 3424 10056
rect 3379 10016 3424 10044
rect 3418 10004 3424 10016
rect 3476 10004 3482 10056
rect 4985 10047 5043 10053
rect 4985 10013 4997 10047
rect 5031 10013 5043 10047
rect 4985 10007 5043 10013
rect 3145 9979 3203 9985
rect 3145 9945 3157 9979
rect 3191 9976 3203 9979
rect 3234 9976 3240 9988
rect 3191 9948 3240 9976
rect 3191 9945 3203 9948
rect 3145 9939 3203 9945
rect 3234 9936 3240 9948
rect 3292 9936 3298 9988
rect 1670 9908 1676 9920
rect 1631 9880 1676 9908
rect 1670 9868 1676 9880
rect 1728 9868 1734 9920
rect 5000 9908 5028 10007
rect 5074 10004 5080 10056
rect 5132 10044 5138 10056
rect 5350 10053 5356 10056
rect 5307 10047 5356 10053
rect 5132 10016 5177 10044
rect 5132 10004 5138 10016
rect 5307 10013 5319 10047
rect 5353 10013 5356 10047
rect 5307 10007 5356 10013
rect 5350 10004 5356 10007
rect 5408 10004 5414 10056
rect 5445 10047 5503 10053
rect 5445 10013 5457 10047
rect 5491 10044 5503 10047
rect 5534 10044 5540 10056
rect 5491 10016 5540 10044
rect 5491 10013 5503 10016
rect 5445 10007 5503 10013
rect 5534 10004 5540 10016
rect 5592 10044 5598 10056
rect 6178 10044 6184 10056
rect 5592 10016 6184 10044
rect 5592 10004 5598 10016
rect 6178 10004 6184 10016
rect 6236 10004 6242 10056
rect 6457 10047 6515 10053
rect 6457 10013 6469 10047
rect 6503 10013 6515 10047
rect 6457 10007 6515 10013
rect 6549 10047 6607 10053
rect 6549 10013 6561 10047
rect 6595 10044 6607 10047
rect 7190 10044 7196 10056
rect 6595 10016 7196 10044
rect 6595 10013 6607 10016
rect 6549 10007 6607 10013
rect 5169 9979 5227 9985
rect 5169 9945 5181 9979
rect 5215 9945 5227 9979
rect 5994 9976 6000 9988
rect 5169 9939 5227 9945
rect 5460 9948 6000 9976
rect 5074 9908 5080 9920
rect 5000 9880 5080 9908
rect 5074 9868 5080 9880
rect 5132 9868 5138 9920
rect 5184 9908 5212 9939
rect 5460 9908 5488 9948
rect 5994 9936 6000 9948
rect 6052 9936 6058 9988
rect 6472 9976 6500 10007
rect 7190 10004 7196 10016
rect 7248 10044 7254 10056
rect 7834 10044 7840 10056
rect 7248 10016 7840 10044
rect 7248 10004 7254 10016
rect 7834 10004 7840 10016
rect 7892 10004 7898 10056
rect 9122 10044 9128 10056
rect 9083 10016 9128 10044
rect 9122 10004 9128 10016
rect 9180 10004 9186 10056
rect 9306 10004 9312 10056
rect 9364 10044 9370 10056
rect 9769 10047 9827 10053
rect 9769 10044 9781 10047
rect 9364 10016 9781 10044
rect 9364 10004 9370 10016
rect 9769 10013 9781 10016
rect 9815 10013 9827 10047
rect 9769 10007 9827 10013
rect 10042 10004 10048 10056
rect 10100 10044 10106 10056
rect 11072 10053 11100 10084
rect 12897 10081 12909 10115
rect 12943 10112 12955 10115
rect 13722 10112 13728 10124
rect 12943 10084 13728 10112
rect 12943 10081 12955 10084
rect 12897 10075 12955 10081
rect 13722 10072 13728 10084
rect 13780 10072 13786 10124
rect 10689 10047 10747 10053
rect 10689 10044 10701 10047
rect 10100 10016 10701 10044
rect 10100 10004 10106 10016
rect 10689 10013 10701 10016
rect 10735 10013 10747 10047
rect 10689 10007 10747 10013
rect 11057 10047 11115 10053
rect 11057 10013 11069 10047
rect 11103 10013 11115 10047
rect 11057 10007 11115 10013
rect 12437 10047 12495 10053
rect 12437 10013 12449 10047
rect 12483 10013 12495 10047
rect 12437 10007 12495 10013
rect 7650 9976 7656 9988
rect 6472 9948 7656 9976
rect 7650 9936 7656 9948
rect 7708 9936 7714 9988
rect 9585 9979 9643 9985
rect 9585 9945 9597 9979
rect 9631 9976 9643 9979
rect 10594 9976 10600 9988
rect 9631 9948 10600 9976
rect 9631 9945 9643 9948
rect 9585 9939 9643 9945
rect 10594 9936 10600 9948
rect 10652 9936 10658 9988
rect 10781 9979 10839 9985
rect 10781 9945 10793 9979
rect 10827 9945 10839 9979
rect 10781 9939 10839 9945
rect 10873 9979 10931 9985
rect 10873 9945 10885 9979
rect 10919 9945 10931 9979
rect 12452 9976 12480 10007
rect 12710 10004 12716 10056
rect 12768 10044 12774 10056
rect 12805 10047 12863 10053
rect 12805 10044 12817 10047
rect 12768 10016 12817 10044
rect 12768 10004 12774 10016
rect 12805 10013 12817 10016
rect 12851 10044 12863 10047
rect 12986 10044 12992 10056
rect 12851 10016 12992 10044
rect 12851 10013 12863 10016
rect 12805 10007 12863 10013
rect 12986 10004 12992 10016
rect 13044 10004 13050 10056
rect 14734 10004 14740 10056
rect 14792 10044 14798 10056
rect 15212 10053 15240 10152
rect 15654 10140 15660 10152
rect 15712 10180 15718 10192
rect 17788 10180 17816 10220
rect 18506 10208 18512 10220
rect 18564 10208 18570 10260
rect 21637 10251 21695 10257
rect 21637 10217 21649 10251
rect 21683 10248 21695 10251
rect 22094 10248 22100 10260
rect 21683 10220 22100 10248
rect 21683 10217 21695 10220
rect 21637 10211 21695 10217
rect 22094 10208 22100 10220
rect 22152 10208 22158 10260
rect 15712 10152 17816 10180
rect 15712 10140 15718 10152
rect 17862 10140 17868 10192
rect 17920 10180 17926 10192
rect 19429 10183 19487 10189
rect 19429 10180 19441 10183
rect 17920 10152 19441 10180
rect 17920 10140 17926 10152
rect 19429 10149 19441 10152
rect 19475 10149 19487 10183
rect 19429 10143 19487 10149
rect 20625 10183 20683 10189
rect 20625 10149 20637 10183
rect 20671 10180 20683 10183
rect 22002 10180 22008 10192
rect 20671 10152 22008 10180
rect 20671 10149 20683 10152
rect 20625 10143 20683 10149
rect 22002 10140 22008 10152
rect 22060 10140 22066 10192
rect 22738 10180 22744 10192
rect 22113 10152 22744 10180
rect 16390 10112 16396 10124
rect 15396 10084 16396 10112
rect 15396 10053 15424 10084
rect 16390 10072 16396 10084
rect 16448 10072 16454 10124
rect 18874 10112 18880 10124
rect 17236 10084 18880 10112
rect 15105 10047 15163 10053
rect 15105 10044 15117 10047
rect 14792 10016 15117 10044
rect 14792 10004 14798 10016
rect 15105 10013 15117 10016
rect 15151 10013 15163 10047
rect 15105 10007 15163 10013
rect 15197 10047 15255 10053
rect 15197 10013 15209 10047
rect 15243 10013 15255 10047
rect 15197 10007 15255 10013
rect 15381 10047 15439 10053
rect 15381 10013 15393 10047
rect 15427 10013 15439 10047
rect 15381 10007 15439 10013
rect 15473 10047 15531 10053
rect 15473 10013 15485 10047
rect 15519 10013 15531 10047
rect 15473 10007 15531 10013
rect 13262 9976 13268 9988
rect 12452 9948 13268 9976
rect 10873 9939 10931 9945
rect 5184 9880 5488 9908
rect 5810 9868 5816 9920
rect 5868 9908 5874 9920
rect 6822 9908 6828 9920
rect 5868 9880 6828 9908
rect 5868 9868 5874 9880
rect 6822 9868 6828 9880
rect 6880 9868 6886 9920
rect 7374 9908 7380 9920
rect 7335 9880 7380 9908
rect 7374 9868 7380 9880
rect 7432 9868 7438 9920
rect 7558 9868 7564 9920
rect 7616 9908 7622 9920
rect 7926 9908 7932 9920
rect 7616 9880 7932 9908
rect 7616 9868 7622 9880
rect 7926 9868 7932 9880
rect 7984 9908 7990 9920
rect 8205 9911 8263 9917
rect 8205 9908 8217 9911
rect 7984 9880 8217 9908
rect 7984 9868 7990 9880
rect 8205 9877 8217 9880
rect 8251 9877 8263 9911
rect 8205 9871 8263 9877
rect 10502 9868 10508 9920
rect 10560 9908 10566 9920
rect 10796 9908 10824 9939
rect 10560 9880 10824 9908
rect 10888 9908 10916 9939
rect 13262 9936 13268 9948
rect 13320 9936 13326 9988
rect 14458 9936 14464 9988
rect 14516 9976 14522 9988
rect 15010 9976 15016 9988
rect 14516 9948 15016 9976
rect 14516 9936 14522 9948
rect 15010 9936 15016 9948
rect 15068 9976 15074 9988
rect 15488 9976 15516 10007
rect 16022 10004 16028 10056
rect 16080 10044 16086 10056
rect 16117 10047 16175 10053
rect 16117 10044 16129 10047
rect 16080 10016 16129 10044
rect 16080 10004 16086 10016
rect 16117 10013 16129 10016
rect 16163 10013 16175 10047
rect 16117 10007 16175 10013
rect 16301 10047 16359 10053
rect 16301 10013 16313 10047
rect 16347 10013 16359 10047
rect 16301 10007 16359 10013
rect 15068 9948 15516 9976
rect 15068 9936 15074 9948
rect 12710 9908 12716 9920
rect 10888 9880 12716 9908
rect 10560 9868 10566 9880
rect 12710 9868 12716 9880
rect 12768 9868 12774 9920
rect 14642 9868 14648 9920
rect 14700 9908 14706 9920
rect 15562 9908 15568 9920
rect 14700 9880 15568 9908
rect 14700 9868 14706 9880
rect 15562 9868 15568 9880
rect 15620 9868 15626 9920
rect 16316 9908 16344 10007
rect 16758 10004 16764 10056
rect 16816 10044 16822 10056
rect 17236 10053 17264 10084
rect 18874 10072 18880 10084
rect 18932 10072 18938 10124
rect 20438 10112 20444 10124
rect 20180 10084 20444 10112
rect 17129 10047 17187 10053
rect 17129 10044 17141 10047
rect 16816 10016 17141 10044
rect 16816 10004 16822 10016
rect 17129 10013 17141 10016
rect 17175 10013 17187 10047
rect 17129 10007 17187 10013
rect 17221 10047 17279 10053
rect 17221 10013 17233 10047
rect 17267 10013 17279 10047
rect 17402 10044 17408 10056
rect 17363 10016 17408 10044
rect 17221 10007 17279 10013
rect 17402 10004 17408 10016
rect 17460 10004 17466 10056
rect 17494 10004 17500 10056
rect 17552 10044 17558 10056
rect 18138 10044 18144 10056
rect 17552 10016 17597 10044
rect 18099 10016 18144 10044
rect 17552 10004 17558 10016
rect 18138 10004 18144 10016
rect 18196 10004 18202 10056
rect 18233 10047 18291 10053
rect 18233 10013 18245 10047
rect 18279 10013 18291 10047
rect 18233 10007 18291 10013
rect 16666 9976 16672 9988
rect 16627 9948 16672 9976
rect 16666 9936 16672 9948
rect 16724 9936 16730 9988
rect 16942 9976 16948 9988
rect 16776 9948 16948 9976
rect 16776 9908 16804 9948
rect 16942 9936 16948 9948
rect 17000 9976 17006 9988
rect 17862 9976 17868 9988
rect 17000 9948 17868 9976
rect 17000 9936 17006 9948
rect 17862 9936 17868 9948
rect 17920 9936 17926 9988
rect 18248 9976 18276 10007
rect 18322 10004 18328 10056
rect 18380 10044 18386 10056
rect 18417 10047 18475 10053
rect 18417 10044 18429 10047
rect 18380 10016 18429 10044
rect 18380 10004 18386 10016
rect 18417 10013 18429 10016
rect 18463 10044 18475 10047
rect 19150 10044 19156 10056
rect 18463 10016 19156 10044
rect 18463 10013 18475 10016
rect 18417 10007 18475 10013
rect 19150 10004 19156 10016
rect 19208 10004 19214 10056
rect 19981 10047 20039 10053
rect 19981 10013 19993 10047
rect 20027 10044 20039 10047
rect 20070 10044 20076 10056
rect 20027 10016 20076 10044
rect 20027 10013 20039 10016
rect 19981 10007 20039 10013
rect 20070 10004 20076 10016
rect 20128 10004 20134 10056
rect 20180 10053 20208 10084
rect 20438 10072 20444 10084
rect 20496 10072 20502 10124
rect 22113 10056 22141 10152
rect 22738 10140 22744 10152
rect 22796 10140 22802 10192
rect 22186 10072 22192 10124
rect 22244 10112 22250 10124
rect 22649 10115 22707 10121
rect 22649 10112 22661 10115
rect 22244 10084 22661 10112
rect 22244 10072 22250 10084
rect 22649 10081 22661 10084
rect 22695 10081 22707 10115
rect 22649 10075 22707 10081
rect 20165 10047 20223 10053
rect 20165 10013 20177 10047
rect 20211 10013 20223 10047
rect 20165 10007 20223 10013
rect 20257 10047 20315 10053
rect 20257 10013 20269 10047
rect 20303 10013 20315 10047
rect 20257 10007 20315 10013
rect 18690 9976 18696 9988
rect 18248 9948 18696 9976
rect 18690 9936 18696 9948
rect 18748 9936 18754 9988
rect 20180 9976 20208 10007
rect 19904 9948 20208 9976
rect 16316 9880 16804 9908
rect 17218 9868 17224 9920
rect 17276 9908 17282 9920
rect 17586 9908 17592 9920
rect 17276 9880 17592 9908
rect 17276 9868 17282 9880
rect 17586 9868 17592 9880
rect 17644 9908 17650 9920
rect 19904 9908 19932 9948
rect 17644 9880 19932 9908
rect 17644 9868 17650 9880
rect 19978 9868 19984 9920
rect 20036 9908 20042 9920
rect 20272 9908 20300 10007
rect 20346 10004 20352 10056
rect 20404 10044 20410 10056
rect 21174 10044 21180 10056
rect 20404 10016 21180 10044
rect 20404 10004 20410 10016
rect 21174 10004 21180 10016
rect 21232 10004 21238 10056
rect 21542 10044 21548 10056
rect 21503 10016 21548 10044
rect 21542 10004 21548 10016
rect 21600 10004 21606 10056
rect 22094 10044 22100 10056
rect 22008 10016 22100 10044
rect 22094 10004 22100 10016
rect 22152 10044 22158 10056
rect 22373 10047 22431 10053
rect 22373 10044 22385 10047
rect 22152 10016 22385 10044
rect 22152 10004 22158 10016
rect 22373 10013 22385 10016
rect 22419 10013 22431 10047
rect 22373 10007 22431 10013
rect 22465 10047 22523 10053
rect 22465 10013 22477 10047
rect 22511 10013 22523 10047
rect 22465 10007 22523 10013
rect 22557 10047 22615 10053
rect 22557 10013 22569 10047
rect 22603 10044 22615 10047
rect 23014 10044 23020 10056
rect 22603 10016 23020 10044
rect 22603 10013 22615 10016
rect 22557 10007 22615 10013
rect 20036 9880 20300 9908
rect 20036 9868 20042 9880
rect 21450 9868 21456 9920
rect 21508 9908 21514 9920
rect 22189 9911 22247 9917
rect 22189 9908 22201 9911
rect 21508 9880 22201 9908
rect 21508 9868 21514 9880
rect 22189 9877 22201 9880
rect 22235 9877 22247 9911
rect 22480 9908 22508 10007
rect 23014 10004 23020 10016
rect 23072 10004 23078 10056
rect 22646 9908 22652 9920
rect 22480 9880 22652 9908
rect 22189 9871 22247 9877
rect 22646 9868 22652 9880
rect 22704 9868 22710 9920
rect 23198 9908 23204 9920
rect 23159 9880 23204 9908
rect 23198 9868 23204 9880
rect 23256 9868 23262 9920
rect 1104 9818 23987 9840
rect 1104 9766 6630 9818
rect 6682 9766 6694 9818
rect 6746 9766 6758 9818
rect 6810 9766 6822 9818
rect 6874 9766 6886 9818
rect 6938 9766 12311 9818
rect 12363 9766 12375 9818
rect 12427 9766 12439 9818
rect 12491 9766 12503 9818
rect 12555 9766 12567 9818
rect 12619 9766 17992 9818
rect 18044 9766 18056 9818
rect 18108 9766 18120 9818
rect 18172 9766 18184 9818
rect 18236 9766 18248 9818
rect 18300 9766 23673 9818
rect 23725 9766 23737 9818
rect 23789 9766 23801 9818
rect 23853 9766 23865 9818
rect 23917 9766 23929 9818
rect 23981 9766 23987 9818
rect 1104 9744 23987 9766
rect 7282 9704 7288 9716
rect 5368 9676 7288 9704
rect 1673 9639 1731 9645
rect 1673 9605 1685 9639
rect 1719 9636 1731 9639
rect 2774 9636 2780 9648
rect 1719 9608 2780 9636
rect 1719 9605 1731 9608
rect 1673 9599 1731 9605
rect 2774 9596 2780 9608
rect 2832 9596 2838 9648
rect 2869 9639 2927 9645
rect 2869 9605 2881 9639
rect 2915 9636 2927 9639
rect 3142 9636 3148 9648
rect 2915 9608 3148 9636
rect 2915 9605 2927 9608
rect 2869 9599 2927 9605
rect 3142 9596 3148 9608
rect 3200 9596 3206 9648
rect 4246 9596 4252 9648
rect 4304 9636 4310 9648
rect 4816 9646 5028 9674
rect 5368 9648 5396 9676
rect 7282 9664 7288 9676
rect 7340 9664 7346 9716
rect 7558 9664 7564 9716
rect 7616 9704 7622 9716
rect 7834 9704 7840 9716
rect 7616 9676 7840 9704
rect 7616 9664 7622 9676
rect 7834 9664 7840 9676
rect 7892 9704 7898 9716
rect 9033 9707 9091 9713
rect 9033 9704 9045 9707
rect 7892 9676 9045 9704
rect 7892 9664 7898 9676
rect 4617 9639 4675 9645
rect 4617 9636 4629 9639
rect 4304 9608 4629 9636
rect 4304 9596 4310 9608
rect 4617 9605 4629 9608
rect 4663 9636 4675 9639
rect 4816 9636 4844 9646
rect 4663 9608 4844 9636
rect 5000 9636 5028 9646
rect 5074 9636 5080 9648
rect 5000 9608 5080 9636
rect 4663 9605 4675 9608
rect 4617 9599 4675 9605
rect 5074 9596 5080 9608
rect 5132 9596 5138 9648
rect 5350 9596 5356 9648
rect 5408 9596 5414 9648
rect 5902 9636 5908 9648
rect 5863 9608 5908 9636
rect 5902 9596 5908 9608
rect 5960 9596 5966 9648
rect 7006 9596 7012 9648
rect 7064 9636 7070 9648
rect 7064 9608 7880 9636
rect 7064 9596 7070 9608
rect 1857 9571 1915 9577
rect 1857 9537 1869 9571
rect 1903 9537 1915 9571
rect 1857 9531 1915 9537
rect 2041 9571 2099 9577
rect 2041 9537 2053 9571
rect 2087 9568 2099 9571
rect 2222 9568 2228 9580
rect 2087 9540 2228 9568
rect 2087 9537 2099 9540
rect 2041 9531 2099 9537
rect 1872 9500 1900 9531
rect 2222 9528 2228 9540
rect 2280 9528 2286 9580
rect 3418 9568 3424 9580
rect 2792 9540 3424 9568
rect 1946 9500 1952 9512
rect 1859 9472 1952 9500
rect 1946 9460 1952 9472
rect 2004 9500 2010 9512
rect 2792 9500 2820 9540
rect 3418 9528 3424 9540
rect 3476 9568 3482 9580
rect 3697 9571 3755 9577
rect 3476 9566 3556 9568
rect 3697 9566 3709 9571
rect 3476 9540 3709 9566
rect 3476 9528 3482 9540
rect 3528 9538 3709 9540
rect 3697 9537 3709 9538
rect 3743 9537 3755 9571
rect 3697 9531 3755 9537
rect 3789 9571 3847 9577
rect 3789 9537 3801 9571
rect 3835 9566 3847 9571
rect 4154 9568 4160 9580
rect 3896 9566 4160 9568
rect 3835 9540 4160 9566
rect 3835 9538 3924 9540
rect 3835 9537 3847 9538
rect 3789 9531 3847 9537
rect 4154 9528 4160 9540
rect 4212 9528 4218 9580
rect 4801 9571 4859 9577
rect 4724 9568 4813 9571
rect 4632 9543 4813 9568
rect 4632 9540 4752 9543
rect 4632 9512 4660 9540
rect 4801 9537 4813 9543
rect 4847 9537 4859 9571
rect 4801 9531 4859 9537
rect 4893 9571 4951 9577
rect 4893 9537 4905 9571
rect 4939 9537 4951 9571
rect 4893 9531 4951 9537
rect 5445 9571 5503 9577
rect 5445 9537 5457 9571
rect 5491 9568 5503 9571
rect 7466 9568 7472 9580
rect 5491 9540 7472 9568
rect 5491 9537 5503 9540
rect 5445 9531 5503 9537
rect 2004 9472 2820 9500
rect 2004 9460 2010 9472
rect 2240 9444 2268 9472
rect 3326 9460 3332 9512
rect 3384 9500 3390 9512
rect 3512 9503 3570 9509
rect 3512 9500 3524 9503
rect 3384 9472 3524 9500
rect 3384 9460 3390 9472
rect 3512 9469 3524 9472
rect 3558 9469 3570 9503
rect 3512 9463 3570 9469
rect 3605 9503 3663 9509
rect 3605 9469 3617 9503
rect 3651 9469 3663 9503
rect 3605 9463 3663 9469
rect 2222 9392 2228 9444
rect 2280 9392 2286 9444
rect 2685 9435 2743 9441
rect 2685 9401 2697 9435
rect 2731 9432 2743 9435
rect 2866 9432 2872 9444
rect 2731 9404 2872 9432
rect 2731 9401 2743 9404
rect 2685 9395 2743 9401
rect 2866 9392 2872 9404
rect 2924 9392 2930 9444
rect 3234 9392 3240 9444
rect 3292 9432 3298 9444
rect 3620 9432 3648 9463
rect 4614 9460 4620 9512
rect 4672 9460 4678 9512
rect 3292 9404 3648 9432
rect 3292 9392 3298 9404
rect 3786 9324 3792 9376
rect 3844 9364 3850 9376
rect 3973 9367 4031 9373
rect 3973 9364 3985 9367
rect 3844 9336 3985 9364
rect 3844 9324 3850 9336
rect 3973 9333 3985 9336
rect 4019 9333 4031 9367
rect 4706 9364 4712 9376
rect 4667 9336 4712 9364
rect 3973 9327 4031 9333
rect 4706 9324 4712 9336
rect 4764 9324 4770 9376
rect 4908 9364 4936 9531
rect 7466 9528 7472 9540
rect 7524 9528 7530 9580
rect 7650 9568 7656 9580
rect 7611 9540 7656 9568
rect 7650 9528 7656 9540
rect 7708 9528 7714 9580
rect 7852 9577 7880 9608
rect 8036 9577 8064 9676
rect 9033 9673 9045 9676
rect 9079 9673 9091 9707
rect 9033 9667 9091 9673
rect 14461 9707 14519 9713
rect 14461 9673 14473 9707
rect 14507 9704 14519 9707
rect 15470 9704 15476 9716
rect 14507 9676 15476 9704
rect 14507 9673 14519 9676
rect 14461 9667 14519 9673
rect 15470 9664 15476 9676
rect 15528 9664 15534 9716
rect 15562 9664 15568 9716
rect 15620 9704 15626 9716
rect 23198 9704 23204 9716
rect 15620 9676 23204 9704
rect 15620 9664 15626 9676
rect 8297 9639 8355 9645
rect 8297 9605 8309 9639
rect 8343 9636 8355 9639
rect 9674 9636 9680 9648
rect 8343 9608 9680 9636
rect 8343 9605 8355 9608
rect 8297 9599 8355 9605
rect 9674 9596 9680 9608
rect 9732 9596 9738 9648
rect 12161 9639 12219 9645
rect 12161 9605 12173 9639
rect 12207 9636 12219 9639
rect 12986 9636 12992 9648
rect 12207 9608 12992 9636
rect 12207 9605 12219 9608
rect 12161 9599 12219 9605
rect 12986 9596 12992 9608
rect 13044 9596 13050 9648
rect 16132 9645 16160 9676
rect 23198 9664 23204 9676
rect 23256 9664 23262 9716
rect 16117 9639 16175 9645
rect 16117 9605 16129 9639
rect 16163 9605 16175 9639
rect 16117 9599 16175 9605
rect 16482 9596 16488 9648
rect 16540 9636 16546 9648
rect 16540 9608 17044 9636
rect 16540 9596 16546 9608
rect 7837 9571 7895 9577
rect 7837 9537 7849 9571
rect 7883 9537 7895 9571
rect 7837 9531 7895 9537
rect 7929 9571 7987 9577
rect 7929 9537 7941 9571
rect 7975 9537 7987 9571
rect 7929 9531 7987 9537
rect 8021 9571 8079 9577
rect 8021 9537 8033 9571
rect 8067 9537 8079 9571
rect 8021 9531 8079 9537
rect 8849 9571 8907 9577
rect 8849 9537 8861 9571
rect 8895 9568 8907 9571
rect 9122 9568 9128 9580
rect 8895 9540 9128 9568
rect 8895 9537 8907 9540
rect 8849 9531 8907 9537
rect 5718 9460 5724 9512
rect 5776 9500 5782 9512
rect 5813 9503 5871 9509
rect 5813 9500 5825 9503
rect 5776 9472 5825 9500
rect 5776 9460 5782 9472
rect 5813 9469 5825 9472
rect 5859 9469 5871 9503
rect 5813 9463 5871 9469
rect 7742 9460 7748 9512
rect 7800 9500 7806 9512
rect 7944 9500 7972 9531
rect 7800 9472 7972 9500
rect 7800 9460 7806 9472
rect 5902 9392 5908 9444
rect 5960 9432 5966 9444
rect 8864 9432 8892 9531
rect 9122 9528 9128 9540
rect 9180 9528 9186 9580
rect 9950 9528 9956 9580
rect 10008 9568 10014 9580
rect 10045 9571 10103 9577
rect 10045 9568 10057 9571
rect 10008 9540 10057 9568
rect 10008 9528 10014 9540
rect 10045 9537 10057 9540
rect 10091 9537 10103 9571
rect 10962 9568 10968 9580
rect 10923 9540 10968 9568
rect 10045 9531 10103 9537
rect 10962 9528 10968 9540
rect 11020 9528 11026 9580
rect 11054 9528 11060 9580
rect 11112 9568 11118 9580
rect 13630 9568 13636 9580
rect 11112 9540 13492 9568
rect 13591 9540 13636 9568
rect 11112 9528 11118 9540
rect 9306 9460 9312 9512
rect 9364 9500 9370 9512
rect 9364 9472 9457 9500
rect 9364 9460 9370 9472
rect 9490 9460 9496 9512
rect 9548 9500 9554 9512
rect 10229 9503 10287 9509
rect 10229 9500 10241 9503
rect 9548 9472 10241 9500
rect 9548 9460 9554 9472
rect 10229 9469 10241 9472
rect 10275 9500 10287 9503
rect 11606 9500 11612 9512
rect 10275 9472 11612 9500
rect 10275 9469 10287 9472
rect 10229 9463 10287 9469
rect 11606 9460 11612 9472
rect 11664 9460 11670 9512
rect 12529 9503 12587 9509
rect 12529 9500 12541 9503
rect 12406 9472 12541 9500
rect 9324 9432 9352 9460
rect 12066 9432 12072 9444
rect 5960 9404 8892 9432
rect 9232 9404 9352 9432
rect 9692 9404 12072 9432
rect 5960 9392 5966 9404
rect 6362 9364 6368 9376
rect 4908 9336 6368 9364
rect 6362 9324 6368 9336
rect 6420 9324 6426 9376
rect 6641 9367 6699 9373
rect 6641 9333 6653 9367
rect 6687 9364 6699 9367
rect 7190 9364 7196 9376
rect 6687 9336 7196 9364
rect 6687 9333 6699 9336
rect 6641 9327 6699 9333
rect 7190 9324 7196 9336
rect 7248 9324 7254 9376
rect 7466 9324 7472 9376
rect 7524 9364 7530 9376
rect 9232 9364 9260 9404
rect 7524 9336 9260 9364
rect 7524 9324 7530 9336
rect 9306 9324 9312 9376
rect 9364 9364 9370 9376
rect 9692 9364 9720 9404
rect 12066 9392 12072 9404
rect 12124 9432 12130 9444
rect 12406 9432 12434 9472
rect 12529 9469 12541 9472
rect 12575 9469 12587 9503
rect 13464 9500 13492 9540
rect 13630 9528 13636 9540
rect 13688 9528 13694 9580
rect 13909 9571 13967 9577
rect 13909 9537 13921 9571
rect 13955 9568 13967 9571
rect 14366 9568 14372 9580
rect 13955 9540 14372 9568
rect 13955 9537 13967 9540
rect 13909 9531 13967 9537
rect 14366 9528 14372 9540
rect 14424 9568 14430 9580
rect 14642 9568 14648 9580
rect 14424 9540 14648 9568
rect 14424 9528 14430 9540
rect 14642 9528 14648 9540
rect 14700 9528 14706 9580
rect 15565 9571 15623 9577
rect 15565 9537 15577 9571
rect 15611 9568 15623 9571
rect 16666 9568 16672 9580
rect 15611 9540 16672 9568
rect 15611 9537 15623 9540
rect 15565 9531 15623 9537
rect 16666 9528 16672 9540
rect 16724 9528 16730 9580
rect 16758 9528 16764 9580
rect 16816 9568 16822 9580
rect 16853 9571 16911 9577
rect 16853 9568 16865 9571
rect 16816 9540 16865 9568
rect 16816 9528 16822 9540
rect 16853 9537 16865 9540
rect 16899 9537 16911 9571
rect 17016 9568 17044 9608
rect 17126 9596 17132 9648
rect 17184 9636 17190 9648
rect 18509 9639 18567 9645
rect 18509 9636 18521 9639
rect 17184 9608 18521 9636
rect 17184 9596 17190 9608
rect 18509 9605 18521 9608
rect 18555 9605 18567 9639
rect 18509 9599 18567 9605
rect 18693 9639 18751 9645
rect 18693 9605 18705 9639
rect 18739 9636 18751 9639
rect 19794 9636 19800 9648
rect 18739 9608 19800 9636
rect 18739 9605 18751 9608
rect 18693 9599 18751 9605
rect 19794 9596 19800 9608
rect 19852 9596 19858 9648
rect 20364 9608 21312 9636
rect 17586 9568 17592 9580
rect 17016 9540 17356 9568
rect 17547 9540 17592 9568
rect 16853 9531 16911 9537
rect 15838 9500 15844 9512
rect 13464 9472 15844 9500
rect 12529 9463 12587 9469
rect 15838 9460 15844 9472
rect 15896 9460 15902 9512
rect 17221 9503 17279 9509
rect 17221 9500 17233 9503
rect 16500 9472 17233 9500
rect 12802 9432 12808 9444
rect 12124 9404 12434 9432
rect 12636 9404 12808 9432
rect 12124 9392 12130 9404
rect 12636 9376 12664 9404
rect 12802 9392 12808 9404
rect 12860 9392 12866 9444
rect 13081 9435 13139 9441
rect 13081 9401 13093 9435
rect 13127 9432 13139 9435
rect 13633 9435 13691 9441
rect 13633 9432 13645 9435
rect 13127 9404 13645 9432
rect 13127 9401 13139 9404
rect 13081 9395 13139 9401
rect 13633 9401 13645 9404
rect 13679 9432 13691 9435
rect 15746 9432 15752 9444
rect 13679 9404 15752 9432
rect 13679 9401 13691 9404
rect 13633 9395 13691 9401
rect 15746 9392 15752 9404
rect 15804 9392 15810 9444
rect 9858 9364 9864 9376
rect 9364 9336 9720 9364
rect 9819 9336 9864 9364
rect 9364 9324 9370 9336
rect 9858 9324 9864 9336
rect 9916 9324 9922 9376
rect 11054 9364 11060 9376
rect 11015 9336 11060 9364
rect 11054 9324 11060 9336
rect 11112 9324 11118 9376
rect 12618 9364 12624 9376
rect 12579 9336 12624 9364
rect 12618 9324 12624 9336
rect 12676 9324 12682 9376
rect 12713 9367 12771 9373
rect 12713 9333 12725 9367
rect 12759 9364 12771 9367
rect 12894 9364 12900 9376
rect 12759 9336 12900 9364
rect 12759 9333 12771 9336
rect 12713 9327 12771 9333
rect 12894 9324 12900 9336
rect 12952 9364 12958 9376
rect 14090 9364 14096 9376
rect 12952 9336 14096 9364
rect 12952 9324 12958 9336
rect 14090 9324 14096 9336
rect 14148 9324 14154 9376
rect 14642 9324 14648 9376
rect 14700 9364 14706 9376
rect 14921 9367 14979 9373
rect 14921 9364 14933 9367
rect 14700 9336 14933 9364
rect 14700 9324 14706 9336
rect 14921 9333 14933 9336
rect 14967 9333 14979 9367
rect 14921 9327 14979 9333
rect 15654 9324 15660 9376
rect 15712 9364 15718 9376
rect 16114 9364 16120 9376
rect 15712 9336 16120 9364
rect 15712 9324 15718 9336
rect 16114 9324 16120 9336
rect 16172 9364 16178 9376
rect 16500 9364 16528 9472
rect 17221 9469 17233 9472
rect 17267 9469 17279 9503
rect 17328 9500 17356 9540
rect 17586 9528 17592 9540
rect 17644 9528 17650 9580
rect 18233 9571 18291 9577
rect 18233 9537 18245 9571
rect 18279 9568 18291 9571
rect 18322 9568 18328 9580
rect 18279 9540 18328 9568
rect 18279 9537 18291 9540
rect 18233 9531 18291 9537
rect 18322 9528 18328 9540
rect 18380 9528 18386 9580
rect 18414 9528 18420 9580
rect 18472 9568 18478 9580
rect 19245 9571 19303 9577
rect 19245 9568 19257 9571
rect 18472 9540 19257 9568
rect 18472 9528 18478 9540
rect 19245 9537 19257 9540
rect 19291 9537 19303 9571
rect 19518 9568 19524 9580
rect 19479 9540 19524 9568
rect 19245 9531 19303 9537
rect 19518 9528 19524 9540
rect 19576 9568 19582 9580
rect 20254 9568 20260 9580
rect 19576 9540 20260 9568
rect 19576 9528 19582 9540
rect 20254 9528 20260 9540
rect 20312 9528 20318 9580
rect 20364 9577 20392 9608
rect 20349 9571 20407 9577
rect 20349 9537 20361 9571
rect 20395 9537 20407 9571
rect 20349 9531 20407 9537
rect 20441 9571 20499 9577
rect 20441 9537 20453 9571
rect 20487 9537 20499 9571
rect 20622 9568 20628 9580
rect 20583 9540 20628 9568
rect 20441 9531 20499 9537
rect 20165 9503 20223 9509
rect 20165 9500 20177 9503
rect 17328 9472 20177 9500
rect 17221 9463 17279 9469
rect 20165 9469 20177 9472
rect 20211 9469 20223 9503
rect 20165 9463 20223 9469
rect 16850 9392 16856 9444
rect 16908 9432 16914 9444
rect 17129 9435 17187 9441
rect 17129 9432 17141 9435
rect 16908 9404 17141 9432
rect 16908 9392 16914 9404
rect 17129 9401 17141 9404
rect 17175 9401 17187 9435
rect 17129 9395 17187 9401
rect 19337 9435 19395 9441
rect 19337 9401 19349 9435
rect 19383 9432 19395 9435
rect 19610 9432 19616 9444
rect 19383 9404 19616 9432
rect 19383 9401 19395 9404
rect 19337 9395 19395 9401
rect 19610 9392 19616 9404
rect 19668 9392 19674 9444
rect 20456 9432 20484 9531
rect 20622 9528 20628 9540
rect 20680 9528 20686 9580
rect 20714 9528 20720 9580
rect 20772 9568 20778 9580
rect 21174 9568 21180 9580
rect 20772 9540 21180 9568
rect 20772 9528 20778 9540
rect 21174 9528 21180 9540
rect 21232 9528 21238 9580
rect 21284 9500 21312 9608
rect 21542 9596 21548 9648
rect 21600 9636 21606 9648
rect 21910 9636 21916 9648
rect 21600 9608 21916 9636
rect 21600 9596 21606 9608
rect 21910 9596 21916 9608
rect 21968 9636 21974 9648
rect 22189 9639 22247 9645
rect 22189 9636 22201 9639
rect 21968 9608 22201 9636
rect 21968 9596 21974 9608
rect 22189 9605 22201 9608
rect 22235 9605 22247 9639
rect 23106 9636 23112 9648
rect 23067 9608 23112 9636
rect 22189 9599 22247 9605
rect 23106 9596 23112 9608
rect 23164 9596 23170 9648
rect 21634 9528 21640 9580
rect 21692 9568 21698 9580
rect 22097 9571 22155 9577
rect 22097 9568 22109 9571
rect 21692 9540 22109 9568
rect 21692 9528 21698 9540
rect 22097 9537 22109 9540
rect 22143 9537 22155 9571
rect 22097 9531 22155 9537
rect 22278 9528 22284 9580
rect 22336 9568 22342 9580
rect 22373 9571 22431 9577
rect 22373 9568 22385 9571
rect 22336 9540 22385 9568
rect 22336 9528 22342 9540
rect 22373 9537 22385 9540
rect 22419 9537 22431 9571
rect 22373 9531 22431 9537
rect 22922 9500 22928 9512
rect 21284 9472 22928 9500
rect 22922 9460 22928 9472
rect 22980 9460 22986 9512
rect 20714 9432 20720 9444
rect 20456 9404 20720 9432
rect 20714 9392 20720 9404
rect 20772 9432 20778 9444
rect 22370 9432 22376 9444
rect 20772 9404 22376 9432
rect 20772 9392 20778 9404
rect 22370 9392 22376 9404
rect 22428 9392 22434 9444
rect 22646 9432 22652 9444
rect 22480 9404 22652 9432
rect 16172 9336 16528 9364
rect 16172 9324 16178 9336
rect 16574 9324 16580 9376
rect 16632 9364 16638 9376
rect 16991 9367 17049 9373
rect 16991 9364 17003 9367
rect 16632 9336 17003 9364
rect 16632 9324 16638 9336
rect 16991 9333 17003 9336
rect 17037 9333 17049 9367
rect 16991 9327 17049 9333
rect 17586 9324 17592 9376
rect 17644 9364 17650 9376
rect 18509 9367 18567 9373
rect 18509 9364 18521 9367
rect 17644 9336 18521 9364
rect 17644 9324 17650 9336
rect 18509 9333 18521 9336
rect 18555 9333 18567 9367
rect 19702 9364 19708 9376
rect 19663 9336 19708 9364
rect 18509 9327 18567 9333
rect 19702 9324 19708 9336
rect 19760 9324 19766 9376
rect 21082 9324 21088 9376
rect 21140 9364 21146 9376
rect 21177 9367 21235 9373
rect 21177 9364 21189 9367
rect 21140 9336 21189 9364
rect 21140 9324 21146 9336
rect 21177 9333 21189 9336
rect 21223 9333 21235 9367
rect 21177 9327 21235 9333
rect 21358 9324 21364 9376
rect 21416 9364 21422 9376
rect 22186 9364 22192 9376
rect 21416 9336 22192 9364
rect 21416 9324 21422 9336
rect 22186 9324 22192 9336
rect 22244 9364 22250 9376
rect 22480 9364 22508 9404
rect 22646 9392 22652 9404
rect 22704 9392 22710 9444
rect 22244 9336 22508 9364
rect 22557 9367 22615 9373
rect 22244 9324 22250 9336
rect 22557 9333 22569 9367
rect 22603 9364 22615 9367
rect 22738 9364 22744 9376
rect 22603 9336 22744 9364
rect 22603 9333 22615 9336
rect 22557 9327 22615 9333
rect 22738 9324 22744 9336
rect 22796 9324 22802 9376
rect 1104 9274 23828 9296
rect 1104 9222 3790 9274
rect 3842 9222 3854 9274
rect 3906 9222 3918 9274
rect 3970 9222 3982 9274
rect 4034 9222 4046 9274
rect 4098 9222 9471 9274
rect 9523 9222 9535 9274
rect 9587 9222 9599 9274
rect 9651 9222 9663 9274
rect 9715 9222 9727 9274
rect 9779 9222 15152 9274
rect 15204 9222 15216 9274
rect 15268 9222 15280 9274
rect 15332 9222 15344 9274
rect 15396 9222 15408 9274
rect 15460 9222 20833 9274
rect 20885 9222 20897 9274
rect 20949 9222 20961 9274
rect 21013 9222 21025 9274
rect 21077 9222 21089 9274
rect 21141 9222 23828 9274
rect 1104 9200 23828 9222
rect 1670 9120 1676 9172
rect 1728 9160 1734 9172
rect 2133 9163 2191 9169
rect 2133 9160 2145 9163
rect 1728 9132 2145 9160
rect 1728 9120 1734 9132
rect 2133 9129 2145 9132
rect 2179 9160 2191 9163
rect 3418 9160 3424 9172
rect 2179 9132 3424 9160
rect 2179 9129 2191 9132
rect 2133 9123 2191 9129
rect 3418 9120 3424 9132
rect 3476 9160 3482 9172
rect 4154 9160 4160 9172
rect 3476 9132 4160 9160
rect 3476 9120 3482 9132
rect 4154 9120 4160 9132
rect 4212 9120 4218 9172
rect 6270 9120 6276 9172
rect 6328 9160 6334 9172
rect 6825 9163 6883 9169
rect 6825 9160 6837 9163
rect 6328 9132 6837 9160
rect 6328 9120 6334 9132
rect 6825 9129 6837 9132
rect 6871 9129 6883 9163
rect 6825 9123 6883 9129
rect 7098 9120 7104 9172
rect 7156 9160 7162 9172
rect 9306 9160 9312 9172
rect 7156 9132 9312 9160
rect 7156 9120 7162 9132
rect 9306 9120 9312 9132
rect 9364 9120 9370 9172
rect 9858 9160 9864 9172
rect 9819 9132 9864 9160
rect 9858 9120 9864 9132
rect 9916 9120 9922 9172
rect 13170 9160 13176 9172
rect 11348 9132 13176 9160
rect 2314 9052 2320 9104
rect 2372 9092 2378 9104
rect 2372 9064 4016 9092
rect 2372 9052 2378 9064
rect 2590 9024 2596 9036
rect 2551 8996 2596 9024
rect 2590 8984 2596 8996
rect 2648 8984 2654 9036
rect 2130 8916 2136 8968
rect 2188 8956 2194 8968
rect 2317 8959 2375 8965
rect 2317 8956 2329 8959
rect 2188 8928 2329 8956
rect 2188 8916 2194 8928
rect 2317 8925 2329 8928
rect 2363 8925 2375 8959
rect 3237 8959 3295 8965
rect 3237 8956 3249 8959
rect 2317 8919 2375 8925
rect 2424 8928 3249 8956
rect 2424 8897 2452 8928
rect 3237 8925 3249 8928
rect 3283 8925 3295 8959
rect 3237 8919 3295 8925
rect 3421 8959 3479 8965
rect 3421 8925 3433 8959
rect 3467 8956 3479 8959
rect 3878 8956 3884 8968
rect 3467 8928 3884 8956
rect 3467 8925 3479 8928
rect 3421 8919 3479 8925
rect 2409 8891 2467 8897
rect 2409 8857 2421 8891
rect 2455 8857 2467 8891
rect 3050 8888 3056 8900
rect 3011 8860 3056 8888
rect 2409 8851 2467 8857
rect 3050 8848 3056 8860
rect 3108 8848 3114 8900
rect 3252 8888 3280 8919
rect 3878 8916 3884 8928
rect 3936 8916 3942 8968
rect 3988 8965 4016 9064
rect 4890 9052 4896 9104
rect 4948 9092 4954 9104
rect 9677 9095 9735 9101
rect 9677 9092 9689 9095
rect 4948 9064 9689 9092
rect 4948 9052 4954 9064
rect 9677 9061 9689 9064
rect 9723 9061 9735 9095
rect 9677 9055 9735 9061
rect 6270 8984 6276 9036
rect 6328 9024 6334 9036
rect 6456 9027 6514 9033
rect 6456 9024 6468 9027
rect 6328 8996 6468 9024
rect 6328 8984 6334 8996
rect 6456 8993 6468 8996
rect 6502 8993 6514 9027
rect 6456 8987 6514 8993
rect 9217 9027 9275 9033
rect 9217 8993 9229 9027
rect 9263 9024 9275 9027
rect 9263 8996 11100 9024
rect 9263 8993 9275 8996
rect 9217 8987 9275 8993
rect 3973 8959 4031 8965
rect 3973 8925 3985 8959
rect 4019 8925 4031 8959
rect 3973 8919 4031 8925
rect 4614 8916 4620 8968
rect 4672 8956 4678 8968
rect 5353 8959 5411 8965
rect 5353 8956 5365 8959
rect 4672 8928 5365 8956
rect 4672 8916 4678 8928
rect 5353 8925 5365 8928
rect 5399 8925 5411 8959
rect 5353 8919 5411 8925
rect 4246 8888 4252 8900
rect 3252 8860 4252 8888
rect 4246 8848 4252 8860
rect 4304 8848 4310 8900
rect 4982 8848 4988 8900
rect 5040 8888 5046 8900
rect 5077 8891 5135 8897
rect 5077 8888 5089 8891
rect 5040 8860 5089 8888
rect 5040 8848 5046 8860
rect 5077 8857 5089 8860
rect 5123 8857 5135 8891
rect 5077 8851 5135 8857
rect 2590 8780 2596 8832
rect 2648 8820 2654 8832
rect 4890 8820 4896 8832
rect 2648 8792 4896 8820
rect 2648 8780 2654 8792
rect 4890 8780 4896 8792
rect 4948 8780 4954 8832
rect 5368 8820 5396 8919
rect 5994 8916 6000 8968
rect 6052 8956 6058 8968
rect 6371 8959 6429 8965
rect 6371 8956 6383 8959
rect 6052 8928 6383 8956
rect 6052 8916 6058 8928
rect 6371 8925 6383 8928
rect 6417 8925 6429 8959
rect 6371 8919 6429 8925
rect 6548 8959 6606 8965
rect 6548 8925 6560 8959
rect 6594 8925 6606 8959
rect 6548 8919 6606 8925
rect 6564 8888 6592 8919
rect 6638 8916 6644 8968
rect 6696 8956 6702 8968
rect 6696 8928 6741 8956
rect 6696 8916 6702 8928
rect 9766 8916 9772 8968
rect 9824 8956 9830 8968
rect 9861 8959 9919 8965
rect 9861 8956 9873 8959
rect 9824 8928 9873 8956
rect 9824 8916 9830 8928
rect 9861 8925 9873 8928
rect 9907 8925 9919 8959
rect 9861 8919 9919 8925
rect 10042 8916 10048 8968
rect 10100 8956 10106 8968
rect 11072 8965 11100 8996
rect 11057 8959 11115 8965
rect 10100 8928 10145 8956
rect 10100 8916 10106 8928
rect 11057 8925 11069 8959
rect 11103 8956 11115 8959
rect 11348 8956 11376 9132
rect 13170 9120 13176 9132
rect 13228 9120 13234 9172
rect 14090 9120 14096 9172
rect 14148 9160 14154 9172
rect 14277 9163 14335 9169
rect 14277 9160 14289 9163
rect 14148 9132 14289 9160
rect 14148 9120 14154 9132
rect 14277 9129 14289 9132
rect 14323 9129 14335 9163
rect 17034 9160 17040 9172
rect 14277 9123 14335 9129
rect 14568 9132 17040 9160
rect 11793 9095 11851 9101
rect 11793 9061 11805 9095
rect 11839 9092 11851 9095
rect 13078 9092 13084 9104
rect 11839 9064 13084 9092
rect 11839 9061 11851 9064
rect 11793 9055 11851 9061
rect 13078 9052 13084 9064
rect 13136 9052 13142 9104
rect 13265 9095 13323 9101
rect 13265 9061 13277 9095
rect 13311 9092 13323 9095
rect 14568 9092 14596 9132
rect 17034 9120 17040 9132
rect 17092 9120 17098 9172
rect 17221 9163 17279 9169
rect 17221 9129 17233 9163
rect 17267 9160 17279 9163
rect 21358 9160 21364 9172
rect 17267 9132 21364 9160
rect 17267 9129 17279 9132
rect 17221 9123 17279 9129
rect 21358 9120 21364 9132
rect 21416 9120 21422 9172
rect 22002 9120 22008 9172
rect 22060 9160 22066 9172
rect 22741 9163 22799 9169
rect 22741 9160 22753 9163
rect 22060 9132 22753 9160
rect 22060 9120 22066 9132
rect 22741 9129 22753 9132
rect 22787 9160 22799 9163
rect 22830 9160 22836 9172
rect 22787 9132 22836 9160
rect 22787 9129 22799 9132
rect 22741 9123 22799 9129
rect 22830 9120 22836 9132
rect 22888 9120 22894 9172
rect 13311 9064 14596 9092
rect 14645 9095 14703 9101
rect 13311 9061 13323 9064
rect 13265 9055 13323 9061
rect 14645 9061 14657 9095
rect 14691 9092 14703 9095
rect 16298 9092 16304 9104
rect 14691 9064 16304 9092
rect 14691 9061 14703 9064
rect 14645 9055 14703 9061
rect 16298 9052 16304 9064
rect 16356 9052 16362 9104
rect 16850 9052 16856 9104
rect 16908 9092 16914 9104
rect 16908 9064 16953 9092
rect 16908 9052 16914 9064
rect 19702 9052 19708 9104
rect 19760 9092 19766 9104
rect 21269 9095 21327 9101
rect 21269 9092 21281 9095
rect 19760 9064 21281 9092
rect 19760 9052 19766 9064
rect 21269 9061 21281 9064
rect 21315 9061 21327 9095
rect 21269 9055 21327 9061
rect 12618 8984 12624 9036
rect 12676 9024 12682 9036
rect 15838 9024 15844 9036
rect 12676 8996 14412 9024
rect 12676 8984 12682 8996
rect 11514 8956 11520 8968
rect 11103 8928 11376 8956
rect 11475 8928 11520 8956
rect 11103 8925 11115 8928
rect 11057 8919 11115 8925
rect 11514 8916 11520 8928
rect 11572 8916 11578 8968
rect 11606 8916 11612 8968
rect 11664 8956 11670 8968
rect 12820 8965 12848 8996
rect 14384 8968 14412 8996
rect 15488 8996 15844 9024
rect 12713 8959 12771 8965
rect 11664 8928 11709 8956
rect 11664 8916 11670 8928
rect 12713 8925 12725 8959
rect 12759 8925 12771 8959
rect 12713 8919 12771 8925
rect 12805 8959 12863 8965
rect 12805 8925 12817 8959
rect 12851 8925 12863 8959
rect 12805 8919 12863 8925
rect 12989 8959 13047 8965
rect 12989 8925 13001 8959
rect 13035 8925 13047 8959
rect 12989 8919 13047 8925
rect 7006 8888 7012 8900
rect 6564 8860 7012 8888
rect 7006 8848 7012 8860
rect 7064 8848 7070 8900
rect 11698 8848 11704 8900
rect 11756 8888 11762 8900
rect 11793 8891 11851 8897
rect 11793 8888 11805 8891
rect 11756 8860 11805 8888
rect 11756 8848 11762 8860
rect 11793 8857 11805 8860
rect 11839 8857 11851 8891
rect 12728 8888 12756 8919
rect 12894 8888 12900 8900
rect 12728 8860 12900 8888
rect 11793 8851 11851 8857
rect 8662 8820 8668 8832
rect 5368 8792 8668 8820
rect 8662 8780 8668 8792
rect 8720 8780 8726 8832
rect 10962 8820 10968 8832
rect 10923 8792 10968 8820
rect 10962 8780 10968 8792
rect 11020 8780 11026 8832
rect 11808 8820 11836 8851
rect 12894 8848 12900 8860
rect 12952 8848 12958 8900
rect 13004 8888 13032 8919
rect 13078 8916 13084 8968
rect 13136 8956 13142 8968
rect 13136 8928 13181 8956
rect 13136 8916 13142 8928
rect 13630 8916 13636 8968
rect 13688 8956 13694 8968
rect 14277 8959 14335 8965
rect 14277 8956 14289 8959
rect 13688 8928 14289 8956
rect 13688 8916 13694 8928
rect 14277 8925 14289 8928
rect 14323 8925 14335 8959
rect 14277 8919 14335 8925
rect 14366 8916 14372 8968
rect 14424 8956 14430 8968
rect 15488 8965 15516 8996
rect 15838 8984 15844 8996
rect 15896 8984 15902 9036
rect 16574 8984 16580 9036
rect 16632 9024 16638 9036
rect 16724 9027 16782 9033
rect 16724 9024 16736 9027
rect 16632 8996 16736 9024
rect 16632 8984 16638 8996
rect 16724 8993 16736 8996
rect 16770 8993 16782 9027
rect 16942 9024 16948 9036
rect 16903 8996 16948 9024
rect 16724 8987 16782 8993
rect 16942 8984 16948 8996
rect 17000 8984 17006 9036
rect 18877 9027 18935 9033
rect 18877 8993 18889 9027
rect 18923 9024 18935 9027
rect 22370 9024 22376 9036
rect 18923 8996 22376 9024
rect 18923 8993 18935 8996
rect 18877 8987 18935 8993
rect 22370 8984 22376 8996
rect 22428 9024 22434 9036
rect 23106 9024 23112 9036
rect 22428 8996 23112 9024
rect 22428 8984 22434 8996
rect 23106 8984 23112 8996
rect 23164 8984 23170 9036
rect 15488 8959 15571 8965
rect 14424 8928 14469 8956
rect 15488 8928 15525 8959
rect 14424 8916 14430 8928
rect 15513 8925 15525 8928
rect 15559 8925 15571 8959
rect 15513 8919 15571 8925
rect 18233 8959 18291 8965
rect 18233 8925 18245 8959
rect 18279 8956 18291 8959
rect 18322 8956 18328 8968
rect 18279 8928 18328 8956
rect 18279 8925 18291 8928
rect 18233 8919 18291 8925
rect 18322 8916 18328 8928
rect 18380 8916 18386 8968
rect 19886 8956 19892 8968
rect 19847 8928 19892 8956
rect 19886 8916 19892 8928
rect 19944 8916 19950 8968
rect 21174 8956 21180 8968
rect 21135 8928 21180 8956
rect 21174 8916 21180 8928
rect 21232 8916 21238 8968
rect 21358 8956 21364 8968
rect 21319 8928 21364 8956
rect 21358 8916 21364 8928
rect 21416 8916 21422 8968
rect 21450 8916 21456 8968
rect 21508 8956 21514 8968
rect 21637 8959 21695 8965
rect 21508 8928 21553 8956
rect 21508 8916 21514 8928
rect 21637 8925 21649 8959
rect 21683 8956 21695 8959
rect 21910 8956 21916 8968
rect 21683 8928 21916 8956
rect 21683 8925 21695 8928
rect 21637 8919 21695 8925
rect 21910 8916 21916 8928
rect 21968 8916 21974 8968
rect 13648 8888 13676 8916
rect 13004 8860 13676 8888
rect 13722 8848 13728 8900
rect 13780 8888 13786 8900
rect 15105 8891 15163 8897
rect 15105 8888 15117 8891
rect 13780 8860 15117 8888
rect 13780 8848 13786 8860
rect 15105 8857 15117 8860
rect 15151 8857 15163 8891
rect 15105 8851 15163 8857
rect 15289 8891 15347 8897
rect 15289 8857 15301 8891
rect 15335 8888 15347 8891
rect 15335 8860 15608 8888
rect 15335 8857 15347 8860
rect 15289 8851 15347 8857
rect 14550 8820 14556 8832
rect 11808 8792 14556 8820
rect 14550 8780 14556 8792
rect 14608 8780 14614 8832
rect 15378 8820 15384 8832
rect 15339 8792 15384 8820
rect 15378 8780 15384 8792
rect 15436 8780 15442 8832
rect 15580 8820 15608 8860
rect 15654 8848 15660 8900
rect 15712 8888 15718 8900
rect 16577 8891 16635 8897
rect 15712 8860 15757 8888
rect 15712 8848 15718 8860
rect 16577 8857 16589 8891
rect 16623 8888 16635 8891
rect 16758 8888 16764 8900
rect 16623 8860 16764 8888
rect 16623 8857 16635 8860
rect 16577 8851 16635 8857
rect 16758 8848 16764 8860
rect 16816 8848 16822 8900
rect 19610 8848 19616 8900
rect 19668 8888 19674 8900
rect 20254 8888 20260 8900
rect 19668 8860 20260 8888
rect 19668 8848 19674 8860
rect 20254 8848 20260 8860
rect 20312 8848 20318 8900
rect 15746 8820 15752 8832
rect 15580 8792 15752 8820
rect 15746 8780 15752 8792
rect 15804 8820 15810 8832
rect 17494 8820 17500 8832
rect 15804 8792 17500 8820
rect 15804 8780 15810 8792
rect 17494 8780 17500 8792
rect 17552 8780 17558 8832
rect 17957 8823 18015 8829
rect 17957 8789 17969 8823
rect 18003 8820 18015 8823
rect 18874 8820 18880 8832
rect 18003 8792 18880 8820
rect 18003 8789 18015 8792
rect 17957 8783 18015 8789
rect 18874 8780 18880 8792
rect 18932 8780 18938 8832
rect 19426 8780 19432 8832
rect 19484 8820 19490 8832
rect 20993 8823 21051 8829
rect 20993 8820 21005 8823
rect 19484 8792 21005 8820
rect 19484 8780 19490 8792
rect 20993 8789 21005 8792
rect 21039 8789 21051 8823
rect 22186 8820 22192 8832
rect 22147 8792 22192 8820
rect 20993 8783 21051 8789
rect 22186 8780 22192 8792
rect 22244 8780 22250 8832
rect 23198 8820 23204 8832
rect 23159 8792 23204 8820
rect 23198 8780 23204 8792
rect 23256 8780 23262 8832
rect 1104 8730 23987 8752
rect 1104 8678 6630 8730
rect 6682 8678 6694 8730
rect 6746 8678 6758 8730
rect 6810 8678 6822 8730
rect 6874 8678 6886 8730
rect 6938 8678 12311 8730
rect 12363 8678 12375 8730
rect 12427 8678 12439 8730
rect 12491 8678 12503 8730
rect 12555 8678 12567 8730
rect 12619 8678 17992 8730
rect 18044 8678 18056 8730
rect 18108 8678 18120 8730
rect 18172 8678 18184 8730
rect 18236 8678 18248 8730
rect 18300 8678 23673 8730
rect 23725 8678 23737 8730
rect 23789 8678 23801 8730
rect 23853 8678 23865 8730
rect 23917 8678 23929 8730
rect 23981 8678 23987 8730
rect 1104 8656 23987 8678
rect 3789 8619 3847 8625
rect 3789 8585 3801 8619
rect 3835 8616 3847 8619
rect 7650 8616 7656 8628
rect 3835 8588 7656 8616
rect 3835 8585 3847 8588
rect 3789 8579 3847 8585
rect 7650 8576 7656 8588
rect 7708 8576 7714 8628
rect 9122 8616 9128 8628
rect 9083 8588 9128 8616
rect 9122 8576 9128 8588
rect 9180 8616 9186 8628
rect 9585 8619 9643 8625
rect 9585 8616 9597 8619
rect 9180 8588 9597 8616
rect 9180 8576 9186 8588
rect 9585 8585 9597 8588
rect 9631 8585 9643 8619
rect 9585 8579 9643 8585
rect 10870 8576 10876 8628
rect 10928 8616 10934 8628
rect 11701 8619 11759 8625
rect 11701 8616 11713 8619
rect 10928 8588 11713 8616
rect 10928 8576 10934 8588
rect 11701 8585 11713 8588
rect 11747 8585 11759 8619
rect 11701 8579 11759 8585
rect 12066 8576 12072 8628
rect 12124 8616 12130 8628
rect 12802 8616 12808 8628
rect 12124 8588 12808 8616
rect 12124 8576 12130 8588
rect 12802 8576 12808 8588
rect 12860 8576 12866 8628
rect 16301 8619 16359 8625
rect 16301 8585 16313 8619
rect 16347 8616 16359 8619
rect 16850 8616 16856 8628
rect 16347 8588 16856 8616
rect 16347 8585 16359 8588
rect 16301 8579 16359 8585
rect 16850 8576 16856 8588
rect 16908 8576 16914 8628
rect 17310 8576 17316 8628
rect 17368 8616 17374 8628
rect 17368 8588 19656 8616
rect 17368 8576 17374 8588
rect 19628 8560 19656 8588
rect 19886 8576 19892 8628
rect 19944 8616 19950 8628
rect 23198 8616 23204 8628
rect 19944 8588 23204 8616
rect 19944 8576 19950 8588
rect 23198 8576 23204 8588
rect 23256 8576 23262 8628
rect 1946 8548 1952 8560
rect 1859 8520 1952 8548
rect 1872 8489 1900 8520
rect 1946 8508 1952 8520
rect 2004 8548 2010 8560
rect 3234 8548 3240 8560
rect 2004 8520 3240 8548
rect 2004 8508 2010 8520
rect 3234 8508 3240 8520
rect 3292 8508 3298 8560
rect 7006 8548 7012 8560
rect 6967 8520 7012 8548
rect 7006 8508 7012 8520
rect 7064 8548 7070 8560
rect 8294 8548 8300 8560
rect 7064 8520 8300 8548
rect 7064 8508 7070 8520
rect 8294 8508 8300 8520
rect 8352 8508 8358 8560
rect 9030 8548 9036 8560
rect 8680 8520 9036 8548
rect 8680 8492 8708 8520
rect 9030 8508 9036 8520
rect 9088 8508 9094 8560
rect 10226 8508 10232 8560
rect 10284 8548 10290 8560
rect 13081 8551 13139 8557
rect 10284 8520 12388 8548
rect 10284 8508 10290 8520
rect 1673 8483 1731 8489
rect 1673 8449 1685 8483
rect 1719 8449 1731 8483
rect 1673 8443 1731 8449
rect 1857 8483 1915 8489
rect 1857 8449 1869 8483
rect 1903 8449 1915 8483
rect 2774 8480 2780 8492
rect 2735 8452 2780 8480
rect 1857 8443 1915 8449
rect 1688 8412 1716 8443
rect 2774 8440 2780 8452
rect 2832 8440 2838 8492
rect 3326 8480 3332 8492
rect 3287 8452 3332 8480
rect 3326 8440 3332 8452
rect 3384 8440 3390 8492
rect 3605 8483 3663 8489
rect 3605 8449 3617 8483
rect 3651 8480 3663 8483
rect 4246 8480 4252 8492
rect 3651 8452 4252 8480
rect 3651 8449 3663 8452
rect 3605 8443 3663 8449
rect 4246 8440 4252 8452
rect 4304 8440 4310 8492
rect 4890 8480 4896 8492
rect 4851 8452 4896 8480
rect 4890 8440 4896 8452
rect 4948 8440 4954 8492
rect 5902 8440 5908 8492
rect 5960 8480 5966 8492
rect 6549 8483 6607 8489
rect 6549 8480 6561 8483
rect 5960 8452 6561 8480
rect 5960 8440 5966 8452
rect 6549 8449 6561 8452
rect 6595 8449 6607 8483
rect 7466 8480 7472 8492
rect 7427 8452 7472 8480
rect 6549 8443 6607 8449
rect 7466 8440 7472 8452
rect 7524 8440 7530 8492
rect 7834 8440 7840 8492
rect 7892 8480 7898 8492
rect 8113 8483 8171 8489
rect 8113 8480 8125 8483
rect 7892 8452 8125 8480
rect 7892 8440 7898 8452
rect 8113 8449 8125 8452
rect 8159 8449 8171 8483
rect 8113 8443 8171 8449
rect 8573 8483 8631 8489
rect 8573 8449 8585 8483
rect 8619 8480 8631 8483
rect 8662 8480 8668 8492
rect 8619 8452 8668 8480
rect 8619 8449 8631 8452
rect 8573 8443 8631 8449
rect 8662 8440 8668 8452
rect 8720 8440 8726 8492
rect 8938 8440 8944 8492
rect 8996 8480 9002 8492
rect 10137 8483 10195 8489
rect 10137 8480 10149 8483
rect 8996 8452 10149 8480
rect 8996 8440 9002 8452
rect 10137 8449 10149 8452
rect 10183 8449 10195 8483
rect 10137 8443 10195 8449
rect 10321 8483 10379 8489
rect 10321 8449 10333 8483
rect 10367 8449 10379 8483
rect 10321 8443 10379 8449
rect 2130 8412 2136 8424
rect 1688 8384 2136 8412
rect 2130 8372 2136 8384
rect 2188 8372 2194 8424
rect 2317 8415 2375 8421
rect 2317 8381 2329 8415
rect 2363 8412 2375 8415
rect 2406 8412 2412 8424
rect 2363 8384 2412 8412
rect 2363 8381 2375 8384
rect 2317 8375 2375 8381
rect 2406 8372 2412 8384
rect 2464 8412 2470 8424
rect 2682 8412 2688 8424
rect 2464 8384 2688 8412
rect 2464 8372 2470 8384
rect 2682 8372 2688 8384
rect 2740 8372 2746 8424
rect 2869 8415 2927 8421
rect 2869 8381 2881 8415
rect 2915 8412 2927 8415
rect 2958 8412 2964 8424
rect 2915 8384 2964 8412
rect 2915 8381 2927 8384
rect 2869 8375 2927 8381
rect 2958 8372 2964 8384
rect 3016 8372 3022 8424
rect 3510 8412 3516 8424
rect 3471 8384 3516 8412
rect 3510 8372 3516 8384
rect 3568 8372 3574 8424
rect 4430 8372 4436 8424
rect 4488 8412 4494 8424
rect 5169 8415 5227 8421
rect 5169 8412 5181 8415
rect 4488 8384 5181 8412
rect 4488 8372 4494 8384
rect 5169 8381 5181 8384
rect 5215 8381 5227 8415
rect 5169 8375 5227 8381
rect 6362 8372 6368 8424
rect 6420 8412 6426 8424
rect 8297 8415 8355 8421
rect 8297 8412 8309 8415
rect 6420 8384 8309 8412
rect 6420 8372 6426 8384
rect 8297 8381 8309 8384
rect 8343 8381 8355 8415
rect 8297 8375 8355 8381
rect 9306 8372 9312 8424
rect 9364 8412 9370 8424
rect 10336 8412 10364 8443
rect 10686 8440 10692 8492
rect 10744 8480 10750 8492
rect 11057 8483 11115 8489
rect 11057 8480 11069 8483
rect 10744 8452 11069 8480
rect 10744 8440 10750 8452
rect 11057 8449 11069 8452
rect 11103 8480 11115 8483
rect 11698 8480 11704 8492
rect 11103 8452 11704 8480
rect 11103 8449 11115 8452
rect 11057 8443 11115 8449
rect 11698 8440 11704 8452
rect 11756 8440 11762 8492
rect 11882 8480 11888 8492
rect 11843 8452 11888 8480
rect 11882 8440 11888 8452
rect 11940 8440 11946 8492
rect 11977 8483 12035 8489
rect 11977 8449 11989 8483
rect 12023 8449 12035 8483
rect 12158 8480 12164 8492
rect 12119 8452 12164 8480
rect 11977 8443 12035 8449
rect 9364 8384 10364 8412
rect 9364 8372 9370 8384
rect 11606 8372 11612 8424
rect 11664 8412 11670 8424
rect 11992 8412 12020 8443
rect 12158 8440 12164 8452
rect 12216 8440 12222 8492
rect 12253 8483 12311 8489
rect 12253 8449 12265 8483
rect 12299 8449 12311 8483
rect 12360 8480 12388 8520
rect 13081 8517 13093 8551
rect 13127 8548 13139 8551
rect 13262 8548 13268 8560
rect 13127 8520 13268 8548
rect 13127 8517 13139 8520
rect 13081 8511 13139 8517
rect 13262 8508 13268 8520
rect 13320 8548 13326 8560
rect 13320 8520 15608 8548
rect 13320 8508 13326 8520
rect 14185 8483 14243 8489
rect 14185 8480 14197 8483
rect 12360 8452 14197 8480
rect 12253 8443 12311 8449
rect 14185 8449 14197 8452
rect 14231 8449 14243 8483
rect 14185 8443 14243 8449
rect 14461 8483 14519 8489
rect 14461 8449 14473 8483
rect 14507 8449 14519 8483
rect 14461 8443 14519 8449
rect 11664 8384 12020 8412
rect 11664 8372 11670 8384
rect 1857 8347 1915 8353
rect 1857 8313 1869 8347
rect 1903 8344 1915 8347
rect 1903 8316 2774 8344
rect 1903 8313 1915 8316
rect 1857 8307 1915 8313
rect 2746 8276 2774 8316
rect 3234 8304 3240 8356
rect 3292 8344 3298 8356
rect 4338 8344 4344 8356
rect 3292 8316 4344 8344
rect 3292 8304 3298 8316
rect 4338 8304 4344 8316
rect 4396 8344 4402 8356
rect 6270 8344 6276 8356
rect 4396 8316 6276 8344
rect 4396 8304 4402 8316
rect 6270 8304 6276 8316
rect 6328 8344 6334 8356
rect 6328 8316 8156 8344
rect 6328 8304 6334 8316
rect 8128 8288 8156 8316
rect 9858 8304 9864 8356
rect 9916 8344 9922 8356
rect 10321 8347 10379 8353
rect 10321 8344 10333 8347
rect 9916 8316 10333 8344
rect 9916 8304 9922 8316
rect 10321 8313 10333 8316
rect 10367 8344 10379 8347
rect 10502 8344 10508 8356
rect 10367 8316 10508 8344
rect 10367 8313 10379 8316
rect 10321 8307 10379 8313
rect 10502 8304 10508 8316
rect 10560 8304 10566 8356
rect 3329 8279 3387 8285
rect 3329 8276 3341 8279
rect 2746 8248 3341 8276
rect 3329 8245 3341 8248
rect 3375 8245 3387 8279
rect 7926 8276 7932 8288
rect 7887 8248 7932 8276
rect 3329 8239 3387 8245
rect 7926 8236 7932 8248
rect 7984 8236 7990 8288
rect 8110 8276 8116 8288
rect 8071 8248 8116 8276
rect 8110 8236 8116 8248
rect 8168 8236 8174 8288
rect 9214 8236 9220 8288
rect 9272 8276 9278 8288
rect 9766 8276 9772 8288
rect 9272 8248 9772 8276
rect 9272 8236 9278 8248
rect 9766 8236 9772 8248
rect 9824 8276 9830 8288
rect 10778 8276 10784 8288
rect 9824 8248 10784 8276
rect 9824 8236 9830 8248
rect 10778 8236 10784 8248
rect 10836 8276 10842 8288
rect 12268 8276 12296 8443
rect 14090 8412 14096 8424
rect 14051 8384 14096 8412
rect 14090 8372 14096 8384
rect 14148 8372 14154 8424
rect 13630 8304 13636 8356
rect 13688 8344 13694 8356
rect 14476 8344 14504 8443
rect 14642 8412 14648 8424
rect 14603 8384 14648 8412
rect 14642 8372 14648 8384
rect 14700 8372 14706 8424
rect 15197 8415 15255 8421
rect 15197 8381 15209 8415
rect 15243 8381 15255 8415
rect 15580 8412 15608 8520
rect 15838 8508 15844 8560
rect 15896 8548 15902 8560
rect 15933 8551 15991 8557
rect 15933 8548 15945 8551
rect 15896 8520 15945 8548
rect 15896 8508 15902 8520
rect 15933 8517 15945 8520
rect 15979 8517 15991 8551
rect 15933 8511 15991 8517
rect 16022 8508 16028 8560
rect 16080 8548 16086 8560
rect 16133 8551 16191 8557
rect 16133 8548 16145 8551
rect 16080 8520 16145 8548
rect 16080 8508 16086 8520
rect 16133 8517 16145 8520
rect 16179 8517 16191 8551
rect 16133 8511 16191 8517
rect 16574 8508 16580 8560
rect 16632 8548 16638 8560
rect 19610 8548 19616 8560
rect 16632 8520 18828 8548
rect 19523 8520 19616 8548
rect 16632 8508 16638 8520
rect 17497 8483 17555 8489
rect 17497 8449 17509 8483
rect 17543 8449 17555 8483
rect 17497 8443 17555 8449
rect 17310 8412 17316 8424
rect 15580 8384 17316 8412
rect 15197 8375 15255 8381
rect 13688 8316 14504 8344
rect 15212 8344 15240 8375
rect 17310 8372 17316 8384
rect 17368 8372 17374 8424
rect 17512 8412 17540 8443
rect 18230 8440 18236 8492
rect 18288 8480 18294 8492
rect 18800 8489 18828 8520
rect 19610 8508 19616 8520
rect 19668 8548 19674 8560
rect 20346 8548 20352 8560
rect 19668 8520 20352 8548
rect 19668 8508 19674 8520
rect 20346 8508 20352 8520
rect 20404 8508 20410 8560
rect 20714 8508 20720 8560
rect 20772 8548 20778 8560
rect 21085 8551 21143 8557
rect 21085 8548 21097 8551
rect 20772 8520 21097 8548
rect 20772 8508 20778 8520
rect 21085 8517 21097 8520
rect 21131 8517 21143 8551
rect 21085 8511 21143 8517
rect 21269 8551 21327 8557
rect 21269 8517 21281 8551
rect 21315 8548 21327 8551
rect 21726 8548 21732 8560
rect 21315 8520 21732 8548
rect 21315 8517 21327 8520
rect 21269 8511 21327 8517
rect 21726 8508 21732 8520
rect 21784 8508 21790 8560
rect 18325 8483 18383 8489
rect 18325 8480 18337 8483
rect 18288 8452 18337 8480
rect 18288 8440 18294 8452
rect 18325 8449 18337 8452
rect 18371 8449 18383 8483
rect 18325 8443 18383 8449
rect 18785 8483 18843 8489
rect 18785 8449 18797 8483
rect 18831 8449 18843 8483
rect 18785 8443 18843 8449
rect 17678 8412 17684 8424
rect 17512 8384 17684 8412
rect 17678 8372 17684 8384
rect 17736 8372 17742 8424
rect 17773 8415 17831 8421
rect 17773 8381 17785 8415
rect 17819 8381 17831 8415
rect 18340 8412 18368 8443
rect 18874 8440 18880 8492
rect 18932 8480 18938 8492
rect 21361 8483 21419 8489
rect 18932 8452 20760 8480
rect 18932 8440 18938 8452
rect 20732 8424 20760 8452
rect 21361 8449 21373 8483
rect 21407 8480 21419 8483
rect 21542 8480 21548 8492
rect 21407 8452 21548 8480
rect 21407 8449 21419 8452
rect 21361 8443 21419 8449
rect 21542 8440 21548 8452
rect 21600 8440 21606 8492
rect 21634 8440 21640 8492
rect 21692 8480 21698 8492
rect 22465 8483 22523 8489
rect 22465 8480 22477 8483
rect 21692 8452 22477 8480
rect 21692 8440 21698 8452
rect 22465 8449 22477 8452
rect 22511 8449 22523 8483
rect 22465 8443 22523 8449
rect 22554 8440 22560 8492
rect 22612 8480 22618 8492
rect 22830 8480 22836 8492
rect 22612 8452 22657 8480
rect 22791 8452 22836 8480
rect 22612 8440 22618 8452
rect 22830 8440 22836 8452
rect 22888 8440 22894 8492
rect 19518 8412 19524 8424
rect 18340 8384 19524 8412
rect 17773 8375 17831 8381
rect 17126 8344 17132 8356
rect 15212 8316 17132 8344
rect 13688 8304 13694 8316
rect 17126 8304 17132 8316
rect 17184 8304 17190 8356
rect 17788 8344 17816 8375
rect 19518 8372 19524 8384
rect 19576 8372 19582 8424
rect 20714 8372 20720 8424
rect 20772 8372 20778 8424
rect 22738 8412 22744 8424
rect 22699 8384 22744 8412
rect 22738 8372 22744 8384
rect 22796 8372 22802 8424
rect 19334 8344 19340 8356
rect 17788 8316 19340 8344
rect 19334 8304 19340 8316
rect 19392 8304 19398 8356
rect 20622 8304 20628 8356
rect 20680 8344 20686 8356
rect 21085 8347 21143 8353
rect 21085 8344 21097 8347
rect 20680 8316 21097 8344
rect 20680 8304 20686 8316
rect 21085 8313 21097 8316
rect 21131 8313 21143 8347
rect 22278 8344 22284 8356
rect 22239 8316 22284 8344
rect 21085 8307 21143 8313
rect 22278 8304 22284 8316
rect 22336 8304 22342 8356
rect 12894 8276 12900 8288
rect 10836 8248 12900 8276
rect 10836 8236 10842 8248
rect 12894 8236 12900 8248
rect 12952 8236 12958 8288
rect 15010 8236 15016 8288
rect 15068 8276 15074 8288
rect 15378 8276 15384 8288
rect 15068 8248 15384 8276
rect 15068 8236 15074 8248
rect 15378 8236 15384 8248
rect 15436 8276 15442 8288
rect 16117 8279 16175 8285
rect 16117 8276 16129 8279
rect 15436 8248 16129 8276
rect 15436 8236 15442 8248
rect 16117 8245 16129 8248
rect 16163 8245 16175 8279
rect 16117 8239 16175 8245
rect 1104 8186 23828 8208
rect 1104 8134 3790 8186
rect 3842 8134 3854 8186
rect 3906 8134 3918 8186
rect 3970 8134 3982 8186
rect 4034 8134 4046 8186
rect 4098 8134 9471 8186
rect 9523 8134 9535 8186
rect 9587 8134 9599 8186
rect 9651 8134 9663 8186
rect 9715 8134 9727 8186
rect 9779 8134 15152 8186
rect 15204 8134 15216 8186
rect 15268 8134 15280 8186
rect 15332 8134 15344 8186
rect 15396 8134 15408 8186
rect 15460 8134 20833 8186
rect 20885 8134 20897 8186
rect 20949 8134 20961 8186
rect 21013 8134 21025 8186
rect 21077 8134 21089 8186
rect 21141 8134 23828 8186
rect 1104 8112 23828 8134
rect 2409 8075 2467 8081
rect 2409 8041 2421 8075
rect 2455 8072 2467 8075
rect 3326 8072 3332 8084
rect 2455 8044 3332 8072
rect 2455 8041 2467 8044
rect 2409 8035 2467 8041
rect 3326 8032 3332 8044
rect 3384 8032 3390 8084
rect 4154 8032 4160 8084
rect 4212 8072 4218 8084
rect 4525 8075 4583 8081
rect 4525 8072 4537 8075
rect 4212 8044 4537 8072
rect 4212 8032 4218 8044
rect 4525 8041 4537 8044
rect 4571 8072 4583 8075
rect 4982 8072 4988 8084
rect 4571 8044 4988 8072
rect 4571 8041 4583 8044
rect 4525 8035 4583 8041
rect 4982 8032 4988 8044
rect 5040 8032 5046 8084
rect 5721 8075 5779 8081
rect 5721 8041 5733 8075
rect 5767 8072 5779 8075
rect 6086 8072 6092 8084
rect 5767 8044 6092 8072
rect 5767 8041 5779 8044
rect 5721 8035 5779 8041
rect 6086 8032 6092 8044
rect 6144 8032 6150 8084
rect 7742 8072 7748 8084
rect 7703 8044 7748 8072
rect 7742 8032 7748 8044
rect 7800 8032 7806 8084
rect 8113 8075 8171 8081
rect 8113 8041 8125 8075
rect 8159 8072 8171 8075
rect 8938 8072 8944 8084
rect 8159 8044 8944 8072
rect 8159 8041 8171 8044
rect 8113 8035 8171 8041
rect 2774 7964 2780 8016
rect 2832 8004 2838 8016
rect 3234 8004 3240 8016
rect 2832 7976 3240 8004
rect 2832 7964 2838 7976
rect 3160 7945 3188 7976
rect 3234 7964 3240 7976
rect 3292 8004 3298 8016
rect 3292 7976 4660 8004
rect 3292 7964 3298 7976
rect 3145 7939 3203 7945
rect 3145 7905 3157 7939
rect 3191 7905 3203 7939
rect 4522 7936 4528 7948
rect 3145 7899 3203 7905
rect 3344 7908 4528 7936
rect 1946 7868 1952 7880
rect 1907 7840 1952 7868
rect 1946 7828 1952 7840
rect 2004 7828 2010 7880
rect 2222 7868 2228 7880
rect 2183 7840 2228 7868
rect 2222 7828 2228 7840
rect 2280 7828 2286 7880
rect 3344 7877 3372 7908
rect 4522 7896 4528 7908
rect 4580 7896 4586 7948
rect 4632 7936 4660 7976
rect 5810 7964 5816 8016
rect 5868 8004 5874 8016
rect 7374 8004 7380 8016
rect 5868 7976 7380 8004
rect 5868 7964 5874 7976
rect 7374 7964 7380 7976
rect 7432 8004 7438 8016
rect 8128 8004 8156 8035
rect 8938 8032 8944 8044
rect 8996 8032 9002 8084
rect 10505 8075 10563 8081
rect 10505 8041 10517 8075
rect 10551 8072 10563 8075
rect 11146 8072 11152 8084
rect 10551 8044 11152 8072
rect 10551 8041 10563 8044
rect 10505 8035 10563 8041
rect 11146 8032 11152 8044
rect 11204 8032 11210 8084
rect 13630 8072 13636 8084
rect 13591 8044 13636 8072
rect 13630 8032 13636 8044
rect 13688 8032 13694 8084
rect 17678 8032 17684 8084
rect 17736 8072 17742 8084
rect 18509 8075 18567 8081
rect 18509 8072 18521 8075
rect 17736 8044 18521 8072
rect 17736 8032 17742 8044
rect 18509 8041 18521 8044
rect 18555 8072 18567 8075
rect 19978 8072 19984 8084
rect 18555 8044 19984 8072
rect 18555 8041 18567 8044
rect 18509 8035 18567 8041
rect 11698 8004 11704 8016
rect 7432 7976 8156 8004
rect 9600 7976 11704 8004
rect 7432 7964 7438 7976
rect 4632 7908 6960 7936
rect 3329 7871 3387 7877
rect 3329 7837 3341 7871
rect 3375 7837 3387 7871
rect 4338 7868 4344 7880
rect 4299 7840 4344 7868
rect 3329 7831 3387 7837
rect 4338 7828 4344 7840
rect 4396 7828 4402 7880
rect 4430 7828 4436 7880
rect 4488 7868 4494 7880
rect 5537 7871 5595 7877
rect 5537 7868 5549 7871
rect 4488 7840 4533 7868
rect 4632 7840 5549 7868
rect 4488 7828 4494 7840
rect 4522 7760 4528 7812
rect 4580 7800 4586 7812
rect 4632 7800 4660 7840
rect 5537 7837 5549 7840
rect 5583 7837 5595 7871
rect 5537 7831 5595 7837
rect 5721 7871 5779 7877
rect 5721 7837 5733 7871
rect 5767 7868 5779 7871
rect 5810 7868 5816 7880
rect 5767 7840 5816 7868
rect 5767 7837 5779 7840
rect 5721 7831 5779 7837
rect 5810 7828 5816 7840
rect 5868 7828 5874 7880
rect 6546 7868 6552 7880
rect 6507 7840 6552 7868
rect 6546 7828 6552 7840
rect 6604 7828 6610 7880
rect 6825 7871 6883 7877
rect 6825 7868 6837 7871
rect 6656 7840 6837 7868
rect 5261 7803 5319 7809
rect 5261 7800 5273 7803
rect 4580 7772 4660 7800
rect 4724 7772 5273 7800
rect 4580 7760 4586 7772
rect 2041 7735 2099 7741
rect 2041 7701 2053 7735
rect 2087 7732 2099 7735
rect 2130 7732 2136 7744
rect 2087 7704 2136 7732
rect 2087 7701 2099 7704
rect 2041 7695 2099 7701
rect 2130 7692 2136 7704
rect 2188 7692 2194 7744
rect 4724 7741 4752 7772
rect 5261 7769 5273 7772
rect 5307 7800 5319 7803
rect 6454 7800 6460 7812
rect 5307 7772 6460 7800
rect 5307 7769 5319 7772
rect 5261 7763 5319 7769
rect 6454 7760 6460 7772
rect 6512 7800 6518 7812
rect 6656 7800 6684 7840
rect 6825 7837 6837 7840
rect 6871 7837 6883 7871
rect 6825 7831 6883 7837
rect 6512 7772 6684 7800
rect 6733 7803 6791 7809
rect 6512 7760 6518 7772
rect 6733 7769 6745 7803
rect 6779 7769 6791 7803
rect 6733 7763 6791 7769
rect 4709 7735 4767 7741
rect 4709 7701 4721 7735
rect 4755 7701 4767 7735
rect 4709 7695 4767 7701
rect 5810 7692 5816 7744
rect 5868 7732 5874 7744
rect 5905 7735 5963 7741
rect 5905 7732 5917 7735
rect 5868 7704 5917 7732
rect 5868 7692 5874 7704
rect 5905 7701 5917 7704
rect 5951 7701 5963 7735
rect 5905 7695 5963 7701
rect 6362 7692 6368 7744
rect 6420 7732 6426 7744
rect 6748 7732 6776 7763
rect 6420 7704 6776 7732
rect 6932 7732 6960 7908
rect 7926 7896 7932 7948
rect 7984 7936 7990 7948
rect 7984 7908 8156 7936
rect 7984 7896 7990 7908
rect 8018 7868 8024 7880
rect 7979 7840 8024 7868
rect 8018 7828 8024 7840
rect 8076 7828 8082 7880
rect 8128 7877 8156 7908
rect 9306 7896 9312 7948
rect 9364 7936 9370 7948
rect 9401 7939 9459 7945
rect 9401 7936 9413 7939
rect 9364 7908 9413 7936
rect 9364 7896 9370 7908
rect 9401 7905 9413 7908
rect 9447 7905 9459 7939
rect 9401 7899 9459 7905
rect 9600 7877 9628 7976
rect 11698 7964 11704 7976
rect 11756 7964 11762 8016
rect 14090 7964 14096 8016
rect 14148 8004 14154 8016
rect 19426 8004 19432 8016
rect 14148 7976 19432 8004
rect 14148 7964 14154 7976
rect 9674 7896 9680 7948
rect 9732 7936 9738 7948
rect 10413 7939 10471 7945
rect 9732 7908 10088 7936
rect 9732 7896 9738 7908
rect 8113 7871 8171 7877
rect 8113 7837 8125 7871
rect 8159 7837 8171 7871
rect 9585 7871 9643 7877
rect 9585 7868 9597 7871
rect 8113 7831 8171 7837
rect 8496 7840 9597 7868
rect 7282 7800 7288 7812
rect 7243 7772 7288 7800
rect 7282 7760 7288 7772
rect 7340 7760 7346 7812
rect 8496 7732 8524 7840
rect 9585 7837 9597 7840
rect 9631 7837 9643 7871
rect 9585 7831 9643 7837
rect 9953 7871 10011 7877
rect 9953 7837 9965 7871
rect 9999 7837 10011 7871
rect 9953 7831 10011 7837
rect 9030 7760 9036 7812
rect 9088 7800 9094 7812
rect 9968 7800 9996 7831
rect 9088 7772 9996 7800
rect 10060 7800 10088 7908
rect 10413 7905 10425 7939
rect 10459 7936 10471 7939
rect 11793 7939 11851 7945
rect 11793 7936 11805 7939
rect 10459 7908 11805 7936
rect 10459 7905 10471 7908
rect 10413 7899 10471 7905
rect 11793 7905 11805 7908
rect 11839 7905 11851 7939
rect 14366 7936 14372 7948
rect 14327 7908 14372 7936
rect 11793 7899 11851 7905
rect 14366 7896 14372 7908
rect 14424 7896 14430 7948
rect 10594 7828 10600 7880
rect 10652 7868 10658 7880
rect 10778 7868 10784 7880
rect 10652 7840 10784 7868
rect 10652 7828 10658 7840
rect 10778 7828 10784 7840
rect 10836 7868 10842 7880
rect 10873 7871 10931 7877
rect 10873 7868 10885 7871
rect 10836 7840 10885 7868
rect 10836 7828 10842 7840
rect 10873 7837 10885 7840
rect 10919 7837 10931 7871
rect 10873 7831 10931 7837
rect 11885 7871 11943 7877
rect 11885 7837 11897 7871
rect 11931 7868 11943 7871
rect 11974 7868 11980 7880
rect 11931 7840 11980 7868
rect 11931 7837 11943 7840
rect 11885 7831 11943 7837
rect 11974 7828 11980 7840
rect 12032 7828 12038 7880
rect 13170 7828 13176 7880
rect 13228 7868 13234 7880
rect 13538 7868 13544 7880
rect 13228 7840 13544 7868
rect 13228 7828 13234 7840
rect 13538 7828 13544 7840
rect 13596 7828 13602 7880
rect 13725 7871 13783 7877
rect 13725 7837 13737 7871
rect 13771 7837 13783 7871
rect 14458 7868 14464 7880
rect 14419 7840 14464 7868
rect 13725 7831 13783 7837
rect 10060 7772 10732 7800
rect 9088 7760 9094 7772
rect 9858 7732 9864 7744
rect 6932 7704 8524 7732
rect 9819 7704 9864 7732
rect 6420 7692 6426 7704
rect 9858 7692 9864 7704
rect 9916 7692 9922 7744
rect 10704 7741 10732 7772
rect 10962 7760 10968 7812
rect 11020 7800 11026 7812
rect 13740 7800 13768 7831
rect 14458 7828 14464 7840
rect 14516 7828 14522 7880
rect 14752 7877 14780 7976
rect 19426 7964 19432 7976
rect 19484 7964 19490 8016
rect 16298 7896 16304 7948
rect 16356 7936 16362 7948
rect 16356 7908 17356 7936
rect 16356 7896 16362 7908
rect 14737 7871 14795 7877
rect 14737 7837 14749 7871
rect 14783 7837 14795 7871
rect 14737 7831 14795 7837
rect 14826 7828 14832 7880
rect 14884 7868 14890 7880
rect 15933 7871 15991 7877
rect 15933 7868 15945 7871
rect 14884 7840 15945 7868
rect 14884 7828 14890 7840
rect 15933 7837 15945 7840
rect 15979 7837 15991 7871
rect 16574 7868 16580 7880
rect 16535 7840 16580 7868
rect 15933 7831 15991 7837
rect 16574 7828 16580 7840
rect 16632 7828 16638 7880
rect 16945 7871 17003 7877
rect 16945 7837 16957 7871
rect 16991 7837 17003 7871
rect 17126 7868 17132 7880
rect 17087 7840 17132 7868
rect 16945 7831 17003 7837
rect 15473 7803 15531 7809
rect 11020 7772 13676 7800
rect 13740 7772 14780 7800
rect 11020 7760 11026 7772
rect 10689 7735 10747 7741
rect 10689 7701 10701 7735
rect 10735 7701 10747 7735
rect 10689 7695 10747 7701
rect 10781 7735 10839 7741
rect 10781 7701 10793 7735
rect 10827 7732 10839 7735
rect 10870 7732 10876 7744
rect 10827 7704 10876 7732
rect 10827 7701 10839 7704
rect 10781 7695 10839 7701
rect 10870 7692 10876 7704
rect 10928 7692 10934 7744
rect 11146 7732 11152 7744
rect 11107 7704 11152 7732
rect 11146 7692 11152 7704
rect 11204 7692 11210 7744
rect 12437 7735 12495 7741
rect 12437 7701 12449 7735
rect 12483 7732 12495 7735
rect 12802 7732 12808 7744
rect 12483 7704 12808 7732
rect 12483 7701 12495 7704
rect 12437 7695 12495 7701
rect 12802 7692 12808 7704
rect 12860 7692 12866 7744
rect 13648 7732 13676 7772
rect 14752 7744 14780 7772
rect 15473 7769 15485 7803
rect 15519 7800 15531 7803
rect 16758 7800 16764 7812
rect 15519 7772 16764 7800
rect 15519 7769 15531 7772
rect 15473 7763 15531 7769
rect 16758 7760 16764 7772
rect 16816 7760 16822 7812
rect 16960 7800 16988 7831
rect 17126 7828 17132 7840
rect 17184 7828 17190 7880
rect 17328 7877 17356 7908
rect 17313 7871 17371 7877
rect 17313 7837 17325 7871
rect 17359 7837 17371 7871
rect 17586 7868 17592 7880
rect 17547 7840 17592 7868
rect 17313 7831 17371 7837
rect 17586 7828 17592 7840
rect 17644 7828 17650 7880
rect 18049 7871 18107 7877
rect 18049 7837 18061 7871
rect 18095 7868 18107 7871
rect 18598 7868 18604 7880
rect 18095 7840 18604 7868
rect 18095 7837 18107 7840
rect 18049 7831 18107 7837
rect 18598 7828 18604 7840
rect 18656 7828 18662 7880
rect 19429 7871 19487 7877
rect 19429 7837 19441 7871
rect 19475 7837 19487 7871
rect 19536 7868 19564 8044
rect 19978 8032 19984 8044
rect 20036 8032 20042 8084
rect 20993 8075 21051 8081
rect 20993 8041 21005 8075
rect 21039 8072 21051 8075
rect 21542 8072 21548 8084
rect 21039 8044 21548 8072
rect 21039 8041 21051 8044
rect 20993 8035 21051 8041
rect 21542 8032 21548 8044
rect 21600 8032 21606 8084
rect 21818 8032 21824 8084
rect 21876 8072 21882 8084
rect 22373 8075 22431 8081
rect 22373 8072 22385 8075
rect 21876 8044 22385 8072
rect 21876 8032 21882 8044
rect 22373 8041 22385 8044
rect 22419 8041 22431 8075
rect 22373 8035 22431 8041
rect 19613 8007 19671 8013
rect 19613 7973 19625 8007
rect 19659 8004 19671 8007
rect 21266 8004 21272 8016
rect 19659 7976 21272 8004
rect 19659 7973 19671 7976
rect 19613 7967 19671 7973
rect 21266 7964 21272 7976
rect 21324 7964 21330 8016
rect 22278 7964 22284 8016
rect 22336 8004 22342 8016
rect 22336 7976 22876 8004
rect 22336 7964 22342 7976
rect 20162 7896 20168 7948
rect 20220 7936 20226 7948
rect 22370 7936 22376 7948
rect 20220 7908 22376 7936
rect 20220 7896 20226 7908
rect 22370 7896 22376 7908
rect 22428 7936 22434 7948
rect 22428 7908 22784 7936
rect 22428 7896 22434 7908
rect 19613 7871 19671 7877
rect 19613 7868 19625 7871
rect 19536 7840 19625 7868
rect 19429 7831 19487 7837
rect 19613 7837 19625 7840
rect 19659 7837 19671 7871
rect 20533 7871 20591 7877
rect 20533 7868 20545 7871
rect 19613 7831 19671 7837
rect 19904 7840 20545 7868
rect 18414 7800 18420 7812
rect 16960 7772 18420 7800
rect 18414 7760 18420 7772
rect 18472 7760 18478 7812
rect 19444 7800 19472 7831
rect 19518 7800 19524 7812
rect 19444 7772 19524 7800
rect 19518 7760 19524 7772
rect 19576 7760 19582 7812
rect 14458 7732 14464 7744
rect 13648 7704 14464 7732
rect 14458 7692 14464 7704
rect 14516 7692 14522 7744
rect 14734 7692 14740 7744
rect 14792 7732 14798 7744
rect 16025 7735 16083 7741
rect 16025 7732 16037 7735
rect 14792 7704 16037 7732
rect 14792 7692 14798 7704
rect 16025 7701 16037 7704
rect 16071 7701 16083 7735
rect 16025 7695 16083 7701
rect 18690 7692 18696 7744
rect 18748 7732 18754 7744
rect 18966 7732 18972 7744
rect 18748 7704 18972 7732
rect 18748 7692 18754 7704
rect 18966 7692 18972 7704
rect 19024 7732 19030 7744
rect 19904 7732 19932 7840
rect 20533 7837 20545 7840
rect 20579 7837 20591 7871
rect 20533 7831 20591 7837
rect 20809 7871 20867 7877
rect 20809 7837 20821 7871
rect 20855 7868 20867 7871
rect 21450 7868 21456 7880
rect 20855 7840 21456 7868
rect 20855 7837 20867 7840
rect 20809 7831 20867 7837
rect 21450 7828 21456 7840
rect 21508 7868 21514 7880
rect 22002 7868 22008 7880
rect 21508 7840 22008 7868
rect 21508 7828 21514 7840
rect 22002 7828 22008 7840
rect 22060 7828 22066 7880
rect 22756 7877 22784 7908
rect 22848 7877 22876 7976
rect 22649 7871 22707 7877
rect 22649 7868 22661 7871
rect 22572 7840 22661 7868
rect 20070 7760 20076 7812
rect 20128 7800 20134 7812
rect 20622 7800 20628 7812
rect 20128 7772 20628 7800
rect 20128 7760 20134 7772
rect 20622 7760 20628 7772
rect 20680 7760 20686 7812
rect 22572 7800 22600 7840
rect 22649 7837 22661 7840
rect 22695 7837 22707 7871
rect 22649 7831 22707 7837
rect 22741 7871 22799 7877
rect 22741 7837 22753 7871
rect 22787 7837 22799 7871
rect 22741 7831 22799 7837
rect 22833 7871 22891 7877
rect 22833 7837 22845 7871
rect 22879 7837 22891 7871
rect 23014 7868 23020 7880
rect 22975 7840 23020 7868
rect 22833 7831 22891 7837
rect 23014 7828 23020 7840
rect 23072 7828 23078 7880
rect 22922 7800 22928 7812
rect 22572 7772 22928 7800
rect 22922 7760 22928 7772
rect 22980 7760 22986 7812
rect 19024 7704 19932 7732
rect 19024 7692 19030 7704
rect 19978 7692 19984 7744
rect 20036 7732 20042 7744
rect 21453 7735 21511 7741
rect 21453 7732 21465 7735
rect 20036 7704 21465 7732
rect 20036 7692 20042 7704
rect 21453 7701 21465 7704
rect 21499 7732 21511 7735
rect 22462 7732 22468 7744
rect 21499 7704 22468 7732
rect 21499 7701 21511 7704
rect 21453 7695 21511 7701
rect 22462 7692 22468 7704
rect 22520 7692 22526 7744
rect 1104 7642 23987 7664
rect 1104 7590 6630 7642
rect 6682 7590 6694 7642
rect 6746 7590 6758 7642
rect 6810 7590 6822 7642
rect 6874 7590 6886 7642
rect 6938 7590 12311 7642
rect 12363 7590 12375 7642
rect 12427 7590 12439 7642
rect 12491 7590 12503 7642
rect 12555 7590 12567 7642
rect 12619 7590 17992 7642
rect 18044 7590 18056 7642
rect 18108 7590 18120 7642
rect 18172 7590 18184 7642
rect 18236 7590 18248 7642
rect 18300 7590 23673 7642
rect 23725 7590 23737 7642
rect 23789 7590 23801 7642
rect 23853 7590 23865 7642
rect 23917 7590 23929 7642
rect 23981 7590 23987 7642
rect 1104 7568 23987 7590
rect 2866 7488 2872 7540
rect 2924 7528 2930 7540
rect 8570 7528 8576 7540
rect 2924 7500 4568 7528
rect 2924 7488 2930 7500
rect 4430 7460 4436 7472
rect 1780 7432 4436 7460
rect 1780 7404 1808 7432
rect 4430 7420 4436 7432
rect 4488 7420 4494 7472
rect 4540 7460 4568 7500
rect 4724 7500 8576 7528
rect 4724 7460 4752 7500
rect 8570 7488 8576 7500
rect 8628 7528 8634 7540
rect 9030 7528 9036 7540
rect 8628 7500 9036 7528
rect 8628 7488 8634 7500
rect 9030 7488 9036 7500
rect 9088 7488 9094 7540
rect 9953 7531 10011 7537
rect 9953 7528 9965 7531
rect 9140 7500 9965 7528
rect 4540 7432 4752 7460
rect 4798 7420 4804 7472
rect 4856 7460 4862 7472
rect 9140 7469 9168 7500
rect 9953 7497 9965 7500
rect 9999 7497 10011 7531
rect 11238 7528 11244 7540
rect 9953 7491 10011 7497
rect 10152 7500 11244 7528
rect 9125 7463 9183 7469
rect 4856 7432 8248 7460
rect 4856 7420 4862 7432
rect 8220 7404 8248 7432
rect 9125 7429 9137 7463
rect 9171 7429 9183 7463
rect 9125 7423 9183 7429
rect 9217 7463 9275 7469
rect 9217 7429 9229 7463
rect 9263 7460 9275 7463
rect 9766 7460 9772 7472
rect 9263 7432 9772 7460
rect 9263 7429 9275 7432
rect 9217 7423 9275 7429
rect 9766 7420 9772 7432
rect 9824 7420 9830 7472
rect 1762 7392 1768 7404
rect 1675 7364 1768 7392
rect 1762 7352 1768 7364
rect 1820 7352 1826 7404
rect 1946 7401 1952 7404
rect 1919 7395 1952 7401
rect 1919 7361 1931 7395
rect 2004 7392 2010 7404
rect 2314 7392 2320 7404
rect 2004 7364 2320 7392
rect 1919 7355 1952 7361
rect 1946 7352 1952 7355
rect 2004 7352 2010 7364
rect 2314 7352 2320 7364
rect 2372 7352 2378 7404
rect 2866 7392 2872 7404
rect 2827 7364 2872 7392
rect 2866 7352 2872 7364
rect 2924 7352 2930 7404
rect 3881 7395 3939 7401
rect 3881 7361 3893 7395
rect 3927 7361 3939 7395
rect 3881 7355 3939 7361
rect 4341 7395 4399 7401
rect 4341 7361 4353 7395
rect 4387 7392 4399 7395
rect 4890 7392 4896 7404
rect 4387 7364 4896 7392
rect 4387 7361 4399 7364
rect 4341 7355 4399 7361
rect 3896 7324 3924 7355
rect 4890 7352 4896 7364
rect 4948 7352 4954 7404
rect 5074 7352 5080 7404
rect 5132 7392 5138 7404
rect 5537 7395 5595 7401
rect 5132 7364 5488 7392
rect 5132 7352 5138 7364
rect 4617 7327 4675 7333
rect 4617 7324 4629 7327
rect 3896 7296 4629 7324
rect 4617 7293 4629 7296
rect 4663 7293 4675 7327
rect 4617 7287 4675 7293
rect 5353 7327 5411 7333
rect 5353 7293 5365 7327
rect 5399 7293 5411 7327
rect 5460 7324 5488 7364
rect 5537 7361 5549 7395
rect 5583 7392 5595 7395
rect 5902 7392 5908 7404
rect 5583 7364 5908 7392
rect 5583 7361 5595 7364
rect 5537 7355 5595 7361
rect 5902 7352 5908 7364
rect 5960 7352 5966 7404
rect 6641 7395 6699 7401
rect 6641 7361 6653 7395
rect 6687 7361 6699 7395
rect 6641 7355 6699 7361
rect 6656 7324 6684 7355
rect 7926 7352 7932 7404
rect 7984 7392 7990 7404
rect 8113 7395 8171 7401
rect 8113 7392 8125 7395
rect 7984 7364 8125 7392
rect 7984 7352 7990 7364
rect 8113 7361 8125 7364
rect 8159 7361 8171 7395
rect 8113 7355 8171 7361
rect 8202 7352 8208 7404
rect 8260 7392 8266 7404
rect 8938 7392 8944 7404
rect 8260 7364 8353 7392
rect 8899 7364 8944 7392
rect 8260 7352 8266 7364
rect 8938 7352 8944 7364
rect 8996 7352 9002 7404
rect 9309 7395 9367 7401
rect 9309 7361 9321 7395
rect 9355 7392 9367 7395
rect 10152 7392 10180 7500
rect 11238 7488 11244 7500
rect 11296 7488 11302 7540
rect 11701 7531 11759 7537
rect 11701 7497 11713 7531
rect 11747 7528 11759 7531
rect 11882 7528 11888 7540
rect 11747 7500 11888 7528
rect 11747 7497 11759 7500
rect 11701 7491 11759 7497
rect 11882 7488 11888 7500
rect 11940 7488 11946 7540
rect 12066 7488 12072 7540
rect 12124 7488 12130 7540
rect 12710 7528 12716 7540
rect 12671 7500 12716 7528
rect 12710 7488 12716 7500
rect 12768 7488 12774 7540
rect 14921 7531 14979 7537
rect 14921 7497 14933 7531
rect 14967 7497 14979 7531
rect 14921 7491 14979 7497
rect 15013 7531 15071 7537
rect 15013 7497 15025 7531
rect 15059 7528 15071 7531
rect 15470 7528 15476 7540
rect 15059 7500 15476 7528
rect 15059 7497 15071 7500
rect 15013 7491 15071 7497
rect 10962 7460 10968 7472
rect 10520 7432 10968 7460
rect 10318 7392 10324 7404
rect 9355 7364 10180 7392
rect 10279 7364 10324 7392
rect 9355 7361 9367 7364
rect 9309 7355 9367 7361
rect 10318 7352 10324 7364
rect 10376 7352 10382 7404
rect 5460 7296 6684 7324
rect 6825 7327 6883 7333
rect 5353 7287 5411 7293
rect 6825 7293 6837 7327
rect 6871 7324 6883 7327
rect 7834 7324 7840 7336
rect 6871 7296 7840 7324
rect 6871 7293 6883 7296
rect 6825 7287 6883 7293
rect 2133 7259 2191 7265
rect 2133 7225 2145 7259
rect 2179 7256 2191 7259
rect 2406 7256 2412 7268
rect 2179 7228 2412 7256
rect 2179 7225 2191 7228
rect 2133 7219 2191 7225
rect 2406 7216 2412 7228
rect 2464 7216 2470 7268
rect 4522 7256 4528 7268
rect 4483 7228 4528 7256
rect 4522 7216 4528 7228
rect 4580 7216 4586 7268
rect 2958 7188 2964 7200
rect 2919 7160 2964 7188
rect 2958 7148 2964 7160
rect 3016 7148 3022 7200
rect 3789 7191 3847 7197
rect 3789 7157 3801 7191
rect 3835 7188 3847 7191
rect 4154 7188 4160 7200
rect 3835 7160 4160 7188
rect 3835 7157 3847 7160
rect 3789 7151 3847 7157
rect 4154 7148 4160 7160
rect 4212 7148 4218 7200
rect 4246 7148 4252 7200
rect 4304 7188 4310 7200
rect 4433 7191 4491 7197
rect 4433 7188 4445 7191
rect 4304 7160 4445 7188
rect 4304 7148 4310 7160
rect 4433 7157 4445 7160
rect 4479 7157 4491 7191
rect 4632 7188 4660 7287
rect 5368 7256 5396 7287
rect 5534 7256 5540 7268
rect 5368 7228 5540 7256
rect 5534 7216 5540 7228
rect 5592 7216 5598 7268
rect 5902 7216 5908 7268
rect 5960 7256 5966 7268
rect 6546 7256 6552 7268
rect 5960 7228 6552 7256
rect 5960 7216 5966 7228
rect 6546 7216 6552 7228
rect 6604 7256 6610 7268
rect 6840 7256 6868 7287
rect 7834 7284 7840 7296
rect 7892 7284 7898 7336
rect 8021 7327 8079 7333
rect 8021 7324 8033 7327
rect 7944 7296 8033 7324
rect 6604 7228 6868 7256
rect 6604 7216 6610 7228
rect 7558 7216 7564 7268
rect 7616 7256 7622 7268
rect 7944 7256 7972 7296
rect 8021 7293 8033 7296
rect 8067 7293 8079 7327
rect 8021 7287 8079 7293
rect 8297 7327 8355 7333
rect 8297 7293 8309 7327
rect 8343 7293 8355 7327
rect 8297 7287 8355 7293
rect 8481 7327 8539 7333
rect 8481 7293 8493 7327
rect 8527 7324 8539 7327
rect 10134 7324 10140 7336
rect 8527 7296 10140 7324
rect 8527 7293 8539 7296
rect 8481 7287 8539 7293
rect 8312 7256 8340 7287
rect 10134 7284 10140 7296
rect 10192 7284 10198 7336
rect 10229 7327 10287 7333
rect 10229 7293 10241 7327
rect 10275 7324 10287 7327
rect 10520 7324 10548 7432
rect 10962 7420 10968 7432
rect 11020 7420 11026 7472
rect 11057 7463 11115 7469
rect 11057 7429 11069 7463
rect 11103 7460 11115 7463
rect 11606 7460 11612 7472
rect 11103 7432 11612 7460
rect 11103 7429 11115 7432
rect 11057 7423 11115 7429
rect 11606 7420 11612 7432
rect 11664 7420 11670 7472
rect 12084 7401 12112 7488
rect 14734 7460 14740 7472
rect 14695 7432 14740 7460
rect 14734 7420 14740 7432
rect 14792 7420 14798 7472
rect 14936 7460 14964 7491
rect 15470 7488 15476 7500
rect 15528 7528 15534 7540
rect 15838 7528 15844 7540
rect 15528 7500 15844 7528
rect 15528 7488 15534 7500
rect 15838 7488 15844 7500
rect 15896 7488 15902 7540
rect 17126 7488 17132 7540
rect 17184 7528 17190 7540
rect 17184 7500 17816 7528
rect 17184 7488 17190 7500
rect 15289 7463 15347 7469
rect 14936 7432 15240 7460
rect 12069 7395 12127 7401
rect 12069 7361 12081 7395
rect 12115 7361 12127 7395
rect 12894 7392 12900 7404
rect 12855 7364 12900 7392
rect 12069 7355 12127 7361
rect 12894 7352 12900 7364
rect 12952 7352 12958 7404
rect 13170 7392 13176 7404
rect 13131 7364 13176 7392
rect 13170 7352 13176 7364
rect 13228 7352 13234 7404
rect 15010 7352 15016 7404
rect 15068 7392 15074 7404
rect 15105 7395 15163 7401
rect 15105 7392 15117 7395
rect 15068 7364 15117 7392
rect 15068 7352 15074 7364
rect 15105 7361 15117 7364
rect 15151 7361 15163 7395
rect 15212 7392 15240 7432
rect 15289 7429 15301 7463
rect 15335 7460 15347 7463
rect 15335 7432 17540 7460
rect 15335 7429 15347 7432
rect 15289 7423 15347 7429
rect 15746 7392 15752 7404
rect 15212 7364 15752 7392
rect 15105 7355 15163 7361
rect 15746 7352 15752 7364
rect 15804 7352 15810 7404
rect 15933 7395 15991 7401
rect 15933 7361 15945 7395
rect 15979 7392 15991 7395
rect 16390 7392 16396 7404
rect 15979 7364 16396 7392
rect 15979 7361 15991 7364
rect 15933 7355 15991 7361
rect 16390 7352 16396 7364
rect 16448 7392 16454 7404
rect 16942 7392 16948 7404
rect 16448 7364 16948 7392
rect 16448 7352 16454 7364
rect 16942 7352 16948 7364
rect 17000 7352 17006 7404
rect 17034 7352 17040 7404
rect 17092 7392 17098 7404
rect 17512 7401 17540 7432
rect 17313 7395 17371 7401
rect 17313 7392 17325 7395
rect 17092 7364 17325 7392
rect 17092 7352 17098 7364
rect 17313 7361 17325 7364
rect 17359 7361 17371 7395
rect 17313 7355 17371 7361
rect 17497 7395 17555 7401
rect 17497 7361 17509 7395
rect 17543 7392 17555 7395
rect 17586 7392 17592 7404
rect 17543 7364 17592 7392
rect 17543 7361 17555 7364
rect 17497 7355 17555 7361
rect 17586 7352 17592 7364
rect 17644 7352 17650 7404
rect 17788 7392 17816 7500
rect 22830 7488 22836 7540
rect 22888 7528 22894 7540
rect 23017 7531 23075 7537
rect 23017 7528 23029 7531
rect 22888 7500 23029 7528
rect 22888 7488 22894 7500
rect 23017 7497 23029 7500
rect 23063 7497 23075 7531
rect 23017 7491 23075 7497
rect 20257 7463 20315 7469
rect 20257 7429 20269 7463
rect 20303 7460 20315 7463
rect 20303 7432 22094 7460
rect 20303 7429 20315 7432
rect 20257 7423 20315 7429
rect 17862 7392 17868 7404
rect 17775 7364 17868 7392
rect 17862 7352 17868 7364
rect 17920 7392 17926 7404
rect 18049 7395 18107 7401
rect 18049 7392 18061 7395
rect 17920 7364 18061 7392
rect 17920 7352 17926 7364
rect 18049 7361 18061 7364
rect 18095 7361 18107 7395
rect 18049 7355 18107 7361
rect 18233 7395 18291 7401
rect 18233 7361 18245 7395
rect 18279 7392 18291 7395
rect 18506 7392 18512 7404
rect 18279 7364 18512 7392
rect 18279 7361 18291 7364
rect 18233 7355 18291 7361
rect 18506 7352 18512 7364
rect 18564 7352 18570 7404
rect 19518 7392 19524 7404
rect 19479 7364 19524 7392
rect 19518 7352 19524 7364
rect 19576 7352 19582 7404
rect 19794 7392 19800 7404
rect 19755 7364 19800 7392
rect 19794 7352 19800 7364
rect 19852 7352 19858 7404
rect 20622 7352 20628 7404
rect 20680 7392 20686 7404
rect 20809 7395 20867 7401
rect 20809 7392 20821 7395
rect 20680 7364 20821 7392
rect 20680 7352 20686 7364
rect 20809 7361 20821 7364
rect 20855 7361 20867 7395
rect 20809 7355 20867 7361
rect 20993 7395 21051 7401
rect 20993 7361 21005 7395
rect 21039 7361 21051 7395
rect 20993 7355 21051 7361
rect 10275 7296 10548 7324
rect 10275 7293 10287 7296
rect 10229 7287 10287 7293
rect 8386 7256 8392 7268
rect 7616 7228 7972 7256
rect 8299 7228 8392 7256
rect 7616 7216 7622 7228
rect 5920 7188 5948 7216
rect 7852 7200 7880 7228
rect 8386 7216 8392 7228
rect 8444 7256 8450 7268
rect 9306 7256 9312 7268
rect 8444 7228 9312 7256
rect 8444 7216 8450 7228
rect 9306 7216 9312 7228
rect 9364 7216 9370 7268
rect 9493 7259 9551 7265
rect 9493 7225 9505 7259
rect 9539 7256 9551 7259
rect 9674 7256 9680 7268
rect 9539 7228 9680 7256
rect 9539 7225 9551 7228
rect 9493 7219 9551 7225
rect 9674 7216 9680 7228
rect 9732 7216 9738 7268
rect 4632 7160 5948 7188
rect 4433 7151 4491 7157
rect 7834 7148 7840 7200
rect 7892 7148 7898 7200
rect 7926 7148 7932 7200
rect 7984 7188 7990 7200
rect 10244 7188 10272 7287
rect 11054 7284 11060 7336
rect 11112 7324 11118 7336
rect 11877 7327 11935 7333
rect 11877 7324 11889 7327
rect 11112 7296 11889 7324
rect 11112 7284 11118 7296
rect 11877 7293 11889 7296
rect 11923 7293 11935 7327
rect 11877 7287 11935 7293
rect 11977 7327 12035 7333
rect 11977 7293 11989 7327
rect 12023 7293 12035 7327
rect 11977 7287 12035 7293
rect 10594 7216 10600 7268
rect 10652 7256 10658 7268
rect 11993 7256 12021 7287
rect 12158 7284 12164 7336
rect 12216 7324 12222 7336
rect 13081 7327 13139 7333
rect 12216 7296 12261 7324
rect 12216 7284 12222 7296
rect 13081 7293 13093 7327
rect 13127 7324 13139 7327
rect 14918 7324 14924 7336
rect 13127 7296 14924 7324
rect 13127 7293 13139 7296
rect 13081 7287 13139 7293
rect 14918 7284 14924 7296
rect 14976 7284 14982 7336
rect 20254 7284 20260 7336
rect 20312 7324 20318 7336
rect 21008 7324 21036 7355
rect 21174 7324 21180 7336
rect 20312 7296 21180 7324
rect 20312 7284 20318 7296
rect 21174 7284 21180 7296
rect 21232 7284 21238 7336
rect 22066 7324 22094 7432
rect 22373 7395 22431 7401
rect 22373 7361 22385 7395
rect 22419 7392 22431 7395
rect 22462 7392 22468 7404
rect 22419 7364 22468 7392
rect 22419 7361 22431 7364
rect 22373 7355 22431 7361
rect 22462 7352 22468 7364
rect 22520 7352 22526 7404
rect 22557 7395 22615 7401
rect 22557 7361 22569 7395
rect 22603 7361 22615 7395
rect 22557 7355 22615 7361
rect 22649 7395 22707 7401
rect 22649 7361 22661 7395
rect 22695 7361 22707 7395
rect 22649 7355 22707 7361
rect 22787 7395 22845 7401
rect 22787 7361 22799 7395
rect 22833 7392 22845 7395
rect 22922 7392 22928 7404
rect 22833 7364 22928 7392
rect 22833 7361 22845 7364
rect 22787 7355 22845 7361
rect 22278 7324 22284 7336
rect 22066 7296 22284 7324
rect 22278 7284 22284 7296
rect 22336 7324 22342 7336
rect 22572 7324 22600 7355
rect 22336 7296 22600 7324
rect 22336 7284 22342 7296
rect 12710 7256 12716 7268
rect 10652 7228 12716 7256
rect 10652 7216 10658 7228
rect 12710 7216 12716 7228
rect 12768 7216 12774 7268
rect 16758 7216 16764 7268
rect 16816 7256 16822 7268
rect 19242 7256 19248 7268
rect 16816 7228 19248 7256
rect 16816 7216 16822 7228
rect 19242 7216 19248 7228
rect 19300 7256 19306 7268
rect 19613 7259 19671 7265
rect 19613 7256 19625 7259
rect 19300 7228 19625 7256
rect 19300 7216 19306 7228
rect 19613 7225 19625 7228
rect 19659 7225 19671 7259
rect 19613 7219 19671 7225
rect 20993 7259 21051 7265
rect 20993 7225 21005 7259
rect 21039 7256 21051 7259
rect 22094 7256 22100 7268
rect 21039 7228 22100 7256
rect 21039 7225 21051 7228
rect 20993 7219 21051 7225
rect 22094 7216 22100 7228
rect 22152 7216 22158 7268
rect 22664 7200 22692 7355
rect 22922 7352 22928 7364
rect 22980 7352 22986 7404
rect 7984 7160 10272 7188
rect 7984 7148 7990 7160
rect 10318 7148 10324 7200
rect 10376 7188 10382 7200
rect 10376 7160 10421 7188
rect 10376 7148 10382 7160
rect 11698 7148 11704 7200
rect 11756 7188 11762 7200
rect 12066 7188 12072 7200
rect 11756 7160 12072 7188
rect 11756 7148 11762 7160
rect 12066 7148 12072 7160
rect 12124 7148 12130 7200
rect 12894 7188 12900 7200
rect 12855 7160 12900 7188
rect 12894 7148 12900 7160
rect 12952 7148 12958 7200
rect 13814 7188 13820 7200
rect 13775 7160 13820 7188
rect 13814 7148 13820 7160
rect 13872 7188 13878 7200
rect 14642 7188 14648 7200
rect 13872 7160 14648 7188
rect 13872 7148 13878 7160
rect 14642 7148 14648 7160
rect 14700 7148 14706 7200
rect 15654 7148 15660 7200
rect 15712 7188 15718 7200
rect 15933 7191 15991 7197
rect 15933 7188 15945 7191
rect 15712 7160 15945 7188
rect 15712 7148 15718 7160
rect 15933 7157 15945 7160
rect 15979 7188 15991 7191
rect 16022 7188 16028 7200
rect 15979 7160 16028 7188
rect 15979 7157 15991 7160
rect 15933 7151 15991 7157
rect 16022 7148 16028 7160
rect 16080 7148 16086 7200
rect 18509 7191 18567 7197
rect 18509 7157 18521 7191
rect 18555 7188 18567 7191
rect 18690 7188 18696 7200
rect 18555 7160 18696 7188
rect 18555 7157 18567 7160
rect 18509 7151 18567 7157
rect 18690 7148 18696 7160
rect 18748 7148 18754 7200
rect 22370 7148 22376 7200
rect 22428 7188 22434 7200
rect 22646 7188 22652 7200
rect 22428 7160 22652 7188
rect 22428 7148 22434 7160
rect 22646 7148 22652 7160
rect 22704 7148 22710 7200
rect 1104 7098 23828 7120
rect 1104 7046 3790 7098
rect 3842 7046 3854 7098
rect 3906 7046 3918 7098
rect 3970 7046 3982 7098
rect 4034 7046 4046 7098
rect 4098 7046 9471 7098
rect 9523 7046 9535 7098
rect 9587 7046 9599 7098
rect 9651 7046 9663 7098
rect 9715 7046 9727 7098
rect 9779 7046 15152 7098
rect 15204 7046 15216 7098
rect 15268 7046 15280 7098
rect 15332 7046 15344 7098
rect 15396 7046 15408 7098
rect 15460 7046 20833 7098
rect 20885 7046 20897 7098
rect 20949 7046 20961 7098
rect 21013 7046 21025 7098
rect 21077 7046 21089 7098
rect 21141 7046 23828 7098
rect 1104 7024 23828 7046
rect 2409 6987 2467 6993
rect 2409 6953 2421 6987
rect 2455 6984 2467 6987
rect 3234 6984 3240 6996
rect 2455 6956 3240 6984
rect 2455 6953 2467 6956
rect 2409 6947 2467 6953
rect 3234 6944 3240 6956
rect 3292 6944 3298 6996
rect 7282 6944 7288 6996
rect 7340 6984 7346 6996
rect 8386 6984 8392 6996
rect 7340 6956 8392 6984
rect 7340 6944 7346 6956
rect 8386 6944 8392 6956
rect 8444 6944 8450 6996
rect 8481 6987 8539 6993
rect 8481 6953 8493 6987
rect 8527 6984 8539 6987
rect 11238 6984 11244 6996
rect 8527 6956 11244 6984
rect 8527 6953 8539 6956
rect 8481 6947 8539 6953
rect 11238 6944 11244 6956
rect 11296 6944 11302 6996
rect 12342 6984 12348 6996
rect 11348 6956 12348 6984
rect 5534 6916 5540 6928
rect 2056 6888 5540 6916
rect 2056 6792 2084 6888
rect 5534 6876 5540 6888
rect 5592 6876 5598 6928
rect 9858 6916 9864 6928
rect 5644 6888 6132 6916
rect 3421 6851 3479 6857
rect 3421 6817 3433 6851
rect 3467 6848 3479 6851
rect 4798 6848 4804 6860
rect 3467 6820 4804 6848
rect 3467 6817 3479 6820
rect 3421 6811 3479 6817
rect 4798 6808 4804 6820
rect 4856 6808 4862 6860
rect 5350 6848 5356 6860
rect 5311 6820 5356 6848
rect 5350 6808 5356 6820
rect 5408 6808 5414 6860
rect 2038 6780 2044 6792
rect 1951 6752 2044 6780
rect 2038 6740 2044 6752
rect 2096 6740 2102 6792
rect 2409 6783 2467 6789
rect 2409 6749 2421 6783
rect 2455 6780 2467 6783
rect 2958 6780 2964 6792
rect 2455 6752 2964 6780
rect 2455 6749 2467 6752
rect 2409 6743 2467 6749
rect 2958 6740 2964 6752
rect 3016 6780 3022 6792
rect 3053 6783 3111 6789
rect 3053 6780 3065 6783
rect 3016 6752 3065 6780
rect 3016 6740 3022 6752
rect 3053 6749 3065 6752
rect 3099 6749 3111 6783
rect 3053 6743 3111 6749
rect 2590 6644 2596 6656
rect 2551 6616 2596 6644
rect 2590 6604 2596 6616
rect 2648 6604 2654 6656
rect 3068 6644 3096 6743
rect 3234 6740 3240 6792
rect 3292 6780 3298 6792
rect 4617 6783 4675 6789
rect 3292 6752 3337 6780
rect 3292 6740 3298 6752
rect 4617 6749 4629 6783
rect 4663 6749 4675 6783
rect 4617 6743 4675 6749
rect 4338 6712 4344 6724
rect 4299 6684 4344 6712
rect 4338 6672 4344 6684
rect 4396 6672 4402 6724
rect 4632 6644 4660 6743
rect 5074 6740 5080 6792
rect 5132 6780 5138 6792
rect 5644 6780 5672 6888
rect 5810 6848 5816 6860
rect 5771 6820 5816 6848
rect 5810 6808 5816 6820
rect 5868 6808 5874 6860
rect 5994 6848 6000 6860
rect 5920 6820 6000 6848
rect 5132 6752 5672 6780
rect 5721 6783 5779 6789
rect 5132 6740 5138 6752
rect 5721 6749 5733 6783
rect 5767 6780 5779 6783
rect 5920 6780 5948 6820
rect 5994 6808 6000 6820
rect 6052 6808 6058 6860
rect 6104 6848 6132 6888
rect 7208 6888 8524 6916
rect 7208 6848 7236 6888
rect 6104 6820 7236 6848
rect 8496 6848 8524 6888
rect 9692 6888 9864 6916
rect 9214 6848 9220 6860
rect 8496 6820 9220 6848
rect 9214 6808 9220 6820
rect 9272 6808 9278 6860
rect 9692 6857 9720 6888
rect 9858 6876 9864 6888
rect 9916 6916 9922 6928
rect 10505 6919 10563 6925
rect 9916 6888 10088 6916
rect 9916 6876 9922 6888
rect 9585 6851 9643 6857
rect 9585 6848 9597 6851
rect 9416 6820 9597 6848
rect 6086 6780 6092 6792
rect 5767 6752 5948 6780
rect 6047 6752 6092 6780
rect 5767 6749 5779 6752
rect 5721 6743 5779 6749
rect 6086 6740 6092 6752
rect 6144 6740 6150 6792
rect 6270 6780 6276 6792
rect 6231 6752 6276 6780
rect 6270 6740 6276 6752
rect 6328 6740 6334 6792
rect 7193 6783 7251 6789
rect 7193 6749 7205 6783
rect 7239 6780 7251 6783
rect 7282 6780 7288 6792
rect 7239 6752 7288 6780
rect 7239 6749 7251 6752
rect 7193 6743 7251 6749
rect 7282 6740 7288 6752
rect 7340 6740 7346 6792
rect 7374 6740 7380 6792
rect 7432 6780 7438 6792
rect 7653 6783 7711 6789
rect 7432 6752 7477 6780
rect 7432 6740 7438 6752
rect 7653 6749 7665 6783
rect 7699 6749 7711 6783
rect 7653 6743 7711 6749
rect 5810 6672 5816 6724
rect 5868 6712 5874 6724
rect 7668 6712 7696 6743
rect 7742 6740 7748 6792
rect 7800 6780 7806 6792
rect 8294 6780 8300 6792
rect 7800 6752 7845 6780
rect 8255 6752 8300 6780
rect 7800 6740 7806 6752
rect 8294 6740 8300 6752
rect 8352 6780 8358 6792
rect 9306 6780 9312 6792
rect 8352 6752 9312 6780
rect 8352 6740 8358 6752
rect 9306 6740 9312 6752
rect 9364 6740 9370 6792
rect 5868 6684 7696 6712
rect 5868 6672 5874 6684
rect 9214 6672 9220 6724
rect 9272 6712 9278 6724
rect 9416 6712 9444 6820
rect 9585 6817 9597 6820
rect 9631 6817 9643 6851
rect 9585 6811 9643 6817
rect 9677 6851 9735 6857
rect 9677 6817 9689 6851
rect 9723 6817 9735 6851
rect 9950 6848 9956 6860
rect 9911 6820 9956 6848
rect 9677 6811 9735 6817
rect 9950 6808 9956 6820
rect 10008 6808 10014 6860
rect 10060 6848 10088 6888
rect 10505 6885 10517 6919
rect 10551 6916 10563 6919
rect 11146 6916 11152 6928
rect 10551 6888 11152 6916
rect 10551 6885 10563 6888
rect 10505 6879 10563 6885
rect 11146 6876 11152 6888
rect 11204 6916 11210 6928
rect 11348 6925 11376 6956
rect 12342 6944 12348 6956
rect 12400 6944 12406 6996
rect 12802 6944 12808 6996
rect 12860 6984 12866 6996
rect 15657 6987 15715 6993
rect 15657 6984 15669 6987
rect 12860 6956 15669 6984
rect 12860 6944 12866 6956
rect 15657 6953 15669 6956
rect 15703 6984 15715 6987
rect 16390 6984 16396 6996
rect 15703 6956 16396 6984
rect 15703 6953 15715 6956
rect 15657 6947 15715 6953
rect 16390 6944 16396 6956
rect 16448 6944 16454 6996
rect 22465 6987 22523 6993
rect 22465 6953 22477 6987
rect 22511 6984 22523 6987
rect 22922 6984 22928 6996
rect 22511 6956 22928 6984
rect 22511 6953 22523 6956
rect 22465 6947 22523 6953
rect 22922 6944 22928 6956
rect 22980 6944 22986 6996
rect 11333 6919 11391 6925
rect 11333 6916 11345 6919
rect 11204 6888 11345 6916
rect 11204 6876 11210 6888
rect 11333 6885 11345 6888
rect 11379 6885 11391 6919
rect 11333 6879 11391 6885
rect 11606 6876 11612 6928
rect 11664 6916 11670 6928
rect 13078 6916 13084 6928
rect 11664 6888 13084 6916
rect 11664 6876 11670 6888
rect 13078 6876 13084 6888
rect 13136 6876 13142 6928
rect 13265 6919 13323 6925
rect 13265 6885 13277 6919
rect 13311 6916 13323 6919
rect 13538 6916 13544 6928
rect 13311 6888 13544 6916
rect 13311 6885 13323 6888
rect 13265 6879 13323 6885
rect 10594 6848 10600 6860
rect 10060 6820 10600 6848
rect 10594 6808 10600 6820
rect 10652 6808 10658 6860
rect 12158 6808 12164 6860
rect 12216 6848 12222 6860
rect 12802 6848 12808 6860
rect 12216 6820 12808 6848
rect 12216 6808 12222 6820
rect 12802 6808 12808 6820
rect 12860 6808 12866 6860
rect 9493 6783 9551 6789
rect 9493 6749 9505 6783
rect 9539 6749 9551 6783
rect 9766 6780 9772 6792
rect 9679 6752 9772 6780
rect 9493 6743 9551 6749
rect 9272 6684 9444 6712
rect 9508 6712 9536 6743
rect 9766 6740 9772 6752
rect 9824 6780 9830 6792
rect 10410 6780 10416 6792
rect 9824 6752 10416 6780
rect 9824 6740 9830 6752
rect 10410 6740 10416 6752
rect 10468 6740 10474 6792
rect 11146 6740 11152 6792
rect 11204 6780 11210 6792
rect 13280 6780 13308 6879
rect 13538 6876 13544 6888
rect 13596 6916 13602 6928
rect 14461 6919 14519 6925
rect 14461 6916 14473 6919
rect 13596 6888 14473 6916
rect 13596 6876 13602 6888
rect 14461 6885 14473 6888
rect 14507 6916 14519 6919
rect 15746 6916 15752 6928
rect 14507 6888 15752 6916
rect 14507 6885 14519 6888
rect 14461 6879 14519 6885
rect 15746 6876 15752 6888
rect 15804 6876 15810 6928
rect 19058 6876 19064 6928
rect 19116 6916 19122 6928
rect 22373 6919 22431 6925
rect 19116 6888 19748 6916
rect 19116 6876 19122 6888
rect 14826 6808 14832 6860
rect 14884 6848 14890 6860
rect 14884 6820 15148 6848
rect 14884 6808 14890 6820
rect 11204 6752 13308 6780
rect 11204 6740 11210 6752
rect 14458 6740 14464 6792
rect 14516 6780 14522 6792
rect 15120 6789 15148 6820
rect 16666 6808 16672 6860
rect 16724 6848 16730 6860
rect 17037 6851 17095 6857
rect 17037 6848 17049 6851
rect 16724 6820 17049 6848
rect 16724 6808 16730 6820
rect 17037 6817 17049 6820
rect 17083 6817 17095 6851
rect 17037 6811 17095 6817
rect 17310 6808 17316 6860
rect 17368 6848 17374 6860
rect 17589 6851 17647 6857
rect 17589 6848 17601 6851
rect 17368 6820 17601 6848
rect 17368 6808 17374 6820
rect 17589 6817 17601 6820
rect 17635 6817 17647 6851
rect 18230 6848 18236 6860
rect 18191 6820 18236 6848
rect 17589 6811 17647 6817
rect 18230 6808 18236 6820
rect 18288 6808 18294 6860
rect 19518 6848 19524 6860
rect 18340 6820 19524 6848
rect 18340 6792 18368 6820
rect 19518 6808 19524 6820
rect 19576 6848 19582 6860
rect 19720 6848 19748 6888
rect 22373 6885 22385 6919
rect 22419 6916 22431 6919
rect 23014 6916 23020 6928
rect 22419 6888 23020 6916
rect 22419 6885 22431 6888
rect 22373 6879 22431 6885
rect 20349 6851 20407 6857
rect 20349 6848 20361 6851
rect 19576 6820 19656 6848
rect 19720 6820 20361 6848
rect 19576 6808 19582 6820
rect 14921 6783 14979 6789
rect 14921 6780 14933 6783
rect 14516 6752 14933 6780
rect 14516 6740 14522 6752
rect 14921 6749 14933 6752
rect 14967 6749 14979 6783
rect 14921 6743 14979 6749
rect 15105 6783 15163 6789
rect 15105 6749 15117 6783
rect 15151 6749 15163 6783
rect 18322 6780 18328 6792
rect 18283 6752 18328 6780
rect 15105 6743 15163 6749
rect 10962 6712 10968 6724
rect 9508 6684 10968 6712
rect 9272 6672 9278 6684
rect 10962 6672 10968 6684
rect 11020 6672 11026 6724
rect 11514 6712 11520 6724
rect 11072 6684 11520 6712
rect 6546 6644 6552 6656
rect 3068 6616 6552 6644
rect 6546 6604 6552 6616
rect 6604 6604 6610 6656
rect 7742 6604 7748 6656
rect 7800 6644 7806 6656
rect 10226 6644 10232 6656
rect 7800 6616 10232 6644
rect 7800 6604 7806 6616
rect 10226 6604 10232 6616
rect 10284 6604 10290 6656
rect 10594 6604 10600 6656
rect 10652 6644 10658 6656
rect 11072 6644 11100 6684
rect 11514 6672 11520 6684
rect 11572 6712 11578 6724
rect 14182 6712 14188 6724
rect 11572 6684 12112 6712
rect 11572 6672 11578 6684
rect 10652 6616 11100 6644
rect 10652 6604 10658 6616
rect 11330 6604 11336 6656
rect 11388 6644 11394 6656
rect 11606 6644 11612 6656
rect 11388 6616 11612 6644
rect 11388 6604 11394 6616
rect 11606 6604 11612 6616
rect 11664 6604 11670 6656
rect 11698 6604 11704 6656
rect 11756 6644 11762 6656
rect 11793 6647 11851 6653
rect 11793 6644 11805 6647
rect 11756 6616 11805 6644
rect 11756 6604 11762 6616
rect 11793 6613 11805 6616
rect 11839 6613 11851 6647
rect 12084 6644 12112 6684
rect 12268 6684 14188 6712
rect 12268 6644 12296 6684
rect 14182 6672 14188 6684
rect 14240 6672 14246 6724
rect 12084 6616 12296 6644
rect 11793 6607 11851 6613
rect 12342 6604 12348 6656
rect 12400 6644 12406 6656
rect 14090 6644 14096 6656
rect 12400 6616 14096 6644
rect 12400 6604 12406 6616
rect 14090 6604 14096 6616
rect 14148 6604 14154 6656
rect 14936 6644 14964 6743
rect 18322 6740 18328 6752
rect 18380 6740 18386 6792
rect 18877 6783 18935 6789
rect 18877 6749 18889 6783
rect 18923 6780 18935 6783
rect 19242 6780 19248 6792
rect 18923 6752 19248 6780
rect 18923 6749 18935 6752
rect 18877 6743 18935 6749
rect 19242 6740 19248 6752
rect 19300 6780 19306 6792
rect 19628 6789 19656 6820
rect 20349 6817 20361 6820
rect 20395 6817 20407 6851
rect 20349 6811 20407 6817
rect 21542 6808 21548 6860
rect 21600 6848 21606 6860
rect 22281 6851 22339 6857
rect 22281 6848 22293 6851
rect 21600 6820 22293 6848
rect 21600 6808 21606 6820
rect 22281 6817 22293 6820
rect 22327 6817 22339 6851
rect 22281 6811 22339 6817
rect 19429 6783 19487 6789
rect 19429 6780 19441 6783
rect 19300 6752 19441 6780
rect 19300 6740 19306 6752
rect 19429 6749 19441 6752
rect 19475 6749 19487 6783
rect 19429 6743 19487 6749
rect 19613 6783 19671 6789
rect 19613 6749 19625 6783
rect 19659 6749 19671 6783
rect 19613 6743 19671 6749
rect 19981 6783 20039 6789
rect 19981 6749 19993 6783
rect 20027 6749 20039 6783
rect 19981 6743 20039 6749
rect 20165 6783 20223 6789
rect 20165 6749 20177 6783
rect 20211 6749 20223 6783
rect 20165 6743 20223 6749
rect 15013 6715 15071 6721
rect 15013 6681 15025 6715
rect 15059 6712 15071 6715
rect 15930 6712 15936 6724
rect 15059 6684 15936 6712
rect 15059 6681 15071 6684
rect 15013 6675 15071 6681
rect 15930 6672 15936 6684
rect 15988 6672 15994 6724
rect 16666 6672 16672 6724
rect 16724 6712 16730 6724
rect 16724 6684 17816 6712
rect 16724 6672 16730 6684
rect 17788 6656 17816 6684
rect 18506 6672 18512 6724
rect 18564 6712 18570 6724
rect 19996 6712 20024 6743
rect 18564 6684 20024 6712
rect 18564 6672 18570 6684
rect 17494 6644 17500 6656
rect 14936 6616 17500 6644
rect 17494 6604 17500 6616
rect 17552 6604 17558 6656
rect 17770 6604 17776 6656
rect 17828 6644 17834 6656
rect 18782 6644 18788 6656
rect 17828 6616 18788 6644
rect 17828 6604 17834 6616
rect 18782 6604 18788 6616
rect 18840 6604 18846 6656
rect 19150 6604 19156 6656
rect 19208 6644 19214 6656
rect 20180 6644 20208 6743
rect 21266 6740 21272 6792
rect 21324 6780 21330 6792
rect 21361 6783 21419 6789
rect 21361 6780 21373 6783
rect 21324 6752 21373 6780
rect 21324 6740 21330 6752
rect 21361 6749 21373 6752
rect 21407 6749 21419 6783
rect 21361 6743 21419 6749
rect 21637 6715 21695 6721
rect 21637 6681 21649 6715
rect 21683 6712 21695 6715
rect 22186 6712 22192 6724
rect 21683 6684 22192 6712
rect 21683 6681 21695 6684
rect 21637 6675 21695 6681
rect 22186 6672 22192 6684
rect 22244 6712 22250 6724
rect 22388 6712 22416 6879
rect 23014 6876 23020 6888
rect 23072 6876 23078 6928
rect 23198 6848 23204 6860
rect 23159 6820 23204 6848
rect 23198 6808 23204 6820
rect 23256 6808 23262 6860
rect 22646 6780 22652 6792
rect 22607 6752 22652 6780
rect 22646 6740 22652 6752
rect 22704 6740 22710 6792
rect 22244 6684 22416 6712
rect 22244 6672 22250 6684
rect 19208 6616 20208 6644
rect 19208 6604 19214 6616
rect 21910 6604 21916 6656
rect 21968 6644 21974 6656
rect 22557 6647 22615 6653
rect 22557 6644 22569 6647
rect 21968 6616 22569 6644
rect 21968 6604 21974 6616
rect 22557 6613 22569 6616
rect 22603 6613 22615 6647
rect 22557 6607 22615 6613
rect 1104 6554 23987 6576
rect 1104 6502 6630 6554
rect 6682 6502 6694 6554
rect 6746 6502 6758 6554
rect 6810 6502 6822 6554
rect 6874 6502 6886 6554
rect 6938 6502 12311 6554
rect 12363 6502 12375 6554
rect 12427 6502 12439 6554
rect 12491 6502 12503 6554
rect 12555 6502 12567 6554
rect 12619 6502 17992 6554
rect 18044 6502 18056 6554
rect 18108 6502 18120 6554
rect 18172 6502 18184 6554
rect 18236 6502 18248 6554
rect 18300 6502 23673 6554
rect 23725 6502 23737 6554
rect 23789 6502 23801 6554
rect 23853 6502 23865 6554
rect 23917 6502 23929 6554
rect 23981 6502 23987 6554
rect 1104 6480 23987 6502
rect 3421 6443 3479 6449
rect 3421 6409 3433 6443
rect 3467 6440 3479 6443
rect 3467 6412 6316 6440
rect 3467 6409 3479 6412
rect 3421 6403 3479 6409
rect 4154 6372 4160 6384
rect 4115 6344 4160 6372
rect 4154 6332 4160 6344
rect 4212 6332 4218 6384
rect 4617 6375 4675 6381
rect 4617 6341 4629 6375
rect 4663 6372 4675 6375
rect 5074 6372 5080 6384
rect 4663 6344 5080 6372
rect 4663 6341 4675 6344
rect 4617 6335 4675 6341
rect 5074 6332 5080 6344
rect 5132 6332 5138 6384
rect 5994 6372 6000 6384
rect 5955 6344 6000 6372
rect 5994 6332 6000 6344
rect 6052 6332 6058 6384
rect 2225 6307 2283 6313
rect 2225 6273 2237 6307
rect 2271 6273 2283 6307
rect 2406 6304 2412 6316
rect 2367 6276 2412 6304
rect 2225 6267 2283 6273
rect 2240 6236 2268 6267
rect 2406 6264 2412 6276
rect 2464 6264 2470 6316
rect 2590 6264 2596 6316
rect 2648 6304 2654 6316
rect 2685 6307 2743 6313
rect 2685 6304 2697 6307
rect 2648 6276 2697 6304
rect 2648 6264 2654 6276
rect 2685 6273 2697 6276
rect 2731 6273 2743 6307
rect 2685 6267 2743 6273
rect 2774 6264 2780 6316
rect 2832 6304 2838 6316
rect 3050 6304 3056 6316
rect 2832 6276 2877 6304
rect 3011 6276 3056 6304
rect 2832 6264 2838 6276
rect 3050 6264 3056 6276
rect 3108 6264 3114 6316
rect 4249 6307 4307 6313
rect 4249 6273 4261 6307
rect 4295 6304 4307 6307
rect 4798 6304 4804 6316
rect 4295 6276 4804 6304
rect 4295 6273 4307 6276
rect 4249 6267 4307 6273
rect 4798 6264 4804 6276
rect 4856 6264 4862 6316
rect 5261 6307 5319 6313
rect 5261 6273 5273 6307
rect 5307 6273 5319 6307
rect 5534 6304 5540 6316
rect 5495 6276 5540 6304
rect 5261 6267 5319 6273
rect 3694 6236 3700 6248
rect 2240 6208 3700 6236
rect 3694 6196 3700 6208
rect 3752 6196 3758 6248
rect 4709 6239 4767 6245
rect 4709 6205 4721 6239
rect 4755 6236 4767 6239
rect 5276 6236 5304 6267
rect 5534 6264 5540 6276
rect 5592 6264 5598 6316
rect 4755 6208 5304 6236
rect 5353 6239 5411 6245
rect 4755 6205 4767 6208
rect 4709 6199 4767 6205
rect 5353 6205 5365 6239
rect 5399 6236 5411 6239
rect 5718 6236 5724 6248
rect 5399 6208 5724 6236
rect 5399 6205 5411 6208
rect 5353 6199 5411 6205
rect 2958 6128 2964 6180
rect 3016 6168 3022 6180
rect 4724 6168 4752 6199
rect 5718 6196 5724 6208
rect 5776 6196 5782 6248
rect 6288 6236 6316 6412
rect 6362 6400 6368 6452
rect 6420 6440 6426 6452
rect 6733 6443 6791 6449
rect 6733 6440 6745 6443
rect 6420 6412 6745 6440
rect 6420 6400 6426 6412
rect 6733 6409 6745 6412
rect 6779 6409 6791 6443
rect 6733 6403 6791 6409
rect 6825 6443 6883 6449
rect 6825 6409 6837 6443
rect 6871 6440 6883 6443
rect 7006 6440 7012 6452
rect 6871 6412 7012 6440
rect 6871 6409 6883 6412
rect 6825 6403 6883 6409
rect 7006 6400 7012 6412
rect 7064 6400 7070 6452
rect 8386 6440 8392 6452
rect 7116 6412 8392 6440
rect 6454 6332 6460 6384
rect 6512 6372 6518 6384
rect 7116 6381 7144 6412
rect 8386 6400 8392 6412
rect 8444 6400 8450 6452
rect 8478 6400 8484 6452
rect 8536 6440 8542 6452
rect 8536 6412 8616 6440
rect 8536 6400 8542 6412
rect 6917 6375 6975 6381
rect 6917 6372 6929 6375
rect 6512 6344 6929 6372
rect 6512 6332 6518 6344
rect 6917 6341 6929 6344
rect 6963 6341 6975 6375
rect 6917 6335 6975 6341
rect 7101 6375 7159 6381
rect 7101 6341 7113 6375
rect 7147 6341 7159 6375
rect 7101 6335 7159 6341
rect 8294 6332 8300 6384
rect 8352 6372 8358 6384
rect 8352 6344 8397 6372
rect 8352 6332 8358 6344
rect 6546 6304 6552 6316
rect 6507 6276 6552 6304
rect 6546 6264 6552 6276
rect 6604 6264 6610 6316
rect 8018 6304 8024 6316
rect 7979 6276 8024 6304
rect 8018 6264 8024 6276
rect 8076 6264 8082 6316
rect 8114 6307 8172 6313
rect 8114 6273 8126 6307
rect 8160 6273 8172 6307
rect 8114 6267 8172 6273
rect 6914 6236 6920 6248
rect 6288 6208 6920 6236
rect 6914 6196 6920 6208
rect 6972 6196 6978 6248
rect 3016 6140 4752 6168
rect 3016 6128 3022 6140
rect 6270 6128 6276 6180
rect 6328 6168 6334 6180
rect 7650 6168 7656 6180
rect 6328 6140 7656 6168
rect 6328 6128 6334 6140
rect 7650 6128 7656 6140
rect 7708 6168 7714 6180
rect 8128 6168 8156 6267
rect 8202 6264 8208 6316
rect 8260 6304 8266 6316
rect 8386 6307 8444 6313
rect 8386 6304 8398 6307
rect 8260 6276 8398 6304
rect 8260 6264 8266 6276
rect 8386 6273 8398 6276
rect 8432 6273 8444 6307
rect 8386 6267 8444 6273
rect 8486 6307 8544 6313
rect 8486 6273 8498 6307
rect 8532 6304 8544 6307
rect 8588 6304 8616 6412
rect 8938 6400 8944 6452
rect 8996 6440 9002 6452
rect 9674 6440 9680 6452
rect 8996 6412 9680 6440
rect 8996 6400 9002 6412
rect 9674 6400 9680 6412
rect 9732 6400 9738 6452
rect 9769 6443 9827 6449
rect 9769 6409 9781 6443
rect 9815 6440 9827 6443
rect 10042 6440 10048 6452
rect 9815 6412 10048 6440
rect 9815 6409 9827 6412
rect 9769 6403 9827 6409
rect 10042 6400 10048 6412
rect 10100 6400 10106 6452
rect 11054 6440 11060 6452
rect 11015 6412 11060 6440
rect 11054 6400 11060 6412
rect 11112 6400 11118 6452
rect 12986 6440 12992 6452
rect 12912 6412 12992 6440
rect 8846 6332 8852 6384
rect 8904 6372 8910 6384
rect 9950 6372 9956 6384
rect 8904 6344 9956 6372
rect 8904 6332 8910 6344
rect 9950 6332 9956 6344
rect 10008 6332 10014 6384
rect 11238 6332 11244 6384
rect 11296 6372 11302 6384
rect 12912 6381 12940 6412
rect 12986 6400 12992 6412
rect 13044 6400 13050 6452
rect 13170 6400 13176 6452
rect 13228 6440 13234 6452
rect 13725 6443 13783 6449
rect 13725 6440 13737 6443
rect 13228 6412 13737 6440
rect 13228 6400 13234 6412
rect 13725 6409 13737 6412
rect 13771 6409 13783 6443
rect 13725 6403 13783 6409
rect 16022 6400 16028 6452
rect 16080 6440 16086 6452
rect 18138 6440 18144 6452
rect 16080 6412 18144 6440
rect 16080 6400 16086 6412
rect 18138 6400 18144 6412
rect 18196 6400 18202 6452
rect 18325 6443 18383 6449
rect 18325 6409 18337 6443
rect 18371 6440 18383 6443
rect 19334 6440 19340 6452
rect 18371 6412 19340 6440
rect 18371 6409 18383 6412
rect 18325 6403 18383 6409
rect 19334 6400 19340 6412
rect 19392 6400 19398 6452
rect 21358 6400 21364 6452
rect 21416 6440 21422 6452
rect 22005 6443 22063 6449
rect 22005 6440 22017 6443
rect 21416 6412 22017 6440
rect 21416 6400 21422 6412
rect 22005 6409 22017 6412
rect 22051 6409 22063 6443
rect 22005 6403 22063 6409
rect 22922 6400 22928 6452
rect 22980 6440 22986 6452
rect 23017 6443 23075 6449
rect 23017 6440 23029 6443
rect 22980 6412 23029 6440
rect 22980 6400 22986 6412
rect 23017 6409 23029 6412
rect 23063 6409 23075 6443
rect 23017 6403 23075 6409
rect 12897 6375 12955 6381
rect 11296 6344 12434 6372
rect 11296 6332 11302 6344
rect 9122 6304 9128 6316
rect 8532 6276 8616 6304
rect 9083 6276 9128 6304
rect 8532 6273 8544 6276
rect 8486 6267 8544 6273
rect 9122 6264 9128 6276
rect 9180 6264 9186 6316
rect 9309 6307 9367 6313
rect 9309 6273 9321 6307
rect 9355 6273 9367 6307
rect 9309 6267 9367 6273
rect 9401 6307 9459 6313
rect 9401 6273 9413 6307
rect 9447 6273 9459 6307
rect 9401 6267 9459 6273
rect 9324 6236 9352 6267
rect 8680 6208 9352 6236
rect 9416 6236 9444 6267
rect 9490 6264 9496 6316
rect 9548 6304 9554 6316
rect 10134 6304 10140 6316
rect 9548 6276 10140 6304
rect 9548 6264 9554 6276
rect 10134 6264 10140 6276
rect 10192 6264 10198 6316
rect 10226 6264 10232 6316
rect 10284 6304 10290 6316
rect 10873 6307 10931 6313
rect 10873 6304 10885 6307
rect 10284 6276 10885 6304
rect 10284 6264 10290 6276
rect 10873 6273 10885 6276
rect 10919 6273 10931 6307
rect 10873 6267 10931 6273
rect 11149 6307 11207 6313
rect 11149 6273 11161 6307
rect 11195 6304 11207 6307
rect 11701 6307 11759 6313
rect 11701 6304 11713 6307
rect 11195 6276 11713 6304
rect 11195 6273 11207 6276
rect 11149 6267 11207 6273
rect 11701 6273 11713 6276
rect 11747 6273 11759 6307
rect 11701 6267 11759 6273
rect 11885 6307 11943 6313
rect 11885 6273 11897 6307
rect 11931 6273 11943 6307
rect 11885 6267 11943 6273
rect 10042 6236 10048 6248
rect 9416 6208 10048 6236
rect 8680 6177 8708 6208
rect 10042 6196 10048 6208
rect 10100 6196 10106 6248
rect 10502 6196 10508 6248
rect 10560 6236 10566 6248
rect 11900 6236 11928 6267
rect 11974 6264 11980 6316
rect 12032 6304 12038 6316
rect 12069 6307 12127 6313
rect 12069 6304 12081 6307
rect 12032 6276 12081 6304
rect 12032 6264 12038 6276
rect 12069 6273 12081 6276
rect 12115 6273 12127 6307
rect 12069 6267 12127 6273
rect 12158 6264 12164 6316
rect 12216 6304 12222 6316
rect 12406 6304 12434 6344
rect 12897 6341 12909 6375
rect 12943 6341 12955 6375
rect 12897 6335 12955 6341
rect 15010 6332 15016 6384
rect 15068 6372 15074 6384
rect 15105 6375 15163 6381
rect 15105 6372 15117 6375
rect 15068 6344 15117 6372
rect 15068 6332 15074 6344
rect 15105 6341 15117 6344
rect 15151 6372 15163 6375
rect 15657 6375 15715 6381
rect 15151 6344 15608 6372
rect 15151 6341 15163 6344
rect 15105 6335 15163 6341
rect 12805 6307 12863 6313
rect 12805 6304 12817 6307
rect 12216 6276 12261 6304
rect 12406 6276 12817 6304
rect 12216 6264 12222 6276
rect 12805 6273 12817 6276
rect 12851 6273 12863 6307
rect 12986 6304 12992 6316
rect 12947 6276 12992 6304
rect 12805 6267 12863 6273
rect 12986 6264 12992 6276
rect 13044 6264 13050 6316
rect 13127 6307 13185 6313
rect 13127 6273 13139 6307
rect 13173 6304 13185 6307
rect 13906 6304 13912 6316
rect 13173 6276 13912 6304
rect 13173 6273 13185 6276
rect 13127 6267 13185 6273
rect 13906 6264 13912 6276
rect 13964 6264 13970 6316
rect 14182 6304 14188 6316
rect 14143 6276 14188 6304
rect 14182 6264 14188 6276
rect 14240 6264 14246 6316
rect 15197 6307 15255 6313
rect 15197 6273 15209 6307
rect 15243 6273 15255 6307
rect 15580 6304 15608 6344
rect 15657 6341 15669 6375
rect 15703 6372 15715 6375
rect 16574 6372 16580 6384
rect 15703 6344 16580 6372
rect 15703 6341 15715 6344
rect 15657 6335 15715 6341
rect 16574 6332 16580 6344
rect 16632 6332 16638 6384
rect 20714 6332 20720 6384
rect 20772 6372 20778 6384
rect 21269 6375 21327 6381
rect 20772 6344 21220 6372
rect 20772 6332 20778 6344
rect 17310 6304 17316 6316
rect 15580 6276 17316 6304
rect 15197 6267 15255 6273
rect 10560 6208 11928 6236
rect 10560 6196 10566 6208
rect 12710 6196 12716 6248
rect 12768 6236 12774 6248
rect 13265 6239 13323 6245
rect 13265 6236 13277 6239
rect 12768 6208 13277 6236
rect 12768 6196 12774 6208
rect 13265 6205 13277 6208
rect 13311 6205 13323 6239
rect 14090 6236 14096 6248
rect 14051 6208 14096 6236
rect 13265 6199 13323 6205
rect 14090 6196 14096 6208
rect 14148 6196 14154 6248
rect 15010 6196 15016 6248
rect 15068 6236 15074 6248
rect 15212 6236 15240 6267
rect 17310 6264 17316 6276
rect 17368 6264 17374 6316
rect 17865 6307 17923 6313
rect 17865 6273 17877 6307
rect 17911 6273 17923 6307
rect 17865 6267 17923 6273
rect 15068 6208 15240 6236
rect 17880 6236 17908 6267
rect 17954 6264 17960 6316
rect 18012 6304 18018 6316
rect 18138 6304 18144 6316
rect 18012 6276 18057 6304
rect 18099 6276 18144 6304
rect 18012 6264 18018 6276
rect 18138 6264 18144 6276
rect 18196 6264 18202 6316
rect 18506 6304 18512 6316
rect 18248 6276 18512 6304
rect 18248 6248 18276 6276
rect 18506 6264 18512 6276
rect 18564 6264 18570 6316
rect 19150 6264 19156 6316
rect 19208 6304 19214 6316
rect 19245 6307 19303 6313
rect 19245 6304 19257 6307
rect 19208 6276 19257 6304
rect 19208 6264 19214 6276
rect 19245 6273 19257 6276
rect 19291 6273 19303 6307
rect 19245 6267 19303 6273
rect 19797 6307 19855 6313
rect 19797 6273 19809 6307
rect 19843 6273 19855 6307
rect 19797 6267 19855 6273
rect 18230 6236 18236 6248
rect 17880 6208 18236 6236
rect 15068 6196 15074 6208
rect 18230 6196 18236 6208
rect 18288 6196 18294 6248
rect 18524 6236 18552 6264
rect 19812 6236 19840 6267
rect 19886 6264 19892 6316
rect 19944 6304 19950 6316
rect 20530 6304 20536 6316
rect 19944 6276 20536 6304
rect 19944 6264 19950 6276
rect 20530 6264 20536 6276
rect 20588 6304 20594 6316
rect 21192 6313 21220 6344
rect 21269 6341 21281 6375
rect 21315 6372 21327 6375
rect 21542 6372 21548 6384
rect 21315 6344 21548 6372
rect 21315 6341 21327 6344
rect 21269 6335 21327 6341
rect 21542 6332 21548 6344
rect 21600 6332 21606 6384
rect 22940 6372 22968 6400
rect 22572 6344 22968 6372
rect 20901 6307 20959 6313
rect 20901 6304 20913 6307
rect 20588 6276 20913 6304
rect 20588 6264 20594 6276
rect 20901 6273 20913 6276
rect 20947 6273 20959 6307
rect 20901 6267 20959 6273
rect 21177 6307 21235 6313
rect 21177 6273 21189 6307
rect 21223 6304 21235 6307
rect 21818 6304 21824 6316
rect 21223 6276 21824 6304
rect 21223 6273 21235 6276
rect 21177 6267 21235 6273
rect 21818 6264 21824 6276
rect 21876 6264 21882 6316
rect 22186 6304 22192 6316
rect 22147 6276 22192 6304
rect 22186 6264 22192 6276
rect 22244 6264 22250 6316
rect 22370 6264 22376 6316
rect 22428 6304 22434 6316
rect 22428 6276 22473 6304
rect 22428 6264 22434 6276
rect 20346 6236 20352 6248
rect 18524 6208 19840 6236
rect 20307 6208 20352 6236
rect 20346 6196 20352 6208
rect 20404 6196 20410 6248
rect 22465 6239 22523 6245
rect 22465 6205 22477 6239
rect 22511 6236 22523 6239
rect 22572 6236 22600 6344
rect 22922 6304 22928 6316
rect 22511 6208 22600 6236
rect 22664 6276 22928 6304
rect 22511 6205 22523 6208
rect 22465 6199 22523 6205
rect 7708 6140 8156 6168
rect 8665 6171 8723 6177
rect 7708 6128 7714 6140
rect 8665 6137 8677 6171
rect 8711 6137 8723 6171
rect 8665 6131 8723 6137
rect 9122 6128 9128 6180
rect 9180 6168 9186 6180
rect 10778 6168 10784 6180
rect 9180 6140 10784 6168
rect 9180 6128 9186 6140
rect 10778 6128 10784 6140
rect 10836 6168 10842 6180
rect 10836 6140 10916 6168
rect 10836 6128 10842 6140
rect 4798 6060 4804 6112
rect 4856 6100 4862 6112
rect 7742 6100 7748 6112
rect 4856 6072 7748 6100
rect 4856 6060 4862 6072
rect 7742 6060 7748 6072
rect 7800 6060 7806 6112
rect 8386 6060 8392 6112
rect 8444 6100 8450 6112
rect 10594 6100 10600 6112
rect 8444 6072 10600 6100
rect 8444 6060 8450 6072
rect 10594 6060 10600 6072
rect 10652 6060 10658 6112
rect 10686 6060 10692 6112
rect 10744 6100 10750 6112
rect 10888 6100 10916 6140
rect 10962 6128 10968 6180
rect 11020 6168 11026 6180
rect 12618 6168 12624 6180
rect 11020 6140 12434 6168
rect 12579 6140 12624 6168
rect 11020 6128 11026 6140
rect 12250 6100 12256 6112
rect 10744 6072 10789 6100
rect 10888 6072 12256 6100
rect 10744 6060 10750 6072
rect 12250 6060 12256 6072
rect 12308 6060 12314 6112
rect 12406 6100 12434 6140
rect 12618 6128 12624 6140
rect 12676 6128 12682 6180
rect 14734 6168 14740 6180
rect 13372 6140 14740 6168
rect 12802 6100 12808 6112
rect 12406 6072 12808 6100
rect 12802 6060 12808 6072
rect 12860 6100 12866 6112
rect 13372 6100 13400 6140
rect 14734 6128 14740 6140
rect 14792 6128 14798 6180
rect 14921 6171 14979 6177
rect 14921 6137 14933 6171
rect 14967 6168 14979 6171
rect 15470 6168 15476 6180
rect 14967 6140 15476 6168
rect 14967 6137 14979 6140
rect 14921 6131 14979 6137
rect 15470 6128 15476 6140
rect 15528 6128 15534 6180
rect 18506 6168 18512 6180
rect 15580 6140 18512 6168
rect 12860 6072 13400 6100
rect 12860 6060 12866 6072
rect 13814 6060 13820 6112
rect 13872 6100 13878 6112
rect 15580 6100 15608 6140
rect 18506 6128 18512 6140
rect 18564 6128 18570 6180
rect 18598 6128 18604 6180
rect 18656 6168 18662 6180
rect 22664 6168 22692 6276
rect 22922 6264 22928 6276
rect 22980 6264 22986 6316
rect 23106 6304 23112 6316
rect 23067 6276 23112 6304
rect 23106 6264 23112 6276
rect 23164 6264 23170 6316
rect 18656 6140 22692 6168
rect 18656 6128 18662 6140
rect 13872 6072 15608 6100
rect 13872 6060 13878 6072
rect 16022 6060 16028 6112
rect 16080 6100 16086 6112
rect 16117 6103 16175 6109
rect 16117 6100 16129 6103
rect 16080 6072 16129 6100
rect 16080 6060 16086 6072
rect 16117 6069 16129 6072
rect 16163 6069 16175 6103
rect 16117 6063 16175 6069
rect 16206 6060 16212 6112
rect 16264 6100 16270 6112
rect 16853 6103 16911 6109
rect 16853 6100 16865 6103
rect 16264 6072 16865 6100
rect 16264 6060 16270 6072
rect 16853 6069 16865 6072
rect 16899 6100 16911 6103
rect 19610 6100 19616 6112
rect 16899 6072 19616 6100
rect 16899 6069 16911 6072
rect 16853 6063 16911 6069
rect 19610 6060 19616 6072
rect 19668 6060 19674 6112
rect 1104 6010 23828 6032
rect 1104 5958 3790 6010
rect 3842 5958 3854 6010
rect 3906 5958 3918 6010
rect 3970 5958 3982 6010
rect 4034 5958 4046 6010
rect 4098 5958 9471 6010
rect 9523 5958 9535 6010
rect 9587 5958 9599 6010
rect 9651 5958 9663 6010
rect 9715 5958 9727 6010
rect 9779 5958 15152 6010
rect 15204 5958 15216 6010
rect 15268 5958 15280 6010
rect 15332 5958 15344 6010
rect 15396 5958 15408 6010
rect 15460 5958 20833 6010
rect 20885 5958 20897 6010
rect 20949 5958 20961 6010
rect 21013 5958 21025 6010
rect 21077 5958 21089 6010
rect 21141 5958 23828 6010
rect 1104 5936 23828 5958
rect 2038 5896 2044 5908
rect 1999 5868 2044 5896
rect 2038 5856 2044 5868
rect 2096 5856 2102 5908
rect 3694 5856 3700 5908
rect 3752 5896 3758 5908
rect 3973 5899 4031 5905
rect 3973 5896 3985 5899
rect 3752 5868 3985 5896
rect 3752 5856 3758 5868
rect 3973 5865 3985 5868
rect 4019 5865 4031 5899
rect 3973 5859 4031 5865
rect 4356 5868 6408 5896
rect 2317 5831 2375 5837
rect 2317 5797 2329 5831
rect 2363 5828 2375 5831
rect 3510 5828 3516 5840
rect 2363 5800 3516 5828
rect 2363 5797 2375 5800
rect 2317 5791 2375 5797
rect 3510 5788 3516 5800
rect 3568 5828 3574 5840
rect 4356 5828 4384 5868
rect 6270 5828 6276 5840
rect 3568 5800 4384 5828
rect 6231 5800 6276 5828
rect 3568 5788 3574 5800
rect 6270 5788 6276 5800
rect 6328 5788 6334 5840
rect 6380 5760 6408 5868
rect 6914 5856 6920 5908
rect 6972 5896 6978 5908
rect 9214 5896 9220 5908
rect 6972 5868 9220 5896
rect 6972 5856 6978 5868
rect 9214 5856 9220 5868
rect 9272 5896 9278 5908
rect 11698 5896 11704 5908
rect 9272 5868 11704 5896
rect 9272 5856 9278 5868
rect 11698 5856 11704 5868
rect 11756 5856 11762 5908
rect 12066 5856 12072 5908
rect 12124 5896 12130 5908
rect 12345 5899 12403 5905
rect 12345 5896 12357 5899
rect 12124 5868 12357 5896
rect 12124 5856 12130 5868
rect 12345 5865 12357 5868
rect 12391 5865 12403 5899
rect 16758 5896 16764 5908
rect 12345 5859 12403 5865
rect 13096 5868 16764 5896
rect 11241 5831 11299 5837
rect 11241 5828 11253 5831
rect 10428 5800 11253 5828
rect 7834 5760 7840 5772
rect 3252 5746 5658 5760
rect 3252 5732 5672 5746
rect 6380 5732 7052 5760
rect 1762 5652 1768 5704
rect 1820 5692 1826 5704
rect 1857 5695 1915 5701
rect 1857 5692 1869 5695
rect 1820 5664 1869 5692
rect 1820 5652 1826 5664
rect 1857 5661 1869 5664
rect 1903 5661 1915 5695
rect 1857 5655 1915 5661
rect 1946 5652 1952 5704
rect 2004 5692 2010 5704
rect 2041 5695 2099 5701
rect 2041 5692 2053 5695
rect 2004 5664 2053 5692
rect 2004 5652 2010 5664
rect 2041 5661 2053 5664
rect 2087 5661 2099 5695
rect 2041 5655 2099 5661
rect 2133 5695 2191 5701
rect 2133 5661 2145 5695
rect 2179 5692 2191 5695
rect 3145 5695 3203 5701
rect 3145 5692 3157 5695
rect 2179 5664 3157 5692
rect 2179 5661 2191 5664
rect 2133 5655 2191 5661
rect 3145 5661 3157 5664
rect 3191 5661 3203 5695
rect 3145 5655 3203 5661
rect 2148 5624 2176 5655
rect 2866 5624 2872 5636
rect 1872 5596 2176 5624
rect 2827 5596 2872 5624
rect 1872 5568 1900 5596
rect 2866 5584 2872 5596
rect 2924 5624 2930 5636
rect 3252 5624 3280 5732
rect 3329 5695 3387 5701
rect 3329 5661 3341 5695
rect 3375 5692 3387 5695
rect 4798 5692 4804 5704
rect 3375 5664 4804 5692
rect 3375 5661 3387 5664
rect 3329 5655 3387 5661
rect 4798 5652 4804 5664
rect 4856 5652 4862 5704
rect 5074 5692 5080 5704
rect 5035 5664 5080 5692
rect 5074 5652 5080 5664
rect 5132 5652 5138 5704
rect 5258 5692 5264 5704
rect 5219 5664 5264 5692
rect 5258 5652 5264 5664
rect 5316 5652 5322 5704
rect 2924 5596 3280 5624
rect 4157 5627 4215 5633
rect 2924 5584 2930 5596
rect 4157 5593 4169 5627
rect 4203 5593 4215 5627
rect 4157 5587 4215 5593
rect 4341 5627 4399 5633
rect 4341 5593 4353 5627
rect 4387 5624 4399 5627
rect 4982 5624 4988 5636
rect 4387 5596 4988 5624
rect 4387 5593 4399 5596
rect 4341 5587 4399 5593
rect 1854 5516 1860 5568
rect 1912 5516 1918 5568
rect 2958 5556 2964 5568
rect 2919 5528 2964 5556
rect 2958 5516 2964 5528
rect 3016 5516 3022 5568
rect 4172 5556 4200 5587
rect 4982 5584 4988 5596
rect 5040 5584 5046 5636
rect 4246 5556 4252 5568
rect 4159 5528 4252 5556
rect 4246 5516 4252 5528
rect 4304 5556 4310 5568
rect 4890 5556 4896 5568
rect 4304 5528 4896 5556
rect 4304 5516 4310 5528
rect 4890 5516 4896 5528
rect 4948 5516 4954 5568
rect 5644 5556 5672 5732
rect 6089 5695 6147 5701
rect 6089 5661 6101 5695
rect 6135 5692 6147 5695
rect 6546 5692 6552 5704
rect 6135 5664 6552 5692
rect 6135 5661 6147 5664
rect 6089 5655 6147 5661
rect 6546 5652 6552 5664
rect 6604 5652 6610 5704
rect 7024 5701 7052 5732
rect 7208 5732 7840 5760
rect 7208 5701 7236 5732
rect 7834 5720 7840 5732
rect 7892 5720 7898 5772
rect 8021 5763 8079 5769
rect 8021 5729 8033 5763
rect 8067 5760 8079 5763
rect 8754 5760 8760 5772
rect 8067 5732 8760 5760
rect 8067 5729 8079 5732
rect 8021 5723 8079 5729
rect 8754 5720 8760 5732
rect 8812 5720 8818 5772
rect 7009 5695 7067 5701
rect 7009 5661 7021 5695
rect 7055 5661 7067 5695
rect 7009 5655 7067 5661
rect 7193 5695 7251 5701
rect 7193 5661 7205 5695
rect 7239 5661 7251 5695
rect 7742 5692 7748 5704
rect 7703 5664 7748 5692
rect 7193 5655 7251 5661
rect 7742 5652 7748 5664
rect 7800 5652 7806 5704
rect 7926 5692 7932 5704
rect 7887 5664 7932 5692
rect 7926 5652 7932 5664
rect 7984 5652 7990 5704
rect 8110 5692 8116 5704
rect 8071 5664 8116 5692
rect 8110 5652 8116 5664
rect 8168 5652 8174 5704
rect 8297 5695 8355 5701
rect 8297 5661 8309 5695
rect 8343 5692 8355 5695
rect 8662 5692 8668 5704
rect 8343 5664 8668 5692
rect 8343 5661 8355 5664
rect 8297 5655 8355 5661
rect 8662 5652 8668 5664
rect 8720 5652 8726 5704
rect 10134 5692 10140 5704
rect 10095 5664 10140 5692
rect 10134 5652 10140 5664
rect 10192 5652 10198 5704
rect 10226 5652 10232 5704
rect 10284 5692 10290 5704
rect 10428 5701 10456 5800
rect 11241 5797 11253 5800
rect 11287 5828 11299 5831
rect 11422 5828 11428 5840
rect 11287 5800 11428 5828
rect 11287 5797 11299 5800
rect 11241 5791 11299 5797
rect 11422 5788 11428 5800
rect 11480 5788 11486 5840
rect 11606 5788 11612 5840
rect 11664 5828 11670 5840
rect 12805 5831 12863 5837
rect 12805 5828 12817 5831
rect 11664 5800 12817 5828
rect 11664 5788 11670 5800
rect 12805 5797 12817 5800
rect 12851 5797 12863 5831
rect 12805 5791 12863 5797
rect 13096 5769 13124 5868
rect 16758 5856 16764 5868
rect 16816 5856 16822 5908
rect 18414 5896 18420 5908
rect 18375 5868 18420 5896
rect 18414 5856 18420 5868
rect 18472 5856 18478 5908
rect 18601 5899 18659 5905
rect 18601 5865 18613 5899
rect 18647 5865 18659 5899
rect 18601 5859 18659 5865
rect 14458 5788 14464 5840
rect 14516 5828 14522 5840
rect 14645 5831 14703 5837
rect 14645 5828 14657 5831
rect 14516 5800 14657 5828
rect 14516 5788 14522 5800
rect 14645 5797 14657 5800
rect 14691 5797 14703 5831
rect 14645 5791 14703 5797
rect 14734 5788 14740 5840
rect 14792 5828 14798 5840
rect 15197 5831 15255 5837
rect 15197 5828 15209 5831
rect 14792 5800 15209 5828
rect 14792 5788 14798 5800
rect 15197 5797 15209 5800
rect 15243 5797 15255 5831
rect 15197 5791 15255 5797
rect 15470 5788 15476 5840
rect 15528 5828 15534 5840
rect 15528 5800 17264 5828
rect 15528 5788 15534 5800
rect 10689 5763 10747 5769
rect 10689 5729 10701 5763
rect 10735 5760 10747 5763
rect 12989 5763 13047 5769
rect 12989 5760 13001 5763
rect 10735 5732 13001 5760
rect 10735 5729 10747 5732
rect 10689 5723 10747 5729
rect 12989 5729 13001 5732
rect 13035 5729 13047 5763
rect 12989 5723 13047 5729
rect 13081 5763 13139 5769
rect 13081 5729 13093 5763
rect 13127 5729 13139 5763
rect 13081 5723 13139 5729
rect 13906 5720 13912 5772
rect 13964 5760 13970 5772
rect 15841 5763 15899 5769
rect 15841 5760 15853 5763
rect 13964 5732 15853 5760
rect 13964 5720 13970 5732
rect 10413 5695 10471 5701
rect 10284 5664 10329 5692
rect 10284 5652 10290 5664
rect 10413 5661 10425 5695
rect 10459 5661 10471 5695
rect 10413 5655 10471 5661
rect 10502 5652 10508 5704
rect 10560 5692 10566 5704
rect 10560 5664 10605 5692
rect 10560 5652 10566 5664
rect 10778 5652 10784 5704
rect 10836 5692 10842 5704
rect 11701 5695 11759 5701
rect 11701 5692 11713 5695
rect 10836 5664 11713 5692
rect 10836 5652 10842 5664
rect 11701 5661 11713 5664
rect 11747 5661 11759 5695
rect 11885 5695 11943 5701
rect 11885 5690 11897 5695
rect 11701 5655 11759 5661
rect 11808 5662 11897 5690
rect 7101 5627 7159 5633
rect 7101 5593 7113 5627
rect 7147 5624 7159 5627
rect 11606 5624 11612 5636
rect 7147 5596 11612 5624
rect 7147 5593 7159 5596
rect 7101 5587 7159 5593
rect 11606 5584 11612 5596
rect 11664 5584 11670 5636
rect 7006 5556 7012 5568
rect 5644 5528 7012 5556
rect 7006 5516 7012 5528
rect 7064 5516 7070 5568
rect 8478 5556 8484 5568
rect 8439 5528 8484 5556
rect 8478 5516 8484 5528
rect 8536 5516 8542 5568
rect 10686 5516 10692 5568
rect 10744 5556 10750 5568
rect 11808 5556 11836 5662
rect 11885 5661 11897 5662
rect 11931 5661 11943 5695
rect 11885 5655 11943 5661
rect 11977 5695 12035 5701
rect 11977 5661 11989 5695
rect 12023 5661 12035 5695
rect 11977 5655 12035 5661
rect 12069 5695 12127 5701
rect 12069 5661 12081 5695
rect 12115 5661 12127 5695
rect 12069 5655 12127 5661
rect 11992 5568 12020 5655
rect 12084 5624 12112 5655
rect 12342 5652 12348 5704
rect 12400 5692 12406 5704
rect 14476 5701 14504 5732
rect 15841 5729 15853 5732
rect 15887 5729 15899 5763
rect 15841 5723 15899 5729
rect 15930 5720 15936 5772
rect 15988 5760 15994 5772
rect 17236 5769 17264 5800
rect 17862 5788 17868 5840
rect 17920 5828 17926 5840
rect 18616 5828 18644 5859
rect 18782 5856 18788 5908
rect 18840 5896 18846 5908
rect 20346 5896 20352 5908
rect 18840 5868 20352 5896
rect 18840 5856 18846 5868
rect 20346 5856 20352 5868
rect 20404 5856 20410 5908
rect 21634 5896 21640 5908
rect 21595 5868 21640 5896
rect 21634 5856 21640 5868
rect 21692 5856 21698 5908
rect 22370 5856 22376 5908
rect 22428 5896 22434 5908
rect 22557 5899 22615 5905
rect 22557 5896 22569 5899
rect 22428 5868 22569 5896
rect 22428 5856 22434 5868
rect 22557 5865 22569 5868
rect 22603 5865 22615 5899
rect 22557 5859 22615 5865
rect 17920 5800 18644 5828
rect 17920 5788 17926 5800
rect 19242 5788 19248 5840
rect 19300 5828 19306 5840
rect 19889 5831 19947 5837
rect 19889 5828 19901 5831
rect 19300 5800 19901 5828
rect 19300 5788 19306 5800
rect 19889 5797 19901 5800
rect 19935 5797 19947 5831
rect 19889 5791 19947 5797
rect 21174 5788 21180 5840
rect 21232 5828 21238 5840
rect 21232 5800 22324 5828
rect 21232 5788 21238 5800
rect 16761 5763 16819 5769
rect 16761 5760 16773 5763
rect 15988 5732 16773 5760
rect 15988 5720 15994 5732
rect 16761 5729 16773 5732
rect 16807 5729 16819 5763
rect 16761 5723 16819 5729
rect 17221 5763 17279 5769
rect 17221 5729 17233 5763
rect 17267 5760 17279 5763
rect 17678 5760 17684 5772
rect 17267 5732 17684 5760
rect 17267 5729 17279 5732
rect 17221 5723 17279 5729
rect 17678 5720 17684 5732
rect 17736 5720 17742 5772
rect 17957 5763 18015 5769
rect 17957 5729 17969 5763
rect 18003 5760 18015 5763
rect 18322 5760 18328 5772
rect 18003 5732 18328 5760
rect 18003 5729 18015 5732
rect 17957 5723 18015 5729
rect 18322 5720 18328 5732
rect 18380 5720 18386 5772
rect 18506 5720 18512 5772
rect 18564 5760 18570 5772
rect 20533 5763 20591 5769
rect 18564 5732 20116 5760
rect 18564 5720 18570 5732
rect 13173 5695 13231 5701
rect 13173 5692 13185 5695
rect 12400 5664 13185 5692
rect 12400 5652 12406 5664
rect 13173 5661 13185 5664
rect 13219 5661 13231 5695
rect 13173 5655 13231 5661
rect 13265 5695 13323 5701
rect 13265 5661 13277 5695
rect 13311 5692 13323 5695
rect 14277 5695 14335 5701
rect 14277 5692 14289 5695
rect 13311 5664 14289 5692
rect 13311 5661 13323 5664
rect 13265 5655 13323 5661
rect 14277 5661 14289 5664
rect 14323 5661 14335 5695
rect 14277 5655 14335 5661
rect 14461 5695 14519 5701
rect 14461 5661 14473 5695
rect 14507 5661 14519 5695
rect 14461 5655 14519 5661
rect 14737 5695 14795 5701
rect 14737 5661 14749 5695
rect 14783 5661 14795 5695
rect 14737 5655 14795 5661
rect 12250 5624 12256 5636
rect 12084 5596 12256 5624
rect 12250 5584 12256 5596
rect 12308 5624 12314 5636
rect 12308 5596 12940 5624
rect 12308 5584 12314 5596
rect 10744 5528 11836 5556
rect 10744 5516 10750 5528
rect 11974 5516 11980 5568
rect 12032 5516 12038 5568
rect 12912 5556 12940 5596
rect 12986 5584 12992 5636
rect 13044 5624 13050 5636
rect 13188 5624 13216 5655
rect 13044 5596 13216 5624
rect 13044 5584 13050 5596
rect 13078 5556 13084 5568
rect 12912 5528 13084 5556
rect 13078 5516 13084 5528
rect 13136 5516 13142 5568
rect 13188 5556 13216 5596
rect 14182 5584 14188 5636
rect 14240 5624 14246 5636
rect 14642 5624 14648 5636
rect 14240 5596 14648 5624
rect 14240 5584 14246 5596
rect 14642 5584 14648 5596
rect 14700 5624 14706 5636
rect 14752 5624 14780 5655
rect 14826 5652 14832 5704
rect 14884 5692 14890 5704
rect 15197 5695 15255 5701
rect 15197 5692 15209 5695
rect 14884 5664 15209 5692
rect 14884 5652 14890 5664
rect 15197 5661 15209 5664
rect 15243 5661 15255 5695
rect 15197 5655 15255 5661
rect 15381 5695 15439 5701
rect 15381 5661 15393 5695
rect 15427 5692 15439 5695
rect 15746 5692 15752 5704
rect 15427 5664 15752 5692
rect 15427 5661 15439 5664
rect 15381 5655 15439 5661
rect 15746 5652 15752 5664
rect 15804 5652 15810 5704
rect 16022 5692 16028 5704
rect 15983 5664 16028 5692
rect 16022 5652 16028 5664
rect 16080 5652 16086 5704
rect 16206 5692 16212 5704
rect 16167 5664 16212 5692
rect 16206 5652 16212 5664
rect 16264 5652 16270 5704
rect 16945 5695 17003 5701
rect 16945 5661 16957 5695
rect 16991 5661 17003 5695
rect 17310 5692 17316 5704
rect 17223 5664 17316 5692
rect 16945 5655 17003 5661
rect 14700 5596 14780 5624
rect 14700 5584 14706 5596
rect 15286 5584 15292 5636
rect 15344 5624 15350 5636
rect 16960 5624 16988 5655
rect 17310 5652 17316 5664
rect 17368 5692 17374 5704
rect 17862 5692 17868 5704
rect 17368 5664 17868 5692
rect 17368 5652 17374 5664
rect 17862 5652 17868 5664
rect 17920 5652 17926 5704
rect 18340 5692 18368 5720
rect 20088 5701 20116 5732
rect 20533 5729 20545 5763
rect 20579 5760 20591 5763
rect 20622 5760 20628 5772
rect 20579 5732 20628 5760
rect 20579 5729 20591 5732
rect 20533 5723 20591 5729
rect 20622 5720 20628 5732
rect 20680 5760 20686 5772
rect 22186 5760 22192 5772
rect 20680 5732 21036 5760
rect 20680 5720 20686 5732
rect 19797 5695 19855 5701
rect 19797 5692 19809 5695
rect 18340 5664 19809 5692
rect 19797 5661 19809 5664
rect 19843 5661 19855 5695
rect 19797 5655 19855 5661
rect 20073 5695 20131 5701
rect 20073 5661 20085 5695
rect 20119 5692 20131 5695
rect 20438 5692 20444 5704
rect 20119 5664 20444 5692
rect 20119 5661 20131 5664
rect 20073 5655 20131 5661
rect 20438 5652 20444 5664
rect 20496 5652 20502 5704
rect 21008 5701 21036 5732
rect 21192 5732 22192 5760
rect 21192 5701 21220 5732
rect 22186 5720 22192 5732
rect 22244 5720 22250 5772
rect 20993 5695 21051 5701
rect 20993 5661 21005 5695
rect 21039 5661 21051 5695
rect 20993 5655 21051 5661
rect 21177 5695 21235 5701
rect 21177 5661 21189 5695
rect 21223 5661 21235 5695
rect 21177 5655 21235 5661
rect 21266 5652 21272 5704
rect 21324 5692 21330 5704
rect 21450 5701 21456 5704
rect 21407 5695 21456 5701
rect 21324 5664 21369 5692
rect 21324 5652 21330 5664
rect 21407 5661 21419 5695
rect 21453 5661 21456 5695
rect 21407 5655 21456 5661
rect 21450 5652 21456 5655
rect 21508 5652 21514 5704
rect 22296 5692 22324 5800
rect 22922 5760 22928 5772
rect 22883 5732 22928 5760
rect 22922 5720 22928 5732
rect 22980 5720 22986 5772
rect 22741 5695 22799 5701
rect 22741 5692 22753 5695
rect 22296 5664 22753 5692
rect 22741 5661 22753 5664
rect 22787 5692 22799 5695
rect 23106 5692 23112 5704
rect 22787 5664 23112 5692
rect 22787 5661 22799 5664
rect 22741 5655 22799 5661
rect 23106 5652 23112 5664
rect 23164 5652 23170 5704
rect 17402 5624 17408 5636
rect 15344 5596 17408 5624
rect 15344 5584 15350 5596
rect 17402 5584 17408 5596
rect 17460 5584 17466 5636
rect 17512 5596 18736 5624
rect 17512 5556 17540 5596
rect 13188 5528 17540 5556
rect 17586 5516 17592 5568
rect 17644 5556 17650 5568
rect 18575 5559 18633 5565
rect 18575 5556 18587 5559
rect 17644 5528 18587 5556
rect 17644 5516 17650 5528
rect 18575 5525 18587 5528
rect 18621 5525 18633 5559
rect 18708 5556 18736 5596
rect 18782 5584 18788 5636
rect 18840 5624 18846 5636
rect 18840 5596 18885 5624
rect 18840 5584 18846 5596
rect 19426 5556 19432 5568
rect 18708 5528 19432 5556
rect 18575 5519 18633 5525
rect 19426 5516 19432 5528
rect 19484 5516 19490 5568
rect 20346 5516 20352 5568
rect 20404 5556 20410 5568
rect 22370 5556 22376 5568
rect 20404 5528 22376 5556
rect 20404 5516 20410 5528
rect 22370 5516 22376 5528
rect 22428 5516 22434 5568
rect 1104 5466 23987 5488
rect 1104 5414 6630 5466
rect 6682 5414 6694 5466
rect 6746 5414 6758 5466
rect 6810 5414 6822 5466
rect 6874 5414 6886 5466
rect 6938 5414 12311 5466
rect 12363 5414 12375 5466
rect 12427 5414 12439 5466
rect 12491 5414 12503 5466
rect 12555 5414 12567 5466
rect 12619 5414 17992 5466
rect 18044 5414 18056 5466
rect 18108 5414 18120 5466
rect 18172 5414 18184 5466
rect 18236 5414 18248 5466
rect 18300 5414 23673 5466
rect 23725 5414 23737 5466
rect 23789 5414 23801 5466
rect 23853 5414 23865 5466
rect 23917 5414 23929 5466
rect 23981 5414 23987 5466
rect 1104 5392 23987 5414
rect 2501 5355 2559 5361
rect 2501 5321 2513 5355
rect 2547 5352 2559 5355
rect 2958 5352 2964 5364
rect 2547 5324 2964 5352
rect 2547 5321 2559 5324
rect 2501 5315 2559 5321
rect 2958 5312 2964 5324
rect 3016 5312 3022 5364
rect 3234 5312 3240 5364
rect 3292 5352 3298 5364
rect 5810 5352 5816 5364
rect 3292 5324 4384 5352
rect 5771 5324 5816 5352
rect 3292 5312 3298 5324
rect 4246 5284 4252 5296
rect 1964 5256 4252 5284
rect 1964 5225 1992 5256
rect 4246 5244 4252 5256
rect 4304 5244 4310 5296
rect 4356 5293 4384 5324
rect 5810 5312 5816 5324
rect 5868 5312 5874 5364
rect 6825 5355 6883 5361
rect 6825 5321 6837 5355
rect 6871 5352 6883 5355
rect 7374 5352 7380 5364
rect 6871 5324 7380 5352
rect 6871 5321 6883 5324
rect 6825 5315 6883 5321
rect 7374 5312 7380 5324
rect 7432 5312 7438 5364
rect 11606 5312 11612 5364
rect 11664 5352 11670 5364
rect 12526 5352 12532 5364
rect 11664 5324 12532 5352
rect 11664 5312 11670 5324
rect 12526 5312 12532 5324
rect 12584 5312 12590 5364
rect 13170 5312 13176 5364
rect 13228 5352 13234 5364
rect 14366 5352 14372 5364
rect 13228 5324 14372 5352
rect 13228 5312 13234 5324
rect 14366 5312 14372 5324
rect 14424 5352 14430 5364
rect 14737 5355 14795 5361
rect 14737 5352 14749 5355
rect 14424 5324 14749 5352
rect 14424 5312 14430 5324
rect 14737 5321 14749 5324
rect 14783 5352 14795 5355
rect 15657 5355 15715 5361
rect 14783 5324 15608 5352
rect 14783 5321 14795 5324
rect 14737 5315 14795 5321
rect 4341 5287 4399 5293
rect 4341 5253 4353 5287
rect 4387 5253 4399 5287
rect 4341 5247 4399 5253
rect 6362 5244 6368 5296
rect 6420 5284 6426 5296
rect 12437 5287 12495 5293
rect 6420 5256 7972 5284
rect 6420 5244 6426 5256
rect 1949 5219 2007 5225
rect 1949 5185 1961 5219
rect 1995 5185 2007 5219
rect 1949 5179 2007 5185
rect 2041 5219 2099 5225
rect 2041 5185 2053 5219
rect 2087 5185 2099 5219
rect 2041 5179 2099 5185
rect 1762 5108 1768 5160
rect 1820 5148 1826 5160
rect 2056 5148 2084 5179
rect 2130 5176 2136 5228
rect 2188 5216 2194 5228
rect 2225 5219 2283 5225
rect 2225 5216 2237 5219
rect 2188 5188 2237 5216
rect 2188 5176 2194 5188
rect 2225 5185 2237 5188
rect 2271 5185 2283 5219
rect 2225 5179 2283 5185
rect 1820 5120 2084 5148
rect 1820 5108 1826 5120
rect 2240 5080 2268 5179
rect 2314 5176 2320 5228
rect 2372 5216 2378 5228
rect 3421 5219 3479 5225
rect 2372 5188 2417 5216
rect 2372 5176 2378 5188
rect 3421 5185 3433 5219
rect 3467 5216 3479 5219
rect 3602 5216 3608 5228
rect 3467 5188 3608 5216
rect 3467 5185 3479 5188
rect 3421 5179 3479 5185
rect 3602 5176 3608 5188
rect 3660 5176 3666 5228
rect 5721 5219 5779 5225
rect 5721 5185 5733 5219
rect 5767 5216 5779 5219
rect 6549 5219 6607 5225
rect 6549 5216 6561 5219
rect 5767 5188 6561 5216
rect 5767 5185 5779 5188
rect 5721 5179 5779 5185
rect 6549 5185 6561 5188
rect 6595 5216 6607 5219
rect 6638 5216 6644 5228
rect 6595 5188 6644 5216
rect 6595 5185 6607 5188
rect 6549 5179 6607 5185
rect 3142 5148 3148 5160
rect 3103 5120 3148 5148
rect 3142 5108 3148 5120
rect 3200 5108 3206 5160
rect 4246 5108 4252 5160
rect 4304 5148 4310 5160
rect 5077 5151 5135 5157
rect 5077 5148 5089 5151
rect 4304 5120 5089 5148
rect 4304 5108 4310 5120
rect 5077 5117 5089 5120
rect 5123 5148 5135 5151
rect 5258 5148 5264 5160
rect 5123 5120 5264 5148
rect 5123 5117 5135 5120
rect 5077 5111 5135 5117
rect 5258 5108 5264 5120
rect 5316 5148 5322 5160
rect 5736 5148 5764 5179
rect 6638 5176 6644 5188
rect 6696 5176 6702 5228
rect 6730 5176 6736 5228
rect 6788 5216 6794 5228
rect 6788 5188 6833 5216
rect 6788 5176 6794 5188
rect 7006 5176 7012 5228
rect 7064 5216 7070 5228
rect 7653 5219 7711 5225
rect 7653 5216 7665 5219
rect 7064 5188 7665 5216
rect 7064 5176 7070 5188
rect 7653 5185 7665 5188
rect 7699 5216 7711 5219
rect 7742 5216 7748 5228
rect 7699 5188 7748 5216
rect 7699 5185 7711 5188
rect 7653 5179 7711 5185
rect 7742 5176 7748 5188
rect 7800 5176 7806 5228
rect 7944 5225 7972 5256
rect 12437 5253 12449 5287
rect 12483 5284 12495 5287
rect 13633 5287 13691 5293
rect 12483 5256 13584 5284
rect 12483 5253 12495 5256
rect 12437 5247 12495 5253
rect 7929 5219 7987 5225
rect 7929 5185 7941 5219
rect 7975 5185 7987 5219
rect 8570 5216 8576 5228
rect 8531 5188 8576 5216
rect 7929 5179 7987 5185
rect 8570 5176 8576 5188
rect 8628 5176 8634 5228
rect 11054 5176 11060 5228
rect 11112 5216 11118 5228
rect 13354 5216 13360 5228
rect 11112 5188 13360 5216
rect 11112 5176 11118 5188
rect 13354 5176 13360 5188
rect 13412 5176 13418 5228
rect 13556 5216 13584 5256
rect 13633 5253 13645 5287
rect 13679 5284 13691 5287
rect 14090 5284 14096 5296
rect 13679 5256 14096 5284
rect 13679 5253 13691 5256
rect 13633 5247 13691 5253
rect 14090 5244 14096 5256
rect 14148 5244 14154 5296
rect 14642 5284 14648 5296
rect 14603 5256 14648 5284
rect 14642 5244 14648 5256
rect 14700 5244 14706 5296
rect 14826 5244 14832 5296
rect 14884 5284 14890 5296
rect 15105 5287 15163 5293
rect 14884 5256 15056 5284
rect 14884 5244 14890 5256
rect 14274 5216 14280 5228
rect 13556 5188 14280 5216
rect 14274 5176 14280 5188
rect 14332 5176 14338 5228
rect 14921 5219 14979 5225
rect 14921 5185 14933 5219
rect 14967 5216 14979 5219
rect 15028 5216 15056 5256
rect 15105 5253 15117 5287
rect 15151 5284 15163 5287
rect 15286 5284 15292 5296
rect 15151 5256 15292 5284
rect 15151 5253 15163 5256
rect 15105 5247 15163 5253
rect 15286 5244 15292 5256
rect 15344 5244 15350 5296
rect 15580 5284 15608 5324
rect 15657 5321 15669 5355
rect 15703 5352 15715 5355
rect 16114 5352 16120 5364
rect 15703 5324 16120 5352
rect 15703 5321 15715 5324
rect 15657 5315 15715 5321
rect 16114 5312 16120 5324
rect 16172 5312 16178 5364
rect 16206 5312 16212 5364
rect 16264 5312 16270 5364
rect 17678 5312 17684 5364
rect 17736 5352 17742 5364
rect 18782 5352 18788 5364
rect 17736 5324 18788 5352
rect 17736 5312 17742 5324
rect 18782 5312 18788 5324
rect 18840 5312 18846 5364
rect 21358 5352 21364 5364
rect 21319 5324 21364 5352
rect 21358 5312 21364 5324
rect 21416 5312 21422 5364
rect 22094 5312 22100 5364
rect 22152 5352 22158 5364
rect 22152 5324 22197 5352
rect 22152 5312 22158 5324
rect 16224 5284 16252 5312
rect 15580 5256 16252 5284
rect 16301 5287 16359 5293
rect 16301 5253 16313 5287
rect 16347 5284 16359 5287
rect 18506 5284 18512 5296
rect 16347 5256 18512 5284
rect 16347 5253 16359 5256
rect 16301 5247 16359 5253
rect 18506 5244 18512 5256
rect 18564 5244 18570 5296
rect 19518 5284 19524 5296
rect 19479 5256 19524 5284
rect 19518 5244 19524 5256
rect 19576 5244 19582 5296
rect 19610 5244 19616 5296
rect 19668 5284 19674 5296
rect 20717 5287 20775 5293
rect 20717 5284 20729 5287
rect 19668 5256 20729 5284
rect 19668 5244 19674 5256
rect 20717 5253 20729 5256
rect 20763 5253 20775 5287
rect 22554 5284 22560 5296
rect 22515 5256 22560 5284
rect 20717 5247 20775 5253
rect 22554 5244 22560 5256
rect 22612 5244 22618 5296
rect 22922 5284 22928 5296
rect 22756 5256 22928 5284
rect 15933 5219 15991 5225
rect 15933 5216 15945 5219
rect 14967 5188 15056 5216
rect 15672 5188 15945 5216
rect 14967 5185 14979 5188
rect 14921 5179 14979 5185
rect 5316 5120 5764 5148
rect 5316 5108 5322 5120
rect 6454 5108 6460 5160
rect 6512 5148 6518 5160
rect 9674 5148 9680 5160
rect 6512 5120 9076 5148
rect 9635 5120 9680 5148
rect 6512 5108 6518 5120
rect 4982 5080 4988 5092
rect 2240 5052 4988 5080
rect 4982 5040 4988 5052
rect 5040 5040 5046 5092
rect 8570 5080 8576 5092
rect 8531 5052 8576 5080
rect 8570 5040 8576 5052
rect 8628 5040 8634 5092
rect 9048 5080 9076 5120
rect 9674 5108 9680 5120
rect 9732 5108 9738 5160
rect 12066 5108 12072 5160
rect 12124 5148 12130 5160
rect 15672 5148 15700 5188
rect 15933 5185 15945 5188
rect 15979 5185 15991 5219
rect 15933 5179 15991 5185
rect 16209 5219 16267 5225
rect 16209 5185 16221 5219
rect 16255 5216 16267 5219
rect 16850 5216 16856 5228
rect 16255 5188 16856 5216
rect 16255 5185 16267 5188
rect 16209 5179 16267 5185
rect 12124 5120 15700 5148
rect 12124 5108 12130 5120
rect 15746 5108 15752 5160
rect 15804 5148 15810 5160
rect 15842 5151 15900 5157
rect 15842 5148 15854 5151
rect 15804 5120 15854 5148
rect 15804 5108 15810 5120
rect 15842 5117 15854 5120
rect 15888 5117 15900 5151
rect 15948 5148 15976 5179
rect 16850 5176 16856 5188
rect 16908 5176 16914 5228
rect 17402 5216 17408 5228
rect 17363 5188 17408 5216
rect 17402 5176 17408 5188
rect 17460 5176 17466 5228
rect 17773 5219 17831 5225
rect 17773 5185 17785 5219
rect 17819 5216 17831 5219
rect 17862 5216 17868 5228
rect 17819 5188 17868 5216
rect 17819 5185 17831 5188
rect 17773 5179 17831 5185
rect 17862 5176 17868 5188
rect 17920 5176 17926 5228
rect 19426 5216 19432 5228
rect 19387 5188 19432 5216
rect 19426 5176 19432 5188
rect 19484 5176 19490 5228
rect 22756 5225 22784 5256
rect 22922 5244 22928 5256
rect 22980 5244 22986 5296
rect 20533 5219 20591 5225
rect 20533 5216 20545 5219
rect 19628 5188 20545 5216
rect 17221 5151 17279 5157
rect 15948 5120 17172 5148
rect 15842 5111 15900 5117
rect 13722 5080 13728 5092
rect 9048 5052 13728 5080
rect 13722 5040 13728 5052
rect 13780 5040 13786 5092
rect 17144 5080 17172 5120
rect 17221 5117 17233 5151
rect 17267 5148 17279 5151
rect 17586 5148 17592 5160
rect 17267 5120 17592 5148
rect 17267 5117 17279 5120
rect 17221 5111 17279 5117
rect 17586 5108 17592 5120
rect 17644 5108 17650 5160
rect 17678 5108 17684 5160
rect 17736 5148 17742 5160
rect 18322 5148 18328 5160
rect 17736 5120 17781 5148
rect 18283 5120 18328 5148
rect 17736 5108 17742 5120
rect 18322 5108 18328 5120
rect 18380 5108 18386 5160
rect 18414 5108 18420 5160
rect 18472 5148 18478 5160
rect 19521 5151 19579 5157
rect 19521 5148 19533 5151
rect 18472 5120 19533 5148
rect 18472 5108 18478 5120
rect 19521 5117 19533 5120
rect 19567 5117 19579 5151
rect 19521 5111 19579 5117
rect 18874 5080 18880 5092
rect 14108 5052 17080 5080
rect 17144 5052 18880 5080
rect 3510 4972 3516 5024
rect 3568 5012 3574 5024
rect 9122 5012 9128 5024
rect 3568 4984 9128 5012
rect 3568 4972 3574 4984
rect 9122 4972 9128 4984
rect 9180 4972 9186 5024
rect 13081 5015 13139 5021
rect 13081 4981 13093 5015
rect 13127 5012 13139 5015
rect 14108 5012 14136 5052
rect 13127 4984 14136 5012
rect 14185 5015 14243 5021
rect 13127 4981 13139 4984
rect 13081 4975 13139 4981
rect 14185 4981 14197 5015
rect 14231 5012 14243 5015
rect 14458 5012 14464 5024
rect 14231 4984 14464 5012
rect 14231 4981 14243 4984
rect 14185 4975 14243 4981
rect 14458 4972 14464 4984
rect 14516 4972 14522 5024
rect 17052 5012 17080 5052
rect 18874 5040 18880 5052
rect 18932 5080 18938 5092
rect 19628 5080 19656 5188
rect 20533 5185 20545 5188
rect 20579 5185 20591 5219
rect 20533 5179 20591 5185
rect 22741 5219 22799 5225
rect 22741 5185 22753 5219
rect 22787 5185 22799 5219
rect 22741 5179 22799 5185
rect 22833 5219 22891 5225
rect 22833 5185 22845 5219
rect 22879 5216 22891 5219
rect 23106 5216 23112 5228
rect 22879 5188 23112 5216
rect 22879 5185 22891 5188
rect 22833 5179 22891 5185
rect 23106 5176 23112 5188
rect 23164 5176 23170 5228
rect 18932 5052 19656 5080
rect 19720 5052 20944 5080
rect 18932 5040 18938 5052
rect 18690 5012 18696 5024
rect 17052 4984 18696 5012
rect 18690 4972 18696 4984
rect 18748 4972 18754 5024
rect 19426 4972 19432 5024
rect 19484 5012 19490 5024
rect 19720 5012 19748 5052
rect 19484 4984 19748 5012
rect 19981 5015 20039 5021
rect 19484 4972 19490 4984
rect 19981 4981 19993 5015
rect 20027 5012 20039 5015
rect 20162 5012 20168 5024
rect 20027 4984 20168 5012
rect 20027 4981 20039 4984
rect 19981 4975 20039 4981
rect 20162 4972 20168 4984
rect 20220 4972 20226 5024
rect 20916 5021 20944 5052
rect 20901 5015 20959 5021
rect 20901 4981 20913 5015
rect 20947 4981 20959 5015
rect 20901 4975 20959 4981
rect 1104 4922 23828 4944
rect 1104 4870 3790 4922
rect 3842 4870 3854 4922
rect 3906 4870 3918 4922
rect 3970 4870 3982 4922
rect 4034 4870 4046 4922
rect 4098 4870 9471 4922
rect 9523 4870 9535 4922
rect 9587 4870 9599 4922
rect 9651 4870 9663 4922
rect 9715 4870 9727 4922
rect 9779 4870 15152 4922
rect 15204 4870 15216 4922
rect 15268 4870 15280 4922
rect 15332 4870 15344 4922
rect 15396 4870 15408 4922
rect 15460 4870 20833 4922
rect 20885 4870 20897 4922
rect 20949 4870 20961 4922
rect 21013 4870 21025 4922
rect 21077 4870 21089 4922
rect 21141 4870 23828 4922
rect 1104 4848 23828 4870
rect 1857 4811 1915 4817
rect 1857 4777 1869 4811
rect 1903 4808 1915 4811
rect 2222 4808 2228 4820
rect 1903 4780 2228 4808
rect 1903 4777 1915 4780
rect 1857 4771 1915 4777
rect 2222 4768 2228 4780
rect 2280 4768 2286 4820
rect 2685 4811 2743 4817
rect 2685 4777 2697 4811
rect 2731 4808 2743 4811
rect 2774 4808 2780 4820
rect 2731 4780 2780 4808
rect 2731 4777 2743 4780
rect 2685 4771 2743 4777
rect 2774 4768 2780 4780
rect 2832 4768 2838 4820
rect 7190 4768 7196 4820
rect 7248 4808 7254 4820
rect 9122 4808 9128 4820
rect 7248 4780 9128 4808
rect 7248 4768 7254 4780
rect 9122 4768 9128 4780
rect 9180 4768 9186 4820
rect 9585 4811 9643 4817
rect 9585 4777 9597 4811
rect 9631 4808 9643 4811
rect 10134 4808 10140 4820
rect 9631 4780 10140 4808
rect 9631 4777 9643 4780
rect 9585 4771 9643 4777
rect 10134 4768 10140 4780
rect 10192 4768 10198 4820
rect 10778 4768 10784 4820
rect 10836 4808 10842 4820
rect 11146 4808 11152 4820
rect 10836 4780 11152 4808
rect 10836 4768 10842 4780
rect 11146 4768 11152 4780
rect 11204 4808 11210 4820
rect 11241 4811 11299 4817
rect 11241 4808 11253 4811
rect 11204 4780 11253 4808
rect 11204 4768 11210 4780
rect 11241 4777 11253 4780
rect 11287 4777 11299 4811
rect 11241 4771 11299 4777
rect 12713 4811 12771 4817
rect 12713 4777 12725 4811
rect 12759 4808 12771 4811
rect 12894 4808 12900 4820
rect 12759 4780 12900 4808
rect 12759 4777 12771 4780
rect 12713 4771 12771 4777
rect 12894 4768 12900 4780
rect 12952 4768 12958 4820
rect 13078 4768 13084 4820
rect 13136 4808 13142 4820
rect 16206 4808 16212 4820
rect 13136 4780 16212 4808
rect 13136 4768 13142 4780
rect 16206 4768 16212 4780
rect 16264 4768 16270 4820
rect 16758 4768 16764 4820
rect 16816 4808 16822 4820
rect 16853 4811 16911 4817
rect 16853 4808 16865 4811
rect 16816 4780 16865 4808
rect 16816 4768 16822 4780
rect 16853 4777 16865 4780
rect 16899 4777 16911 4811
rect 16853 4771 16911 4777
rect 18690 4768 18696 4820
rect 18748 4808 18754 4820
rect 20530 4808 20536 4820
rect 18748 4780 20392 4808
rect 20491 4780 20536 4808
rect 18748 4768 18754 4780
rect 4338 4700 4344 4752
rect 4396 4740 4402 4752
rect 5258 4740 5264 4752
rect 4396 4712 5264 4740
rect 4396 4700 4402 4712
rect 5258 4700 5264 4712
rect 5316 4740 5322 4752
rect 6546 4740 6552 4752
rect 5316 4712 6552 4740
rect 5316 4700 5322 4712
rect 5810 4672 5816 4684
rect 4540 4644 5816 4672
rect 1762 4564 1768 4616
rect 1820 4604 1826 4616
rect 2314 4604 2320 4616
rect 1820 4576 2320 4604
rect 1820 4564 1826 4576
rect 2314 4564 2320 4576
rect 2372 4564 2378 4616
rect 2406 4564 2412 4616
rect 2464 4604 2470 4616
rect 2777 4607 2835 4613
rect 2777 4604 2789 4607
rect 2464 4576 2789 4604
rect 2464 4564 2470 4576
rect 2777 4573 2789 4576
rect 2823 4573 2835 4607
rect 2777 4567 2835 4573
rect 4154 4564 4160 4616
rect 4212 4604 4218 4616
rect 4540 4613 4568 4644
rect 5810 4632 5816 4644
rect 5868 4632 5874 4684
rect 4433 4607 4491 4613
rect 4433 4604 4445 4607
rect 4212 4576 4445 4604
rect 4212 4564 4218 4576
rect 4433 4573 4445 4576
rect 4479 4573 4491 4607
rect 4433 4567 4491 4573
rect 4525 4607 4583 4613
rect 4525 4573 4537 4607
rect 4571 4573 4583 4607
rect 4525 4567 4583 4573
rect 4985 4607 5043 4613
rect 4985 4573 4997 4607
rect 5031 4604 5043 4607
rect 5534 4604 5540 4616
rect 5031 4576 5540 4604
rect 5031 4573 5043 4576
rect 4985 4567 5043 4573
rect 5534 4564 5540 4576
rect 5592 4564 5598 4616
rect 5718 4604 5724 4616
rect 5679 4576 5724 4604
rect 5718 4564 5724 4576
rect 5776 4564 5782 4616
rect 5920 4613 5948 4712
rect 6546 4700 6552 4712
rect 6604 4740 6610 4752
rect 6730 4740 6736 4752
rect 6604 4712 6736 4740
rect 6604 4700 6610 4712
rect 6730 4700 6736 4712
rect 6788 4740 6794 4752
rect 10042 4740 10048 4752
rect 6788 4712 6960 4740
rect 10003 4712 10048 4740
rect 6788 4700 6794 4712
rect 6086 4632 6092 4684
rect 6144 4672 6150 4684
rect 6144 4644 6592 4672
rect 6144 4632 6150 4644
rect 6564 4613 6592 4644
rect 6638 4632 6644 4684
rect 6696 4672 6702 4684
rect 6825 4675 6883 4681
rect 6825 4672 6837 4675
rect 6696 4644 6837 4672
rect 6696 4632 6702 4644
rect 6825 4641 6837 4644
rect 6871 4641 6883 4675
rect 6825 4635 6883 4641
rect 6932 4613 6960 4712
rect 10042 4700 10048 4712
rect 10100 4700 10106 4752
rect 12268 4712 12434 4740
rect 7374 4632 7380 4684
rect 7432 4672 7438 4684
rect 7432 4644 8156 4672
rect 7432 4632 7438 4644
rect 5905 4607 5963 4613
rect 5905 4573 5917 4607
rect 5951 4573 5963 4607
rect 5905 4567 5963 4573
rect 6365 4607 6423 4613
rect 6365 4573 6377 4607
rect 6411 4573 6423 4607
rect 6365 4567 6423 4573
rect 6549 4607 6607 4613
rect 6549 4573 6561 4607
rect 6595 4573 6607 4607
rect 6549 4567 6607 4573
rect 6917 4607 6975 4613
rect 6917 4573 6929 4607
rect 6963 4573 6975 4607
rect 6917 4567 6975 4573
rect 4249 4539 4307 4545
rect 4249 4505 4261 4539
rect 4295 4536 4307 4539
rect 4338 4536 4344 4548
rect 4295 4508 4344 4536
rect 4295 4505 4307 4508
rect 4249 4499 4307 4505
rect 3418 4468 3424 4480
rect 3379 4440 3424 4468
rect 3418 4428 3424 4440
rect 3476 4428 3482 4480
rect 4154 4428 4160 4480
rect 4212 4468 4218 4480
rect 4264 4468 4292 4499
rect 4338 4496 4344 4508
rect 4396 4496 4402 4548
rect 4617 4539 4675 4545
rect 4617 4536 4629 4539
rect 4448 4508 4629 4536
rect 4448 4480 4476 4508
rect 4617 4505 4629 4508
rect 4663 4536 4675 4539
rect 5074 4536 5080 4548
rect 4663 4508 5080 4536
rect 4663 4505 4675 4508
rect 4617 4499 4675 4505
rect 5074 4496 5080 4508
rect 5132 4496 5138 4548
rect 5350 4496 5356 4548
rect 5408 4536 5414 4548
rect 6380 4536 6408 4567
rect 7926 4564 7932 4616
rect 7984 4604 7990 4616
rect 8021 4607 8079 4613
rect 8021 4604 8033 4607
rect 7984 4576 8033 4604
rect 7984 4564 7990 4576
rect 8021 4573 8033 4576
rect 8067 4573 8079 4607
rect 8128 4604 8156 4644
rect 8478 4632 8484 4684
rect 8536 4672 8542 4684
rect 9125 4675 9183 4681
rect 9125 4672 9137 4675
rect 8536 4644 9137 4672
rect 8536 4632 8542 4644
rect 9125 4641 9137 4644
rect 9171 4641 9183 4675
rect 9125 4635 9183 4641
rect 9217 4675 9275 4681
rect 9217 4641 9229 4675
rect 9263 4672 9275 4675
rect 9858 4672 9864 4684
rect 9263 4644 9864 4672
rect 9263 4641 9275 4644
rect 9217 4635 9275 4641
rect 9858 4632 9864 4644
rect 9916 4632 9922 4684
rect 10410 4632 10416 4684
rect 10468 4672 10474 4684
rect 10689 4675 10747 4681
rect 10689 4672 10701 4675
rect 10468 4644 10701 4672
rect 10468 4632 10474 4644
rect 10689 4641 10701 4644
rect 10735 4641 10747 4675
rect 10689 4635 10747 4641
rect 9401 4607 9459 4613
rect 9401 4604 9413 4607
rect 8128 4576 9413 4604
rect 8021 4567 8079 4573
rect 9401 4573 9413 4576
rect 9447 4573 9459 4607
rect 9401 4567 9459 4573
rect 10229 4607 10287 4613
rect 10229 4573 10241 4607
rect 10275 4573 10287 4607
rect 10229 4567 10287 4573
rect 7558 4536 7564 4548
rect 5408 4508 6408 4536
rect 7519 4508 7564 4536
rect 5408 4496 5414 4508
rect 7558 4496 7564 4508
rect 7616 4496 7622 4548
rect 10244 4536 10272 4567
rect 10318 4564 10324 4616
rect 10376 4604 10382 4616
rect 10597 4607 10655 4613
rect 10376 4576 10421 4604
rect 10376 4564 10382 4576
rect 10597 4573 10609 4607
rect 10643 4604 10655 4607
rect 11698 4604 11704 4616
rect 10643 4576 11704 4604
rect 10643 4573 10655 4576
rect 10597 4567 10655 4573
rect 11698 4564 11704 4576
rect 11756 4564 11762 4616
rect 12268 4613 12296 4712
rect 12406 4672 12434 4712
rect 12526 4700 12532 4752
rect 12584 4740 12590 4752
rect 20364 4740 20392 4780
rect 20530 4768 20536 4780
rect 20588 4768 20594 4820
rect 21085 4743 21143 4749
rect 21085 4740 21097 4743
rect 12584 4712 19748 4740
rect 20364 4712 21097 4740
rect 12584 4700 12590 4712
rect 13446 4672 13452 4684
rect 12406 4644 13452 4672
rect 13446 4632 13452 4644
rect 13504 4632 13510 4684
rect 13556 4644 16436 4672
rect 12253 4607 12311 4613
rect 12253 4573 12265 4607
rect 12299 4573 12311 4607
rect 12253 4567 12311 4573
rect 12526 4564 12532 4616
rect 12584 4604 12590 4616
rect 13354 4604 13360 4616
rect 12584 4576 12629 4604
rect 13315 4576 13360 4604
rect 12584 4564 12590 4576
rect 13354 4564 13360 4576
rect 13412 4564 13418 4616
rect 13556 4604 13584 4644
rect 13722 4604 13728 4616
rect 13464 4576 13584 4604
rect 13683 4576 13728 4604
rect 9324 4508 10272 4536
rect 9324 4480 9352 4508
rect 12066 4496 12072 4548
rect 12124 4536 12130 4548
rect 12345 4539 12403 4545
rect 12345 4536 12357 4539
rect 12124 4508 12357 4536
rect 12124 4496 12130 4508
rect 12345 4505 12357 4508
rect 12391 4505 12403 4539
rect 12345 4499 12403 4505
rect 12802 4496 12808 4548
rect 12860 4536 12866 4548
rect 13464 4545 13492 4576
rect 13722 4564 13728 4576
rect 13780 4564 13786 4616
rect 14366 4604 14372 4616
rect 14327 4576 14372 4604
rect 14366 4564 14372 4576
rect 14424 4564 14430 4616
rect 15473 4607 15531 4613
rect 15473 4573 15485 4607
rect 15519 4604 15531 4607
rect 16022 4604 16028 4616
rect 15519 4576 16028 4604
rect 15519 4573 15531 4576
rect 15473 4567 15531 4573
rect 16022 4564 16028 4576
rect 16080 4564 16086 4616
rect 16206 4604 16212 4616
rect 16167 4576 16212 4604
rect 16206 4564 16212 4576
rect 16264 4564 16270 4616
rect 16302 4607 16360 4613
rect 16302 4573 16314 4607
rect 16348 4573 16360 4607
rect 16302 4567 16360 4573
rect 13449 4539 13507 4545
rect 13449 4536 13461 4539
rect 12860 4508 13461 4536
rect 12860 4496 12866 4508
rect 13449 4505 13461 4508
rect 13495 4505 13507 4539
rect 13449 4499 13507 4505
rect 13538 4496 13544 4548
rect 13596 4536 13602 4548
rect 13740 4536 13768 4564
rect 15838 4536 15844 4548
rect 13596 4508 13641 4536
rect 13740 4508 15844 4536
rect 13596 4496 13602 4508
rect 15838 4496 15844 4508
rect 15896 4536 15902 4548
rect 16316 4536 16344 4567
rect 15896 4508 16344 4536
rect 16408 4536 16436 4644
rect 16482 4564 16488 4616
rect 16540 4604 16546 4616
rect 16715 4607 16773 4613
rect 16540 4576 16585 4604
rect 16540 4564 16546 4576
rect 16715 4573 16727 4607
rect 16761 4604 16773 4607
rect 17310 4604 17316 4616
rect 16761 4576 17316 4604
rect 16761 4573 16773 4576
rect 16715 4567 16773 4573
rect 17310 4564 17316 4576
rect 17368 4604 17374 4616
rect 17865 4607 17923 4613
rect 17865 4604 17877 4607
rect 17368 4576 17877 4604
rect 17368 4564 17374 4576
rect 17865 4573 17877 4576
rect 17911 4573 17923 4607
rect 19426 4604 19432 4616
rect 19387 4576 19432 4604
rect 17865 4567 17923 4573
rect 19426 4564 19432 4576
rect 19484 4564 19490 4616
rect 19720 4613 19748 4712
rect 21085 4709 21097 4712
rect 21131 4740 21143 4743
rect 21450 4740 21456 4752
rect 21131 4712 21456 4740
rect 21131 4709 21143 4712
rect 21085 4703 21143 4709
rect 21450 4700 21456 4712
rect 21508 4700 21514 4752
rect 22094 4632 22100 4684
rect 22152 4672 22158 4684
rect 22152 4644 22197 4672
rect 22152 4632 22158 4644
rect 22370 4632 22376 4684
rect 22428 4672 22434 4684
rect 22428 4644 22692 4672
rect 22428 4632 22434 4644
rect 19705 4607 19763 4613
rect 19705 4573 19717 4607
rect 19751 4573 19763 4607
rect 20438 4604 20444 4616
rect 19705 4567 19763 4573
rect 19812 4576 20444 4604
rect 16574 4536 16580 4548
rect 16408 4508 16580 4536
rect 15896 4496 15902 4508
rect 16574 4496 16580 4508
rect 16632 4496 16638 4548
rect 16942 4496 16948 4548
rect 17000 4536 17006 4548
rect 19521 4539 19579 4545
rect 19521 4536 19533 4539
rect 17000 4508 19533 4536
rect 17000 4496 17006 4508
rect 19521 4505 19533 4508
rect 19567 4505 19579 4539
rect 19521 4499 19579 4505
rect 4212 4440 4292 4468
rect 4212 4428 4218 4440
rect 4430 4428 4436 4480
rect 4488 4428 4494 4480
rect 5813 4471 5871 4477
rect 5813 4437 5825 4471
rect 5859 4468 5871 4471
rect 9306 4468 9312 4480
rect 5859 4440 9312 4468
rect 5859 4437 5871 4440
rect 5813 4431 5871 4437
rect 9306 4428 9312 4440
rect 9364 4428 9370 4480
rect 11974 4428 11980 4480
rect 12032 4468 12038 4480
rect 13173 4471 13231 4477
rect 13173 4468 13185 4471
rect 12032 4440 13185 4468
rect 12032 4428 12038 4440
rect 13173 4437 13185 4440
rect 13219 4437 13231 4471
rect 13173 4431 13231 4437
rect 14921 4471 14979 4477
rect 14921 4437 14933 4471
rect 14967 4468 14979 4471
rect 15746 4468 15752 4480
rect 14967 4440 15752 4468
rect 14967 4437 14979 4440
rect 14921 4431 14979 4437
rect 15746 4428 15752 4440
rect 15804 4468 15810 4480
rect 17405 4471 17463 4477
rect 17405 4468 17417 4471
rect 15804 4440 17417 4468
rect 15804 4428 15810 4440
rect 17405 4437 17417 4440
rect 17451 4468 17463 4471
rect 18598 4468 18604 4480
rect 17451 4440 18604 4468
rect 17451 4437 17463 4440
rect 17405 4431 17463 4437
rect 18598 4428 18604 4440
rect 18656 4428 18662 4480
rect 18877 4471 18935 4477
rect 18877 4437 18889 4471
rect 18923 4468 18935 4471
rect 19812 4468 19840 4576
rect 20438 4564 20444 4576
rect 20496 4564 20502 4616
rect 22664 4613 22692 4644
rect 22649 4607 22707 4613
rect 22649 4573 22661 4607
rect 22695 4573 22707 4607
rect 22649 4567 22707 4573
rect 23017 4607 23075 4613
rect 23017 4573 23029 4607
rect 23063 4604 23075 4607
rect 23106 4604 23112 4616
rect 23063 4576 23112 4604
rect 23063 4573 23075 4576
rect 23017 4567 23075 4573
rect 23106 4564 23112 4576
rect 23164 4564 23170 4616
rect 19889 4539 19947 4545
rect 19889 4505 19901 4539
rect 19935 4536 19947 4539
rect 20806 4536 20812 4548
rect 19935 4508 20812 4536
rect 19935 4505 19947 4508
rect 19889 4499 19947 4505
rect 20806 4496 20812 4508
rect 20864 4496 20870 4548
rect 18923 4440 19840 4468
rect 18923 4437 18935 4440
rect 18877 4431 18935 4437
rect 1104 4378 23987 4400
rect 1104 4326 6630 4378
rect 6682 4326 6694 4378
rect 6746 4326 6758 4378
rect 6810 4326 6822 4378
rect 6874 4326 6886 4378
rect 6938 4326 12311 4378
rect 12363 4326 12375 4378
rect 12427 4326 12439 4378
rect 12491 4326 12503 4378
rect 12555 4326 12567 4378
rect 12619 4326 17992 4378
rect 18044 4326 18056 4378
rect 18108 4326 18120 4378
rect 18172 4326 18184 4378
rect 18236 4326 18248 4378
rect 18300 4326 23673 4378
rect 23725 4326 23737 4378
rect 23789 4326 23801 4378
rect 23853 4326 23865 4378
rect 23917 4326 23929 4378
rect 23981 4326 23987 4378
rect 1104 4304 23987 4326
rect 6733 4267 6791 4273
rect 6733 4233 6745 4267
rect 6779 4264 6791 4267
rect 7006 4264 7012 4276
rect 6779 4236 7012 4264
rect 6779 4233 6791 4236
rect 6733 4227 6791 4233
rect 7006 4224 7012 4236
rect 7064 4224 7070 4276
rect 8478 4264 8484 4276
rect 8439 4236 8484 4264
rect 8478 4224 8484 4236
rect 8536 4224 8542 4276
rect 10318 4224 10324 4276
rect 10376 4264 10382 4276
rect 10873 4267 10931 4273
rect 10873 4264 10885 4267
rect 10376 4236 10885 4264
rect 10376 4224 10382 4236
rect 10873 4233 10885 4236
rect 10919 4233 10931 4267
rect 12066 4264 12072 4276
rect 11979 4236 12072 4264
rect 10873 4227 10931 4233
rect 12066 4224 12072 4236
rect 12124 4224 12130 4276
rect 14001 4267 14059 4273
rect 14001 4233 14013 4267
rect 14047 4264 14059 4267
rect 14366 4264 14372 4276
rect 14047 4236 14372 4264
rect 14047 4233 14059 4236
rect 14001 4227 14059 4233
rect 14366 4224 14372 4236
rect 14424 4224 14430 4276
rect 14550 4264 14556 4276
rect 14511 4236 14556 4264
rect 14550 4224 14556 4236
rect 14608 4224 14614 4276
rect 16022 4224 16028 4276
rect 16080 4264 16086 4276
rect 17957 4267 18015 4273
rect 17957 4264 17969 4267
rect 16080 4236 17969 4264
rect 16080 4224 16086 4236
rect 17957 4233 17969 4236
rect 18003 4264 18015 4267
rect 18322 4264 18328 4276
rect 18003 4236 18328 4264
rect 18003 4233 18015 4236
rect 17957 4227 18015 4233
rect 18322 4224 18328 4236
rect 18380 4224 18386 4276
rect 18506 4264 18512 4276
rect 18467 4236 18512 4264
rect 18506 4224 18512 4236
rect 18564 4224 18570 4276
rect 2314 4156 2320 4208
rect 2372 4196 2378 4208
rect 4430 4196 4436 4208
rect 2372 4168 4436 4196
rect 2372 4156 2378 4168
rect 4430 4156 4436 4168
rect 4488 4196 4494 4208
rect 5721 4199 5779 4205
rect 4488 4168 5396 4196
rect 4488 4156 4494 4168
rect 5368 4140 5396 4168
rect 5721 4165 5733 4199
rect 5767 4196 5779 4199
rect 6362 4196 6368 4208
rect 5767 4168 6368 4196
rect 5767 4165 5779 4168
rect 5721 4159 5779 4165
rect 6362 4156 6368 4168
rect 6420 4156 6426 4208
rect 6546 4156 6552 4208
rect 6604 4196 6610 4208
rect 6641 4199 6699 4205
rect 6641 4196 6653 4199
rect 6604 4168 6653 4196
rect 6604 4156 6610 4168
rect 6641 4165 6653 4168
rect 6687 4165 6699 4199
rect 6641 4159 6699 4165
rect 6748 4168 7420 4196
rect 1854 4128 1860 4140
rect 1815 4100 1860 4128
rect 1854 4088 1860 4100
rect 1912 4088 1918 4140
rect 2038 4088 2044 4140
rect 2096 4128 2102 4140
rect 2133 4131 2191 4137
rect 2133 4128 2145 4131
rect 2096 4100 2145 4128
rect 2096 4088 2102 4100
rect 2133 4097 2145 4100
rect 2179 4128 2191 4131
rect 2590 4128 2596 4140
rect 2179 4100 2596 4128
rect 2179 4097 2191 4100
rect 2133 4091 2191 4097
rect 2590 4088 2596 4100
rect 2648 4088 2654 4140
rect 2685 4131 2743 4137
rect 2685 4097 2697 4131
rect 2731 4128 2743 4131
rect 4246 4128 4252 4140
rect 2731 4100 4252 4128
rect 2731 4097 2743 4100
rect 2685 4091 2743 4097
rect 2700 4060 2728 4091
rect 4246 4088 4252 4100
rect 4304 4088 4310 4140
rect 4617 4131 4675 4137
rect 4617 4097 4629 4131
rect 4663 4097 4675 4131
rect 4617 4091 4675 4097
rect 2056 4032 2728 4060
rect 1946 3952 1952 4004
rect 2004 3992 2010 4004
rect 2056 4001 2084 4032
rect 3694 4020 3700 4072
rect 3752 4060 3758 4072
rect 4341 4063 4399 4069
rect 4341 4060 4353 4063
rect 3752 4032 4353 4060
rect 3752 4020 3758 4032
rect 4341 4029 4353 4032
rect 4387 4029 4399 4063
rect 4632 4060 4660 4091
rect 4890 4088 4896 4140
rect 4948 4128 4954 4140
rect 5169 4131 5227 4137
rect 5169 4128 5181 4131
rect 4948 4100 5181 4128
rect 4948 4088 4954 4100
rect 5169 4097 5181 4100
rect 5215 4097 5227 4131
rect 5169 4091 5227 4097
rect 5350 4088 5356 4140
rect 5408 4128 5414 4140
rect 6380 4128 6408 4156
rect 6748 4128 6776 4168
rect 7392 4137 7420 4168
rect 7558 4156 7564 4208
rect 7616 4196 7622 4208
rect 9030 4196 9036 4208
rect 7616 4168 9036 4196
rect 7616 4156 7622 4168
rect 9030 4156 9036 4168
rect 9088 4196 9094 4208
rect 12084 4196 12112 4224
rect 13814 4196 13820 4208
rect 9088 4168 12112 4196
rect 13096 4168 13820 4196
rect 9088 4156 9094 4168
rect 5408 4100 5501 4128
rect 6380 4100 6776 4128
rect 6825 4131 6883 4137
rect 5408 4088 5414 4100
rect 6825 4097 6837 4131
rect 6871 4097 6883 4131
rect 6825 4091 6883 4097
rect 7377 4131 7435 4137
rect 7377 4097 7389 4131
rect 7423 4097 7435 4131
rect 7377 4091 7435 4097
rect 5442 4060 5448 4072
rect 4632 4032 5448 4060
rect 4341 4023 4399 4029
rect 5442 4020 5448 4032
rect 5500 4020 5506 4072
rect 2041 3995 2099 4001
rect 2041 3992 2053 3995
rect 2004 3964 2053 3992
rect 2004 3952 2010 3964
rect 2041 3961 2053 3964
rect 2087 3961 2099 3995
rect 4154 3992 4160 4004
rect 2041 3955 2099 3961
rect 2700 3964 4160 3992
rect 1670 3924 1676 3936
rect 1631 3896 1676 3924
rect 1670 3884 1676 3896
rect 1728 3884 1734 3936
rect 1854 3884 1860 3936
rect 1912 3924 1918 3936
rect 2700 3924 2728 3964
rect 4154 3952 4160 3964
rect 4212 3952 4218 4004
rect 4982 3952 4988 4004
rect 5040 3992 5046 4004
rect 6840 3992 6868 4091
rect 8294 4088 8300 4140
rect 8352 4128 8358 4140
rect 8389 4131 8447 4137
rect 8389 4128 8401 4131
rect 8352 4100 8401 4128
rect 8352 4088 8358 4100
rect 8389 4097 8401 4100
rect 8435 4097 8447 4131
rect 8389 4091 8447 4097
rect 8573 4131 8631 4137
rect 8573 4097 8585 4131
rect 8619 4128 8631 4131
rect 8662 4128 8668 4140
rect 8619 4100 8668 4128
rect 8619 4097 8631 4100
rect 8573 4091 8631 4097
rect 8662 4088 8668 4100
rect 8720 4088 8726 4140
rect 10686 4128 10692 4140
rect 8864 4100 10692 4128
rect 7190 4060 7196 4072
rect 7151 4032 7196 4060
rect 7190 4020 7196 4032
rect 7248 4020 7254 4072
rect 8202 4020 8208 4072
rect 8260 4060 8266 4072
rect 8864 4060 8892 4100
rect 10686 4088 10692 4100
rect 10744 4088 10750 4140
rect 10778 4088 10784 4140
rect 10836 4128 10842 4140
rect 11698 4128 11704 4140
rect 10836 4100 10881 4128
rect 11659 4100 11704 4128
rect 10836 4088 10842 4100
rect 11698 4088 11704 4100
rect 11756 4088 11762 4140
rect 11977 4131 12035 4137
rect 11977 4097 11989 4131
rect 12023 4128 12035 4131
rect 12897 4131 12955 4137
rect 12023 4100 12112 4128
rect 12023 4097 12035 4100
rect 11977 4091 12035 4097
rect 12084 4072 12112 4100
rect 12897 4097 12909 4131
rect 12943 4128 12955 4131
rect 13096 4128 13124 4168
rect 13814 4156 13820 4168
rect 13872 4156 13878 4208
rect 17972 4168 18828 4196
rect 12943 4100 13124 4128
rect 12943 4097 12955 4100
rect 12897 4091 12955 4097
rect 14090 4088 14096 4140
rect 14148 4128 14154 4140
rect 15746 4128 15752 4140
rect 14148 4100 15608 4128
rect 15707 4100 15752 4128
rect 14148 4088 14154 4100
rect 8260 4032 8892 4060
rect 8260 4020 8266 4032
rect 8938 4020 8944 4072
rect 8996 4060 9002 4072
rect 10962 4060 10968 4072
rect 8996 4032 10968 4060
rect 8996 4020 9002 4032
rect 10962 4020 10968 4032
rect 11020 4060 11026 4072
rect 11149 4063 11207 4069
rect 11149 4060 11161 4063
rect 11020 4032 11161 4060
rect 11020 4020 11026 4032
rect 11149 4029 11161 4032
rect 11195 4029 11207 4063
rect 11873 4063 11931 4069
rect 11873 4060 11885 4063
rect 11149 4023 11207 4029
rect 11808 4032 11885 4060
rect 5040 3964 6868 3992
rect 5040 3952 5046 3964
rect 7282 3952 7288 4004
rect 7340 3992 7346 4004
rect 9033 3995 9091 4001
rect 9033 3992 9045 3995
rect 7340 3964 9045 3992
rect 7340 3952 7346 3964
rect 9033 3961 9045 3964
rect 9079 3961 9091 3995
rect 9033 3955 9091 3961
rect 9214 3952 9220 4004
rect 9272 3992 9278 4004
rect 11808 3992 11836 4032
rect 11873 4029 11885 4032
rect 11919 4029 11931 4063
rect 11873 4023 11931 4029
rect 12066 4020 12072 4072
rect 12124 4020 12130 4072
rect 12253 4063 12311 4069
rect 12253 4029 12265 4063
rect 12299 4029 12311 4063
rect 12253 4023 12311 4029
rect 12345 4063 12403 4069
rect 12345 4029 12357 4063
rect 12391 4060 12403 4063
rect 14734 4060 14740 4072
rect 12391 4032 14740 4060
rect 12391 4029 12403 4032
rect 12345 4023 12403 4029
rect 9272 3964 11836 3992
rect 9272 3952 9278 3964
rect 2866 3924 2872 3936
rect 1912 3896 2728 3924
rect 2827 3896 2872 3924
rect 1912 3884 1918 3896
rect 2866 3884 2872 3896
rect 2924 3884 2930 3936
rect 3418 3884 3424 3936
rect 3476 3924 3482 3936
rect 3697 3927 3755 3933
rect 3697 3924 3709 3927
rect 3476 3896 3709 3924
rect 3476 3884 3482 3896
rect 3697 3893 3709 3896
rect 3743 3924 3755 3927
rect 4338 3924 4344 3936
rect 3743 3896 4344 3924
rect 3743 3893 3755 3896
rect 3697 3887 3755 3893
rect 4338 3884 4344 3896
rect 4396 3884 4402 3936
rect 7006 3884 7012 3936
rect 7064 3924 7070 3936
rect 7837 3927 7895 3933
rect 7837 3924 7849 3927
rect 7064 3896 7849 3924
rect 7064 3884 7070 3896
rect 7837 3893 7849 3896
rect 7883 3893 7895 3927
rect 7837 3887 7895 3893
rect 9122 3884 9128 3936
rect 9180 3924 9186 3936
rect 9677 3927 9735 3933
rect 9677 3924 9689 3927
rect 9180 3896 9689 3924
rect 9180 3884 9186 3896
rect 9677 3893 9689 3896
rect 9723 3893 9735 3927
rect 11808 3924 11836 3964
rect 12158 3952 12164 4004
rect 12216 3992 12222 4004
rect 12268 3992 12296 4023
rect 14734 4020 14740 4032
rect 14792 4020 14798 4072
rect 14918 4020 14924 4072
rect 14976 4060 14982 4072
rect 15473 4063 15531 4069
rect 15473 4060 15485 4063
rect 14976 4032 15485 4060
rect 14976 4020 14982 4032
rect 15473 4029 15485 4032
rect 15519 4029 15531 4063
rect 15580 4060 15608 4100
rect 15746 4088 15752 4100
rect 15804 4088 15810 4140
rect 15841 4131 15899 4137
rect 15841 4097 15853 4131
rect 15887 4097 15899 4131
rect 15841 4091 15899 4097
rect 15856 4060 15884 4091
rect 15930 4088 15936 4140
rect 15988 4128 15994 4140
rect 15988 4100 16033 4128
rect 15988 4088 15994 4100
rect 16114 4088 16120 4140
rect 16172 4128 16178 4140
rect 16853 4131 16911 4137
rect 16172 4100 16217 4128
rect 16172 4088 16178 4100
rect 16853 4097 16865 4131
rect 16899 4128 16911 4131
rect 17405 4131 17463 4137
rect 17405 4128 17417 4131
rect 16899 4100 17417 4128
rect 16899 4097 16911 4100
rect 16853 4091 16911 4097
rect 17405 4097 17417 4100
rect 17451 4097 17463 4131
rect 17405 4091 17463 4097
rect 16868 4060 16896 4091
rect 15580 4032 16896 4060
rect 17420 4060 17448 4091
rect 17494 4088 17500 4140
rect 17552 4128 17558 4140
rect 17972 4128 18000 4168
rect 17552 4100 18000 4128
rect 17552 4088 17558 4100
rect 18046 4088 18052 4140
rect 18104 4128 18110 4140
rect 18800 4137 18828 4168
rect 18874 4156 18880 4208
rect 18932 4196 18938 4208
rect 18932 4168 18977 4196
rect 18932 4156 18938 4168
rect 18693 4131 18751 4137
rect 18693 4128 18705 4131
rect 18104 4100 18705 4128
rect 18104 4088 18110 4100
rect 18693 4097 18705 4100
rect 18739 4097 18751 4131
rect 18693 4091 18751 4097
rect 18785 4131 18843 4137
rect 18785 4097 18797 4131
rect 18831 4097 18843 4131
rect 19058 4128 19064 4140
rect 19019 4100 19064 4128
rect 18785 4091 18843 4097
rect 19058 4088 19064 4100
rect 19116 4088 19122 4140
rect 19978 4128 19984 4140
rect 19939 4100 19984 4128
rect 19978 4088 19984 4100
rect 20036 4088 20042 4140
rect 20162 4128 20168 4140
rect 20123 4100 20168 4128
rect 20162 4088 20168 4100
rect 20220 4088 20226 4140
rect 20346 4128 20352 4140
rect 20307 4100 20352 4128
rect 20346 4088 20352 4100
rect 20404 4088 20410 4140
rect 20530 4128 20536 4140
rect 20491 4100 20536 4128
rect 20530 4088 20536 4100
rect 20588 4088 20594 4140
rect 20806 4128 20812 4140
rect 20767 4100 20812 4128
rect 20806 4088 20812 4100
rect 20864 4128 20870 4140
rect 21174 4128 21180 4140
rect 20864 4100 21180 4128
rect 20864 4088 20870 4100
rect 21174 4088 21180 4100
rect 21232 4088 21238 4140
rect 22462 4088 22468 4140
rect 22520 4128 22526 4140
rect 22741 4131 22799 4137
rect 22741 4128 22753 4131
rect 22520 4100 22753 4128
rect 22520 4088 22526 4100
rect 22741 4097 22753 4100
rect 22787 4097 22799 4131
rect 22741 4091 22799 4097
rect 18506 4060 18512 4072
rect 17420 4032 18512 4060
rect 15473 4023 15531 4029
rect 18506 4020 18512 4032
rect 18564 4020 18570 4072
rect 19521 4063 19579 4069
rect 19521 4029 19533 4063
rect 19567 4029 19579 4063
rect 19521 4023 19579 4029
rect 16942 3992 16948 4004
rect 12216 3964 16948 3992
rect 12216 3952 12222 3964
rect 16942 3952 16948 3964
rect 17000 3952 17006 4004
rect 17862 3952 17868 4004
rect 17920 3992 17926 4004
rect 19536 3992 19564 4023
rect 17920 3964 19564 3992
rect 17920 3952 17926 3964
rect 12802 3924 12808 3936
rect 11808 3896 12808 3924
rect 9677 3887 9735 3893
rect 12802 3884 12808 3896
rect 12860 3884 12866 3936
rect 13449 3927 13507 3933
rect 13449 3893 13461 3927
rect 13495 3924 13507 3927
rect 13630 3924 13636 3936
rect 13495 3896 13636 3924
rect 13495 3893 13507 3896
rect 13449 3887 13507 3893
rect 13630 3884 13636 3896
rect 13688 3884 13694 3936
rect 16574 3884 16580 3936
rect 16632 3924 16638 3936
rect 18690 3924 18696 3936
rect 16632 3896 18696 3924
rect 16632 3884 16638 3896
rect 18690 3884 18696 3896
rect 18748 3884 18754 3936
rect 22281 3927 22339 3933
rect 22281 3893 22293 3927
rect 22327 3924 22339 3927
rect 22370 3924 22376 3936
rect 22327 3896 22376 3924
rect 22327 3893 22339 3896
rect 22281 3887 22339 3893
rect 22370 3884 22376 3896
rect 22428 3884 22434 3936
rect 1104 3834 23828 3856
rect 1104 3782 3790 3834
rect 3842 3782 3854 3834
rect 3906 3782 3918 3834
rect 3970 3782 3982 3834
rect 4034 3782 4046 3834
rect 4098 3782 9471 3834
rect 9523 3782 9535 3834
rect 9587 3782 9599 3834
rect 9651 3782 9663 3834
rect 9715 3782 9727 3834
rect 9779 3782 15152 3834
rect 15204 3782 15216 3834
rect 15268 3782 15280 3834
rect 15332 3782 15344 3834
rect 15396 3782 15408 3834
rect 15460 3782 20833 3834
rect 20885 3782 20897 3834
rect 20949 3782 20961 3834
rect 21013 3782 21025 3834
rect 21077 3782 21089 3834
rect 21141 3782 23828 3834
rect 1104 3760 23828 3782
rect 2590 3680 2596 3732
rect 2648 3720 2654 3732
rect 4065 3723 4123 3729
rect 2648 3692 3832 3720
rect 2648 3680 2654 3692
rect 2774 3652 2780 3664
rect 2746 3612 2780 3652
rect 2832 3612 2838 3664
rect 2746 3584 2774 3612
rect 2424 3556 2774 3584
rect 1670 3476 1676 3528
rect 1728 3516 1734 3528
rect 2424 3525 2452 3556
rect 2041 3519 2099 3525
rect 2041 3516 2053 3519
rect 1728 3488 2053 3516
rect 1728 3476 1734 3488
rect 2041 3485 2053 3488
rect 2087 3485 2099 3519
rect 2041 3479 2099 3485
rect 2409 3519 2467 3525
rect 2409 3485 2421 3519
rect 2455 3485 2467 3519
rect 2409 3479 2467 3485
rect 2501 3519 2559 3525
rect 2501 3485 2513 3519
rect 2547 3516 2559 3519
rect 2590 3516 2596 3528
rect 2547 3488 2596 3516
rect 2547 3485 2559 3488
rect 2501 3479 2559 3485
rect 2590 3476 2596 3488
rect 2648 3476 2654 3528
rect 2682 3476 2688 3528
rect 2740 3516 2746 3528
rect 2849 3519 2907 3525
rect 2740 3488 2785 3516
rect 2740 3476 2746 3488
rect 2849 3485 2861 3519
rect 2895 3516 2907 3519
rect 3418 3516 3424 3528
rect 2895 3488 3424 3516
rect 2895 3485 2907 3488
rect 2849 3479 2907 3485
rect 3418 3476 3424 3488
rect 3476 3476 3482 3528
rect 3804 3516 3832 3692
rect 4065 3689 4077 3723
rect 4111 3720 4123 3723
rect 4338 3720 4344 3732
rect 4111 3692 4344 3720
rect 4111 3689 4123 3692
rect 4065 3683 4123 3689
rect 4338 3680 4344 3692
rect 4396 3680 4402 3732
rect 7377 3723 7435 3729
rect 7377 3689 7389 3723
rect 7423 3720 7435 3723
rect 9214 3720 9220 3732
rect 7423 3692 9220 3720
rect 7423 3689 7435 3692
rect 7377 3683 7435 3689
rect 9214 3680 9220 3692
rect 9272 3680 9278 3732
rect 9306 3680 9312 3732
rect 9364 3720 9370 3732
rect 9401 3723 9459 3729
rect 9401 3720 9413 3723
rect 9364 3692 9413 3720
rect 9364 3680 9370 3692
rect 9401 3689 9413 3692
rect 9447 3689 9459 3723
rect 9401 3683 9459 3689
rect 9582 3680 9588 3732
rect 9640 3720 9646 3732
rect 13354 3720 13360 3732
rect 9640 3692 13360 3720
rect 9640 3680 9646 3692
rect 13354 3680 13360 3692
rect 13412 3680 13418 3732
rect 13538 3680 13544 3732
rect 13596 3720 13602 3732
rect 13725 3723 13783 3729
rect 13725 3720 13737 3723
rect 13596 3692 13737 3720
rect 13596 3680 13602 3692
rect 13725 3689 13737 3692
rect 13771 3689 13783 3723
rect 13725 3683 13783 3689
rect 14550 3680 14556 3732
rect 14608 3720 14614 3732
rect 15197 3723 15255 3729
rect 15197 3720 15209 3723
rect 14608 3692 15209 3720
rect 14608 3680 14614 3692
rect 15197 3689 15209 3692
rect 15243 3689 15255 3723
rect 15197 3683 15255 3689
rect 5721 3655 5779 3661
rect 5721 3621 5733 3655
rect 5767 3652 5779 3655
rect 6454 3652 6460 3664
rect 5767 3624 6460 3652
rect 5767 3621 5779 3624
rect 5721 3615 5779 3621
rect 6454 3612 6460 3624
rect 6512 3612 6518 3664
rect 8478 3612 8484 3664
rect 8536 3652 8542 3664
rect 9493 3655 9551 3661
rect 9493 3652 9505 3655
rect 8536 3624 9505 3652
rect 8536 3612 8542 3624
rect 9493 3621 9505 3624
rect 9539 3652 9551 3655
rect 14277 3655 14335 3661
rect 14277 3652 14289 3655
rect 9539 3624 14289 3652
rect 9539 3621 9551 3624
rect 9493 3615 9551 3621
rect 14277 3621 14289 3624
rect 14323 3621 14335 3655
rect 15212 3652 15240 3683
rect 15930 3680 15936 3732
rect 15988 3720 15994 3732
rect 18049 3723 18107 3729
rect 18049 3720 18061 3723
rect 15988 3692 18061 3720
rect 15988 3680 15994 3692
rect 18049 3689 18061 3692
rect 18095 3689 18107 3723
rect 18049 3683 18107 3689
rect 18138 3680 18144 3732
rect 18196 3720 18202 3732
rect 21818 3720 21824 3732
rect 18196 3692 18920 3720
rect 21779 3692 21824 3720
rect 18196 3680 18202 3692
rect 18782 3652 18788 3664
rect 15212 3624 18788 3652
rect 14277 3615 14335 3621
rect 18782 3612 18788 3624
rect 18840 3612 18846 3664
rect 4982 3584 4988 3596
rect 4943 3556 4988 3584
rect 4982 3544 4988 3556
rect 5040 3544 5046 3596
rect 5350 3544 5356 3596
rect 5408 3584 5414 3596
rect 5408 3556 6408 3584
rect 5408 3544 5414 3556
rect 3970 3516 3976 3528
rect 3804 3488 3976 3516
rect 3970 3476 3976 3488
rect 4028 3516 4034 3528
rect 4801 3519 4859 3525
rect 4801 3516 4813 3519
rect 4028 3488 4813 3516
rect 4028 3476 4034 3488
rect 4801 3485 4813 3488
rect 4847 3516 4859 3519
rect 5166 3516 5172 3528
rect 4847 3488 5172 3516
rect 4847 3485 4859 3488
rect 4801 3479 4859 3485
rect 5166 3476 5172 3488
rect 5224 3516 5230 3528
rect 6273 3519 6331 3525
rect 6273 3516 6285 3519
rect 5224 3488 6285 3516
rect 5224 3476 5230 3488
rect 6273 3485 6285 3488
rect 6319 3485 6331 3519
rect 6380 3516 6408 3556
rect 6546 3544 6552 3596
rect 6604 3584 6610 3596
rect 10321 3587 10379 3593
rect 10321 3584 10333 3587
rect 6604 3556 10333 3584
rect 6604 3544 6610 3556
rect 10321 3553 10333 3556
rect 10367 3553 10379 3587
rect 10321 3547 10379 3553
rect 10594 3544 10600 3596
rect 10652 3584 10658 3596
rect 12066 3584 12072 3596
rect 10652 3556 11836 3584
rect 12027 3556 12072 3584
rect 10652 3544 10658 3556
rect 6917 3519 6975 3525
rect 6917 3516 6929 3519
rect 6380 3488 6929 3516
rect 6273 3479 6331 3485
rect 6917 3485 6929 3488
rect 6963 3485 6975 3519
rect 6917 3479 6975 3485
rect 7101 3519 7159 3525
rect 7101 3485 7113 3519
rect 7147 3516 7159 3519
rect 7374 3516 7380 3528
rect 7147 3488 7380 3516
rect 7147 3485 7159 3488
rect 7101 3479 7159 3485
rect 7374 3476 7380 3488
rect 7432 3476 7438 3528
rect 8294 3516 8300 3528
rect 8255 3488 8300 3516
rect 8294 3476 8300 3488
rect 8352 3476 8358 3528
rect 8478 3516 8484 3528
rect 8439 3488 8484 3516
rect 8478 3476 8484 3488
rect 8536 3476 8542 3528
rect 8573 3519 8631 3525
rect 8573 3485 8585 3519
rect 8619 3516 8631 3519
rect 8938 3516 8944 3528
rect 8619 3488 8944 3516
rect 8619 3485 8631 3488
rect 8573 3479 8631 3485
rect 8938 3476 8944 3488
rect 8996 3476 9002 3528
rect 9122 3516 9128 3528
rect 9083 3488 9128 3516
rect 9122 3476 9128 3488
rect 9180 3476 9186 3528
rect 9306 3516 9312 3528
rect 9267 3488 9312 3516
rect 9306 3476 9312 3488
rect 9364 3476 9370 3528
rect 9490 3476 9496 3528
rect 9548 3516 9554 3528
rect 9585 3519 9643 3525
rect 9585 3516 9597 3519
rect 9548 3488 9597 3516
rect 9548 3476 9554 3488
rect 9585 3485 9597 3488
rect 9631 3485 9643 3519
rect 11698 3516 11704 3528
rect 11659 3488 11704 3516
rect 9585 3479 9643 3485
rect 11698 3476 11704 3488
rect 11756 3476 11762 3528
rect 11808 3516 11836 3556
rect 12066 3544 12072 3556
rect 12124 3544 12130 3596
rect 12161 3587 12219 3593
rect 12161 3553 12173 3587
rect 12207 3553 12219 3587
rect 12161 3547 12219 3553
rect 12176 3516 12204 3547
rect 12250 3544 12256 3596
rect 12308 3584 12314 3596
rect 15746 3584 15752 3596
rect 12308 3556 12353 3584
rect 14568 3556 15752 3584
rect 12308 3544 12314 3556
rect 13446 3516 13452 3528
rect 11808 3488 12204 3516
rect 13407 3488 13452 3516
rect 13446 3476 13452 3488
rect 13504 3476 13510 3528
rect 13538 3476 13544 3528
rect 13596 3516 13602 3528
rect 14568 3525 14596 3556
rect 15746 3544 15752 3556
rect 15804 3544 15810 3596
rect 18138 3584 18144 3596
rect 17236 3556 18144 3584
rect 14553 3519 14611 3525
rect 13596 3488 13641 3516
rect 13596 3476 13602 3488
rect 14553 3485 14565 3519
rect 14599 3485 14611 3519
rect 14553 3479 14611 3485
rect 14737 3519 14795 3525
rect 14737 3485 14749 3519
rect 14783 3485 14795 3519
rect 15838 3516 15844 3528
rect 15799 3488 15844 3516
rect 14737 3479 14795 3485
rect 3326 3448 3332 3460
rect 3287 3420 3332 3448
rect 3326 3408 3332 3420
rect 3384 3408 3390 3460
rect 4890 3448 4896 3460
rect 4851 3420 4896 3448
rect 4890 3408 4896 3420
rect 4948 3408 4954 3460
rect 5261 3451 5319 3457
rect 5261 3417 5273 3451
rect 5307 3417 5319 3451
rect 5261 3411 5319 3417
rect 5276 3380 5304 3411
rect 5810 3408 5816 3460
rect 5868 3448 5874 3460
rect 8312 3448 8340 3476
rect 5868 3420 8340 3448
rect 9861 3451 9919 3457
rect 5868 3408 5874 3420
rect 9861 3417 9873 3451
rect 9907 3448 9919 3451
rect 13081 3451 13139 3457
rect 13081 3448 13093 3451
rect 9907 3420 13093 3448
rect 9907 3417 9919 3420
rect 9861 3411 9919 3417
rect 13081 3417 13093 3420
rect 13127 3417 13139 3451
rect 13081 3411 13139 3417
rect 13354 3408 13360 3460
rect 13412 3448 13418 3460
rect 14752 3448 14780 3479
rect 15838 3476 15844 3488
rect 15896 3476 15902 3528
rect 16114 3516 16120 3528
rect 16075 3488 16120 3516
rect 16114 3476 16120 3488
rect 16172 3476 16178 3528
rect 16574 3516 16580 3528
rect 16535 3488 16580 3516
rect 16574 3476 16580 3488
rect 16632 3476 16638 3528
rect 16942 3516 16948 3528
rect 16903 3488 16948 3516
rect 16942 3476 16948 3488
rect 17000 3476 17006 3528
rect 13412 3420 14780 3448
rect 15749 3451 15807 3457
rect 13412 3408 13418 3420
rect 15749 3417 15761 3451
rect 15795 3448 15807 3451
rect 17236 3448 17264 3556
rect 18138 3544 18144 3556
rect 18196 3544 18202 3596
rect 18690 3584 18696 3596
rect 18651 3556 18696 3584
rect 18690 3544 18696 3556
rect 18748 3544 18754 3596
rect 18892 3584 18920 3692
rect 21818 3680 21824 3692
rect 21876 3680 21882 3732
rect 22370 3720 22376 3732
rect 22331 3692 22376 3720
rect 22370 3680 22376 3692
rect 22428 3680 22434 3732
rect 19334 3612 19340 3664
rect 19392 3652 19398 3664
rect 19521 3655 19579 3661
rect 19521 3652 19533 3655
rect 19392 3624 19533 3652
rect 19392 3612 19398 3624
rect 19521 3621 19533 3624
rect 19567 3621 19579 3655
rect 19521 3615 19579 3621
rect 20530 3584 20536 3596
rect 18892 3556 20536 3584
rect 20530 3544 20536 3556
rect 20588 3584 20594 3596
rect 20588 3556 20760 3584
rect 20588 3544 20594 3556
rect 17313 3519 17371 3525
rect 17313 3485 17325 3519
rect 17359 3516 17371 3519
rect 18046 3516 18052 3528
rect 17359 3488 18052 3516
rect 17359 3485 17371 3488
rect 17313 3479 17371 3485
rect 15795 3420 17264 3448
rect 15795 3417 15807 3420
rect 15749 3411 15807 3417
rect 7558 3380 7564 3392
rect 5276 3352 7564 3380
rect 7558 3340 7564 3352
rect 7616 3340 7622 3392
rect 7650 3340 7656 3392
rect 7708 3380 7714 3392
rect 11146 3380 11152 3392
rect 7708 3352 11152 3380
rect 7708 3340 7714 3352
rect 11146 3340 11152 3352
rect 11204 3340 11210 3392
rect 11238 3340 11244 3392
rect 11296 3380 11302 3392
rect 12250 3380 12256 3392
rect 11296 3352 12256 3380
rect 11296 3340 11302 3352
rect 12250 3340 12256 3352
rect 12308 3340 12314 3392
rect 13446 3340 13452 3392
rect 13504 3380 13510 3392
rect 14461 3383 14519 3389
rect 14461 3380 14473 3383
rect 13504 3352 14473 3380
rect 13504 3340 13510 3352
rect 14461 3349 14473 3352
rect 14507 3349 14519 3383
rect 14461 3343 14519 3349
rect 14642 3340 14648 3392
rect 14700 3380 14706 3392
rect 17328 3380 17356 3479
rect 18046 3476 18052 3488
rect 18104 3476 18110 3528
rect 18230 3516 18236 3528
rect 18191 3488 18236 3516
rect 18230 3476 18236 3488
rect 18288 3476 18294 3528
rect 18506 3476 18512 3528
rect 18564 3525 18570 3528
rect 18564 3519 18593 3525
rect 18581 3485 18593 3519
rect 18564 3479 18593 3485
rect 18564 3476 18570 3479
rect 18782 3476 18788 3528
rect 18840 3516 18846 3528
rect 19429 3519 19487 3525
rect 19429 3516 19441 3519
rect 18840 3488 19441 3516
rect 18840 3476 18846 3488
rect 19429 3485 19441 3488
rect 19475 3516 19487 3519
rect 19978 3516 19984 3528
rect 19475 3488 19984 3516
rect 19475 3485 19487 3488
rect 19429 3479 19487 3485
rect 19978 3476 19984 3488
rect 20036 3476 20042 3528
rect 20162 3516 20168 3528
rect 20123 3488 20168 3516
rect 20162 3476 20168 3488
rect 20220 3476 20226 3528
rect 20346 3516 20352 3528
rect 20307 3488 20352 3516
rect 20346 3476 20352 3488
rect 20404 3476 20410 3528
rect 20732 3525 20760 3556
rect 20717 3519 20775 3525
rect 20717 3485 20729 3519
rect 20763 3485 20775 3519
rect 21174 3516 21180 3528
rect 21135 3488 21180 3516
rect 20717 3479 20775 3485
rect 21174 3476 21180 3488
rect 21232 3476 21238 3528
rect 23293 3519 23351 3525
rect 23293 3485 23305 3519
rect 23339 3516 23351 3519
rect 23382 3516 23388 3528
rect 23339 3488 23388 3516
rect 23339 3485 23351 3488
rect 23293 3479 23351 3485
rect 23382 3476 23388 3488
rect 23440 3476 23446 3528
rect 17862 3408 17868 3460
rect 17920 3448 17926 3460
rect 18325 3451 18383 3457
rect 18325 3448 18337 3451
rect 17920 3420 18337 3448
rect 17920 3408 17926 3420
rect 18325 3417 18337 3420
rect 18371 3417 18383 3451
rect 18325 3411 18383 3417
rect 18417 3451 18475 3457
rect 18417 3417 18429 3451
rect 18463 3448 18475 3451
rect 18874 3448 18880 3460
rect 18463 3420 18880 3448
rect 18463 3417 18475 3420
rect 18417 3411 18475 3417
rect 18874 3408 18880 3420
rect 18932 3408 18938 3460
rect 14700 3352 17356 3380
rect 14700 3340 14706 3352
rect 1104 3290 23987 3312
rect 1104 3238 6630 3290
rect 6682 3238 6694 3290
rect 6746 3238 6758 3290
rect 6810 3238 6822 3290
rect 6874 3238 6886 3290
rect 6938 3238 12311 3290
rect 12363 3238 12375 3290
rect 12427 3238 12439 3290
rect 12491 3238 12503 3290
rect 12555 3238 12567 3290
rect 12619 3238 17992 3290
rect 18044 3238 18056 3290
rect 18108 3238 18120 3290
rect 18172 3238 18184 3290
rect 18236 3238 18248 3290
rect 18300 3238 23673 3290
rect 23725 3238 23737 3290
rect 23789 3238 23801 3290
rect 23853 3238 23865 3290
rect 23917 3238 23929 3290
rect 23981 3238 23987 3290
rect 1104 3216 23987 3238
rect 1854 3136 1860 3188
rect 1912 3176 1918 3188
rect 2590 3176 2596 3188
rect 1912 3148 2360 3176
rect 2551 3148 2596 3176
rect 1912 3136 1918 3148
rect 1946 3000 1952 3052
rect 2004 3040 2010 3052
rect 2332 3049 2360 3148
rect 2590 3136 2596 3148
rect 2648 3136 2654 3188
rect 5534 3136 5540 3188
rect 5592 3176 5598 3188
rect 8202 3176 8208 3188
rect 5592 3148 8208 3176
rect 5592 3136 5598 3148
rect 8202 3136 8208 3148
rect 8260 3176 8266 3188
rect 8389 3179 8447 3185
rect 8260 3148 8340 3176
rect 8260 3136 8266 3148
rect 5350 3068 5356 3120
rect 5408 3108 5414 3120
rect 6733 3111 6791 3117
rect 6733 3108 6745 3111
rect 5408 3080 6745 3108
rect 5408 3068 5414 3080
rect 6733 3077 6745 3080
rect 6779 3077 6791 3111
rect 6733 3071 6791 3077
rect 2225 3043 2283 3049
rect 2225 3040 2237 3043
rect 2004 3012 2237 3040
rect 2004 3000 2010 3012
rect 2225 3009 2237 3012
rect 2271 3009 2283 3043
rect 2225 3003 2283 3009
rect 2317 3043 2375 3049
rect 2317 3009 2329 3043
rect 2363 3009 2375 3043
rect 2317 3003 2375 3009
rect 2409 3043 2467 3049
rect 2409 3009 2421 3043
rect 2455 3040 2467 3043
rect 2498 3040 2504 3052
rect 2455 3012 2504 3040
rect 2455 3009 2467 3012
rect 2409 3003 2467 3009
rect 2498 3000 2504 3012
rect 2556 3000 2562 3052
rect 3510 3040 3516 3052
rect 3471 3012 3516 3040
rect 3510 3000 3516 3012
rect 3568 3000 3574 3052
rect 3970 3040 3976 3052
rect 3931 3012 3976 3040
rect 3970 3000 3976 3012
rect 4028 3000 4034 3052
rect 4157 3043 4215 3049
rect 4157 3009 4169 3043
rect 4203 3040 4215 3043
rect 4246 3040 4252 3052
rect 4203 3012 4252 3040
rect 4203 3009 4215 3012
rect 4157 3003 4215 3009
rect 4246 3000 4252 3012
rect 4304 3000 4310 3052
rect 4430 3040 4436 3052
rect 4391 3012 4436 3040
rect 4430 3000 4436 3012
rect 4488 3000 4494 3052
rect 4617 3043 4675 3049
rect 4617 3009 4629 3043
rect 4663 3040 4675 3043
rect 5261 3043 5319 3049
rect 5261 3040 5273 3043
rect 4663 3012 5273 3040
rect 4663 3009 4675 3012
rect 4617 3003 4675 3009
rect 5261 3009 5273 3012
rect 5307 3040 5319 3043
rect 5718 3040 5724 3052
rect 5307 3012 5724 3040
rect 5307 3009 5319 3012
rect 5261 3003 5319 3009
rect 5718 3000 5724 3012
rect 5776 3000 5782 3052
rect 5810 3000 5816 3052
rect 5868 3040 5874 3052
rect 7006 3040 7012 3052
rect 5868 3012 5913 3040
rect 6967 3012 7012 3040
rect 5868 3000 5874 3012
rect 7006 3000 7012 3012
rect 7064 3000 7070 3052
rect 8312 3049 8340 3148
rect 8389 3145 8401 3179
rect 8435 3176 8447 3179
rect 9306 3176 9312 3188
rect 8435 3148 9312 3176
rect 8435 3145 8447 3148
rect 8389 3139 8447 3145
rect 9306 3136 9312 3148
rect 9364 3136 9370 3188
rect 9582 3136 9588 3188
rect 9640 3136 9646 3188
rect 9858 3176 9864 3188
rect 9819 3148 9864 3176
rect 9858 3136 9864 3148
rect 9916 3136 9922 3188
rect 11238 3176 11244 3188
rect 10428 3148 11244 3176
rect 8570 3108 8576 3120
rect 8483 3080 8576 3108
rect 8496 3049 8524 3080
rect 8570 3068 8576 3080
rect 8628 3108 8634 3120
rect 9217 3111 9275 3117
rect 9217 3108 9229 3111
rect 8628 3080 9229 3108
rect 8628 3068 8634 3080
rect 9217 3077 9229 3080
rect 9263 3108 9275 3111
rect 9600 3108 9628 3136
rect 10321 3111 10379 3117
rect 10321 3108 10333 3111
rect 9263 3080 9628 3108
rect 10060 3080 10333 3108
rect 9263 3077 9275 3080
rect 9217 3071 9275 3077
rect 8297 3043 8355 3049
rect 8297 3009 8309 3043
rect 8343 3009 8355 3043
rect 8297 3003 8355 3009
rect 8481 3043 8539 3049
rect 8481 3009 8493 3043
rect 8527 3009 8539 3043
rect 8481 3003 8539 3009
rect 9585 3043 9643 3049
rect 9585 3009 9597 3043
rect 9631 3040 9643 3043
rect 10060 3040 10088 3080
rect 10321 3077 10333 3080
rect 10367 3077 10379 3111
rect 10321 3071 10379 3077
rect 10428 3040 10456 3148
rect 11238 3136 11244 3148
rect 11296 3136 11302 3188
rect 11422 3136 11428 3188
rect 11480 3176 11486 3188
rect 11701 3179 11759 3185
rect 11701 3176 11713 3179
rect 11480 3148 11713 3176
rect 11480 3136 11486 3148
rect 11701 3145 11713 3148
rect 11747 3176 11759 3179
rect 12342 3176 12348 3188
rect 11747 3148 12348 3176
rect 11747 3145 11759 3148
rect 11701 3139 11759 3145
rect 12342 3136 12348 3148
rect 12400 3136 12406 3188
rect 12805 3179 12863 3185
rect 12805 3145 12817 3179
rect 12851 3176 12863 3179
rect 13538 3176 13544 3188
rect 12851 3148 13544 3176
rect 12851 3145 12863 3148
rect 12805 3139 12863 3145
rect 13538 3136 13544 3148
rect 13596 3136 13602 3188
rect 13630 3136 13636 3188
rect 13688 3176 13694 3188
rect 14185 3179 14243 3185
rect 13688 3148 13733 3176
rect 13688 3136 13694 3148
rect 14185 3145 14197 3179
rect 14231 3176 14243 3179
rect 14550 3176 14556 3188
rect 14231 3148 14556 3176
rect 14231 3145 14243 3148
rect 14185 3139 14243 3145
rect 14550 3136 14556 3148
rect 14608 3136 14614 3188
rect 14734 3176 14740 3188
rect 14695 3148 14740 3176
rect 14734 3136 14740 3148
rect 14792 3136 14798 3188
rect 16850 3176 16856 3188
rect 16811 3148 16856 3176
rect 16850 3136 16856 3148
rect 16908 3136 16914 3188
rect 18233 3179 18291 3185
rect 18233 3145 18245 3179
rect 18279 3176 18291 3179
rect 18322 3176 18328 3188
rect 18279 3148 18328 3176
rect 18279 3145 18291 3148
rect 18233 3139 18291 3145
rect 18322 3136 18328 3148
rect 18380 3136 18386 3188
rect 19518 3136 19524 3188
rect 19576 3176 19582 3188
rect 20349 3179 20407 3185
rect 20349 3176 20361 3179
rect 19576 3148 20361 3176
rect 19576 3136 19582 3148
rect 20349 3145 20361 3148
rect 20395 3145 20407 3179
rect 20349 3139 20407 3145
rect 10686 3068 10692 3120
rect 10744 3108 10750 3120
rect 14752 3108 14780 3136
rect 17862 3108 17868 3120
rect 10744 3080 14228 3108
rect 14752 3080 14964 3108
rect 10744 3068 10750 3080
rect 10594 3040 10600 3052
rect 9631 3012 10088 3040
rect 10336 3012 10456 3040
rect 10555 3012 10600 3040
rect 9631 3009 9643 3012
rect 9585 3003 9643 3009
rect 3329 2975 3387 2981
rect 3329 2941 3341 2975
rect 3375 2972 3387 2975
rect 3418 2972 3424 2984
rect 3375 2944 3424 2972
rect 3375 2941 3387 2944
rect 3329 2935 3387 2941
rect 3418 2932 3424 2944
rect 3476 2932 3482 2984
rect 5353 2975 5411 2981
rect 5353 2941 5365 2975
rect 5399 2972 5411 2975
rect 5442 2972 5448 2984
rect 5399 2944 5448 2972
rect 5399 2941 5411 2944
rect 5353 2935 5411 2941
rect 5442 2932 5448 2944
rect 5500 2932 5506 2984
rect 5626 2972 5632 2984
rect 5587 2944 5632 2972
rect 5626 2932 5632 2944
rect 5684 2932 5690 2984
rect 10336 2981 10364 3012
rect 10594 3000 10600 3012
rect 10652 3000 10658 3052
rect 11054 3000 11060 3052
rect 11112 3040 11118 3052
rect 12158 3040 12164 3052
rect 11112 3012 12164 3040
rect 11112 3000 11118 3012
rect 12158 3000 12164 3012
rect 12216 3040 12222 3052
rect 12437 3043 12495 3049
rect 12437 3040 12449 3043
rect 12216 3012 12449 3040
rect 12216 3000 12222 3012
rect 12437 3009 12449 3012
rect 12483 3009 12495 3043
rect 12437 3003 12495 3009
rect 12621 3043 12679 3049
rect 12621 3009 12633 3043
rect 12667 3040 12679 3043
rect 13262 3040 13268 3052
rect 12667 3012 13268 3040
rect 12667 3009 12679 3012
rect 12621 3003 12679 3009
rect 13262 3000 13268 3012
rect 13320 3000 13326 3052
rect 14200 3040 14228 3080
rect 14642 3040 14648 3052
rect 14200 3012 14648 3040
rect 14634 3010 14648 3012
rect 14642 3000 14648 3010
rect 14700 3000 14706 3052
rect 14826 3040 14832 3052
rect 14787 3012 14832 3040
rect 14826 3000 14832 3012
rect 14884 3000 14890 3052
rect 14936 3040 14964 3080
rect 17144 3080 17868 3108
rect 15749 3043 15807 3049
rect 14936 3038 15700 3040
rect 15749 3038 15761 3043
rect 14936 3012 15761 3038
rect 15672 3010 15761 3012
rect 15749 3009 15761 3010
rect 15795 3009 15807 3043
rect 15749 3003 15807 3009
rect 15933 3043 15991 3049
rect 15933 3009 15945 3043
rect 15979 3009 15991 3043
rect 17034 3040 17040 3052
rect 16995 3012 17040 3040
rect 15933 3003 15991 3009
rect 9677 2975 9735 2981
rect 9677 2941 9689 2975
rect 9723 2941 9735 2975
rect 9677 2935 9735 2941
rect 10321 2975 10379 2981
rect 10321 2941 10333 2975
rect 10367 2941 10379 2975
rect 11422 2972 11428 2984
rect 10321 2935 10379 2941
rect 10428 2944 11428 2972
rect 2130 2864 2136 2916
rect 2188 2904 2194 2916
rect 3142 2904 3148 2916
rect 2188 2876 3148 2904
rect 2188 2864 2194 2876
rect 3142 2864 3148 2876
rect 3200 2864 3206 2916
rect 4249 2907 4307 2913
rect 4249 2873 4261 2907
rect 4295 2873 4307 2907
rect 4249 2867 4307 2873
rect 4341 2907 4399 2913
rect 4341 2873 4353 2907
rect 4387 2904 4399 2907
rect 4890 2904 4896 2916
rect 4387 2876 4896 2904
rect 4387 2873 4399 2876
rect 4341 2867 4399 2873
rect 1673 2839 1731 2845
rect 1673 2805 1685 2839
rect 1719 2836 1731 2839
rect 4154 2836 4160 2848
rect 1719 2808 4160 2836
rect 1719 2805 1731 2808
rect 1673 2799 1731 2805
rect 4154 2796 4160 2808
rect 4212 2796 4218 2848
rect 4264 2836 4292 2867
rect 4890 2864 4896 2876
rect 4948 2864 4954 2916
rect 7837 2907 7895 2913
rect 7837 2873 7849 2907
rect 7883 2904 7895 2907
rect 8570 2904 8576 2916
rect 7883 2876 8576 2904
rect 7883 2873 7895 2876
rect 7837 2867 7895 2873
rect 8570 2864 8576 2876
rect 8628 2864 8634 2916
rect 9692 2904 9720 2935
rect 10428 2904 10456 2944
rect 11422 2932 11428 2944
rect 11480 2932 11486 2984
rect 12066 2932 12072 2984
rect 12124 2972 12130 2984
rect 15948 2972 15976 3003
rect 17034 3000 17040 3012
rect 17092 3040 17098 3052
rect 17144 3040 17172 3080
rect 17862 3068 17868 3080
rect 17920 3068 17926 3120
rect 18598 3108 18604 3120
rect 18559 3080 18604 3108
rect 18598 3068 18604 3080
rect 18656 3068 18662 3120
rect 20165 3111 20223 3117
rect 20165 3108 20177 3111
rect 19306 3080 20177 3108
rect 17310 3040 17316 3052
rect 17092 3012 17172 3040
rect 17271 3012 17316 3040
rect 17092 3000 17098 3012
rect 17310 3000 17316 3012
rect 17368 3000 17374 3052
rect 18417 3043 18475 3049
rect 18417 3009 18429 3043
rect 18463 3009 18475 3043
rect 18690 3040 18696 3052
rect 18603 3012 18696 3040
rect 18417 3003 18475 3009
rect 18432 2972 18460 3003
rect 18690 3000 18696 3012
rect 18748 3040 18754 3052
rect 19306 3040 19334 3080
rect 20165 3077 20177 3080
rect 20211 3108 20223 3111
rect 20622 3108 20628 3120
rect 20211 3080 20628 3108
rect 20211 3077 20223 3080
rect 20165 3071 20223 3077
rect 20622 3068 20628 3080
rect 20680 3068 20686 3120
rect 18748 3012 19334 3040
rect 19981 3043 20039 3049
rect 18748 3000 18754 3012
rect 19981 3009 19993 3043
rect 20027 3009 20039 3043
rect 19981 3003 20039 3009
rect 19058 2972 19064 2984
rect 12124 2944 19064 2972
rect 12124 2932 12130 2944
rect 19058 2932 19064 2944
rect 19116 2972 19122 2984
rect 19996 2972 20024 3003
rect 19116 2944 20024 2972
rect 19116 2932 19122 2944
rect 9692 2876 10456 2904
rect 10505 2907 10563 2913
rect 10505 2873 10517 2907
rect 10551 2904 10563 2907
rect 11149 2907 11207 2913
rect 11149 2904 11161 2907
rect 10551 2876 11161 2904
rect 10551 2873 10563 2876
rect 10505 2867 10563 2873
rect 11149 2873 11161 2876
rect 11195 2904 11207 2907
rect 11238 2904 11244 2916
rect 11195 2876 11244 2904
rect 11195 2873 11207 2876
rect 11149 2867 11207 2873
rect 11238 2864 11244 2876
rect 11296 2864 11302 2916
rect 17586 2864 17592 2916
rect 17644 2904 17650 2916
rect 19426 2904 19432 2916
rect 17644 2876 19432 2904
rect 17644 2864 17650 2876
rect 19426 2864 19432 2876
rect 19484 2864 19490 2916
rect 20162 2864 20168 2916
rect 20220 2904 20226 2916
rect 20809 2907 20867 2913
rect 20809 2904 20821 2907
rect 20220 2876 20821 2904
rect 20220 2864 20226 2876
rect 20809 2873 20821 2876
rect 20855 2873 20867 2907
rect 20809 2867 20867 2873
rect 4982 2836 4988 2848
rect 4264 2808 4988 2836
rect 4982 2796 4988 2808
rect 5040 2796 5046 2848
rect 6086 2796 6092 2848
rect 6144 2836 6150 2848
rect 10410 2836 10416 2848
rect 6144 2808 10416 2836
rect 6144 2796 6150 2808
rect 10410 2796 10416 2808
rect 10468 2796 10474 2848
rect 15746 2796 15752 2848
rect 15804 2836 15810 2848
rect 15841 2839 15899 2845
rect 15841 2836 15853 2839
rect 15804 2808 15853 2836
rect 15804 2796 15810 2808
rect 15841 2805 15853 2808
rect 15887 2836 15899 2839
rect 17221 2839 17279 2845
rect 17221 2836 17233 2839
rect 15887 2808 17233 2836
rect 15887 2805 15899 2808
rect 15841 2799 15899 2805
rect 17221 2805 17233 2808
rect 17267 2805 17279 2839
rect 17221 2799 17279 2805
rect 18322 2796 18328 2848
rect 18380 2836 18386 2848
rect 19153 2839 19211 2845
rect 19153 2836 19165 2839
rect 18380 2808 19165 2836
rect 18380 2796 18386 2808
rect 19153 2805 19165 2808
rect 19199 2805 19211 2839
rect 19153 2799 19211 2805
rect 21450 2796 21456 2848
rect 21508 2836 21514 2848
rect 22005 2839 22063 2845
rect 22005 2836 22017 2839
rect 21508 2808 22017 2836
rect 21508 2796 21514 2808
rect 22005 2805 22017 2808
rect 22051 2805 22063 2839
rect 22005 2799 22063 2805
rect 22738 2796 22744 2848
rect 22796 2836 22802 2848
rect 22833 2839 22891 2845
rect 22833 2836 22845 2839
rect 22796 2808 22845 2836
rect 22796 2796 22802 2808
rect 22833 2805 22845 2808
rect 22879 2805 22891 2839
rect 22833 2799 22891 2805
rect 1104 2746 23828 2768
rect 1104 2694 3790 2746
rect 3842 2694 3854 2746
rect 3906 2694 3918 2746
rect 3970 2694 3982 2746
rect 4034 2694 4046 2746
rect 4098 2694 9471 2746
rect 9523 2694 9535 2746
rect 9587 2694 9599 2746
rect 9651 2694 9663 2746
rect 9715 2694 9727 2746
rect 9779 2694 15152 2746
rect 15204 2694 15216 2746
rect 15268 2694 15280 2746
rect 15332 2694 15344 2746
rect 15396 2694 15408 2746
rect 15460 2694 20833 2746
rect 20885 2694 20897 2746
rect 20949 2694 20961 2746
rect 21013 2694 21025 2746
rect 21077 2694 21089 2746
rect 21141 2694 23828 2746
rect 1104 2672 23828 2694
rect 4430 2592 4436 2644
rect 4488 2632 4494 2644
rect 5353 2635 5411 2641
rect 4488 2604 5120 2632
rect 4488 2592 4494 2604
rect 4890 2524 4896 2576
rect 4948 2564 4954 2576
rect 5092 2573 5120 2604
rect 5353 2601 5365 2635
rect 5399 2632 5411 2635
rect 5810 2632 5816 2644
rect 5399 2604 5816 2632
rect 5399 2601 5411 2604
rect 5353 2595 5411 2601
rect 5810 2592 5816 2604
rect 5868 2592 5874 2644
rect 5997 2635 6055 2641
rect 5997 2601 6009 2635
rect 6043 2632 6055 2635
rect 6178 2632 6184 2644
rect 6043 2604 6184 2632
rect 6043 2601 6055 2604
rect 5997 2595 6055 2601
rect 6178 2592 6184 2604
rect 6236 2632 6242 2644
rect 6236 2604 7512 2632
rect 6236 2592 6242 2604
rect 4985 2567 5043 2573
rect 4985 2564 4997 2567
rect 4948 2536 4997 2564
rect 4948 2524 4954 2536
rect 4985 2533 4997 2536
rect 5031 2533 5043 2567
rect 4985 2527 5043 2533
rect 5073 2567 5131 2573
rect 5073 2533 5085 2567
rect 5119 2533 5131 2567
rect 5073 2527 5131 2533
rect 4065 2499 4123 2505
rect 4065 2496 4077 2499
rect 2516 2468 4077 2496
rect 2516 2437 2544 2468
rect 4065 2465 4077 2468
rect 4111 2465 4123 2499
rect 4065 2459 4123 2465
rect 4264 2468 6776 2496
rect 2501 2431 2559 2437
rect 2501 2397 2513 2431
rect 2547 2397 2559 2431
rect 2501 2391 2559 2397
rect 3421 2431 3479 2437
rect 3421 2397 3433 2431
rect 3467 2397 3479 2431
rect 3421 2391 3479 2397
rect 2225 2363 2283 2369
rect 2225 2329 2237 2363
rect 2271 2360 2283 2363
rect 2774 2360 2780 2372
rect 2271 2332 2780 2360
rect 2271 2329 2283 2332
rect 2225 2323 2283 2329
rect 2774 2320 2780 2332
rect 2832 2320 2838 2372
rect 3145 2363 3203 2369
rect 3145 2329 3157 2363
rect 3191 2329 3203 2363
rect 3436 2360 3464 2391
rect 4154 2388 4160 2440
rect 4212 2428 4218 2440
rect 4264 2437 4292 2468
rect 4249 2431 4307 2437
rect 4249 2428 4261 2431
rect 4212 2400 4261 2428
rect 4212 2388 4218 2400
rect 4249 2397 4261 2400
rect 4295 2397 4307 2431
rect 4249 2391 4307 2397
rect 4338 2388 4344 2440
rect 4396 2428 4402 2440
rect 4893 2431 4951 2437
rect 4893 2428 4905 2431
rect 4396 2400 4905 2428
rect 4396 2388 4402 2400
rect 4893 2397 4905 2400
rect 4939 2397 4951 2431
rect 5166 2428 5172 2440
rect 5127 2400 5172 2428
rect 4893 2391 4951 2397
rect 5166 2388 5172 2400
rect 5224 2388 5230 2440
rect 6454 2428 6460 2440
rect 5920 2400 6460 2428
rect 5920 2360 5948 2400
rect 6454 2388 6460 2400
rect 6512 2388 6518 2440
rect 6748 2428 6776 2468
rect 7009 2431 7067 2437
rect 7009 2428 7021 2431
rect 6748 2400 7021 2428
rect 7009 2397 7021 2400
rect 7055 2428 7067 2431
rect 7374 2428 7380 2440
rect 7055 2400 7380 2428
rect 7055 2397 7067 2400
rect 7009 2391 7067 2397
rect 7374 2388 7380 2400
rect 7432 2388 7438 2440
rect 7484 2437 7512 2604
rect 12342 2592 12348 2644
rect 12400 2632 12406 2644
rect 14458 2632 14464 2644
rect 12400 2604 14464 2632
rect 12400 2592 12406 2604
rect 14458 2592 14464 2604
rect 14516 2632 14522 2644
rect 16301 2635 16359 2641
rect 16301 2632 16313 2635
rect 14516 2604 16313 2632
rect 14516 2592 14522 2604
rect 16301 2601 16313 2604
rect 16347 2632 16359 2635
rect 17310 2632 17316 2644
rect 16347 2604 17316 2632
rect 16347 2601 16359 2604
rect 16301 2595 16359 2601
rect 17310 2592 17316 2604
rect 17368 2592 17374 2644
rect 18598 2592 18604 2644
rect 18656 2632 18662 2644
rect 18785 2635 18843 2641
rect 18785 2632 18797 2635
rect 18656 2604 18797 2632
rect 18656 2592 18662 2604
rect 18785 2601 18797 2604
rect 18831 2601 18843 2635
rect 19426 2632 19432 2644
rect 19387 2604 19432 2632
rect 18785 2595 18843 2601
rect 19426 2592 19432 2604
rect 19484 2592 19490 2644
rect 20622 2592 20628 2644
rect 20680 2632 20686 2644
rect 21361 2635 21419 2641
rect 21361 2632 21373 2635
rect 20680 2604 21373 2632
rect 20680 2592 20686 2604
rect 21361 2601 21373 2604
rect 21407 2601 21419 2635
rect 21361 2595 21419 2601
rect 7650 2496 7656 2508
rect 7611 2468 7656 2496
rect 7650 2456 7656 2468
rect 7708 2456 7714 2508
rect 16298 2456 16304 2508
rect 16356 2496 16362 2508
rect 17497 2499 17555 2505
rect 17497 2496 17509 2499
rect 16356 2468 17509 2496
rect 16356 2456 16362 2468
rect 17497 2465 17509 2468
rect 17543 2465 17555 2499
rect 17497 2459 17555 2465
rect 18874 2456 18880 2508
rect 18932 2496 18938 2508
rect 20073 2499 20131 2505
rect 20073 2496 20085 2499
rect 18932 2468 20085 2496
rect 18932 2456 18938 2468
rect 20073 2465 20085 2468
rect 20119 2465 20131 2499
rect 20073 2459 20131 2465
rect 7469 2431 7527 2437
rect 7469 2397 7481 2431
rect 7515 2397 7527 2431
rect 7469 2391 7527 2397
rect 8573 2431 8631 2437
rect 8573 2397 8585 2431
rect 8619 2428 8631 2431
rect 9214 2428 9220 2440
rect 8619 2400 9220 2428
rect 8619 2397 8631 2400
rect 8573 2391 8631 2397
rect 9214 2388 9220 2400
rect 9272 2388 9278 2440
rect 9858 2428 9864 2440
rect 9819 2400 9864 2428
rect 9858 2388 9864 2400
rect 9916 2388 9922 2440
rect 10502 2428 10508 2440
rect 10463 2400 10508 2428
rect 10502 2388 10508 2400
rect 10560 2388 10566 2440
rect 11146 2428 11152 2440
rect 11107 2400 11152 2428
rect 11146 2388 11152 2400
rect 11204 2388 11210 2440
rect 11790 2388 11796 2440
rect 11848 2428 11854 2440
rect 11885 2431 11943 2437
rect 11885 2428 11897 2431
rect 11848 2400 11897 2428
rect 11848 2388 11854 2400
rect 11885 2397 11897 2400
rect 11931 2397 11943 2431
rect 11885 2391 11943 2397
rect 12529 2431 12587 2437
rect 12529 2397 12541 2431
rect 12575 2428 12587 2431
rect 12710 2428 12716 2440
rect 12575 2400 12716 2428
rect 12575 2397 12587 2400
rect 12529 2391 12587 2397
rect 12710 2388 12716 2400
rect 12768 2388 12774 2440
rect 13078 2388 13084 2440
rect 13136 2428 13142 2440
rect 13173 2431 13231 2437
rect 13173 2428 13185 2431
rect 13136 2400 13185 2428
rect 13136 2388 13142 2400
rect 13173 2397 13185 2400
rect 13219 2397 13231 2431
rect 13173 2391 13231 2397
rect 13722 2388 13728 2440
rect 13780 2428 13786 2440
rect 14277 2431 14335 2437
rect 14277 2428 14289 2431
rect 13780 2400 14289 2428
rect 13780 2388 13786 2400
rect 14277 2397 14289 2400
rect 14323 2397 14335 2431
rect 14277 2391 14335 2397
rect 14366 2388 14372 2440
rect 14424 2428 14430 2440
rect 14921 2431 14979 2437
rect 14921 2428 14933 2431
rect 14424 2400 14933 2428
rect 14424 2388 14430 2400
rect 14921 2397 14933 2400
rect 14967 2397 14979 2431
rect 14921 2391 14979 2397
rect 15010 2388 15016 2440
rect 15068 2428 15074 2440
rect 15565 2431 15623 2437
rect 15565 2428 15577 2431
rect 15068 2400 15577 2428
rect 15068 2388 15074 2400
rect 15565 2397 15577 2400
rect 15611 2397 15623 2431
rect 15565 2391 15623 2397
rect 15654 2388 15660 2440
rect 15712 2428 15718 2440
rect 16853 2431 16911 2437
rect 16853 2428 16865 2431
rect 15712 2400 16865 2428
rect 15712 2388 15718 2400
rect 16853 2397 16865 2400
rect 16899 2397 16911 2431
rect 16853 2391 16911 2397
rect 16942 2388 16948 2440
rect 17000 2428 17006 2440
rect 18141 2431 18199 2437
rect 18141 2428 18153 2431
rect 17000 2400 18153 2428
rect 17000 2388 17006 2400
rect 18141 2397 18153 2400
rect 18187 2397 18199 2431
rect 18141 2391 18199 2397
rect 19518 2388 19524 2440
rect 19576 2428 19582 2440
rect 20717 2431 20775 2437
rect 20717 2428 20729 2431
rect 19576 2400 20729 2428
rect 19576 2388 19582 2400
rect 20717 2397 20729 2400
rect 20763 2397 20775 2431
rect 20717 2391 20775 2397
rect 20806 2388 20812 2440
rect 20864 2428 20870 2440
rect 22005 2431 22063 2437
rect 22005 2428 22017 2431
rect 20864 2400 22017 2428
rect 20864 2388 20870 2400
rect 22005 2397 22017 2400
rect 22051 2397 22063 2431
rect 22005 2391 22063 2397
rect 22094 2388 22100 2440
rect 22152 2428 22158 2440
rect 22649 2431 22707 2437
rect 22649 2428 22661 2431
rect 22152 2400 22661 2428
rect 22152 2388 22158 2400
rect 22649 2397 22661 2400
rect 22695 2397 22707 2431
rect 22649 2391 22707 2397
rect 3436 2332 5948 2360
rect 3145 2323 3203 2329
rect 3160 2292 3188 2323
rect 5994 2320 6000 2372
rect 6052 2360 6058 2372
rect 6733 2363 6791 2369
rect 6733 2360 6745 2363
rect 6052 2332 6745 2360
rect 6052 2320 6058 2332
rect 6733 2329 6745 2332
rect 6779 2329 6791 2363
rect 7392 2360 7420 2388
rect 9125 2363 9183 2369
rect 9125 2360 9137 2363
rect 7392 2332 9137 2360
rect 6733 2323 6791 2329
rect 9125 2329 9137 2332
rect 9171 2329 9183 2363
rect 9125 2323 9183 2329
rect 4706 2292 4712 2304
rect 3160 2264 4712 2292
rect 4706 2252 4712 2264
rect 4764 2252 4770 2304
rect 1104 2202 23987 2224
rect 1104 2150 6630 2202
rect 6682 2150 6694 2202
rect 6746 2150 6758 2202
rect 6810 2150 6822 2202
rect 6874 2150 6886 2202
rect 6938 2150 12311 2202
rect 12363 2150 12375 2202
rect 12427 2150 12439 2202
rect 12491 2150 12503 2202
rect 12555 2150 12567 2202
rect 12619 2150 17992 2202
rect 18044 2150 18056 2202
rect 18108 2150 18120 2202
rect 18172 2150 18184 2202
rect 18236 2150 18248 2202
rect 18300 2150 23673 2202
rect 23725 2150 23737 2202
rect 23789 2150 23801 2202
rect 23853 2150 23865 2202
rect 23917 2150 23929 2202
rect 23981 2150 23987 2202
rect 1104 2128 23987 2150
rect 1486 1164 1492 1216
rect 1544 1204 1550 1216
rect 7650 1204 7656 1216
rect 1544 1176 7656 1204
rect 1544 1164 1550 1176
rect 7650 1164 7656 1176
rect 7708 1164 7714 1216
<< via1 >>
rect 3790 22278 3842 22330
rect 3854 22278 3906 22330
rect 3918 22278 3970 22330
rect 3982 22278 4034 22330
rect 4046 22278 4098 22330
rect 9471 22278 9523 22330
rect 9535 22278 9587 22330
rect 9599 22278 9651 22330
rect 9663 22278 9715 22330
rect 9727 22278 9779 22330
rect 15152 22278 15204 22330
rect 15216 22278 15268 22330
rect 15280 22278 15332 22330
rect 15344 22278 15396 22330
rect 15408 22278 15460 22330
rect 20833 22278 20885 22330
rect 20897 22278 20949 22330
rect 20961 22278 21013 22330
rect 21025 22278 21077 22330
rect 21089 22278 21141 22330
rect 21180 22040 21232 22092
rect 10508 22015 10560 22024
rect 10508 21981 10517 22015
rect 10517 21981 10551 22015
rect 10551 21981 10560 22015
rect 10508 21972 10560 21981
rect 7472 21904 7524 21956
rect 19984 21972 20036 22024
rect 22376 21972 22428 22024
rect 6276 21836 6328 21888
rect 8944 21836 8996 21888
rect 11336 21836 11388 21888
rect 12440 21836 12492 21888
rect 17408 21904 17460 21956
rect 14004 21836 14056 21888
rect 15108 21836 15160 21888
rect 15660 21879 15712 21888
rect 15660 21845 15669 21879
rect 15669 21845 15703 21879
rect 15703 21845 15712 21879
rect 15660 21836 15712 21845
rect 17684 21879 17736 21888
rect 17684 21845 17693 21879
rect 17693 21845 17727 21879
rect 17727 21845 17736 21879
rect 17684 21836 17736 21845
rect 22376 21836 22428 21888
rect 6630 21734 6682 21786
rect 6694 21734 6746 21786
rect 6758 21734 6810 21786
rect 6822 21734 6874 21786
rect 6886 21734 6938 21786
rect 12311 21734 12363 21786
rect 12375 21734 12427 21786
rect 12439 21734 12491 21786
rect 12503 21734 12555 21786
rect 12567 21734 12619 21786
rect 17992 21734 18044 21786
rect 18056 21734 18108 21786
rect 18120 21734 18172 21786
rect 18184 21734 18236 21786
rect 18248 21734 18300 21786
rect 23673 21734 23725 21786
rect 23737 21734 23789 21786
rect 23801 21734 23853 21786
rect 23865 21734 23917 21786
rect 23929 21734 23981 21786
rect 2504 21632 2556 21684
rect 5816 21632 5868 21684
rect 2044 21428 2096 21480
rect 2780 21539 2832 21548
rect 2780 21505 2814 21539
rect 2814 21505 2832 21539
rect 5356 21564 5408 21616
rect 9128 21564 9180 21616
rect 2780 21496 2832 21505
rect 5448 21496 5500 21548
rect 10508 21496 10560 21548
rect 1860 21292 1912 21344
rect 6184 21292 6236 21344
rect 8852 21292 8904 21344
rect 11336 21292 11388 21344
rect 11796 21292 11848 21344
rect 13820 21564 13872 21616
rect 14556 21564 14608 21616
rect 13084 21539 13136 21548
rect 13084 21505 13093 21539
rect 13093 21505 13127 21539
rect 13127 21505 13136 21539
rect 13084 21496 13136 21505
rect 14004 21496 14056 21548
rect 14096 21496 14148 21548
rect 15108 21539 15160 21548
rect 13268 21428 13320 21480
rect 12900 21360 12952 21412
rect 15108 21505 15117 21539
rect 15117 21505 15151 21539
rect 15151 21505 15160 21539
rect 15108 21496 15160 21505
rect 19156 21632 19208 21684
rect 19984 21675 20036 21684
rect 19984 21641 19993 21675
rect 19993 21641 20027 21675
rect 20027 21641 20036 21675
rect 19984 21632 20036 21641
rect 21180 21632 21232 21684
rect 17040 21496 17092 21548
rect 17684 21496 17736 21548
rect 14924 21471 14976 21480
rect 14924 21437 14933 21471
rect 14933 21437 14967 21471
rect 14967 21437 14976 21471
rect 14924 21428 14976 21437
rect 15016 21471 15068 21480
rect 15016 21437 15025 21471
rect 15025 21437 15059 21471
rect 15059 21437 15068 21471
rect 15016 21428 15068 21437
rect 14372 21360 14424 21412
rect 15752 21403 15804 21412
rect 15752 21369 15761 21403
rect 15761 21369 15795 21403
rect 15795 21369 15804 21403
rect 15752 21360 15804 21369
rect 21272 21539 21324 21548
rect 21272 21505 21281 21539
rect 21281 21505 21315 21539
rect 21315 21505 21324 21539
rect 22376 21539 22428 21548
rect 21272 21496 21324 21505
rect 22376 21505 22385 21539
rect 22385 21505 22419 21539
rect 22419 21505 22428 21539
rect 22376 21496 22428 21505
rect 14648 21292 14700 21344
rect 16488 21292 16540 21344
rect 3790 21190 3842 21242
rect 3854 21190 3906 21242
rect 3918 21190 3970 21242
rect 3982 21190 4034 21242
rect 4046 21190 4098 21242
rect 9471 21190 9523 21242
rect 9535 21190 9587 21242
rect 9599 21190 9651 21242
rect 9663 21190 9715 21242
rect 9727 21190 9779 21242
rect 15152 21190 15204 21242
rect 15216 21190 15268 21242
rect 15280 21190 15332 21242
rect 15344 21190 15396 21242
rect 15408 21190 15460 21242
rect 20833 21190 20885 21242
rect 20897 21190 20949 21242
rect 20961 21190 21013 21242
rect 21025 21190 21077 21242
rect 21089 21190 21141 21242
rect 9404 21088 9456 21140
rect 11336 21088 11388 21140
rect 5356 20995 5408 21004
rect 5356 20961 5365 20995
rect 5365 20961 5399 20995
rect 5399 20961 5408 20995
rect 5356 20952 5408 20961
rect 9128 20995 9180 21004
rect 9128 20961 9137 20995
rect 9137 20961 9171 20995
rect 9171 20961 9180 20995
rect 9128 20952 9180 20961
rect 2044 20927 2096 20936
rect 2044 20893 2053 20927
rect 2053 20893 2087 20927
rect 2087 20893 2096 20927
rect 2044 20884 2096 20893
rect 13452 21063 13504 21072
rect 13452 21029 13461 21063
rect 13461 21029 13495 21063
rect 13495 21029 13504 21063
rect 13452 21020 13504 21029
rect 13636 21020 13688 21072
rect 16488 21088 16540 21140
rect 21272 21131 21324 21140
rect 21272 21097 21281 21131
rect 21281 21097 21315 21131
rect 21315 21097 21324 21131
rect 21272 21088 21324 21097
rect 14464 21020 14516 21072
rect 14556 21063 14608 21072
rect 14556 21029 14565 21063
rect 14565 21029 14599 21063
rect 14599 21029 14608 21063
rect 14556 21020 14608 21029
rect 15568 21020 15620 21072
rect 16212 21063 16264 21072
rect 16212 21029 16221 21063
rect 16221 21029 16255 21063
rect 16255 21029 16264 21063
rect 16212 21020 16264 21029
rect 11796 20927 11848 20936
rect 1676 20816 1728 20868
rect 4712 20816 4764 20868
rect 9404 20859 9456 20868
rect 9404 20825 9438 20859
rect 9438 20825 9456 20859
rect 9404 20816 9456 20825
rect 3148 20748 3200 20800
rect 3516 20748 3568 20800
rect 11244 20816 11296 20868
rect 11336 20816 11388 20868
rect 11796 20893 11805 20927
rect 11805 20893 11839 20927
rect 11839 20893 11848 20927
rect 11796 20884 11848 20893
rect 12716 20884 12768 20936
rect 14280 20884 14332 20936
rect 10048 20748 10100 20800
rect 13360 20816 13412 20868
rect 14832 20816 14884 20868
rect 15476 20884 15528 20936
rect 15660 20884 15712 20936
rect 16120 20884 16172 20936
rect 22100 20952 22152 21004
rect 16672 20927 16724 20936
rect 16672 20893 16681 20927
rect 16681 20893 16715 20927
rect 16715 20893 16724 20927
rect 16672 20884 16724 20893
rect 16948 20927 17000 20936
rect 16948 20893 16957 20927
rect 16957 20893 16991 20927
rect 16991 20893 17000 20927
rect 16948 20884 17000 20893
rect 18328 20884 18380 20936
rect 21180 20927 21232 20936
rect 21180 20893 21189 20927
rect 21189 20893 21223 20927
rect 21223 20893 21232 20927
rect 21180 20884 21232 20893
rect 22376 20884 22428 20936
rect 15292 20816 15344 20868
rect 12716 20748 12768 20800
rect 13268 20748 13320 20800
rect 15384 20791 15436 20800
rect 15384 20757 15393 20791
rect 15393 20757 15427 20791
rect 15427 20757 15436 20791
rect 15384 20748 15436 20757
rect 15476 20748 15528 20800
rect 15660 20748 15712 20800
rect 6630 20646 6682 20698
rect 6694 20646 6746 20698
rect 6758 20646 6810 20698
rect 6822 20646 6874 20698
rect 6886 20646 6938 20698
rect 12311 20646 12363 20698
rect 12375 20646 12427 20698
rect 12439 20646 12491 20698
rect 12503 20646 12555 20698
rect 12567 20646 12619 20698
rect 17992 20646 18044 20698
rect 18056 20646 18108 20698
rect 18120 20646 18172 20698
rect 18184 20646 18236 20698
rect 18248 20646 18300 20698
rect 23673 20646 23725 20698
rect 23737 20646 23789 20698
rect 23801 20646 23853 20698
rect 23865 20646 23917 20698
rect 23929 20646 23981 20698
rect 11060 20544 11112 20596
rect 4344 20451 4396 20460
rect 4344 20417 4353 20451
rect 4353 20417 4387 20451
rect 4387 20417 4396 20451
rect 4344 20408 4396 20417
rect 9036 20408 9088 20460
rect 12072 20408 12124 20460
rect 12164 20451 12216 20460
rect 12164 20417 12173 20451
rect 12173 20417 12207 20451
rect 12207 20417 12216 20451
rect 14924 20544 14976 20596
rect 15752 20544 15804 20596
rect 13636 20476 13688 20528
rect 12164 20408 12216 20417
rect 12716 20408 12768 20460
rect 13176 20451 13228 20460
rect 13176 20417 13185 20451
rect 13185 20417 13219 20451
rect 13219 20417 13228 20451
rect 13176 20408 13228 20417
rect 13544 20451 13596 20460
rect 13544 20417 13553 20451
rect 13553 20417 13587 20451
rect 13587 20417 13596 20451
rect 13544 20408 13596 20417
rect 15384 20476 15436 20528
rect 14740 20408 14792 20460
rect 14924 20408 14976 20460
rect 15568 20408 15620 20460
rect 15752 20408 15804 20460
rect 15936 20408 15988 20460
rect 17316 20544 17368 20596
rect 16304 20451 16356 20460
rect 16304 20417 16313 20451
rect 16313 20417 16347 20451
rect 16347 20417 16356 20451
rect 16304 20408 16356 20417
rect 16948 20408 17000 20460
rect 17868 20544 17920 20596
rect 2044 20340 2096 20392
rect 14832 20340 14884 20392
rect 13636 20272 13688 20324
rect 15476 20272 15528 20324
rect 17684 20451 17736 20460
rect 17684 20417 17693 20451
rect 17693 20417 17727 20451
rect 17727 20417 17736 20451
rect 17684 20408 17736 20417
rect 18604 20451 18656 20460
rect 18604 20417 18613 20451
rect 18613 20417 18647 20451
rect 18647 20417 18656 20451
rect 18604 20408 18656 20417
rect 19432 20544 19484 20596
rect 22100 20587 22152 20596
rect 22100 20553 22109 20587
rect 22109 20553 22143 20587
rect 22143 20553 22152 20587
rect 22100 20544 22152 20553
rect 18972 20451 19024 20460
rect 18972 20417 18981 20451
rect 18981 20417 19015 20451
rect 19015 20417 19024 20451
rect 19432 20451 19484 20460
rect 18972 20408 19024 20417
rect 19432 20417 19441 20451
rect 19441 20417 19475 20451
rect 19475 20417 19484 20451
rect 19432 20408 19484 20417
rect 20168 20408 20220 20460
rect 22192 20451 22244 20460
rect 20076 20340 20128 20392
rect 17684 20272 17736 20324
rect 19340 20272 19392 20324
rect 22192 20417 22201 20451
rect 22201 20417 22235 20451
rect 22235 20417 22244 20451
rect 22192 20408 22244 20417
rect 11336 20204 11388 20256
rect 14648 20204 14700 20256
rect 16304 20204 16356 20256
rect 3790 20102 3842 20154
rect 3854 20102 3906 20154
rect 3918 20102 3970 20154
rect 3982 20102 4034 20154
rect 4046 20102 4098 20154
rect 9471 20102 9523 20154
rect 9535 20102 9587 20154
rect 9599 20102 9651 20154
rect 9663 20102 9715 20154
rect 9727 20102 9779 20154
rect 15152 20102 15204 20154
rect 15216 20102 15268 20154
rect 15280 20102 15332 20154
rect 15344 20102 15396 20154
rect 15408 20102 15460 20154
rect 20833 20102 20885 20154
rect 20897 20102 20949 20154
rect 20961 20102 21013 20154
rect 21025 20102 21077 20154
rect 21089 20102 21141 20154
rect 12072 20000 12124 20052
rect 15016 20000 15068 20052
rect 18972 20000 19024 20052
rect 2044 19907 2096 19916
rect 2044 19873 2053 19907
rect 2053 19873 2087 19907
rect 2087 19873 2096 19907
rect 2044 19864 2096 19873
rect 9128 19907 9180 19916
rect 9128 19873 9137 19907
rect 9137 19873 9171 19907
rect 9171 19873 9180 19907
rect 9128 19864 9180 19873
rect 13268 19932 13320 19984
rect 15292 19932 15344 19984
rect 16304 19932 16356 19984
rect 16488 19975 16540 19984
rect 16488 19941 16497 19975
rect 16497 19941 16531 19975
rect 16531 19941 16540 19975
rect 16488 19932 16540 19941
rect 16764 19932 16816 19984
rect 1584 19728 1636 19780
rect 5724 19728 5776 19780
rect 3608 19660 3660 19712
rect 4436 19660 4488 19712
rect 10784 19660 10836 19712
rect 11336 19660 11388 19712
rect 12164 19864 12216 19916
rect 12900 19864 12952 19916
rect 15016 19864 15068 19916
rect 15384 19907 15436 19916
rect 15384 19873 15393 19907
rect 15393 19873 15427 19907
rect 15427 19873 15436 19907
rect 15384 19864 15436 19873
rect 17684 19864 17736 19916
rect 19432 19864 19484 19916
rect 20444 19864 20496 19916
rect 13452 19796 13504 19848
rect 14648 19839 14700 19848
rect 14648 19805 14657 19839
rect 14657 19805 14691 19839
rect 14691 19805 14700 19839
rect 14648 19796 14700 19805
rect 16028 19796 16080 19848
rect 16396 19839 16448 19848
rect 16396 19805 16405 19839
rect 16405 19805 16439 19839
rect 16439 19805 16448 19839
rect 16396 19796 16448 19805
rect 17040 19796 17092 19848
rect 18696 19796 18748 19848
rect 20996 19796 21048 19848
rect 13084 19728 13136 19780
rect 16856 19728 16908 19780
rect 14924 19660 14976 19712
rect 15936 19660 15988 19712
rect 17868 19660 17920 19712
rect 19892 19660 19944 19712
rect 6630 19558 6682 19610
rect 6694 19558 6746 19610
rect 6758 19558 6810 19610
rect 6822 19558 6874 19610
rect 6886 19558 6938 19610
rect 12311 19558 12363 19610
rect 12375 19558 12427 19610
rect 12439 19558 12491 19610
rect 12503 19558 12555 19610
rect 12567 19558 12619 19610
rect 17992 19558 18044 19610
rect 18056 19558 18108 19610
rect 18120 19558 18172 19610
rect 18184 19558 18236 19610
rect 18248 19558 18300 19610
rect 23673 19558 23725 19610
rect 23737 19558 23789 19610
rect 23801 19558 23853 19610
rect 23865 19558 23917 19610
rect 23929 19558 23981 19610
rect 5172 19456 5224 19508
rect 5908 19456 5960 19508
rect 11980 19456 12032 19508
rect 16488 19456 16540 19508
rect 7564 19388 7616 19440
rect 3424 19320 3476 19372
rect 4344 19320 4396 19372
rect 7472 19320 7524 19372
rect 8024 19363 8076 19372
rect 8024 19329 8033 19363
rect 8033 19329 8067 19363
rect 8067 19329 8076 19363
rect 8024 19320 8076 19329
rect 9036 19320 9088 19372
rect 14556 19320 14608 19372
rect 15752 19388 15804 19440
rect 16672 19388 16724 19440
rect 18696 19388 18748 19440
rect 14740 19320 14792 19372
rect 15200 19320 15252 19372
rect 2780 19252 2832 19304
rect 12992 19252 13044 19304
rect 15936 19320 15988 19372
rect 17132 19320 17184 19372
rect 17316 19363 17368 19372
rect 17316 19329 17325 19363
rect 17325 19329 17359 19363
rect 17359 19329 17368 19363
rect 17316 19320 17368 19329
rect 18512 19320 18564 19372
rect 19340 19363 19392 19372
rect 19340 19329 19349 19363
rect 19349 19329 19383 19363
rect 19383 19329 19392 19363
rect 19340 19320 19392 19329
rect 19524 19363 19576 19372
rect 19524 19329 19533 19363
rect 19533 19329 19567 19363
rect 19567 19329 19576 19363
rect 19524 19320 19576 19329
rect 19616 19363 19668 19372
rect 19616 19329 19625 19363
rect 19625 19329 19659 19363
rect 19659 19329 19668 19363
rect 20260 19363 20312 19372
rect 19616 19320 19668 19329
rect 20260 19329 20269 19363
rect 20269 19329 20303 19363
rect 20303 19329 20312 19363
rect 20260 19320 20312 19329
rect 21180 19320 21232 19372
rect 22100 19320 22152 19372
rect 15660 19252 15712 19304
rect 18972 19252 19024 19304
rect 19156 19295 19208 19304
rect 19156 19261 19165 19295
rect 19165 19261 19199 19295
rect 19199 19261 19208 19295
rect 19156 19252 19208 19261
rect 20076 19295 20128 19304
rect 20076 19261 20085 19295
rect 20085 19261 20119 19295
rect 20119 19261 20128 19295
rect 20076 19252 20128 19261
rect 20996 19295 21048 19304
rect 20996 19261 21005 19295
rect 21005 19261 21039 19295
rect 21039 19261 21048 19295
rect 20996 19252 21048 19261
rect 21364 19252 21416 19304
rect 14188 19184 14240 19236
rect 15200 19184 15252 19236
rect 15568 19184 15620 19236
rect 22376 19184 22428 19236
rect 14464 19116 14516 19168
rect 14832 19116 14884 19168
rect 19708 19116 19760 19168
rect 21732 19116 21784 19168
rect 3790 19014 3842 19066
rect 3854 19014 3906 19066
rect 3918 19014 3970 19066
rect 3982 19014 4034 19066
rect 4046 19014 4098 19066
rect 9471 19014 9523 19066
rect 9535 19014 9587 19066
rect 9599 19014 9651 19066
rect 9663 19014 9715 19066
rect 9727 19014 9779 19066
rect 15152 19014 15204 19066
rect 15216 19014 15268 19066
rect 15280 19014 15332 19066
rect 15344 19014 15396 19066
rect 15408 19014 15460 19066
rect 20833 19014 20885 19066
rect 20897 19014 20949 19066
rect 20961 19014 21013 19066
rect 21025 19014 21077 19066
rect 21089 19014 21141 19066
rect 5816 18955 5868 18964
rect 5816 18921 5825 18955
rect 5825 18921 5859 18955
rect 5859 18921 5868 18955
rect 5816 18912 5868 18921
rect 7472 18912 7524 18964
rect 14280 18955 14332 18964
rect 14280 18921 14289 18955
rect 14289 18921 14323 18955
rect 14323 18921 14332 18955
rect 14280 18912 14332 18921
rect 14556 18912 14608 18964
rect 15292 18912 15344 18964
rect 15660 18912 15712 18964
rect 16028 18955 16080 18964
rect 16028 18921 16037 18955
rect 16037 18921 16071 18955
rect 16071 18921 16080 18955
rect 16028 18912 16080 18921
rect 18328 18955 18380 18964
rect 18328 18921 18337 18955
rect 18337 18921 18371 18955
rect 18371 18921 18380 18955
rect 18328 18912 18380 18921
rect 14832 18844 14884 18896
rect 18880 18912 18932 18964
rect 19616 18912 19668 18964
rect 22376 18955 22428 18964
rect 22376 18921 22385 18955
rect 22385 18921 22419 18955
rect 22419 18921 22428 18955
rect 22376 18912 22428 18921
rect 9128 18819 9180 18828
rect 9128 18785 9137 18819
rect 9137 18785 9171 18819
rect 9171 18785 9180 18819
rect 9128 18776 9180 18785
rect 12900 18776 12952 18828
rect 13268 18819 13320 18828
rect 13268 18785 13277 18819
rect 13277 18785 13311 18819
rect 13311 18785 13320 18819
rect 13268 18776 13320 18785
rect 16580 18776 16632 18828
rect 20720 18844 20772 18896
rect 2780 18708 2832 18760
rect 5816 18708 5868 18760
rect 12992 18708 13044 18760
rect 13360 18751 13412 18760
rect 13360 18717 13369 18751
rect 13369 18717 13403 18751
rect 13403 18717 13412 18751
rect 13360 18708 13412 18717
rect 14464 18751 14516 18760
rect 14464 18717 14473 18751
rect 14473 18717 14507 18751
rect 14507 18717 14516 18751
rect 14464 18708 14516 18717
rect 15752 18751 15804 18760
rect 8300 18640 8352 18692
rect 10876 18640 10928 18692
rect 12072 18640 12124 18692
rect 14372 18640 14424 18692
rect 14556 18683 14608 18692
rect 14556 18649 14565 18683
rect 14565 18649 14599 18683
rect 14599 18649 14608 18683
rect 14556 18640 14608 18649
rect 2596 18572 2648 18624
rect 10600 18572 10652 18624
rect 14464 18572 14516 18624
rect 14740 18683 14792 18692
rect 14740 18649 14775 18683
rect 14775 18649 14792 18683
rect 14740 18640 14792 18649
rect 15292 18640 15344 18692
rect 15752 18717 15761 18751
rect 15761 18717 15795 18751
rect 15795 18717 15804 18751
rect 15752 18708 15804 18717
rect 16488 18708 16540 18760
rect 16672 18751 16724 18760
rect 16672 18717 16681 18751
rect 16681 18717 16715 18751
rect 16715 18717 16724 18751
rect 16672 18708 16724 18717
rect 16948 18751 17000 18760
rect 16948 18717 16957 18751
rect 16957 18717 16991 18751
rect 16991 18717 17000 18751
rect 16948 18708 17000 18717
rect 18880 18776 18932 18828
rect 18512 18751 18564 18760
rect 18512 18717 18521 18751
rect 18521 18717 18555 18751
rect 18555 18717 18564 18751
rect 18512 18708 18564 18717
rect 17132 18640 17184 18692
rect 17776 18640 17828 18692
rect 18788 18751 18840 18760
rect 18788 18717 18797 18751
rect 18797 18717 18831 18751
rect 18831 18717 18840 18751
rect 18788 18708 18840 18717
rect 18972 18708 19024 18760
rect 19708 18751 19760 18760
rect 19708 18717 19717 18751
rect 19717 18717 19751 18751
rect 19751 18717 19760 18751
rect 19708 18708 19760 18717
rect 19892 18751 19944 18760
rect 19892 18717 19937 18751
rect 19937 18717 19944 18751
rect 19892 18708 19944 18717
rect 20076 18751 20128 18760
rect 20076 18717 20085 18751
rect 20085 18717 20119 18751
rect 20119 18717 20128 18751
rect 20076 18708 20128 18717
rect 20260 18708 20312 18760
rect 20444 18708 20496 18760
rect 21180 18708 21232 18760
rect 20628 18640 20680 18692
rect 15660 18572 15712 18624
rect 17408 18572 17460 18624
rect 20904 18615 20956 18624
rect 20904 18581 20913 18615
rect 20913 18581 20947 18615
rect 20947 18581 20956 18615
rect 20904 18572 20956 18581
rect 22100 18572 22152 18624
rect 6630 18470 6682 18522
rect 6694 18470 6746 18522
rect 6758 18470 6810 18522
rect 6822 18470 6874 18522
rect 6886 18470 6938 18522
rect 12311 18470 12363 18522
rect 12375 18470 12427 18522
rect 12439 18470 12491 18522
rect 12503 18470 12555 18522
rect 12567 18470 12619 18522
rect 17992 18470 18044 18522
rect 18056 18470 18108 18522
rect 18120 18470 18172 18522
rect 18184 18470 18236 18522
rect 18248 18470 18300 18522
rect 23673 18470 23725 18522
rect 23737 18470 23789 18522
rect 23801 18470 23853 18522
rect 23865 18470 23917 18522
rect 23929 18470 23981 18522
rect 9128 18411 9180 18420
rect 9128 18377 9137 18411
rect 9137 18377 9171 18411
rect 9171 18377 9180 18411
rect 9128 18368 9180 18377
rect 13544 18411 13596 18420
rect 13544 18377 13553 18411
rect 13553 18377 13587 18411
rect 13587 18377 13596 18411
rect 13544 18368 13596 18377
rect 14740 18368 14792 18420
rect 16488 18368 16540 18420
rect 17224 18368 17276 18420
rect 7472 18300 7524 18352
rect 2320 18232 2372 18284
rect 14004 18300 14056 18352
rect 16120 18300 16172 18352
rect 18788 18368 18840 18420
rect 19892 18368 19944 18420
rect 21456 18368 21508 18420
rect 22192 18368 22244 18420
rect 19248 18300 19300 18352
rect 2780 18164 2832 18216
rect 12900 18164 12952 18216
rect 3332 18028 3384 18080
rect 13268 18028 13320 18080
rect 14832 18232 14884 18284
rect 15476 18164 15528 18216
rect 18696 18232 18748 18284
rect 19708 18232 19760 18284
rect 20352 18300 20404 18352
rect 22376 18368 22428 18420
rect 20165 18275 20217 18284
rect 20165 18241 20192 18275
rect 20192 18241 20217 18275
rect 20165 18232 20217 18241
rect 20260 18275 20312 18284
rect 20260 18241 20274 18275
rect 20274 18241 20308 18275
rect 20308 18241 20312 18275
rect 20260 18232 20312 18241
rect 22284 18275 22336 18284
rect 18420 18164 18472 18216
rect 22284 18241 22293 18275
rect 22293 18241 22327 18275
rect 22327 18241 22336 18275
rect 22284 18232 22336 18241
rect 22468 18275 22520 18284
rect 22468 18241 22477 18275
rect 22477 18241 22511 18275
rect 22511 18241 22520 18275
rect 22652 18275 22704 18284
rect 22468 18232 22520 18241
rect 22652 18241 22661 18275
rect 22661 18241 22695 18275
rect 22695 18241 22704 18275
rect 22652 18232 22704 18241
rect 14464 18096 14516 18148
rect 16856 18096 16908 18148
rect 16028 18028 16080 18080
rect 16120 18028 16172 18080
rect 16948 18071 17000 18080
rect 16948 18037 16957 18071
rect 16957 18037 16991 18071
rect 16991 18037 17000 18071
rect 16948 18028 17000 18037
rect 17316 18028 17368 18080
rect 19892 18028 19944 18080
rect 3790 17926 3842 17978
rect 3854 17926 3906 17978
rect 3918 17926 3970 17978
rect 3982 17926 4034 17978
rect 4046 17926 4098 17978
rect 9471 17926 9523 17978
rect 9535 17926 9587 17978
rect 9599 17926 9651 17978
rect 9663 17926 9715 17978
rect 9727 17926 9779 17978
rect 15152 17926 15204 17978
rect 15216 17926 15268 17978
rect 15280 17926 15332 17978
rect 15344 17926 15396 17978
rect 15408 17926 15460 17978
rect 20833 17926 20885 17978
rect 20897 17926 20949 17978
rect 20961 17926 21013 17978
rect 21025 17926 21077 17978
rect 21089 17926 21141 17978
rect 14556 17824 14608 17876
rect 18512 17824 18564 17876
rect 19800 17867 19852 17876
rect 19800 17833 19809 17867
rect 19809 17833 19843 17867
rect 19843 17833 19852 17867
rect 19800 17824 19852 17833
rect 22652 17867 22704 17876
rect 22652 17833 22661 17867
rect 22661 17833 22695 17867
rect 22695 17833 22704 17867
rect 22652 17824 22704 17833
rect 12164 17756 12216 17808
rect 7104 17731 7156 17740
rect 7104 17697 7113 17731
rect 7113 17697 7147 17731
rect 7147 17697 7156 17731
rect 7104 17688 7156 17697
rect 8024 17688 8076 17740
rect 9128 17731 9180 17740
rect 9128 17697 9137 17731
rect 9137 17697 9171 17731
rect 9171 17697 9180 17731
rect 9128 17688 9180 17697
rect 17776 17688 17828 17740
rect 2688 17620 2740 17672
rect 12072 17620 12124 17672
rect 2412 17552 2464 17604
rect 6368 17552 6420 17604
rect 13268 17552 13320 17604
rect 13820 17620 13872 17672
rect 14464 17663 14516 17672
rect 14464 17629 14473 17663
rect 14473 17629 14507 17663
rect 14507 17629 14516 17663
rect 14464 17620 14516 17629
rect 16304 17620 16356 17672
rect 16488 17663 16540 17672
rect 16488 17629 16497 17663
rect 16497 17629 16531 17663
rect 16531 17629 16540 17663
rect 16488 17620 16540 17629
rect 14832 17552 14884 17604
rect 17316 17552 17368 17604
rect 17500 17620 17552 17672
rect 17868 17620 17920 17672
rect 18328 17620 18380 17672
rect 19708 17731 19760 17740
rect 19708 17697 19717 17731
rect 19717 17697 19751 17731
rect 19751 17697 19760 17731
rect 19708 17688 19760 17697
rect 19984 17620 20036 17672
rect 20076 17620 20128 17672
rect 21824 17663 21876 17672
rect 21824 17629 21833 17663
rect 21833 17629 21867 17663
rect 21867 17629 21876 17663
rect 21824 17620 21876 17629
rect 19340 17552 19392 17604
rect 19432 17552 19484 17604
rect 2964 17484 3016 17536
rect 5540 17484 5592 17536
rect 10416 17484 10468 17536
rect 11796 17484 11848 17536
rect 12900 17527 12952 17536
rect 12900 17493 12909 17527
rect 12909 17493 12943 17527
rect 12943 17493 12952 17527
rect 12900 17484 12952 17493
rect 15844 17484 15896 17536
rect 16396 17527 16448 17536
rect 16396 17493 16405 17527
rect 16405 17493 16439 17527
rect 16439 17493 16448 17527
rect 16396 17484 16448 17493
rect 16580 17484 16632 17536
rect 17592 17484 17644 17536
rect 20812 17484 20864 17536
rect 20904 17484 20956 17536
rect 22008 17527 22060 17536
rect 22008 17493 22017 17527
rect 22017 17493 22051 17527
rect 22051 17493 22060 17527
rect 22008 17484 22060 17493
rect 6630 17382 6682 17434
rect 6694 17382 6746 17434
rect 6758 17382 6810 17434
rect 6822 17382 6874 17434
rect 6886 17382 6938 17434
rect 12311 17382 12363 17434
rect 12375 17382 12427 17434
rect 12439 17382 12491 17434
rect 12503 17382 12555 17434
rect 12567 17382 12619 17434
rect 17992 17382 18044 17434
rect 18056 17382 18108 17434
rect 18120 17382 18172 17434
rect 18184 17382 18236 17434
rect 18248 17382 18300 17434
rect 23673 17382 23725 17434
rect 23737 17382 23789 17434
rect 23801 17382 23853 17434
rect 23865 17382 23917 17434
rect 23929 17382 23981 17434
rect 12164 17323 12216 17332
rect 12164 17289 12173 17323
rect 12173 17289 12207 17323
rect 12207 17289 12216 17323
rect 12164 17280 12216 17289
rect 10876 17212 10928 17264
rect 14004 17323 14056 17332
rect 14004 17289 14013 17323
rect 14013 17289 14047 17323
rect 14047 17289 14056 17323
rect 14004 17280 14056 17289
rect 14096 17280 14148 17332
rect 8024 17144 8076 17196
rect 8208 17144 8260 17196
rect 15016 17212 15068 17264
rect 18880 17280 18932 17332
rect 19524 17280 19576 17332
rect 20720 17323 20772 17332
rect 20720 17289 20729 17323
rect 20729 17289 20763 17323
rect 20763 17289 20772 17323
rect 20720 17280 20772 17289
rect 13176 17187 13228 17196
rect 2688 17119 2740 17128
rect 2688 17085 2697 17119
rect 2697 17085 2731 17119
rect 2731 17085 2740 17119
rect 2688 17076 2740 17085
rect 5080 17076 5132 17128
rect 13176 17153 13185 17187
rect 13185 17153 13219 17187
rect 13219 17153 13228 17187
rect 13176 17144 13228 17153
rect 14556 17144 14608 17196
rect 15936 17144 15988 17196
rect 17316 17212 17368 17264
rect 17040 17144 17092 17196
rect 20076 17212 20128 17264
rect 13636 17076 13688 17128
rect 14096 17076 14148 17128
rect 11888 17008 11940 17060
rect 13084 17051 13136 17060
rect 13084 17017 13093 17051
rect 13093 17017 13127 17051
rect 13127 17017 13136 17051
rect 13084 17008 13136 17017
rect 14280 17008 14332 17060
rect 14464 17119 14516 17128
rect 14464 17085 14473 17119
rect 14473 17085 14507 17119
rect 14507 17085 14516 17119
rect 14464 17076 14516 17085
rect 15108 17076 15160 17128
rect 15292 17119 15344 17128
rect 15292 17085 15301 17119
rect 15301 17085 15335 17119
rect 15335 17085 15344 17119
rect 15292 17076 15344 17085
rect 15752 17076 15804 17128
rect 16396 17076 16448 17128
rect 18420 17144 18472 17196
rect 19248 17144 19300 17196
rect 20904 17187 20956 17196
rect 20904 17153 20913 17187
rect 20913 17153 20947 17187
rect 20947 17153 20956 17187
rect 20904 17144 20956 17153
rect 22284 17144 22336 17196
rect 18788 17076 18840 17128
rect 20720 17119 20772 17128
rect 20720 17085 20729 17119
rect 20729 17085 20763 17119
rect 20763 17085 20772 17119
rect 20720 17076 20772 17085
rect 20812 17076 20864 17128
rect 22376 17076 22428 17128
rect 14740 17008 14792 17060
rect 17132 17051 17184 17060
rect 5356 16940 5408 16992
rect 8392 16983 8444 16992
rect 8392 16949 8401 16983
rect 8401 16949 8435 16983
rect 8435 16949 8444 16983
rect 8392 16940 8444 16949
rect 9220 16940 9272 16992
rect 11704 16940 11756 16992
rect 14372 16940 14424 16992
rect 15292 16940 15344 16992
rect 16028 16983 16080 16992
rect 16028 16949 16037 16983
rect 16037 16949 16071 16983
rect 16071 16949 16080 16983
rect 16028 16940 16080 16949
rect 17132 17017 17141 17051
rect 17141 17017 17175 17051
rect 17175 17017 17184 17051
rect 17132 17008 17184 17017
rect 17868 17008 17920 17060
rect 19708 17008 19760 17060
rect 20352 17008 20404 17060
rect 17592 16940 17644 16992
rect 17776 16940 17828 16992
rect 18052 16983 18104 16992
rect 18052 16949 18061 16983
rect 18061 16949 18095 16983
rect 18095 16949 18104 16983
rect 18052 16940 18104 16949
rect 18972 16940 19024 16992
rect 19248 16983 19300 16992
rect 19248 16949 19257 16983
rect 19257 16949 19291 16983
rect 19291 16949 19300 16983
rect 19248 16940 19300 16949
rect 22744 16940 22796 16992
rect 3790 16838 3842 16890
rect 3854 16838 3906 16890
rect 3918 16838 3970 16890
rect 3982 16838 4034 16890
rect 4046 16838 4098 16890
rect 9471 16838 9523 16890
rect 9535 16838 9587 16890
rect 9599 16838 9651 16890
rect 9663 16838 9715 16890
rect 9727 16838 9779 16890
rect 15152 16838 15204 16890
rect 15216 16838 15268 16890
rect 15280 16838 15332 16890
rect 15344 16838 15396 16890
rect 15408 16838 15460 16890
rect 20833 16838 20885 16890
rect 20897 16838 20949 16890
rect 20961 16838 21013 16890
rect 21025 16838 21077 16890
rect 21089 16838 21141 16890
rect 13268 16736 13320 16788
rect 14280 16736 14332 16788
rect 14832 16736 14884 16788
rect 14924 16736 14976 16788
rect 17316 16736 17368 16788
rect 18512 16736 18564 16788
rect 7104 16643 7156 16652
rect 7104 16609 7113 16643
rect 7113 16609 7147 16643
rect 7147 16609 7156 16643
rect 7104 16600 7156 16609
rect 8208 16600 8260 16652
rect 11796 16600 11848 16652
rect 12716 16600 12768 16652
rect 14096 16668 14148 16720
rect 2688 16532 2740 16584
rect 3056 16532 3108 16584
rect 8392 16532 8444 16584
rect 11888 16575 11940 16584
rect 11888 16541 11897 16575
rect 11897 16541 11931 16575
rect 11931 16541 11940 16575
rect 11888 16532 11940 16541
rect 12164 16532 12216 16584
rect 12992 16575 13044 16584
rect 12992 16541 13016 16575
rect 13016 16541 13044 16575
rect 12992 16532 13044 16541
rect 13084 16575 13136 16584
rect 13084 16541 13105 16575
rect 13105 16541 13136 16575
rect 13084 16532 13136 16541
rect 14188 16532 14240 16584
rect 14372 16575 14424 16584
rect 14372 16541 14381 16575
rect 14381 16541 14415 16575
rect 14415 16541 14424 16575
rect 14372 16532 14424 16541
rect 14740 16668 14792 16720
rect 15752 16668 15804 16720
rect 14648 16600 14700 16652
rect 16028 16668 16080 16720
rect 16304 16668 16356 16720
rect 17040 16668 17092 16720
rect 19248 16668 19300 16720
rect 20536 16668 20588 16720
rect 22376 16736 22428 16788
rect 22284 16668 22336 16720
rect 15660 16575 15712 16584
rect 2780 16464 2832 16516
rect 4896 16396 4948 16448
rect 5264 16439 5316 16448
rect 5264 16405 5273 16439
rect 5273 16405 5307 16439
rect 5307 16405 5316 16439
rect 5264 16396 5316 16405
rect 6460 16396 6512 16448
rect 8484 16439 8536 16448
rect 8484 16405 8493 16439
rect 8493 16405 8527 16439
rect 8527 16405 8536 16439
rect 8484 16396 8536 16405
rect 10692 16439 10744 16448
rect 10692 16405 10701 16439
rect 10701 16405 10735 16439
rect 10735 16405 10744 16439
rect 10692 16396 10744 16405
rect 12072 16439 12124 16448
rect 12072 16405 12081 16439
rect 12081 16405 12115 16439
rect 12115 16405 12124 16439
rect 12072 16396 12124 16405
rect 15660 16541 15669 16575
rect 15669 16541 15703 16575
rect 15703 16541 15712 16575
rect 15660 16532 15712 16541
rect 15844 16532 15896 16584
rect 17040 16532 17092 16584
rect 17408 16600 17460 16652
rect 17776 16643 17828 16652
rect 17776 16609 17785 16643
rect 17785 16609 17819 16643
rect 17819 16609 17828 16643
rect 17776 16600 17828 16609
rect 18328 16600 18380 16652
rect 18512 16600 18564 16652
rect 20352 16643 20404 16652
rect 20352 16609 20361 16643
rect 20361 16609 20395 16643
rect 20395 16609 20404 16643
rect 20352 16600 20404 16609
rect 14372 16396 14424 16448
rect 16948 16464 17000 16516
rect 17408 16507 17460 16516
rect 17408 16473 17417 16507
rect 17417 16473 17451 16507
rect 17451 16473 17460 16507
rect 17408 16464 17460 16473
rect 16672 16396 16724 16448
rect 18328 16464 18380 16516
rect 18788 16464 18840 16516
rect 20444 16532 20496 16584
rect 23296 16464 23348 16516
rect 17868 16396 17920 16448
rect 18880 16439 18932 16448
rect 18880 16405 18889 16439
rect 18889 16405 18923 16439
rect 18923 16405 18932 16439
rect 18880 16396 18932 16405
rect 20168 16396 20220 16448
rect 20996 16439 21048 16448
rect 20996 16405 21005 16439
rect 21005 16405 21039 16439
rect 21039 16405 21048 16439
rect 20996 16396 21048 16405
rect 22284 16396 22336 16448
rect 6630 16294 6682 16346
rect 6694 16294 6746 16346
rect 6758 16294 6810 16346
rect 6822 16294 6874 16346
rect 6886 16294 6938 16346
rect 12311 16294 12363 16346
rect 12375 16294 12427 16346
rect 12439 16294 12491 16346
rect 12503 16294 12555 16346
rect 12567 16294 12619 16346
rect 17992 16294 18044 16346
rect 18056 16294 18108 16346
rect 18120 16294 18172 16346
rect 18184 16294 18236 16346
rect 18248 16294 18300 16346
rect 23673 16294 23725 16346
rect 23737 16294 23789 16346
rect 23801 16294 23853 16346
rect 23865 16294 23917 16346
rect 23929 16294 23981 16346
rect 8208 16192 8260 16244
rect 9220 16192 9272 16244
rect 14740 16192 14792 16244
rect 18328 16235 18380 16244
rect 18328 16201 18337 16235
rect 18337 16201 18371 16235
rect 18371 16201 18380 16235
rect 18328 16192 18380 16201
rect 20260 16192 20312 16244
rect 4344 16167 4396 16176
rect 4344 16133 4353 16167
rect 4353 16133 4387 16167
rect 4387 16133 4396 16167
rect 4344 16124 4396 16133
rect 11704 16099 11756 16108
rect 11704 16065 11713 16099
rect 11713 16065 11747 16099
rect 11747 16065 11756 16099
rect 11704 16056 11756 16065
rect 11980 16099 12032 16108
rect 11980 16065 11989 16099
rect 11989 16065 12023 16099
rect 12023 16065 12032 16099
rect 11980 16056 12032 16065
rect 12164 15988 12216 16040
rect 14096 15988 14148 16040
rect 16488 15988 16540 16040
rect 17132 16124 17184 16176
rect 20168 16124 20220 16176
rect 20996 16192 21048 16244
rect 18420 16056 18472 16108
rect 19432 16056 19484 16108
rect 19616 16099 19668 16108
rect 19616 16065 19625 16099
rect 19625 16065 19659 16099
rect 19659 16065 19668 16099
rect 19616 16056 19668 16065
rect 19800 16099 19852 16108
rect 19800 16065 19809 16099
rect 19809 16065 19843 16099
rect 19843 16065 19852 16099
rect 19800 16056 19852 16065
rect 20812 16167 20864 16176
rect 20812 16133 20821 16167
rect 20821 16133 20855 16167
rect 20855 16133 20864 16167
rect 20812 16124 20864 16133
rect 20996 16099 21048 16108
rect 17592 15988 17644 16040
rect 19156 15988 19208 16040
rect 20996 16065 21005 16099
rect 21005 16065 21039 16099
rect 21039 16065 21048 16099
rect 20996 16056 21048 16065
rect 21824 16056 21876 16108
rect 21916 15988 21968 16040
rect 22560 15988 22612 16040
rect 2688 15920 2740 15972
rect 3148 15920 3200 15972
rect 12072 15920 12124 15972
rect 15568 15920 15620 15972
rect 17040 15920 17092 15972
rect 17776 15920 17828 15972
rect 21180 15920 21232 15972
rect 3056 15895 3108 15904
rect 3056 15861 3065 15895
rect 3065 15861 3099 15895
rect 3099 15861 3108 15895
rect 3056 15852 3108 15861
rect 13084 15852 13136 15904
rect 13912 15852 13964 15904
rect 15660 15895 15712 15904
rect 15660 15861 15669 15895
rect 15669 15861 15703 15895
rect 15703 15861 15712 15895
rect 15660 15852 15712 15861
rect 17132 15895 17184 15904
rect 17132 15861 17141 15895
rect 17141 15861 17175 15895
rect 17175 15861 17184 15895
rect 17132 15852 17184 15861
rect 19708 15852 19760 15904
rect 20996 15852 21048 15904
rect 21272 15852 21324 15904
rect 22652 15895 22704 15904
rect 22652 15861 22661 15895
rect 22661 15861 22695 15895
rect 22695 15861 22704 15895
rect 22652 15852 22704 15861
rect 3790 15750 3842 15802
rect 3854 15750 3906 15802
rect 3918 15750 3970 15802
rect 3982 15750 4034 15802
rect 4046 15750 4098 15802
rect 9471 15750 9523 15802
rect 9535 15750 9587 15802
rect 9599 15750 9651 15802
rect 9663 15750 9715 15802
rect 9727 15750 9779 15802
rect 15152 15750 15204 15802
rect 15216 15750 15268 15802
rect 15280 15750 15332 15802
rect 15344 15750 15396 15802
rect 15408 15750 15460 15802
rect 20833 15750 20885 15802
rect 20897 15750 20949 15802
rect 20961 15750 21013 15802
rect 21025 15750 21077 15802
rect 21089 15750 21141 15802
rect 13268 15648 13320 15700
rect 15016 15648 15068 15700
rect 10692 15580 10744 15632
rect 3056 15512 3108 15564
rect 8208 15512 8260 15564
rect 10140 15512 10192 15564
rect 2504 15487 2556 15496
rect 2504 15453 2513 15487
rect 2513 15453 2547 15487
rect 2547 15453 2556 15487
rect 2504 15444 2556 15453
rect 3700 15444 3752 15496
rect 11244 15487 11296 15496
rect 11244 15453 11253 15487
rect 11253 15453 11287 15487
rect 11287 15453 11296 15487
rect 11244 15444 11296 15453
rect 11428 15512 11480 15564
rect 15016 15512 15068 15564
rect 19248 15648 19300 15700
rect 19616 15648 19668 15700
rect 20352 15648 20404 15700
rect 22008 15648 22060 15700
rect 22744 15691 22796 15700
rect 22744 15657 22753 15691
rect 22753 15657 22787 15691
rect 22787 15657 22796 15691
rect 22744 15648 22796 15657
rect 16856 15580 16908 15632
rect 11796 15444 11848 15496
rect 11888 15444 11940 15496
rect 13544 15444 13596 15496
rect 13912 15444 13964 15496
rect 14740 15444 14792 15496
rect 15200 15444 15252 15496
rect 15660 15444 15712 15496
rect 16212 15444 16264 15496
rect 16672 15487 16724 15496
rect 16672 15453 16681 15487
rect 16681 15453 16715 15487
rect 16715 15453 16724 15487
rect 16672 15444 16724 15453
rect 18972 15580 19024 15632
rect 22560 15580 22612 15632
rect 18788 15512 18840 15564
rect 19892 15512 19944 15564
rect 19524 15444 19576 15496
rect 21364 15444 21416 15496
rect 22652 15444 22704 15496
rect 23020 15444 23072 15496
rect 2688 15376 2740 15428
rect 2228 15308 2280 15360
rect 3148 15308 3200 15360
rect 3332 15419 3384 15428
rect 3332 15385 3341 15419
rect 3341 15385 3375 15419
rect 3375 15385 3384 15419
rect 4252 15419 4304 15428
rect 3332 15376 3384 15385
rect 4252 15385 4261 15419
rect 4261 15385 4295 15419
rect 4295 15385 4304 15419
rect 4252 15376 4304 15385
rect 6552 15376 6604 15428
rect 12900 15419 12952 15428
rect 4528 15308 4580 15360
rect 7932 15308 7984 15360
rect 11152 15308 11204 15360
rect 12900 15385 12909 15419
rect 12909 15385 12943 15419
rect 12943 15385 12952 15419
rect 12900 15376 12952 15385
rect 16580 15376 16632 15428
rect 14740 15308 14792 15360
rect 16120 15308 16172 15360
rect 16396 15308 16448 15360
rect 16488 15308 16540 15360
rect 17408 15376 17460 15428
rect 19064 15376 19116 15428
rect 19800 15376 19852 15428
rect 20812 15419 20864 15428
rect 20812 15385 20821 15419
rect 20821 15385 20855 15419
rect 20855 15385 20864 15419
rect 20812 15376 20864 15385
rect 6630 15206 6682 15258
rect 6694 15206 6746 15258
rect 6758 15206 6810 15258
rect 6822 15206 6874 15258
rect 6886 15206 6938 15258
rect 12311 15206 12363 15258
rect 12375 15206 12427 15258
rect 12439 15206 12491 15258
rect 12503 15206 12555 15258
rect 12567 15206 12619 15258
rect 17992 15206 18044 15258
rect 18056 15206 18108 15258
rect 18120 15206 18172 15258
rect 18184 15206 18236 15258
rect 18248 15206 18300 15258
rect 23673 15206 23725 15258
rect 23737 15206 23789 15258
rect 23801 15206 23853 15258
rect 23865 15206 23917 15258
rect 23929 15206 23981 15258
rect 3240 15104 3292 15156
rect 3424 15104 3476 15156
rect 6276 15104 6328 15156
rect 1860 15079 1912 15088
rect 1860 15045 1869 15079
rect 1869 15045 1903 15079
rect 1903 15045 1912 15079
rect 1860 15036 1912 15045
rect 2136 15036 2188 15088
rect 4160 15036 4212 15088
rect 5264 15036 5316 15088
rect 1768 15011 1820 15020
rect 1768 14977 1777 15011
rect 1777 14977 1811 15011
rect 1811 14977 1820 15011
rect 1768 14968 1820 14977
rect 2320 14968 2372 15020
rect 3056 14968 3108 15020
rect 4988 15011 5040 15020
rect 4988 14977 4997 15011
rect 4997 14977 5031 15011
rect 5031 14977 5040 15011
rect 4988 14968 5040 14977
rect 4620 14900 4672 14952
rect 4988 14832 5040 14884
rect 5632 14968 5684 15020
rect 11888 15104 11940 15156
rect 15476 15104 15528 15156
rect 16488 15104 16540 15156
rect 19248 15104 19300 15156
rect 22468 15104 22520 15156
rect 11796 15036 11848 15088
rect 12900 15036 12952 15088
rect 8208 14968 8260 15020
rect 12624 14968 12676 15020
rect 13084 15011 13136 15020
rect 13084 14977 13093 15011
rect 13093 14977 13127 15011
rect 13127 14977 13136 15011
rect 13084 14968 13136 14977
rect 13268 15011 13320 15020
rect 13268 14977 13277 15011
rect 13277 14977 13311 15011
rect 13311 14977 13320 15011
rect 13268 14968 13320 14977
rect 18512 15036 18564 15088
rect 19340 15079 19392 15088
rect 19340 15045 19349 15079
rect 19349 15045 19383 15079
rect 19383 15045 19392 15079
rect 19340 15036 19392 15045
rect 14924 14968 14976 15020
rect 15568 15011 15620 15020
rect 15568 14977 15577 15011
rect 15577 14977 15611 15011
rect 15611 14977 15620 15011
rect 15568 14968 15620 14977
rect 7840 14900 7892 14952
rect 12900 14900 12952 14952
rect 14188 14900 14240 14952
rect 6184 14832 6236 14884
rect 6644 14832 6696 14884
rect 11796 14832 11848 14884
rect 13544 14832 13596 14884
rect 14832 14875 14884 14884
rect 14832 14841 14841 14875
rect 14841 14841 14875 14875
rect 14875 14841 14884 14875
rect 14832 14832 14884 14841
rect 15200 14900 15252 14952
rect 16948 14968 17000 15020
rect 19248 14968 19300 15020
rect 19800 15011 19852 15020
rect 16580 14900 16632 14952
rect 17316 14900 17368 14952
rect 18328 14900 18380 14952
rect 16304 14832 16356 14884
rect 2872 14764 2924 14816
rect 3148 14764 3200 14816
rect 3424 14764 3476 14816
rect 6000 14764 6052 14816
rect 6092 14764 6144 14816
rect 7656 14764 7708 14816
rect 13360 14764 13412 14816
rect 16212 14764 16264 14816
rect 18788 14764 18840 14816
rect 19800 14977 19809 15011
rect 19809 14977 19843 15011
rect 19843 14977 19852 15011
rect 19800 14968 19852 14977
rect 19892 15011 19944 15020
rect 19892 14977 19901 15011
rect 19901 14977 19935 15011
rect 19935 14977 19944 15011
rect 19892 14968 19944 14977
rect 20260 14968 20312 15020
rect 21180 14968 21232 15020
rect 22008 15011 22060 15020
rect 22008 14977 22017 15011
rect 22017 14977 22051 15011
rect 22051 14977 22060 15011
rect 22008 14968 22060 14977
rect 22100 15011 22152 15020
rect 22100 14977 22110 15011
rect 22110 14977 22144 15011
rect 22144 14977 22152 15011
rect 22284 15011 22336 15020
rect 22100 14968 22152 14977
rect 22284 14977 22293 15011
rect 22293 14977 22327 15011
rect 22327 14977 22336 15011
rect 22284 14968 22336 14977
rect 20812 14900 20864 14952
rect 21364 14832 21416 14884
rect 22284 14832 22336 14884
rect 22836 14968 22888 15020
rect 21824 14764 21876 14816
rect 23112 14807 23164 14816
rect 23112 14773 23121 14807
rect 23121 14773 23155 14807
rect 23155 14773 23164 14807
rect 23112 14764 23164 14773
rect 3790 14662 3842 14714
rect 3854 14662 3906 14714
rect 3918 14662 3970 14714
rect 3982 14662 4034 14714
rect 4046 14662 4098 14714
rect 9471 14662 9523 14714
rect 9535 14662 9587 14714
rect 9599 14662 9651 14714
rect 9663 14662 9715 14714
rect 9727 14662 9779 14714
rect 15152 14662 15204 14714
rect 15216 14662 15268 14714
rect 15280 14662 15332 14714
rect 15344 14662 15396 14714
rect 15408 14662 15460 14714
rect 20833 14662 20885 14714
rect 20897 14662 20949 14714
rect 20961 14662 21013 14714
rect 21025 14662 21077 14714
rect 21089 14662 21141 14714
rect 1676 14560 1728 14612
rect 4712 14603 4764 14612
rect 2228 14399 2280 14408
rect 2228 14365 2237 14399
rect 2237 14365 2271 14399
rect 2271 14365 2280 14399
rect 2228 14356 2280 14365
rect 2320 14356 2372 14408
rect 2688 14356 2740 14408
rect 4252 14492 4304 14544
rect 3240 14424 3292 14476
rect 3516 14424 3568 14476
rect 4712 14569 4721 14603
rect 4721 14569 4755 14603
rect 4755 14569 4764 14603
rect 4712 14560 4764 14569
rect 4620 14492 4672 14544
rect 6552 14560 6604 14612
rect 8300 14560 8352 14612
rect 12808 14560 12860 14612
rect 13820 14560 13872 14612
rect 6000 14492 6052 14544
rect 6092 14424 6144 14476
rect 7196 14492 7248 14544
rect 9312 14492 9364 14544
rect 10508 14492 10560 14544
rect 1952 14288 2004 14340
rect 3240 14331 3292 14340
rect 3240 14297 3249 14331
rect 3249 14297 3283 14331
rect 3283 14297 3292 14331
rect 4620 14356 4672 14408
rect 5264 14356 5316 14408
rect 5448 14356 5500 14408
rect 7288 14424 7340 14476
rect 11888 14492 11940 14544
rect 11060 14467 11112 14476
rect 7012 14399 7064 14408
rect 7012 14365 7021 14399
rect 7021 14365 7055 14399
rect 7055 14365 7064 14399
rect 7012 14356 7064 14365
rect 7380 14399 7432 14408
rect 7380 14365 7389 14399
rect 7389 14365 7423 14399
rect 7423 14365 7432 14399
rect 7380 14356 7432 14365
rect 7932 14399 7984 14408
rect 7932 14365 7941 14399
rect 7941 14365 7975 14399
rect 7975 14365 7984 14399
rect 7932 14356 7984 14365
rect 3240 14288 3292 14297
rect 3516 14288 3568 14340
rect 6092 14331 6144 14340
rect 6092 14297 6101 14331
rect 6101 14297 6135 14331
rect 6135 14297 6144 14331
rect 6092 14288 6144 14297
rect 6184 14331 6236 14340
rect 6184 14297 6193 14331
rect 6193 14297 6227 14331
rect 6227 14297 6236 14331
rect 6184 14288 6236 14297
rect 8300 14288 8352 14340
rect 11060 14433 11069 14467
rect 11069 14433 11103 14467
rect 11103 14433 11112 14467
rect 11060 14424 11112 14433
rect 13360 14492 13412 14544
rect 14924 14560 14976 14612
rect 17408 14560 17460 14612
rect 19340 14560 19392 14612
rect 15200 14492 15252 14544
rect 16396 14492 16448 14544
rect 19708 14492 19760 14544
rect 20352 14560 20404 14612
rect 20720 14560 20772 14612
rect 21272 14492 21324 14544
rect 12348 14467 12400 14476
rect 12348 14433 12357 14467
rect 12357 14433 12391 14467
rect 12391 14433 12400 14467
rect 12348 14424 12400 14433
rect 12716 14424 12768 14476
rect 14188 14424 14240 14476
rect 9312 14399 9364 14408
rect 9312 14365 9321 14399
rect 9321 14365 9355 14399
rect 9355 14365 9364 14399
rect 9312 14356 9364 14365
rect 9680 14399 9732 14408
rect 9680 14365 9689 14399
rect 9689 14365 9723 14399
rect 9723 14365 9732 14399
rect 9680 14356 9732 14365
rect 9404 14331 9456 14340
rect 2872 14263 2924 14272
rect 2872 14229 2881 14263
rect 2881 14229 2915 14263
rect 2915 14229 2924 14263
rect 2872 14220 2924 14229
rect 7012 14220 7064 14272
rect 9404 14297 9413 14331
rect 9413 14297 9447 14331
rect 9447 14297 9456 14331
rect 9404 14288 9456 14297
rect 11152 14331 11204 14340
rect 9220 14220 9272 14272
rect 11152 14297 11161 14331
rect 11161 14297 11195 14331
rect 11195 14297 11204 14331
rect 11152 14288 11204 14297
rect 11796 14288 11848 14340
rect 12808 14356 12860 14408
rect 13544 14356 13596 14408
rect 14280 14399 14332 14408
rect 14280 14365 14289 14399
rect 14289 14365 14323 14399
rect 14323 14365 14332 14399
rect 14280 14356 14332 14365
rect 14556 14399 14608 14408
rect 13360 14288 13412 14340
rect 14004 14288 14056 14340
rect 14188 14288 14240 14340
rect 14556 14365 14565 14399
rect 14565 14365 14599 14399
rect 14599 14365 14608 14399
rect 14556 14356 14608 14365
rect 15384 14424 15436 14476
rect 16212 14467 16264 14476
rect 16212 14433 16221 14467
rect 16221 14433 16255 14467
rect 16255 14433 16264 14467
rect 16212 14424 16264 14433
rect 17132 14424 17184 14476
rect 15936 14356 15988 14408
rect 16764 14356 16816 14408
rect 17316 14399 17368 14408
rect 17316 14365 17325 14399
rect 17325 14365 17359 14399
rect 17359 14365 17368 14399
rect 17316 14356 17368 14365
rect 17408 14399 17460 14408
rect 17408 14365 17417 14399
rect 17417 14365 17451 14399
rect 17451 14365 17460 14399
rect 17408 14356 17460 14365
rect 19340 14356 19392 14408
rect 19616 14399 19668 14408
rect 19616 14365 19625 14399
rect 19625 14365 19659 14399
rect 19659 14365 19668 14399
rect 19616 14356 19668 14365
rect 14648 14331 14700 14340
rect 14648 14297 14657 14331
rect 14657 14297 14691 14331
rect 14691 14297 14700 14331
rect 14648 14288 14700 14297
rect 15476 14288 15528 14340
rect 11336 14220 11388 14272
rect 15384 14220 15436 14272
rect 15660 14263 15712 14272
rect 15660 14229 15669 14263
rect 15669 14229 15703 14263
rect 15703 14229 15712 14263
rect 15660 14220 15712 14229
rect 16120 14263 16172 14272
rect 16120 14229 16129 14263
rect 16129 14229 16163 14263
rect 16163 14229 16172 14263
rect 16120 14220 16172 14229
rect 19156 14288 19208 14340
rect 21456 14356 21508 14408
rect 21732 14399 21784 14408
rect 21732 14365 21741 14399
rect 21741 14365 21775 14399
rect 21775 14365 21784 14399
rect 21732 14356 21784 14365
rect 22100 14356 22152 14408
rect 22836 14399 22888 14408
rect 22836 14365 22845 14399
rect 22845 14365 22879 14399
rect 22879 14365 22888 14399
rect 22836 14356 22888 14365
rect 20076 14288 20128 14340
rect 17224 14220 17276 14272
rect 18696 14220 18748 14272
rect 20260 14220 20312 14272
rect 22468 14220 22520 14272
rect 22928 14220 22980 14272
rect 6630 14118 6682 14170
rect 6694 14118 6746 14170
rect 6758 14118 6810 14170
rect 6822 14118 6874 14170
rect 6886 14118 6938 14170
rect 12311 14118 12363 14170
rect 12375 14118 12427 14170
rect 12439 14118 12491 14170
rect 12503 14118 12555 14170
rect 12567 14118 12619 14170
rect 17992 14118 18044 14170
rect 18056 14118 18108 14170
rect 18120 14118 18172 14170
rect 18184 14118 18236 14170
rect 18248 14118 18300 14170
rect 23673 14118 23725 14170
rect 23737 14118 23789 14170
rect 23801 14118 23853 14170
rect 23865 14118 23917 14170
rect 23929 14118 23981 14170
rect 3056 14016 3108 14068
rect 3700 14016 3752 14068
rect 5080 14059 5132 14068
rect 5080 14025 5089 14059
rect 5089 14025 5123 14059
rect 5123 14025 5132 14059
rect 5080 14016 5132 14025
rect 10140 14016 10192 14068
rect 12808 14059 12860 14068
rect 12808 14025 12817 14059
rect 12817 14025 12851 14059
rect 12851 14025 12860 14059
rect 12808 14016 12860 14025
rect 16120 14016 16172 14068
rect 16948 14016 17000 14068
rect 17408 14016 17460 14068
rect 2872 13991 2924 14000
rect 2872 13957 2906 13991
rect 2906 13957 2924 13991
rect 2872 13948 2924 13957
rect 2504 13880 2556 13932
rect 13084 13948 13136 14000
rect 5448 13923 5500 13932
rect 5448 13889 5457 13923
rect 5457 13889 5491 13923
rect 5491 13889 5500 13923
rect 5448 13880 5500 13889
rect 6184 13880 6236 13932
rect 8208 13923 8260 13932
rect 8208 13889 8217 13923
rect 8217 13889 8251 13923
rect 8251 13889 8260 13923
rect 8208 13880 8260 13889
rect 1860 13855 1912 13864
rect 1860 13821 1869 13855
rect 1869 13821 1903 13855
rect 1903 13821 1912 13855
rect 1860 13812 1912 13821
rect 5356 13812 5408 13864
rect 5908 13812 5960 13864
rect 7840 13812 7892 13864
rect 9680 13880 9732 13932
rect 10048 13923 10100 13932
rect 10048 13889 10057 13923
rect 10057 13889 10091 13923
rect 10091 13889 10100 13923
rect 10048 13880 10100 13889
rect 10692 13880 10744 13932
rect 10784 13880 10836 13932
rect 12716 13880 12768 13932
rect 14464 13880 14516 13932
rect 15200 13948 15252 14000
rect 15844 13991 15896 14000
rect 15844 13957 15853 13991
rect 15853 13957 15887 13991
rect 15887 13957 15896 13991
rect 15844 13948 15896 13957
rect 16028 13948 16080 14000
rect 11796 13855 11848 13864
rect 11796 13821 11805 13855
rect 11805 13821 11839 13855
rect 11839 13821 11848 13855
rect 11796 13812 11848 13821
rect 14280 13812 14332 13864
rect 14924 13923 14976 13932
rect 14924 13889 14933 13923
rect 14933 13889 14967 13923
rect 14967 13889 14976 13923
rect 15752 13923 15804 13932
rect 14924 13880 14976 13889
rect 15752 13889 15761 13923
rect 15761 13889 15795 13923
rect 15795 13889 15804 13923
rect 15752 13880 15804 13889
rect 15936 13923 15988 13932
rect 15936 13889 15945 13923
rect 15945 13889 15979 13923
rect 15979 13889 15988 13923
rect 15936 13880 15988 13889
rect 16948 13880 17000 13932
rect 15660 13812 15712 13864
rect 17960 13923 18012 13932
rect 17960 13889 17969 13923
rect 17969 13889 18003 13923
rect 18003 13889 18012 13923
rect 19800 14016 19852 14068
rect 17960 13880 18012 13889
rect 18236 13923 18288 13932
rect 18236 13889 18245 13923
rect 18245 13889 18279 13923
rect 18279 13889 18288 13923
rect 18236 13880 18288 13889
rect 20260 13880 20312 13932
rect 21456 14016 21508 14068
rect 19156 13812 19208 13864
rect 2320 13744 2372 13796
rect 17684 13787 17736 13796
rect 17684 13753 17693 13787
rect 17693 13753 17727 13787
rect 17727 13753 17736 13787
rect 17684 13744 17736 13753
rect 2044 13719 2096 13728
rect 2044 13685 2053 13719
rect 2053 13685 2087 13719
rect 2087 13685 2096 13719
rect 2044 13676 2096 13685
rect 3700 13676 3752 13728
rect 5724 13676 5776 13728
rect 7012 13676 7064 13728
rect 10324 13676 10376 13728
rect 11612 13676 11664 13728
rect 14096 13719 14148 13728
rect 14096 13685 14105 13719
rect 14105 13685 14139 13719
rect 14139 13685 14148 13719
rect 14096 13676 14148 13685
rect 15476 13676 15528 13728
rect 15660 13676 15712 13728
rect 18880 13676 18932 13728
rect 19524 13855 19576 13864
rect 19524 13821 19533 13855
rect 19533 13821 19567 13855
rect 19567 13821 19576 13855
rect 19524 13812 19576 13821
rect 20812 13889 20821 13898
rect 20821 13889 20855 13898
rect 20855 13889 20864 13898
rect 20812 13846 20864 13889
rect 20996 13923 21048 13932
rect 20996 13889 20999 13923
rect 20999 13889 21033 13923
rect 21033 13889 21048 13923
rect 20996 13880 21048 13889
rect 21640 13880 21692 13932
rect 22744 13948 22796 14000
rect 22284 13923 22336 13932
rect 22284 13889 22293 13923
rect 22293 13889 22327 13923
rect 22327 13889 22336 13923
rect 22284 13880 22336 13889
rect 22560 13923 22612 13932
rect 22560 13889 22569 13923
rect 22569 13889 22603 13923
rect 22603 13889 22612 13923
rect 22560 13880 22612 13889
rect 21824 13744 21876 13796
rect 23112 13880 23164 13932
rect 23388 13744 23440 13796
rect 19984 13676 20036 13728
rect 22284 13676 22336 13728
rect 3790 13574 3842 13626
rect 3854 13574 3906 13626
rect 3918 13574 3970 13626
rect 3982 13574 4034 13626
rect 4046 13574 4098 13626
rect 9471 13574 9523 13626
rect 9535 13574 9587 13626
rect 9599 13574 9651 13626
rect 9663 13574 9715 13626
rect 9727 13574 9779 13626
rect 15152 13574 15204 13626
rect 15216 13574 15268 13626
rect 15280 13574 15332 13626
rect 15344 13574 15396 13626
rect 15408 13574 15460 13626
rect 20833 13574 20885 13626
rect 20897 13574 20949 13626
rect 20961 13574 21013 13626
rect 21025 13574 21077 13626
rect 21089 13574 21141 13626
rect 2504 13472 2556 13524
rect 3700 13404 3752 13456
rect 3516 13336 3568 13388
rect 4252 13336 4304 13388
rect 2320 13311 2372 13320
rect 2320 13277 2329 13311
rect 2329 13277 2363 13311
rect 2363 13277 2372 13311
rect 2320 13268 2372 13277
rect 2688 13268 2740 13320
rect 4620 13515 4672 13524
rect 4620 13481 4629 13515
rect 4629 13481 4663 13515
rect 4663 13481 4672 13515
rect 4620 13472 4672 13481
rect 4988 13472 5040 13524
rect 6184 13472 6236 13524
rect 11336 13472 11388 13524
rect 15752 13472 15804 13524
rect 17316 13472 17368 13524
rect 19616 13472 19668 13524
rect 19708 13472 19760 13524
rect 19800 13472 19852 13524
rect 21456 13515 21508 13524
rect 21456 13481 21465 13515
rect 21465 13481 21499 13515
rect 21499 13481 21508 13515
rect 21456 13472 21508 13481
rect 4528 13404 4580 13456
rect 7104 13404 7156 13456
rect 10048 13404 10100 13456
rect 5448 13336 5500 13388
rect 6276 13336 6328 13388
rect 10324 13379 10376 13388
rect 5172 13311 5224 13320
rect 5172 13277 5181 13311
rect 5181 13277 5215 13311
rect 5215 13277 5224 13311
rect 5172 13268 5224 13277
rect 5264 13268 5316 13320
rect 10324 13345 10333 13379
rect 10333 13345 10367 13379
rect 10367 13345 10376 13379
rect 10324 13336 10376 13345
rect 2780 13200 2832 13252
rect 3516 13200 3568 13252
rect 3976 13200 4028 13252
rect 4252 13243 4304 13252
rect 4252 13209 4261 13243
rect 4261 13209 4295 13243
rect 4295 13209 4304 13243
rect 4252 13200 4304 13209
rect 4344 13200 4396 13252
rect 6552 13200 6604 13252
rect 10140 13200 10192 13252
rect 10692 13311 10744 13320
rect 10692 13277 10701 13311
rect 10701 13277 10735 13311
rect 10735 13277 10744 13311
rect 10692 13268 10744 13277
rect 13360 13404 13412 13456
rect 16028 13404 16080 13456
rect 14740 13336 14792 13388
rect 11704 13268 11756 13320
rect 12072 13268 12124 13320
rect 14280 13311 14332 13320
rect 14280 13277 14289 13311
rect 14289 13277 14323 13311
rect 14323 13277 14332 13311
rect 14280 13268 14332 13277
rect 14464 13268 14516 13320
rect 14648 13268 14700 13320
rect 15292 13311 15344 13320
rect 15292 13277 15301 13311
rect 15301 13277 15335 13311
rect 15335 13277 15344 13311
rect 15292 13268 15344 13277
rect 15476 13311 15528 13320
rect 15476 13277 15485 13311
rect 15485 13277 15519 13311
rect 15519 13277 15528 13311
rect 15476 13268 15528 13277
rect 16948 13336 17000 13388
rect 16856 13268 16908 13320
rect 18420 13404 18472 13456
rect 3332 13132 3384 13184
rect 5264 13132 5316 13184
rect 7196 13175 7248 13184
rect 7196 13141 7205 13175
rect 7205 13141 7239 13175
rect 7239 13141 7248 13175
rect 7196 13132 7248 13141
rect 7748 13132 7800 13184
rect 11888 13132 11940 13184
rect 12992 13200 13044 13252
rect 15844 13200 15896 13252
rect 16580 13200 16632 13252
rect 16764 13200 16816 13252
rect 17960 13336 18012 13388
rect 18788 13336 18840 13388
rect 19524 13336 19576 13388
rect 17592 13268 17644 13320
rect 19248 13268 19300 13320
rect 20904 13336 20956 13388
rect 21548 13336 21600 13388
rect 22100 13336 22152 13388
rect 14004 13132 14056 13184
rect 14556 13132 14608 13184
rect 14648 13175 14700 13184
rect 14648 13141 14657 13175
rect 14657 13141 14691 13175
rect 14691 13141 14700 13175
rect 14648 13132 14700 13141
rect 15292 13132 15344 13184
rect 15476 13132 15528 13184
rect 16120 13132 16172 13184
rect 16304 13132 16356 13184
rect 19156 13200 19208 13252
rect 17776 13132 17828 13184
rect 18880 13175 18932 13184
rect 18880 13141 18889 13175
rect 18889 13141 18923 13175
rect 18923 13141 18932 13175
rect 18880 13132 18932 13141
rect 19616 13200 19668 13252
rect 19984 13200 20036 13252
rect 20352 13200 20404 13252
rect 22468 13268 22520 13320
rect 22928 13200 22980 13252
rect 23112 13200 23164 13252
rect 22652 13132 22704 13184
rect 6630 13030 6682 13082
rect 6694 13030 6746 13082
rect 6758 13030 6810 13082
rect 6822 13030 6874 13082
rect 6886 13030 6938 13082
rect 12311 13030 12363 13082
rect 12375 13030 12427 13082
rect 12439 13030 12491 13082
rect 12503 13030 12555 13082
rect 12567 13030 12619 13082
rect 17992 13030 18044 13082
rect 18056 13030 18108 13082
rect 18120 13030 18172 13082
rect 18184 13030 18236 13082
rect 18248 13030 18300 13082
rect 23673 13030 23725 13082
rect 23737 13030 23789 13082
rect 23801 13030 23853 13082
rect 23865 13030 23917 13082
rect 23929 13030 23981 13082
rect 2044 12928 2096 12980
rect 4344 12928 4396 12980
rect 6552 12928 6604 12980
rect 7840 12928 7892 12980
rect 9220 12928 9272 12980
rect 11888 12928 11940 12980
rect 2596 12903 2648 12912
rect 2596 12869 2605 12903
rect 2605 12869 2639 12903
rect 2639 12869 2648 12903
rect 2596 12860 2648 12869
rect 2780 12860 2832 12912
rect 3976 12903 4028 12912
rect 3976 12869 3985 12903
rect 3985 12869 4019 12903
rect 4019 12869 4028 12903
rect 3976 12860 4028 12869
rect 2688 12792 2740 12844
rect 3332 12792 3384 12844
rect 4988 12860 5040 12912
rect 4252 12792 4304 12844
rect 7748 12860 7800 12912
rect 8668 12860 8720 12912
rect 10140 12860 10192 12912
rect 5264 12835 5316 12844
rect 5264 12801 5273 12835
rect 5273 12801 5307 12835
rect 5307 12801 5316 12835
rect 5264 12792 5316 12801
rect 5632 12792 5684 12844
rect 6000 12792 6052 12844
rect 7564 12835 7616 12844
rect 7564 12801 7573 12835
rect 7573 12801 7607 12835
rect 7607 12801 7616 12835
rect 7564 12792 7616 12801
rect 8116 12835 8168 12844
rect 8116 12801 8125 12835
rect 8125 12801 8159 12835
rect 8159 12801 8168 12835
rect 8116 12792 8168 12801
rect 8300 12835 8352 12844
rect 8300 12801 8309 12835
rect 8309 12801 8343 12835
rect 8343 12801 8352 12835
rect 8300 12792 8352 12801
rect 8944 12835 8996 12844
rect 8944 12801 8953 12835
rect 8953 12801 8987 12835
rect 8987 12801 8996 12835
rect 8944 12792 8996 12801
rect 9036 12835 9088 12844
rect 9036 12801 9045 12835
rect 9045 12801 9079 12835
rect 9079 12801 9088 12835
rect 9312 12835 9364 12844
rect 9036 12792 9088 12801
rect 9312 12801 9321 12835
rect 9321 12801 9355 12835
rect 9355 12801 9364 12835
rect 9312 12792 9364 12801
rect 10416 12835 10468 12844
rect 10416 12801 10425 12835
rect 10425 12801 10459 12835
rect 10459 12801 10468 12835
rect 10416 12792 10468 12801
rect 11704 12860 11756 12912
rect 11796 12792 11848 12844
rect 12072 12860 12124 12912
rect 11980 12792 12032 12844
rect 12716 12860 12768 12912
rect 13360 12860 13412 12912
rect 12900 12792 12952 12844
rect 13176 12792 13228 12844
rect 14740 12860 14792 12912
rect 15660 12860 15712 12912
rect 17224 12903 17276 12912
rect 17224 12869 17233 12903
rect 17233 12869 17267 12903
rect 17267 12869 17276 12903
rect 17224 12860 17276 12869
rect 3424 12656 3476 12708
rect 1952 12588 2004 12640
rect 2596 12588 2648 12640
rect 5448 12656 5500 12708
rect 7104 12699 7156 12708
rect 7104 12665 7113 12699
rect 7113 12665 7147 12699
rect 7147 12665 7156 12699
rect 8852 12724 8904 12776
rect 7104 12656 7156 12665
rect 4252 12588 4304 12640
rect 5724 12588 5776 12640
rect 7012 12588 7064 12640
rect 7840 12656 7892 12708
rect 11152 12767 11204 12776
rect 11152 12733 11161 12767
rect 11161 12733 11195 12767
rect 11195 12733 11204 12767
rect 11152 12724 11204 12733
rect 13728 12767 13780 12776
rect 13728 12733 13737 12767
rect 13737 12733 13771 12767
rect 13771 12733 13780 12767
rect 13728 12724 13780 12733
rect 14096 12724 14148 12776
rect 15660 12724 15712 12776
rect 15936 12767 15988 12776
rect 15936 12733 15945 12767
rect 15945 12733 15979 12767
rect 15979 12733 15988 12767
rect 15936 12724 15988 12733
rect 16120 12767 16172 12776
rect 16120 12733 16129 12767
rect 16129 12733 16163 12767
rect 16163 12733 16172 12767
rect 16948 12835 17000 12844
rect 16948 12801 16958 12835
rect 16958 12801 16992 12835
rect 16992 12801 17000 12835
rect 17132 12835 17184 12844
rect 16948 12792 17000 12801
rect 17132 12801 17141 12835
rect 17141 12801 17175 12835
rect 17175 12801 17184 12835
rect 17132 12792 17184 12801
rect 17684 12928 17736 12980
rect 19340 12928 19392 12980
rect 17592 12860 17644 12912
rect 19984 12928 20036 12980
rect 20260 12928 20312 12980
rect 22284 12971 22336 12980
rect 17868 12792 17920 12844
rect 19340 12792 19392 12844
rect 21364 12860 21416 12912
rect 19892 12835 19944 12844
rect 19892 12801 19901 12835
rect 19901 12801 19935 12835
rect 19935 12801 19944 12835
rect 19892 12792 19944 12801
rect 20260 12792 20312 12844
rect 20352 12792 20404 12844
rect 20628 12792 20680 12844
rect 20720 12792 20772 12844
rect 21272 12792 21324 12844
rect 21732 12860 21784 12912
rect 22284 12937 22293 12971
rect 22293 12937 22327 12971
rect 22327 12937 22336 12971
rect 22284 12928 22336 12937
rect 22744 12903 22796 12912
rect 22744 12869 22779 12903
rect 22779 12869 22796 12903
rect 22744 12860 22796 12869
rect 16120 12724 16172 12733
rect 22100 12724 22152 12776
rect 16672 12656 16724 12708
rect 8024 12588 8076 12640
rect 8760 12631 8812 12640
rect 8760 12597 8769 12631
rect 8769 12597 8803 12631
rect 8803 12597 8812 12631
rect 8760 12588 8812 12597
rect 11796 12588 11848 12640
rect 12532 12588 12584 12640
rect 16856 12588 16908 12640
rect 17592 12588 17644 12640
rect 18512 12656 18564 12708
rect 19800 12699 19852 12708
rect 19800 12665 19809 12699
rect 19809 12665 19843 12699
rect 19843 12665 19852 12699
rect 19800 12656 19852 12665
rect 18604 12631 18656 12640
rect 18604 12597 18613 12631
rect 18613 12597 18647 12631
rect 18647 12597 18656 12631
rect 18604 12588 18656 12597
rect 19340 12588 19392 12640
rect 20628 12588 20680 12640
rect 22652 12835 22704 12844
rect 22652 12801 22661 12835
rect 22661 12801 22695 12835
rect 22695 12801 22704 12835
rect 22928 12835 22980 12844
rect 22652 12792 22704 12801
rect 22928 12801 22937 12835
rect 22937 12801 22971 12835
rect 22971 12801 22980 12835
rect 22928 12792 22980 12801
rect 23020 12656 23072 12708
rect 22744 12588 22796 12640
rect 3790 12486 3842 12538
rect 3854 12486 3906 12538
rect 3918 12486 3970 12538
rect 3982 12486 4034 12538
rect 4046 12486 4098 12538
rect 9471 12486 9523 12538
rect 9535 12486 9587 12538
rect 9599 12486 9651 12538
rect 9663 12486 9715 12538
rect 9727 12486 9779 12538
rect 15152 12486 15204 12538
rect 15216 12486 15268 12538
rect 15280 12486 15332 12538
rect 15344 12486 15396 12538
rect 15408 12486 15460 12538
rect 20833 12486 20885 12538
rect 20897 12486 20949 12538
rect 20961 12486 21013 12538
rect 21025 12486 21077 12538
rect 21089 12486 21141 12538
rect 1584 12384 1636 12436
rect 2044 12316 2096 12368
rect 4160 12384 4212 12436
rect 5632 12384 5684 12436
rect 7196 12384 7248 12436
rect 7380 12427 7432 12436
rect 7380 12393 7389 12427
rect 7389 12393 7423 12427
rect 7423 12393 7432 12427
rect 7380 12384 7432 12393
rect 7564 12384 7616 12436
rect 10692 12384 10744 12436
rect 10968 12384 11020 12436
rect 11980 12427 12032 12436
rect 11980 12393 11989 12427
rect 11989 12393 12023 12427
rect 12023 12393 12032 12427
rect 11980 12384 12032 12393
rect 12164 12384 12216 12436
rect 15476 12384 15528 12436
rect 16304 12427 16356 12436
rect 16304 12393 16313 12427
rect 16313 12393 16347 12427
rect 16347 12393 16356 12427
rect 16304 12384 16356 12393
rect 18972 12384 19024 12436
rect 19156 12384 19208 12436
rect 20352 12384 20404 12436
rect 2136 12180 2188 12232
rect 2320 12180 2372 12232
rect 2596 12248 2648 12300
rect 7288 12316 7340 12368
rect 8208 12316 8260 12368
rect 12532 12359 12584 12368
rect 12532 12325 12541 12359
rect 12541 12325 12575 12359
rect 12575 12325 12584 12359
rect 12532 12316 12584 12325
rect 13176 12316 13228 12368
rect 15568 12316 15620 12368
rect 6276 12248 6328 12300
rect 1952 12112 2004 12164
rect 1676 12044 1728 12096
rect 2228 12044 2280 12096
rect 3700 12180 3752 12232
rect 4160 12223 4212 12232
rect 4160 12189 4169 12223
rect 4169 12189 4203 12223
rect 4203 12189 4212 12223
rect 6552 12223 6604 12232
rect 4160 12180 4212 12189
rect 3332 12112 3384 12164
rect 6552 12189 6561 12223
rect 6561 12189 6595 12223
rect 6595 12189 6604 12223
rect 6552 12180 6604 12189
rect 8300 12248 8352 12300
rect 7196 12223 7248 12232
rect 7196 12189 7205 12223
rect 7205 12189 7239 12223
rect 7239 12189 7248 12223
rect 7196 12180 7248 12189
rect 7012 12112 7064 12164
rect 8208 12180 8260 12232
rect 10784 12248 10836 12300
rect 10508 12180 10560 12232
rect 10692 12223 10744 12232
rect 10692 12189 10701 12223
rect 10701 12189 10735 12223
rect 10735 12189 10744 12223
rect 10692 12180 10744 12189
rect 12072 12248 12124 12300
rect 13268 12248 13320 12300
rect 14372 12248 14424 12300
rect 15016 12248 15068 12300
rect 21272 12316 21324 12368
rect 21640 12316 21692 12368
rect 7840 12112 7892 12164
rect 11888 12112 11940 12164
rect 14004 12180 14056 12232
rect 14280 12223 14332 12232
rect 14280 12189 14289 12223
rect 14289 12189 14323 12223
rect 14323 12189 14332 12223
rect 14280 12180 14332 12189
rect 14740 12180 14792 12232
rect 16028 12112 16080 12164
rect 16120 12155 16172 12164
rect 16120 12121 16129 12155
rect 16129 12121 16163 12155
rect 16163 12121 16172 12155
rect 16856 12180 16908 12232
rect 17960 12248 18012 12300
rect 19708 12248 19760 12300
rect 17684 12223 17736 12232
rect 17684 12189 17693 12223
rect 17693 12189 17727 12223
rect 17727 12189 17736 12223
rect 17868 12223 17920 12232
rect 17684 12180 17736 12189
rect 17868 12189 17877 12223
rect 17877 12189 17911 12223
rect 17911 12189 17920 12223
rect 17868 12180 17920 12189
rect 18420 12180 18472 12232
rect 20812 12223 20864 12232
rect 20812 12189 20821 12223
rect 20821 12189 20855 12223
rect 20855 12189 20864 12223
rect 20812 12180 20864 12189
rect 21640 12180 21692 12232
rect 22836 12316 22888 12368
rect 22284 12248 22336 12300
rect 22928 12248 22980 12300
rect 22008 12223 22060 12232
rect 22008 12189 22017 12223
rect 22017 12189 22051 12223
rect 22051 12189 22060 12223
rect 22008 12180 22060 12189
rect 22192 12180 22244 12232
rect 23204 12180 23256 12232
rect 16120 12112 16172 12121
rect 4344 12044 4396 12096
rect 5908 12044 5960 12096
rect 9312 12044 9364 12096
rect 13360 12044 13412 12096
rect 15752 12044 15804 12096
rect 16948 12112 17000 12164
rect 17408 12044 17460 12096
rect 18604 12112 18656 12164
rect 20168 12112 20220 12164
rect 21272 12112 21324 12164
rect 21548 12155 21600 12164
rect 21548 12121 21557 12155
rect 21557 12121 21591 12155
rect 21591 12121 21600 12155
rect 21548 12112 21600 12121
rect 22376 12112 22428 12164
rect 22652 12112 22704 12164
rect 21180 12044 21232 12096
rect 21456 12044 21508 12096
rect 6630 11942 6682 11994
rect 6694 11942 6746 11994
rect 6758 11942 6810 11994
rect 6822 11942 6874 11994
rect 6886 11942 6938 11994
rect 12311 11942 12363 11994
rect 12375 11942 12427 11994
rect 12439 11942 12491 11994
rect 12503 11942 12555 11994
rect 12567 11942 12619 11994
rect 17992 11942 18044 11994
rect 18056 11942 18108 11994
rect 18120 11942 18172 11994
rect 18184 11942 18236 11994
rect 18248 11942 18300 11994
rect 23673 11942 23725 11994
rect 23737 11942 23789 11994
rect 23801 11942 23853 11994
rect 23865 11942 23917 11994
rect 23929 11942 23981 11994
rect 1768 11840 1820 11892
rect 2504 11883 2556 11892
rect 2504 11849 2513 11883
rect 2513 11849 2547 11883
rect 2547 11849 2556 11883
rect 2504 11840 2556 11849
rect 2688 11883 2740 11892
rect 2688 11849 2697 11883
rect 2697 11849 2731 11883
rect 2731 11849 2740 11883
rect 2688 11840 2740 11849
rect 2964 11840 3016 11892
rect 4896 11840 4948 11892
rect 3332 11772 3384 11824
rect 5172 11815 5224 11824
rect 1676 11747 1728 11756
rect 1676 11713 1685 11747
rect 1685 11713 1719 11747
rect 1719 11713 1728 11747
rect 1676 11704 1728 11713
rect 2964 11704 3016 11756
rect 3516 11704 3568 11756
rect 5172 11781 5181 11815
rect 5181 11781 5215 11815
rect 5215 11781 5224 11815
rect 5172 11772 5224 11781
rect 5632 11840 5684 11892
rect 7012 11840 7064 11892
rect 9220 11840 9272 11892
rect 11612 11840 11664 11892
rect 13176 11840 13228 11892
rect 17500 11840 17552 11892
rect 19156 11840 19208 11892
rect 19800 11840 19852 11892
rect 21364 11883 21416 11892
rect 21364 11849 21373 11883
rect 21373 11849 21407 11883
rect 21407 11849 21416 11883
rect 21364 11840 21416 11849
rect 23020 11883 23072 11892
rect 23020 11849 23029 11883
rect 23029 11849 23063 11883
rect 23063 11849 23072 11883
rect 23020 11840 23072 11849
rect 7196 11772 7248 11824
rect 4988 11747 5040 11756
rect 4988 11713 4997 11747
rect 4997 11713 5031 11747
rect 5031 11713 5040 11747
rect 4988 11704 5040 11713
rect 1860 11679 1912 11688
rect 1860 11645 1869 11679
rect 1869 11645 1903 11679
rect 1903 11645 1912 11679
rect 1860 11636 1912 11645
rect 1952 11636 2004 11688
rect 4620 11636 4672 11688
rect 4896 11636 4948 11688
rect 5448 11747 5500 11756
rect 5448 11713 5457 11747
rect 5457 11713 5491 11747
rect 5491 11713 5500 11747
rect 5448 11704 5500 11713
rect 6276 11704 6328 11756
rect 7840 11747 7892 11756
rect 7840 11713 7849 11747
rect 7849 11713 7883 11747
rect 7883 11713 7892 11747
rect 7840 11704 7892 11713
rect 8668 11747 8720 11756
rect 8668 11713 8677 11747
rect 8677 11713 8711 11747
rect 8711 11713 8720 11747
rect 8668 11704 8720 11713
rect 9128 11704 9180 11756
rect 11060 11772 11112 11824
rect 11704 11815 11756 11824
rect 11704 11781 11713 11815
rect 11713 11781 11747 11815
rect 11747 11781 11756 11815
rect 11704 11772 11756 11781
rect 11980 11772 12032 11824
rect 12716 11772 12768 11824
rect 14188 11772 14240 11824
rect 15108 11772 15160 11824
rect 18788 11772 18840 11824
rect 19524 11772 19576 11824
rect 22928 11772 22980 11824
rect 23296 11772 23348 11824
rect 9312 11704 9364 11756
rect 10232 11704 10284 11756
rect 10508 11704 10560 11756
rect 10784 11704 10836 11756
rect 11244 11704 11296 11756
rect 12072 11704 12124 11756
rect 17408 11747 17460 11756
rect 17408 11713 17417 11747
rect 17417 11713 17451 11747
rect 17451 11713 17460 11747
rect 17408 11704 17460 11713
rect 17592 11747 17644 11756
rect 17592 11713 17601 11747
rect 17601 11713 17635 11747
rect 17635 11713 17644 11747
rect 17592 11704 17644 11713
rect 17776 11704 17828 11756
rect 18972 11704 19024 11756
rect 5632 11636 5684 11688
rect 2136 11500 2188 11552
rect 2780 11500 2832 11552
rect 6552 11500 6604 11552
rect 7196 11679 7248 11688
rect 7196 11645 7205 11679
rect 7205 11645 7239 11679
rect 7239 11645 7248 11679
rect 10048 11679 10100 11688
rect 7196 11636 7248 11645
rect 10048 11645 10057 11679
rect 10057 11645 10091 11679
rect 10091 11645 10100 11679
rect 10048 11636 10100 11645
rect 13452 11636 13504 11688
rect 13728 11636 13780 11688
rect 15660 11636 15712 11688
rect 7656 11568 7708 11620
rect 17316 11636 17368 11688
rect 19340 11636 19392 11688
rect 19984 11704 20036 11756
rect 21364 11704 21416 11756
rect 21732 11704 21784 11756
rect 22100 11747 22152 11756
rect 22100 11713 22109 11747
rect 22109 11713 22143 11747
rect 22143 11713 22152 11747
rect 23020 11747 23072 11756
rect 22100 11704 22152 11713
rect 23020 11713 23029 11747
rect 23029 11713 23063 11747
rect 23063 11713 23072 11747
rect 23020 11704 23072 11713
rect 23112 11704 23164 11756
rect 22652 11636 22704 11688
rect 8116 11500 8168 11552
rect 9864 11500 9916 11552
rect 10968 11500 11020 11552
rect 13544 11500 13596 11552
rect 14372 11500 14424 11552
rect 14740 11543 14792 11552
rect 14740 11509 14749 11543
rect 14749 11509 14783 11543
rect 14783 11509 14792 11543
rect 14740 11500 14792 11509
rect 15568 11500 15620 11552
rect 15936 11543 15988 11552
rect 15936 11509 15945 11543
rect 15945 11509 15979 11543
rect 15979 11509 15988 11543
rect 15936 11500 15988 11509
rect 18420 11543 18472 11552
rect 18420 11509 18429 11543
rect 18429 11509 18463 11543
rect 18463 11509 18472 11543
rect 18420 11500 18472 11509
rect 18788 11500 18840 11552
rect 19984 11500 20036 11552
rect 3790 11398 3842 11450
rect 3854 11398 3906 11450
rect 3918 11398 3970 11450
rect 3982 11398 4034 11450
rect 4046 11398 4098 11450
rect 9471 11398 9523 11450
rect 9535 11398 9587 11450
rect 9599 11398 9651 11450
rect 9663 11398 9715 11450
rect 9727 11398 9779 11450
rect 15152 11398 15204 11450
rect 15216 11398 15268 11450
rect 15280 11398 15332 11450
rect 15344 11398 15396 11450
rect 15408 11398 15460 11450
rect 20833 11398 20885 11450
rect 20897 11398 20949 11450
rect 20961 11398 21013 11450
rect 21025 11398 21077 11450
rect 21089 11398 21141 11450
rect 3240 11296 3292 11348
rect 7472 11296 7524 11348
rect 1860 11228 1912 11280
rect 3884 11228 3936 11280
rect 4344 11228 4396 11280
rect 7932 11228 7984 11280
rect 4068 11203 4120 11212
rect 1584 11135 1636 11144
rect 1584 11101 1593 11135
rect 1593 11101 1627 11135
rect 1627 11101 1636 11135
rect 1584 11092 1636 11101
rect 2412 11135 2464 11144
rect 2412 11101 2421 11135
rect 2421 11101 2455 11135
rect 2455 11101 2464 11135
rect 2412 11092 2464 11101
rect 4068 11169 4077 11203
rect 4077 11169 4111 11203
rect 4111 11169 4120 11203
rect 4068 11160 4120 11169
rect 4160 11160 4212 11212
rect 4620 11160 4672 11212
rect 5724 11160 5776 11212
rect 7840 11160 7892 11212
rect 2872 11092 2924 11144
rect 3516 11092 3568 11144
rect 4344 11135 4396 11144
rect 4344 11101 4353 11135
rect 4353 11101 4387 11135
rect 4387 11101 4396 11135
rect 4344 11092 4396 11101
rect 5908 11092 5960 11144
rect 7288 11092 7340 11144
rect 7472 11092 7524 11144
rect 9220 11092 9272 11144
rect 9864 11160 9916 11212
rect 9772 11135 9824 11144
rect 9772 11101 9781 11135
rect 9781 11101 9815 11135
rect 9815 11101 9824 11135
rect 9772 11092 9824 11101
rect 10600 11135 10652 11144
rect 10600 11101 10609 11135
rect 10609 11101 10643 11135
rect 10643 11101 10652 11135
rect 10600 11092 10652 11101
rect 13084 11296 13136 11348
rect 13544 11296 13596 11348
rect 14648 11296 14700 11348
rect 16028 11296 16080 11348
rect 19616 11339 19668 11348
rect 19616 11305 19625 11339
rect 19625 11305 19659 11339
rect 19659 11305 19668 11339
rect 22284 11339 22336 11348
rect 19616 11296 19668 11305
rect 22284 11305 22293 11339
rect 22293 11305 22327 11339
rect 22327 11305 22336 11339
rect 22284 11296 22336 11305
rect 15016 11228 15068 11280
rect 15568 11228 15620 11280
rect 16856 11228 16908 11280
rect 16948 11228 17000 11280
rect 11888 11135 11940 11144
rect 11888 11101 11897 11135
rect 11897 11101 11931 11135
rect 11931 11101 11940 11135
rect 11888 11092 11940 11101
rect 12624 11135 12676 11144
rect 4252 11024 4304 11076
rect 6092 11024 6144 11076
rect 8576 11024 8628 11076
rect 10048 11024 10100 11076
rect 10968 11024 11020 11076
rect 12624 11101 12633 11135
rect 12633 11101 12667 11135
rect 12667 11101 12676 11135
rect 12624 11092 12676 11101
rect 13084 11135 13136 11144
rect 13084 11101 13093 11135
rect 13093 11101 13127 11135
rect 13127 11101 13136 11135
rect 13084 11092 13136 11101
rect 13452 11135 13504 11144
rect 13452 11101 13461 11135
rect 13461 11101 13495 11135
rect 13495 11101 13504 11135
rect 13452 11092 13504 11101
rect 13820 11092 13872 11144
rect 14280 11135 14332 11144
rect 14280 11101 14289 11135
rect 14289 11101 14323 11135
rect 14323 11101 14332 11135
rect 14280 11092 14332 11101
rect 12992 11024 13044 11076
rect 5816 10956 5868 11008
rect 7380 10956 7432 11008
rect 9772 10956 9824 11008
rect 12164 10956 12216 11008
rect 13360 11067 13412 11076
rect 13360 11033 13369 11067
rect 13369 11033 13403 11067
rect 13403 11033 13412 11067
rect 13360 11024 13412 11033
rect 14188 11024 14240 11076
rect 15384 11160 15436 11212
rect 14924 11092 14976 11144
rect 15752 11203 15804 11212
rect 15752 11169 15761 11203
rect 15761 11169 15795 11203
rect 15795 11169 15804 11203
rect 15752 11160 15804 11169
rect 15936 11160 15988 11212
rect 21180 11228 21232 11280
rect 23388 11228 23440 11280
rect 16120 11092 16172 11144
rect 16856 11135 16908 11144
rect 16856 11101 16865 11135
rect 16865 11101 16899 11135
rect 16899 11101 16908 11135
rect 16856 11092 16908 11101
rect 17776 11092 17828 11144
rect 18236 11092 18288 11144
rect 18604 11135 18656 11144
rect 18604 11101 18613 11135
rect 18613 11101 18647 11135
rect 18647 11101 18656 11135
rect 18604 11092 18656 11101
rect 18788 11092 18840 11144
rect 19708 11135 19760 11144
rect 19708 11101 19717 11135
rect 19717 11101 19751 11135
rect 19751 11101 19760 11135
rect 19708 11092 19760 11101
rect 15108 11024 15160 11076
rect 17868 11024 17920 11076
rect 18880 11067 18932 11076
rect 18880 11033 18889 11067
rect 18889 11033 18923 11067
rect 18923 11033 18932 11067
rect 18880 11024 18932 11033
rect 19616 11024 19668 11076
rect 21456 11092 21508 11144
rect 23020 11160 23072 11212
rect 22652 11024 22704 11076
rect 23296 11024 23348 11076
rect 15660 10956 15712 11008
rect 15752 10956 15804 11008
rect 16488 10956 16540 11008
rect 18420 10956 18472 11008
rect 18788 10956 18840 11008
rect 21364 10999 21416 11008
rect 21364 10965 21373 10999
rect 21373 10965 21407 10999
rect 21407 10965 21416 10999
rect 21364 10956 21416 10965
rect 21732 10956 21784 11008
rect 6630 10854 6682 10906
rect 6694 10854 6746 10906
rect 6758 10854 6810 10906
rect 6822 10854 6874 10906
rect 6886 10854 6938 10906
rect 12311 10854 12363 10906
rect 12375 10854 12427 10906
rect 12439 10854 12491 10906
rect 12503 10854 12555 10906
rect 12567 10854 12619 10906
rect 17992 10854 18044 10906
rect 18056 10854 18108 10906
rect 18120 10854 18172 10906
rect 18184 10854 18236 10906
rect 18248 10854 18300 10906
rect 23673 10854 23725 10906
rect 23737 10854 23789 10906
rect 23801 10854 23853 10906
rect 23865 10854 23917 10906
rect 23929 10854 23981 10906
rect 1584 10752 1636 10804
rect 2964 10752 3016 10804
rect 4252 10752 4304 10804
rect 4344 10752 4396 10804
rect 4712 10752 4764 10804
rect 6368 10752 6420 10804
rect 2044 10684 2096 10736
rect 2320 10548 2372 10600
rect 2596 10480 2648 10532
rect 2780 10616 2832 10668
rect 4068 10684 4120 10736
rect 4620 10684 4672 10736
rect 3332 10548 3384 10600
rect 5724 10616 5776 10668
rect 6552 10616 6604 10668
rect 10876 10752 10928 10804
rect 11888 10752 11940 10804
rect 13360 10752 13412 10804
rect 13636 10795 13688 10804
rect 13636 10761 13645 10795
rect 13645 10761 13679 10795
rect 13679 10761 13688 10795
rect 13636 10752 13688 10761
rect 14832 10752 14884 10804
rect 15752 10795 15804 10804
rect 15752 10761 15761 10795
rect 15761 10761 15795 10795
rect 15795 10761 15804 10795
rect 15752 10752 15804 10761
rect 16212 10752 16264 10804
rect 17592 10752 17644 10804
rect 7012 10727 7064 10736
rect 7012 10693 7021 10727
rect 7021 10693 7055 10727
rect 7055 10693 7064 10727
rect 7012 10684 7064 10693
rect 4620 10548 4672 10600
rect 5356 10548 5408 10600
rect 5632 10548 5684 10600
rect 7932 10659 7984 10668
rect 7932 10625 7941 10659
rect 7941 10625 7975 10659
rect 7975 10625 7984 10659
rect 7932 10616 7984 10625
rect 7288 10591 7340 10600
rect 7288 10557 7297 10591
rect 7297 10557 7331 10591
rect 7331 10557 7340 10591
rect 7288 10548 7340 10557
rect 7748 10548 7800 10600
rect 4160 10480 4212 10532
rect 5540 10480 5592 10532
rect 2136 10455 2188 10464
rect 2136 10421 2145 10455
rect 2145 10421 2179 10455
rect 2179 10421 2188 10455
rect 2136 10412 2188 10421
rect 3516 10412 3568 10464
rect 4804 10412 4856 10464
rect 5816 10412 5868 10464
rect 6828 10480 6880 10532
rect 9128 10684 9180 10736
rect 11704 10684 11756 10736
rect 12900 10684 12952 10736
rect 13912 10684 13964 10736
rect 15476 10684 15528 10736
rect 15568 10727 15620 10736
rect 15568 10693 15577 10727
rect 15577 10693 15611 10727
rect 15611 10693 15620 10727
rect 15568 10684 15620 10693
rect 9312 10616 9364 10668
rect 10048 10548 10100 10600
rect 13084 10616 13136 10668
rect 14648 10616 14700 10668
rect 12808 10548 12860 10600
rect 10232 10480 10284 10532
rect 12900 10480 12952 10532
rect 14924 10659 14976 10668
rect 14924 10625 14933 10659
rect 14933 10625 14967 10659
rect 14967 10625 14976 10659
rect 14924 10616 14976 10625
rect 15016 10548 15068 10600
rect 15384 10616 15436 10668
rect 16396 10684 16448 10736
rect 17132 10684 17184 10736
rect 18052 10659 18104 10668
rect 18052 10625 18061 10659
rect 18061 10625 18095 10659
rect 18095 10625 18104 10659
rect 18052 10616 18104 10625
rect 19156 10752 19208 10804
rect 21640 10752 21692 10804
rect 19156 10659 19208 10702
rect 19156 10650 19187 10659
rect 19187 10650 19208 10659
rect 19984 10684 20036 10736
rect 22560 10752 22612 10804
rect 19708 10616 19760 10668
rect 19800 10616 19852 10668
rect 20076 10659 20128 10668
rect 20076 10625 20085 10659
rect 20085 10625 20119 10659
rect 20119 10625 20128 10659
rect 20076 10616 20128 10625
rect 21548 10616 21600 10668
rect 22836 10684 22888 10736
rect 23112 10752 23164 10804
rect 22652 10616 22704 10668
rect 17592 10591 17644 10600
rect 17592 10557 17601 10591
rect 17601 10557 17635 10591
rect 17635 10557 17644 10591
rect 17592 10548 17644 10557
rect 18604 10548 18656 10600
rect 16672 10480 16724 10532
rect 18052 10480 18104 10532
rect 19616 10548 19668 10600
rect 20536 10548 20588 10600
rect 20720 10548 20772 10600
rect 19064 10523 19116 10532
rect 19064 10489 19073 10523
rect 19073 10489 19107 10523
rect 19107 10489 19116 10523
rect 19064 10480 19116 10489
rect 19248 10480 19300 10532
rect 22468 10548 22520 10600
rect 7288 10412 7340 10464
rect 7656 10412 7708 10464
rect 10508 10412 10560 10464
rect 12256 10412 12308 10464
rect 13452 10412 13504 10464
rect 16488 10412 16540 10464
rect 17408 10412 17460 10464
rect 19524 10412 19576 10464
rect 19800 10412 19852 10464
rect 21548 10412 21600 10464
rect 22376 10412 22428 10464
rect 22560 10455 22612 10464
rect 22560 10421 22569 10455
rect 22569 10421 22603 10455
rect 22603 10421 22612 10455
rect 22560 10412 22612 10421
rect 3790 10310 3842 10362
rect 3854 10310 3906 10362
rect 3918 10310 3970 10362
rect 3982 10310 4034 10362
rect 4046 10310 4098 10362
rect 9471 10310 9523 10362
rect 9535 10310 9587 10362
rect 9599 10310 9651 10362
rect 9663 10310 9715 10362
rect 9727 10310 9779 10362
rect 15152 10310 15204 10362
rect 15216 10310 15268 10362
rect 15280 10310 15332 10362
rect 15344 10310 15396 10362
rect 15408 10310 15460 10362
rect 20833 10310 20885 10362
rect 20897 10310 20949 10362
rect 20961 10310 21013 10362
rect 21025 10310 21077 10362
rect 21089 10310 21141 10362
rect 2504 10208 2556 10260
rect 4988 10208 5040 10260
rect 6460 10208 6512 10260
rect 8576 10251 8628 10260
rect 2688 10140 2740 10192
rect 3056 10140 3108 10192
rect 5540 10140 5592 10192
rect 6276 10140 6328 10192
rect 3332 10072 3384 10124
rect 4160 10072 4212 10124
rect 7104 10140 7156 10192
rect 7564 10140 7616 10192
rect 8576 10217 8585 10251
rect 8585 10217 8619 10251
rect 8619 10217 8628 10251
rect 8576 10208 8628 10217
rect 13544 10251 13596 10260
rect 13544 10217 13553 10251
rect 13553 10217 13587 10251
rect 13587 10217 13596 10251
rect 13544 10208 13596 10217
rect 13912 10208 13964 10260
rect 12256 10183 12308 10192
rect 12256 10149 12265 10183
rect 12265 10149 12299 10183
rect 12299 10149 12308 10183
rect 12256 10140 12308 10149
rect 13360 10140 13412 10192
rect 15752 10208 15804 10260
rect 17684 10251 17736 10260
rect 17684 10217 17693 10251
rect 17693 10217 17727 10251
rect 17727 10217 17736 10251
rect 17684 10208 17736 10217
rect 6828 10072 6880 10124
rect 8024 10072 8076 10124
rect 9680 10072 9732 10124
rect 3056 10004 3108 10056
rect 3424 10047 3476 10056
rect 3424 10013 3433 10047
rect 3433 10013 3467 10047
rect 3467 10013 3476 10047
rect 3424 10004 3476 10013
rect 3240 9936 3292 9988
rect 1676 9911 1728 9920
rect 1676 9877 1685 9911
rect 1685 9877 1719 9911
rect 1719 9877 1728 9911
rect 1676 9868 1728 9877
rect 5080 10047 5132 10056
rect 5080 10013 5089 10047
rect 5089 10013 5123 10047
rect 5123 10013 5132 10047
rect 5080 10004 5132 10013
rect 5356 10004 5408 10056
rect 5540 10004 5592 10056
rect 6184 10004 6236 10056
rect 5080 9868 5132 9920
rect 6000 9936 6052 9988
rect 7196 10004 7248 10056
rect 7840 10004 7892 10056
rect 9128 10047 9180 10056
rect 9128 10013 9137 10047
rect 9137 10013 9171 10047
rect 9171 10013 9180 10047
rect 9128 10004 9180 10013
rect 9312 10004 9364 10056
rect 10048 10004 10100 10056
rect 13728 10072 13780 10124
rect 7656 9936 7708 9988
rect 10600 9936 10652 9988
rect 12716 10004 12768 10056
rect 12992 10004 13044 10056
rect 14740 10004 14792 10056
rect 15660 10140 15712 10192
rect 18512 10208 18564 10260
rect 22100 10208 22152 10260
rect 17868 10140 17920 10192
rect 22008 10140 22060 10192
rect 16396 10072 16448 10124
rect 5816 9868 5868 9920
rect 6828 9868 6880 9920
rect 7380 9911 7432 9920
rect 7380 9877 7389 9911
rect 7389 9877 7423 9911
rect 7423 9877 7432 9911
rect 7380 9868 7432 9877
rect 7564 9868 7616 9920
rect 7932 9868 7984 9920
rect 10508 9868 10560 9920
rect 13268 9936 13320 9988
rect 14464 9936 14516 9988
rect 15016 9936 15068 9988
rect 16028 10004 16080 10056
rect 12716 9868 12768 9920
rect 14648 9868 14700 9920
rect 15568 9868 15620 9920
rect 16764 10004 16816 10056
rect 18880 10072 18932 10124
rect 17408 10047 17460 10056
rect 17408 10013 17417 10047
rect 17417 10013 17451 10047
rect 17451 10013 17460 10047
rect 17408 10004 17460 10013
rect 17500 10047 17552 10056
rect 17500 10013 17509 10047
rect 17509 10013 17543 10047
rect 17543 10013 17552 10047
rect 18144 10047 18196 10056
rect 17500 10004 17552 10013
rect 18144 10013 18153 10047
rect 18153 10013 18187 10047
rect 18187 10013 18196 10047
rect 18144 10004 18196 10013
rect 16672 9979 16724 9988
rect 16672 9945 16681 9979
rect 16681 9945 16715 9979
rect 16715 9945 16724 9979
rect 16672 9936 16724 9945
rect 16948 9936 17000 9988
rect 17868 9936 17920 9988
rect 18328 10004 18380 10056
rect 19156 10004 19208 10056
rect 20076 10004 20128 10056
rect 20444 10072 20496 10124
rect 22744 10140 22796 10192
rect 22192 10072 22244 10124
rect 18696 9936 18748 9988
rect 17224 9868 17276 9920
rect 17592 9868 17644 9920
rect 19984 9868 20036 9920
rect 20352 10047 20404 10056
rect 20352 10013 20361 10047
rect 20361 10013 20395 10047
rect 20395 10013 20404 10047
rect 20352 10004 20404 10013
rect 21180 10004 21232 10056
rect 21548 10047 21600 10056
rect 21548 10013 21557 10047
rect 21557 10013 21591 10047
rect 21591 10013 21600 10047
rect 21548 10004 21600 10013
rect 22100 10004 22152 10056
rect 21456 9868 21508 9920
rect 23020 10004 23072 10056
rect 22652 9868 22704 9920
rect 23204 9911 23256 9920
rect 23204 9877 23213 9911
rect 23213 9877 23247 9911
rect 23247 9877 23256 9911
rect 23204 9868 23256 9877
rect 6630 9766 6682 9818
rect 6694 9766 6746 9818
rect 6758 9766 6810 9818
rect 6822 9766 6874 9818
rect 6886 9766 6938 9818
rect 12311 9766 12363 9818
rect 12375 9766 12427 9818
rect 12439 9766 12491 9818
rect 12503 9766 12555 9818
rect 12567 9766 12619 9818
rect 17992 9766 18044 9818
rect 18056 9766 18108 9818
rect 18120 9766 18172 9818
rect 18184 9766 18236 9818
rect 18248 9766 18300 9818
rect 23673 9766 23725 9818
rect 23737 9766 23789 9818
rect 23801 9766 23853 9818
rect 23865 9766 23917 9818
rect 23929 9766 23981 9818
rect 2780 9596 2832 9648
rect 3148 9596 3200 9648
rect 4252 9596 4304 9648
rect 7288 9664 7340 9716
rect 7564 9664 7616 9716
rect 7840 9664 7892 9716
rect 5080 9596 5132 9648
rect 5356 9596 5408 9648
rect 5908 9639 5960 9648
rect 5908 9605 5917 9639
rect 5917 9605 5951 9639
rect 5951 9605 5960 9639
rect 5908 9596 5960 9605
rect 7012 9596 7064 9648
rect 2228 9528 2280 9580
rect 1952 9460 2004 9512
rect 3424 9528 3476 9580
rect 4160 9528 4212 9580
rect 3332 9460 3384 9512
rect 2228 9392 2280 9444
rect 2872 9392 2924 9444
rect 3240 9392 3292 9444
rect 4620 9460 4672 9512
rect 3792 9324 3844 9376
rect 4712 9367 4764 9376
rect 4712 9333 4721 9367
rect 4721 9333 4755 9367
rect 4755 9333 4764 9367
rect 4712 9324 4764 9333
rect 7472 9528 7524 9580
rect 7656 9571 7708 9580
rect 7656 9537 7665 9571
rect 7665 9537 7699 9571
rect 7699 9537 7708 9571
rect 7656 9528 7708 9537
rect 15476 9664 15528 9716
rect 15568 9664 15620 9716
rect 9680 9596 9732 9648
rect 12992 9596 13044 9648
rect 23204 9664 23256 9716
rect 16488 9596 16540 9648
rect 5724 9460 5776 9512
rect 7748 9460 7800 9512
rect 5908 9392 5960 9444
rect 9128 9528 9180 9580
rect 9956 9528 10008 9580
rect 10968 9571 11020 9580
rect 10968 9537 10977 9571
rect 10977 9537 11011 9571
rect 11011 9537 11020 9571
rect 10968 9528 11020 9537
rect 11060 9528 11112 9580
rect 13636 9571 13688 9580
rect 9312 9503 9364 9512
rect 9312 9469 9321 9503
rect 9321 9469 9355 9503
rect 9355 9469 9364 9503
rect 9312 9460 9364 9469
rect 9496 9460 9548 9512
rect 11612 9460 11664 9512
rect 6368 9324 6420 9376
rect 7196 9367 7248 9376
rect 7196 9333 7205 9367
rect 7205 9333 7239 9367
rect 7239 9333 7248 9367
rect 7196 9324 7248 9333
rect 7472 9324 7524 9376
rect 9312 9324 9364 9376
rect 12072 9392 12124 9444
rect 13636 9537 13645 9571
rect 13645 9537 13679 9571
rect 13679 9537 13688 9571
rect 13636 9528 13688 9537
rect 14372 9528 14424 9580
rect 14648 9528 14700 9580
rect 16672 9528 16724 9580
rect 16764 9528 16816 9580
rect 17132 9596 17184 9648
rect 19800 9596 19852 9648
rect 17592 9571 17644 9580
rect 15844 9460 15896 9512
rect 12808 9392 12860 9444
rect 15752 9392 15804 9444
rect 9864 9367 9916 9376
rect 9864 9333 9873 9367
rect 9873 9333 9907 9367
rect 9907 9333 9916 9367
rect 9864 9324 9916 9333
rect 11060 9367 11112 9376
rect 11060 9333 11069 9367
rect 11069 9333 11103 9367
rect 11103 9333 11112 9367
rect 11060 9324 11112 9333
rect 12624 9367 12676 9376
rect 12624 9333 12633 9367
rect 12633 9333 12667 9367
rect 12667 9333 12676 9367
rect 12624 9324 12676 9333
rect 12900 9324 12952 9376
rect 14096 9324 14148 9376
rect 14648 9324 14700 9376
rect 15660 9324 15712 9376
rect 16120 9324 16172 9376
rect 17592 9537 17601 9571
rect 17601 9537 17635 9571
rect 17635 9537 17644 9571
rect 17592 9528 17644 9537
rect 18328 9528 18380 9580
rect 18420 9528 18472 9580
rect 19524 9571 19576 9580
rect 19524 9537 19533 9571
rect 19533 9537 19567 9571
rect 19567 9537 19576 9571
rect 19524 9528 19576 9537
rect 20260 9528 20312 9580
rect 20628 9571 20680 9580
rect 16856 9392 16908 9444
rect 19616 9392 19668 9444
rect 20628 9537 20637 9571
rect 20637 9537 20671 9571
rect 20671 9537 20680 9571
rect 20628 9528 20680 9537
rect 20720 9571 20772 9580
rect 20720 9537 20729 9571
rect 20729 9537 20763 9571
rect 20763 9537 20772 9571
rect 20720 9528 20772 9537
rect 21180 9528 21232 9580
rect 21548 9596 21600 9648
rect 21916 9596 21968 9648
rect 23112 9639 23164 9648
rect 23112 9605 23121 9639
rect 23121 9605 23155 9639
rect 23155 9605 23164 9639
rect 23112 9596 23164 9605
rect 21640 9528 21692 9580
rect 22284 9528 22336 9580
rect 22928 9460 22980 9512
rect 20720 9392 20772 9444
rect 22376 9392 22428 9444
rect 16580 9324 16632 9376
rect 17592 9324 17644 9376
rect 19708 9367 19760 9376
rect 19708 9333 19717 9367
rect 19717 9333 19751 9367
rect 19751 9333 19760 9367
rect 19708 9324 19760 9333
rect 21088 9324 21140 9376
rect 21364 9324 21416 9376
rect 22192 9324 22244 9376
rect 22652 9392 22704 9444
rect 22744 9324 22796 9376
rect 3790 9222 3842 9274
rect 3854 9222 3906 9274
rect 3918 9222 3970 9274
rect 3982 9222 4034 9274
rect 4046 9222 4098 9274
rect 9471 9222 9523 9274
rect 9535 9222 9587 9274
rect 9599 9222 9651 9274
rect 9663 9222 9715 9274
rect 9727 9222 9779 9274
rect 15152 9222 15204 9274
rect 15216 9222 15268 9274
rect 15280 9222 15332 9274
rect 15344 9222 15396 9274
rect 15408 9222 15460 9274
rect 20833 9222 20885 9274
rect 20897 9222 20949 9274
rect 20961 9222 21013 9274
rect 21025 9222 21077 9274
rect 21089 9222 21141 9274
rect 1676 9120 1728 9172
rect 3424 9120 3476 9172
rect 4160 9120 4212 9172
rect 6276 9120 6328 9172
rect 7104 9120 7156 9172
rect 9312 9120 9364 9172
rect 9864 9163 9916 9172
rect 9864 9129 9873 9163
rect 9873 9129 9907 9163
rect 9907 9129 9916 9163
rect 9864 9120 9916 9129
rect 2320 9052 2372 9104
rect 2596 9027 2648 9036
rect 2596 8993 2605 9027
rect 2605 8993 2639 9027
rect 2639 8993 2648 9027
rect 2596 8984 2648 8993
rect 2136 8916 2188 8968
rect 3056 8891 3108 8900
rect 3056 8857 3065 8891
rect 3065 8857 3099 8891
rect 3099 8857 3108 8891
rect 3056 8848 3108 8857
rect 3884 8916 3936 8968
rect 4896 9052 4948 9104
rect 6276 8984 6328 9036
rect 4620 8916 4672 8968
rect 4252 8891 4304 8900
rect 4252 8857 4261 8891
rect 4261 8857 4295 8891
rect 4295 8857 4304 8891
rect 4252 8848 4304 8857
rect 4988 8848 5040 8900
rect 2596 8780 2648 8832
rect 4896 8780 4948 8832
rect 6000 8916 6052 8968
rect 6644 8959 6696 8968
rect 6644 8925 6653 8959
rect 6653 8925 6687 8959
rect 6687 8925 6696 8959
rect 6644 8916 6696 8925
rect 9772 8916 9824 8968
rect 10048 8959 10100 8968
rect 10048 8925 10057 8959
rect 10057 8925 10091 8959
rect 10091 8925 10100 8959
rect 10048 8916 10100 8925
rect 13176 9120 13228 9172
rect 14096 9120 14148 9172
rect 13084 9052 13136 9104
rect 17040 9120 17092 9172
rect 21364 9120 21416 9172
rect 22008 9120 22060 9172
rect 22836 9120 22888 9172
rect 16304 9052 16356 9104
rect 16856 9095 16908 9104
rect 16856 9061 16865 9095
rect 16865 9061 16899 9095
rect 16899 9061 16908 9095
rect 16856 9052 16908 9061
rect 19708 9052 19760 9104
rect 12624 8984 12676 9036
rect 11520 8959 11572 8968
rect 11520 8925 11529 8959
rect 11529 8925 11563 8959
rect 11563 8925 11572 8959
rect 11520 8916 11572 8925
rect 11612 8959 11664 8968
rect 11612 8925 11621 8959
rect 11621 8925 11655 8959
rect 11655 8925 11664 8959
rect 11612 8916 11664 8925
rect 7012 8848 7064 8900
rect 11704 8848 11756 8900
rect 8668 8780 8720 8832
rect 10968 8823 11020 8832
rect 10968 8789 10977 8823
rect 10977 8789 11011 8823
rect 11011 8789 11020 8823
rect 10968 8780 11020 8789
rect 12900 8848 12952 8900
rect 13084 8959 13136 8968
rect 13084 8925 13093 8959
rect 13093 8925 13127 8959
rect 13127 8925 13136 8959
rect 13084 8916 13136 8925
rect 13636 8916 13688 8968
rect 14372 8959 14424 8968
rect 14372 8925 14381 8959
rect 14381 8925 14415 8959
rect 14415 8925 14424 8959
rect 15844 8984 15896 9036
rect 16580 8984 16632 9036
rect 16948 9027 17000 9036
rect 16948 8993 16957 9027
rect 16957 8993 16991 9027
rect 16991 8993 17000 9027
rect 16948 8984 17000 8993
rect 22376 8984 22428 9036
rect 23112 8984 23164 9036
rect 14372 8916 14424 8925
rect 18328 8916 18380 8968
rect 19892 8959 19944 8968
rect 19892 8925 19901 8959
rect 19901 8925 19935 8959
rect 19935 8925 19944 8959
rect 19892 8916 19944 8925
rect 21180 8959 21232 8968
rect 21180 8925 21189 8959
rect 21189 8925 21223 8959
rect 21223 8925 21232 8959
rect 21180 8916 21232 8925
rect 21364 8959 21416 8968
rect 21364 8925 21373 8959
rect 21373 8925 21407 8959
rect 21407 8925 21416 8959
rect 21364 8916 21416 8925
rect 21456 8959 21508 8968
rect 21456 8925 21465 8959
rect 21465 8925 21499 8959
rect 21499 8925 21508 8959
rect 21456 8916 21508 8925
rect 21916 8916 21968 8968
rect 13728 8848 13780 8900
rect 14556 8780 14608 8832
rect 15384 8823 15436 8832
rect 15384 8789 15393 8823
rect 15393 8789 15427 8823
rect 15427 8789 15436 8823
rect 15384 8780 15436 8789
rect 15660 8891 15712 8900
rect 15660 8857 15669 8891
rect 15669 8857 15703 8891
rect 15703 8857 15712 8891
rect 15660 8848 15712 8857
rect 16764 8848 16816 8900
rect 19616 8848 19668 8900
rect 20260 8891 20312 8900
rect 20260 8857 20269 8891
rect 20269 8857 20303 8891
rect 20303 8857 20312 8891
rect 20260 8848 20312 8857
rect 15752 8780 15804 8832
rect 17500 8780 17552 8832
rect 18880 8780 18932 8832
rect 19432 8780 19484 8832
rect 22192 8823 22244 8832
rect 22192 8789 22201 8823
rect 22201 8789 22235 8823
rect 22235 8789 22244 8823
rect 22192 8780 22244 8789
rect 23204 8823 23256 8832
rect 23204 8789 23213 8823
rect 23213 8789 23247 8823
rect 23247 8789 23256 8823
rect 23204 8780 23256 8789
rect 6630 8678 6682 8730
rect 6694 8678 6746 8730
rect 6758 8678 6810 8730
rect 6822 8678 6874 8730
rect 6886 8678 6938 8730
rect 12311 8678 12363 8730
rect 12375 8678 12427 8730
rect 12439 8678 12491 8730
rect 12503 8678 12555 8730
rect 12567 8678 12619 8730
rect 17992 8678 18044 8730
rect 18056 8678 18108 8730
rect 18120 8678 18172 8730
rect 18184 8678 18236 8730
rect 18248 8678 18300 8730
rect 23673 8678 23725 8730
rect 23737 8678 23789 8730
rect 23801 8678 23853 8730
rect 23865 8678 23917 8730
rect 23929 8678 23981 8730
rect 7656 8576 7708 8628
rect 9128 8619 9180 8628
rect 9128 8585 9137 8619
rect 9137 8585 9171 8619
rect 9171 8585 9180 8619
rect 9128 8576 9180 8585
rect 10876 8576 10928 8628
rect 12072 8576 12124 8628
rect 12808 8576 12860 8628
rect 16856 8576 16908 8628
rect 17316 8576 17368 8628
rect 19892 8576 19944 8628
rect 23204 8576 23256 8628
rect 1952 8508 2004 8560
rect 3240 8508 3292 8560
rect 7012 8551 7064 8560
rect 7012 8517 7021 8551
rect 7021 8517 7055 8551
rect 7055 8517 7064 8551
rect 7012 8508 7064 8517
rect 8300 8508 8352 8560
rect 9036 8508 9088 8560
rect 10232 8508 10284 8560
rect 2780 8483 2832 8492
rect 2780 8449 2789 8483
rect 2789 8449 2823 8483
rect 2823 8449 2832 8483
rect 2780 8440 2832 8449
rect 3332 8483 3384 8492
rect 3332 8449 3341 8483
rect 3341 8449 3375 8483
rect 3375 8449 3384 8483
rect 3332 8440 3384 8449
rect 4252 8440 4304 8492
rect 4896 8483 4948 8492
rect 4896 8449 4905 8483
rect 4905 8449 4939 8483
rect 4939 8449 4948 8483
rect 4896 8440 4948 8449
rect 5908 8440 5960 8492
rect 7472 8483 7524 8492
rect 7472 8449 7481 8483
rect 7481 8449 7515 8483
rect 7515 8449 7524 8483
rect 7472 8440 7524 8449
rect 7840 8440 7892 8492
rect 8668 8440 8720 8492
rect 8944 8440 8996 8492
rect 2136 8372 2188 8424
rect 2412 8372 2464 8424
rect 2688 8372 2740 8424
rect 2964 8372 3016 8424
rect 3516 8415 3568 8424
rect 3516 8381 3525 8415
rect 3525 8381 3559 8415
rect 3559 8381 3568 8415
rect 3516 8372 3568 8381
rect 4436 8372 4488 8424
rect 6368 8372 6420 8424
rect 9312 8372 9364 8424
rect 10692 8440 10744 8492
rect 11704 8440 11756 8492
rect 11888 8483 11940 8492
rect 11888 8449 11897 8483
rect 11897 8449 11931 8483
rect 11931 8449 11940 8483
rect 11888 8440 11940 8449
rect 12164 8483 12216 8492
rect 11612 8372 11664 8424
rect 12164 8449 12173 8483
rect 12173 8449 12207 8483
rect 12207 8449 12216 8483
rect 12164 8440 12216 8449
rect 13268 8508 13320 8560
rect 3240 8304 3292 8356
rect 4344 8304 4396 8356
rect 6276 8304 6328 8356
rect 9864 8304 9916 8356
rect 10508 8304 10560 8356
rect 7932 8279 7984 8288
rect 7932 8245 7941 8279
rect 7941 8245 7975 8279
rect 7975 8245 7984 8279
rect 7932 8236 7984 8245
rect 8116 8279 8168 8288
rect 8116 8245 8125 8279
rect 8125 8245 8159 8279
rect 8159 8245 8168 8279
rect 8116 8236 8168 8245
rect 9220 8236 9272 8288
rect 9772 8236 9824 8288
rect 10784 8236 10836 8288
rect 14096 8415 14148 8424
rect 14096 8381 14105 8415
rect 14105 8381 14139 8415
rect 14139 8381 14148 8415
rect 14096 8372 14148 8381
rect 13636 8304 13688 8356
rect 14648 8415 14700 8424
rect 14648 8381 14657 8415
rect 14657 8381 14691 8415
rect 14691 8381 14700 8415
rect 14648 8372 14700 8381
rect 15844 8508 15896 8560
rect 16028 8508 16080 8560
rect 16580 8508 16632 8560
rect 19616 8551 19668 8560
rect 17316 8415 17368 8424
rect 17316 8381 17325 8415
rect 17325 8381 17359 8415
rect 17359 8381 17368 8415
rect 17316 8372 17368 8381
rect 18236 8440 18288 8492
rect 19616 8517 19625 8551
rect 19625 8517 19659 8551
rect 19659 8517 19668 8551
rect 20352 8551 20404 8560
rect 19616 8508 19668 8517
rect 20352 8517 20361 8551
rect 20361 8517 20395 8551
rect 20395 8517 20404 8551
rect 20352 8508 20404 8517
rect 20720 8508 20772 8560
rect 21732 8508 21784 8560
rect 17684 8372 17736 8424
rect 18880 8440 18932 8492
rect 21548 8440 21600 8492
rect 21640 8440 21692 8492
rect 22560 8483 22612 8492
rect 22560 8449 22569 8483
rect 22569 8449 22603 8483
rect 22603 8449 22612 8483
rect 22836 8483 22888 8492
rect 22560 8440 22612 8449
rect 22836 8449 22845 8483
rect 22845 8449 22879 8483
rect 22879 8449 22888 8483
rect 22836 8440 22888 8449
rect 17132 8304 17184 8356
rect 19524 8372 19576 8424
rect 20720 8372 20772 8424
rect 22744 8415 22796 8424
rect 22744 8381 22753 8415
rect 22753 8381 22787 8415
rect 22787 8381 22796 8415
rect 22744 8372 22796 8381
rect 19340 8304 19392 8356
rect 20628 8304 20680 8356
rect 22284 8347 22336 8356
rect 22284 8313 22293 8347
rect 22293 8313 22327 8347
rect 22327 8313 22336 8347
rect 22284 8304 22336 8313
rect 12900 8236 12952 8288
rect 15016 8236 15068 8288
rect 15384 8236 15436 8288
rect 3790 8134 3842 8186
rect 3854 8134 3906 8186
rect 3918 8134 3970 8186
rect 3982 8134 4034 8186
rect 4046 8134 4098 8186
rect 9471 8134 9523 8186
rect 9535 8134 9587 8186
rect 9599 8134 9651 8186
rect 9663 8134 9715 8186
rect 9727 8134 9779 8186
rect 15152 8134 15204 8186
rect 15216 8134 15268 8186
rect 15280 8134 15332 8186
rect 15344 8134 15396 8186
rect 15408 8134 15460 8186
rect 20833 8134 20885 8186
rect 20897 8134 20949 8186
rect 20961 8134 21013 8186
rect 21025 8134 21077 8186
rect 21089 8134 21141 8186
rect 3332 8032 3384 8084
rect 4160 8032 4212 8084
rect 4988 8032 5040 8084
rect 6092 8032 6144 8084
rect 7748 8075 7800 8084
rect 7748 8041 7757 8075
rect 7757 8041 7791 8075
rect 7791 8041 7800 8075
rect 7748 8032 7800 8041
rect 2780 7964 2832 8016
rect 3240 7964 3292 8016
rect 1952 7871 2004 7880
rect 1952 7837 1961 7871
rect 1961 7837 1995 7871
rect 1995 7837 2004 7871
rect 1952 7828 2004 7837
rect 2228 7871 2280 7880
rect 2228 7837 2237 7871
rect 2237 7837 2271 7871
rect 2271 7837 2280 7871
rect 2228 7828 2280 7837
rect 4528 7896 4580 7948
rect 5816 7964 5868 8016
rect 7380 7964 7432 8016
rect 8944 8032 8996 8084
rect 11152 8032 11204 8084
rect 13636 8075 13688 8084
rect 13636 8041 13645 8075
rect 13645 8041 13679 8075
rect 13679 8041 13688 8075
rect 13636 8032 13688 8041
rect 17684 8032 17736 8084
rect 4344 7871 4396 7880
rect 4344 7837 4353 7871
rect 4353 7837 4387 7871
rect 4387 7837 4396 7871
rect 4344 7828 4396 7837
rect 4436 7871 4488 7880
rect 4436 7837 4445 7871
rect 4445 7837 4479 7871
rect 4479 7837 4488 7871
rect 4436 7828 4488 7837
rect 4528 7760 4580 7812
rect 5816 7828 5868 7880
rect 6552 7871 6604 7880
rect 6552 7837 6561 7871
rect 6561 7837 6595 7871
rect 6595 7837 6604 7871
rect 6552 7828 6604 7837
rect 2136 7692 2188 7744
rect 6460 7760 6512 7812
rect 5816 7692 5868 7744
rect 6368 7692 6420 7744
rect 7932 7896 7984 7948
rect 8024 7871 8076 7880
rect 8024 7837 8033 7871
rect 8033 7837 8067 7871
rect 8067 7837 8076 7871
rect 8024 7828 8076 7837
rect 9312 7896 9364 7948
rect 11704 7964 11756 8016
rect 14096 7964 14148 8016
rect 9680 7896 9732 7948
rect 7288 7803 7340 7812
rect 7288 7769 7297 7803
rect 7297 7769 7331 7803
rect 7331 7769 7340 7803
rect 7288 7760 7340 7769
rect 9036 7760 9088 7812
rect 14372 7939 14424 7948
rect 14372 7905 14381 7939
rect 14381 7905 14415 7939
rect 14415 7905 14424 7939
rect 14372 7896 14424 7905
rect 10600 7828 10652 7880
rect 10784 7828 10836 7880
rect 11980 7828 12032 7880
rect 13176 7828 13228 7880
rect 13544 7871 13596 7880
rect 13544 7837 13553 7871
rect 13553 7837 13587 7871
rect 13587 7837 13596 7871
rect 13544 7828 13596 7837
rect 14464 7871 14516 7880
rect 9864 7735 9916 7744
rect 9864 7701 9873 7735
rect 9873 7701 9907 7735
rect 9907 7701 9916 7735
rect 9864 7692 9916 7701
rect 10968 7760 11020 7812
rect 14464 7837 14473 7871
rect 14473 7837 14507 7871
rect 14507 7837 14516 7871
rect 14464 7828 14516 7837
rect 19432 7964 19484 8016
rect 16304 7896 16356 7948
rect 14832 7871 14884 7880
rect 14832 7837 14841 7871
rect 14841 7837 14875 7871
rect 14875 7837 14884 7871
rect 14832 7828 14884 7837
rect 16580 7871 16632 7880
rect 16580 7837 16589 7871
rect 16589 7837 16623 7871
rect 16623 7837 16632 7871
rect 16580 7828 16632 7837
rect 17132 7871 17184 7880
rect 10876 7692 10928 7744
rect 11152 7735 11204 7744
rect 11152 7701 11161 7735
rect 11161 7701 11195 7735
rect 11195 7701 11204 7735
rect 11152 7692 11204 7701
rect 12808 7692 12860 7744
rect 16764 7760 16816 7812
rect 17132 7837 17141 7871
rect 17141 7837 17175 7871
rect 17175 7837 17184 7871
rect 17132 7828 17184 7837
rect 17592 7871 17644 7880
rect 17592 7837 17601 7871
rect 17601 7837 17635 7871
rect 17635 7837 17644 7871
rect 17592 7828 17644 7837
rect 18604 7828 18656 7880
rect 19984 8032 20036 8084
rect 21548 8032 21600 8084
rect 21824 8032 21876 8084
rect 21272 7964 21324 8016
rect 22284 7964 22336 8016
rect 20168 7896 20220 7948
rect 22376 7896 22428 7948
rect 18420 7760 18472 7812
rect 19524 7760 19576 7812
rect 14464 7692 14516 7744
rect 14740 7692 14792 7744
rect 18696 7692 18748 7744
rect 18972 7692 19024 7744
rect 21456 7828 21508 7880
rect 22008 7828 22060 7880
rect 20076 7760 20128 7812
rect 20628 7803 20680 7812
rect 20628 7769 20637 7803
rect 20637 7769 20671 7803
rect 20671 7769 20680 7803
rect 20628 7760 20680 7769
rect 23020 7871 23072 7880
rect 23020 7837 23029 7871
rect 23029 7837 23063 7871
rect 23063 7837 23072 7871
rect 23020 7828 23072 7837
rect 22928 7760 22980 7812
rect 19984 7692 20036 7744
rect 22468 7692 22520 7744
rect 6630 7590 6682 7642
rect 6694 7590 6746 7642
rect 6758 7590 6810 7642
rect 6822 7590 6874 7642
rect 6886 7590 6938 7642
rect 12311 7590 12363 7642
rect 12375 7590 12427 7642
rect 12439 7590 12491 7642
rect 12503 7590 12555 7642
rect 12567 7590 12619 7642
rect 17992 7590 18044 7642
rect 18056 7590 18108 7642
rect 18120 7590 18172 7642
rect 18184 7590 18236 7642
rect 18248 7590 18300 7642
rect 23673 7590 23725 7642
rect 23737 7590 23789 7642
rect 23801 7590 23853 7642
rect 23865 7590 23917 7642
rect 23929 7590 23981 7642
rect 2872 7488 2924 7540
rect 4436 7420 4488 7472
rect 8576 7488 8628 7540
rect 9036 7488 9088 7540
rect 4804 7420 4856 7472
rect 9772 7420 9824 7472
rect 1768 7395 1820 7404
rect 1768 7361 1777 7395
rect 1777 7361 1811 7395
rect 1811 7361 1820 7395
rect 1768 7352 1820 7361
rect 1952 7395 2004 7404
rect 1952 7361 1965 7395
rect 1965 7361 2004 7395
rect 1952 7352 2004 7361
rect 2320 7352 2372 7404
rect 2872 7395 2924 7404
rect 2872 7361 2881 7395
rect 2881 7361 2915 7395
rect 2915 7361 2924 7395
rect 2872 7352 2924 7361
rect 4896 7352 4948 7404
rect 5080 7352 5132 7404
rect 5908 7352 5960 7404
rect 7932 7352 7984 7404
rect 8208 7395 8260 7404
rect 8208 7361 8217 7395
rect 8217 7361 8251 7395
rect 8251 7361 8260 7395
rect 8944 7395 8996 7404
rect 8208 7352 8260 7361
rect 8944 7361 8953 7395
rect 8953 7361 8987 7395
rect 8987 7361 8996 7395
rect 8944 7352 8996 7361
rect 11244 7488 11296 7540
rect 11888 7488 11940 7540
rect 12072 7488 12124 7540
rect 12716 7531 12768 7540
rect 12716 7497 12725 7531
rect 12725 7497 12759 7531
rect 12759 7497 12768 7531
rect 12716 7488 12768 7497
rect 10324 7395 10376 7404
rect 10324 7361 10333 7395
rect 10333 7361 10367 7395
rect 10367 7361 10376 7395
rect 10324 7352 10376 7361
rect 2412 7216 2464 7268
rect 4528 7259 4580 7268
rect 4528 7225 4537 7259
rect 4537 7225 4571 7259
rect 4571 7225 4580 7259
rect 4528 7216 4580 7225
rect 2964 7191 3016 7200
rect 2964 7157 2973 7191
rect 2973 7157 3007 7191
rect 3007 7157 3016 7191
rect 2964 7148 3016 7157
rect 4160 7148 4212 7200
rect 4252 7148 4304 7200
rect 5540 7216 5592 7268
rect 5908 7216 5960 7268
rect 6552 7216 6604 7268
rect 7840 7284 7892 7336
rect 7564 7216 7616 7268
rect 10140 7284 10192 7336
rect 10968 7420 11020 7472
rect 11612 7420 11664 7472
rect 14740 7463 14792 7472
rect 14740 7429 14749 7463
rect 14749 7429 14783 7463
rect 14783 7429 14792 7463
rect 14740 7420 14792 7429
rect 15476 7488 15528 7540
rect 15844 7488 15896 7540
rect 17132 7488 17184 7540
rect 12900 7395 12952 7404
rect 12900 7361 12909 7395
rect 12909 7361 12943 7395
rect 12943 7361 12952 7395
rect 12900 7352 12952 7361
rect 13176 7395 13228 7404
rect 13176 7361 13185 7395
rect 13185 7361 13219 7395
rect 13219 7361 13228 7395
rect 13176 7352 13228 7361
rect 15016 7352 15068 7404
rect 15752 7352 15804 7404
rect 16396 7352 16448 7404
rect 16948 7352 17000 7404
rect 17040 7352 17092 7404
rect 17592 7352 17644 7404
rect 22836 7488 22888 7540
rect 17868 7352 17920 7404
rect 18512 7352 18564 7404
rect 19524 7395 19576 7404
rect 19524 7361 19533 7395
rect 19533 7361 19567 7395
rect 19567 7361 19576 7395
rect 19524 7352 19576 7361
rect 19800 7395 19852 7404
rect 19800 7361 19809 7395
rect 19809 7361 19843 7395
rect 19843 7361 19852 7395
rect 19800 7352 19852 7361
rect 20628 7352 20680 7404
rect 8392 7216 8444 7268
rect 9312 7216 9364 7268
rect 9680 7216 9732 7268
rect 7840 7148 7892 7200
rect 7932 7148 7984 7200
rect 11060 7284 11112 7336
rect 10600 7216 10652 7268
rect 12164 7327 12216 7336
rect 12164 7293 12173 7327
rect 12173 7293 12207 7327
rect 12207 7293 12216 7327
rect 12164 7284 12216 7293
rect 14924 7284 14976 7336
rect 20260 7284 20312 7336
rect 21180 7284 21232 7336
rect 22468 7352 22520 7404
rect 22284 7284 22336 7336
rect 12716 7216 12768 7268
rect 16764 7216 16816 7268
rect 19248 7216 19300 7268
rect 22100 7216 22152 7268
rect 22928 7352 22980 7404
rect 10324 7191 10376 7200
rect 10324 7157 10333 7191
rect 10333 7157 10367 7191
rect 10367 7157 10376 7191
rect 10324 7148 10376 7157
rect 11704 7148 11756 7200
rect 12072 7148 12124 7200
rect 12900 7191 12952 7200
rect 12900 7157 12909 7191
rect 12909 7157 12943 7191
rect 12943 7157 12952 7191
rect 12900 7148 12952 7157
rect 13820 7191 13872 7200
rect 13820 7157 13829 7191
rect 13829 7157 13863 7191
rect 13863 7157 13872 7191
rect 13820 7148 13872 7157
rect 14648 7148 14700 7200
rect 15660 7148 15712 7200
rect 16028 7148 16080 7200
rect 18696 7148 18748 7200
rect 22376 7148 22428 7200
rect 22652 7148 22704 7200
rect 3790 7046 3842 7098
rect 3854 7046 3906 7098
rect 3918 7046 3970 7098
rect 3982 7046 4034 7098
rect 4046 7046 4098 7098
rect 9471 7046 9523 7098
rect 9535 7046 9587 7098
rect 9599 7046 9651 7098
rect 9663 7046 9715 7098
rect 9727 7046 9779 7098
rect 15152 7046 15204 7098
rect 15216 7046 15268 7098
rect 15280 7046 15332 7098
rect 15344 7046 15396 7098
rect 15408 7046 15460 7098
rect 20833 7046 20885 7098
rect 20897 7046 20949 7098
rect 20961 7046 21013 7098
rect 21025 7046 21077 7098
rect 21089 7046 21141 7098
rect 3240 6944 3292 6996
rect 7288 6944 7340 6996
rect 8392 6944 8444 6996
rect 11244 6944 11296 6996
rect 5540 6876 5592 6928
rect 4804 6808 4856 6860
rect 5356 6851 5408 6860
rect 5356 6817 5365 6851
rect 5365 6817 5399 6851
rect 5399 6817 5408 6851
rect 5356 6808 5408 6817
rect 2044 6783 2096 6792
rect 2044 6749 2053 6783
rect 2053 6749 2087 6783
rect 2087 6749 2096 6783
rect 2044 6740 2096 6749
rect 2964 6740 3016 6792
rect 2596 6647 2648 6656
rect 2596 6613 2605 6647
rect 2605 6613 2639 6647
rect 2639 6613 2648 6647
rect 2596 6604 2648 6613
rect 3240 6783 3292 6792
rect 3240 6749 3249 6783
rect 3249 6749 3283 6783
rect 3283 6749 3292 6783
rect 3240 6740 3292 6749
rect 4344 6715 4396 6724
rect 4344 6681 4353 6715
rect 4353 6681 4387 6715
rect 4387 6681 4396 6715
rect 4344 6672 4396 6681
rect 5080 6740 5132 6792
rect 5816 6851 5868 6860
rect 5816 6817 5825 6851
rect 5825 6817 5859 6851
rect 5859 6817 5868 6851
rect 5816 6808 5868 6817
rect 6000 6808 6052 6860
rect 9220 6808 9272 6860
rect 9864 6876 9916 6928
rect 6092 6783 6144 6792
rect 6092 6749 6101 6783
rect 6101 6749 6135 6783
rect 6135 6749 6144 6783
rect 6092 6740 6144 6749
rect 6276 6783 6328 6792
rect 6276 6749 6285 6783
rect 6285 6749 6319 6783
rect 6319 6749 6328 6783
rect 6276 6740 6328 6749
rect 7288 6740 7340 6792
rect 7380 6783 7432 6792
rect 7380 6749 7389 6783
rect 7389 6749 7423 6783
rect 7423 6749 7432 6783
rect 7380 6740 7432 6749
rect 5816 6672 5868 6724
rect 7748 6783 7800 6792
rect 7748 6749 7757 6783
rect 7757 6749 7791 6783
rect 7791 6749 7800 6783
rect 8300 6783 8352 6792
rect 7748 6740 7800 6749
rect 8300 6749 8309 6783
rect 8309 6749 8343 6783
rect 8343 6749 8352 6783
rect 8300 6740 8352 6749
rect 9312 6740 9364 6792
rect 9220 6672 9272 6724
rect 9956 6851 10008 6860
rect 9956 6817 9965 6851
rect 9965 6817 9999 6851
rect 9999 6817 10008 6851
rect 9956 6808 10008 6817
rect 11152 6876 11204 6928
rect 12348 6944 12400 6996
rect 12808 6944 12860 6996
rect 16396 6987 16448 6996
rect 16396 6953 16405 6987
rect 16405 6953 16439 6987
rect 16439 6953 16448 6987
rect 16396 6944 16448 6953
rect 22928 6944 22980 6996
rect 11612 6876 11664 6928
rect 13084 6876 13136 6928
rect 10600 6808 10652 6860
rect 12164 6808 12216 6860
rect 12808 6808 12860 6860
rect 9772 6783 9824 6792
rect 9772 6749 9781 6783
rect 9781 6749 9815 6783
rect 9815 6749 9824 6783
rect 9772 6740 9824 6749
rect 10416 6740 10468 6792
rect 11152 6740 11204 6792
rect 13544 6876 13596 6928
rect 15752 6876 15804 6928
rect 19064 6876 19116 6928
rect 14832 6808 14884 6860
rect 14464 6740 14516 6792
rect 16672 6808 16724 6860
rect 17316 6808 17368 6860
rect 18236 6851 18288 6860
rect 18236 6817 18245 6851
rect 18245 6817 18279 6851
rect 18279 6817 18288 6851
rect 18236 6808 18288 6817
rect 19524 6808 19576 6860
rect 18328 6783 18380 6792
rect 10968 6672 11020 6724
rect 6552 6604 6604 6656
rect 7748 6604 7800 6656
rect 10232 6604 10284 6656
rect 10600 6604 10652 6656
rect 11520 6672 11572 6724
rect 11336 6604 11388 6656
rect 11612 6604 11664 6656
rect 11704 6604 11756 6656
rect 14188 6672 14240 6724
rect 12348 6604 12400 6656
rect 14096 6604 14148 6656
rect 18328 6749 18337 6783
rect 18337 6749 18371 6783
rect 18371 6749 18380 6783
rect 18328 6740 18380 6749
rect 19248 6740 19300 6792
rect 21548 6808 21600 6860
rect 15936 6672 15988 6724
rect 16672 6672 16724 6724
rect 18512 6672 18564 6724
rect 17500 6604 17552 6656
rect 17776 6604 17828 6656
rect 18788 6604 18840 6656
rect 19156 6604 19208 6656
rect 21272 6740 21324 6792
rect 22192 6672 22244 6724
rect 23020 6876 23072 6928
rect 23204 6851 23256 6860
rect 23204 6817 23213 6851
rect 23213 6817 23247 6851
rect 23247 6817 23256 6851
rect 23204 6808 23256 6817
rect 22652 6783 22704 6792
rect 22652 6749 22661 6783
rect 22661 6749 22695 6783
rect 22695 6749 22704 6783
rect 22652 6740 22704 6749
rect 21916 6604 21968 6656
rect 6630 6502 6682 6554
rect 6694 6502 6746 6554
rect 6758 6502 6810 6554
rect 6822 6502 6874 6554
rect 6886 6502 6938 6554
rect 12311 6502 12363 6554
rect 12375 6502 12427 6554
rect 12439 6502 12491 6554
rect 12503 6502 12555 6554
rect 12567 6502 12619 6554
rect 17992 6502 18044 6554
rect 18056 6502 18108 6554
rect 18120 6502 18172 6554
rect 18184 6502 18236 6554
rect 18248 6502 18300 6554
rect 23673 6502 23725 6554
rect 23737 6502 23789 6554
rect 23801 6502 23853 6554
rect 23865 6502 23917 6554
rect 23929 6502 23981 6554
rect 4160 6375 4212 6384
rect 4160 6341 4169 6375
rect 4169 6341 4203 6375
rect 4203 6341 4212 6375
rect 4160 6332 4212 6341
rect 5080 6332 5132 6384
rect 6000 6375 6052 6384
rect 6000 6341 6009 6375
rect 6009 6341 6043 6375
rect 6043 6341 6052 6375
rect 6000 6332 6052 6341
rect 2412 6307 2464 6316
rect 2412 6273 2421 6307
rect 2421 6273 2455 6307
rect 2455 6273 2464 6307
rect 2412 6264 2464 6273
rect 2596 6264 2648 6316
rect 2780 6307 2832 6316
rect 2780 6273 2789 6307
rect 2789 6273 2823 6307
rect 2823 6273 2832 6307
rect 3056 6307 3108 6316
rect 2780 6264 2832 6273
rect 3056 6273 3065 6307
rect 3065 6273 3099 6307
rect 3099 6273 3108 6307
rect 3056 6264 3108 6273
rect 4804 6264 4856 6316
rect 5540 6307 5592 6316
rect 3700 6196 3752 6248
rect 5540 6273 5549 6307
rect 5549 6273 5583 6307
rect 5583 6273 5592 6307
rect 5540 6264 5592 6273
rect 2964 6128 3016 6180
rect 5724 6196 5776 6248
rect 6368 6400 6420 6452
rect 7012 6400 7064 6452
rect 6460 6332 6512 6384
rect 8392 6400 8444 6452
rect 8484 6400 8536 6452
rect 8300 6375 8352 6384
rect 8300 6341 8309 6375
rect 8309 6341 8343 6375
rect 8343 6341 8352 6375
rect 8300 6332 8352 6341
rect 6552 6307 6604 6316
rect 6552 6273 6561 6307
rect 6561 6273 6595 6307
rect 6595 6273 6604 6307
rect 6552 6264 6604 6273
rect 8024 6307 8076 6316
rect 8024 6273 8033 6307
rect 8033 6273 8067 6307
rect 8067 6273 8076 6307
rect 8024 6264 8076 6273
rect 6920 6196 6972 6248
rect 6276 6128 6328 6180
rect 7656 6128 7708 6180
rect 8208 6264 8260 6316
rect 8944 6400 8996 6452
rect 9680 6400 9732 6452
rect 10048 6400 10100 6452
rect 11060 6443 11112 6452
rect 11060 6409 11069 6443
rect 11069 6409 11103 6443
rect 11103 6409 11112 6443
rect 11060 6400 11112 6409
rect 8852 6332 8904 6384
rect 9956 6332 10008 6384
rect 11244 6332 11296 6384
rect 12992 6400 13044 6452
rect 13176 6400 13228 6452
rect 16028 6400 16080 6452
rect 18144 6400 18196 6452
rect 19340 6400 19392 6452
rect 21364 6400 21416 6452
rect 22928 6400 22980 6452
rect 9128 6307 9180 6316
rect 9128 6273 9137 6307
rect 9137 6273 9171 6307
rect 9171 6273 9180 6307
rect 9128 6264 9180 6273
rect 9496 6307 9548 6316
rect 9496 6273 9505 6307
rect 9505 6273 9539 6307
rect 9539 6273 9548 6307
rect 9496 6264 9548 6273
rect 10140 6264 10192 6316
rect 10232 6264 10284 6316
rect 10048 6196 10100 6248
rect 10508 6196 10560 6248
rect 11980 6264 12032 6316
rect 12164 6307 12216 6316
rect 12164 6273 12173 6307
rect 12173 6273 12207 6307
rect 12207 6273 12216 6307
rect 15016 6332 15068 6384
rect 12164 6264 12216 6273
rect 12992 6307 13044 6316
rect 12992 6273 13001 6307
rect 13001 6273 13035 6307
rect 13035 6273 13044 6307
rect 12992 6264 13044 6273
rect 13912 6307 13964 6316
rect 13912 6273 13921 6307
rect 13921 6273 13955 6307
rect 13955 6273 13964 6307
rect 13912 6264 13964 6273
rect 14188 6307 14240 6316
rect 14188 6273 14197 6307
rect 14197 6273 14231 6307
rect 14231 6273 14240 6307
rect 14188 6264 14240 6273
rect 16580 6332 16632 6384
rect 20720 6332 20772 6384
rect 12716 6196 12768 6248
rect 14096 6239 14148 6248
rect 14096 6205 14105 6239
rect 14105 6205 14139 6239
rect 14139 6205 14148 6239
rect 14096 6196 14148 6205
rect 15016 6196 15068 6248
rect 17316 6264 17368 6316
rect 17960 6307 18012 6316
rect 17960 6273 17969 6307
rect 17969 6273 18003 6307
rect 18003 6273 18012 6307
rect 18144 6307 18196 6316
rect 17960 6264 18012 6273
rect 18144 6273 18153 6307
rect 18153 6273 18187 6307
rect 18187 6273 18196 6307
rect 18144 6264 18196 6273
rect 18512 6264 18564 6316
rect 19156 6264 19208 6316
rect 18236 6196 18288 6248
rect 19892 6264 19944 6316
rect 20536 6264 20588 6316
rect 21548 6332 21600 6384
rect 21824 6264 21876 6316
rect 22192 6307 22244 6316
rect 22192 6273 22201 6307
rect 22201 6273 22235 6307
rect 22235 6273 22244 6307
rect 22192 6264 22244 6273
rect 22376 6307 22428 6316
rect 22376 6273 22385 6307
rect 22385 6273 22419 6307
rect 22419 6273 22428 6307
rect 22376 6264 22428 6273
rect 20352 6239 20404 6248
rect 20352 6205 20361 6239
rect 20361 6205 20395 6239
rect 20395 6205 20404 6239
rect 20352 6196 20404 6205
rect 22928 6307 22980 6316
rect 9128 6128 9180 6180
rect 10784 6128 10836 6180
rect 4804 6060 4856 6112
rect 7748 6060 7800 6112
rect 8392 6060 8444 6112
rect 10600 6060 10652 6112
rect 10692 6103 10744 6112
rect 10692 6069 10701 6103
rect 10701 6069 10735 6103
rect 10735 6069 10744 6103
rect 10968 6128 11020 6180
rect 12624 6171 12676 6180
rect 10692 6060 10744 6069
rect 12256 6060 12308 6112
rect 12624 6137 12633 6171
rect 12633 6137 12667 6171
rect 12667 6137 12676 6171
rect 12624 6128 12676 6137
rect 12808 6060 12860 6112
rect 14740 6128 14792 6180
rect 15476 6128 15528 6180
rect 13820 6060 13872 6112
rect 18512 6128 18564 6180
rect 18604 6128 18656 6180
rect 22928 6273 22937 6307
rect 22937 6273 22971 6307
rect 22971 6273 22980 6307
rect 22928 6264 22980 6273
rect 23112 6307 23164 6316
rect 23112 6273 23121 6307
rect 23121 6273 23155 6307
rect 23155 6273 23164 6307
rect 23112 6264 23164 6273
rect 16028 6060 16080 6112
rect 16212 6060 16264 6112
rect 19616 6060 19668 6112
rect 3790 5958 3842 6010
rect 3854 5958 3906 6010
rect 3918 5958 3970 6010
rect 3982 5958 4034 6010
rect 4046 5958 4098 6010
rect 9471 5958 9523 6010
rect 9535 5958 9587 6010
rect 9599 5958 9651 6010
rect 9663 5958 9715 6010
rect 9727 5958 9779 6010
rect 15152 5958 15204 6010
rect 15216 5958 15268 6010
rect 15280 5958 15332 6010
rect 15344 5958 15396 6010
rect 15408 5958 15460 6010
rect 20833 5958 20885 6010
rect 20897 5958 20949 6010
rect 20961 5958 21013 6010
rect 21025 5958 21077 6010
rect 21089 5958 21141 6010
rect 2044 5899 2096 5908
rect 2044 5865 2053 5899
rect 2053 5865 2087 5899
rect 2087 5865 2096 5899
rect 2044 5856 2096 5865
rect 3700 5856 3752 5908
rect 3516 5788 3568 5840
rect 6276 5831 6328 5840
rect 6276 5797 6285 5831
rect 6285 5797 6319 5831
rect 6319 5797 6328 5831
rect 6276 5788 6328 5797
rect 6920 5856 6972 5908
rect 9220 5899 9272 5908
rect 9220 5865 9229 5899
rect 9229 5865 9263 5899
rect 9263 5865 9272 5899
rect 9220 5856 9272 5865
rect 11704 5856 11756 5908
rect 12072 5856 12124 5908
rect 1768 5652 1820 5704
rect 1952 5652 2004 5704
rect 2872 5627 2924 5636
rect 2872 5593 2881 5627
rect 2881 5593 2915 5627
rect 2915 5593 2924 5627
rect 4804 5652 4856 5704
rect 5080 5695 5132 5704
rect 5080 5661 5089 5695
rect 5089 5661 5123 5695
rect 5123 5661 5132 5695
rect 5080 5652 5132 5661
rect 5264 5695 5316 5704
rect 5264 5661 5273 5695
rect 5273 5661 5307 5695
rect 5307 5661 5316 5695
rect 5264 5652 5316 5661
rect 2872 5584 2924 5593
rect 1860 5516 1912 5568
rect 2964 5559 3016 5568
rect 2964 5525 2973 5559
rect 2973 5525 3007 5559
rect 3007 5525 3016 5559
rect 2964 5516 3016 5525
rect 4988 5584 5040 5636
rect 4252 5516 4304 5568
rect 4896 5516 4948 5568
rect 6552 5652 6604 5704
rect 7840 5720 7892 5772
rect 8760 5720 8812 5772
rect 7748 5695 7800 5704
rect 7748 5661 7757 5695
rect 7757 5661 7791 5695
rect 7791 5661 7800 5695
rect 7748 5652 7800 5661
rect 7932 5695 7984 5704
rect 7932 5661 7941 5695
rect 7941 5661 7975 5695
rect 7975 5661 7984 5695
rect 7932 5652 7984 5661
rect 8116 5695 8168 5704
rect 8116 5661 8125 5695
rect 8125 5661 8159 5695
rect 8159 5661 8168 5695
rect 8116 5652 8168 5661
rect 8668 5652 8720 5704
rect 10140 5695 10192 5704
rect 10140 5661 10149 5695
rect 10149 5661 10183 5695
rect 10183 5661 10192 5695
rect 10140 5652 10192 5661
rect 10232 5695 10284 5704
rect 10232 5661 10241 5695
rect 10241 5661 10275 5695
rect 10275 5661 10284 5695
rect 11428 5788 11480 5840
rect 11612 5788 11664 5840
rect 16764 5856 16816 5908
rect 18420 5899 18472 5908
rect 18420 5865 18429 5899
rect 18429 5865 18463 5899
rect 18463 5865 18472 5899
rect 18420 5856 18472 5865
rect 14464 5788 14516 5840
rect 14740 5788 14792 5840
rect 15476 5788 15528 5840
rect 13912 5720 13964 5772
rect 10232 5652 10284 5661
rect 10508 5695 10560 5704
rect 10508 5661 10517 5695
rect 10517 5661 10551 5695
rect 10551 5661 10560 5695
rect 10508 5652 10560 5661
rect 10784 5652 10836 5704
rect 11612 5584 11664 5636
rect 7012 5516 7064 5568
rect 8484 5559 8536 5568
rect 8484 5525 8493 5559
rect 8493 5525 8527 5559
rect 8527 5525 8536 5559
rect 8484 5516 8536 5525
rect 10692 5516 10744 5568
rect 12348 5652 12400 5704
rect 15936 5720 15988 5772
rect 17868 5788 17920 5840
rect 18788 5856 18840 5908
rect 20352 5856 20404 5908
rect 21640 5899 21692 5908
rect 21640 5865 21649 5899
rect 21649 5865 21683 5899
rect 21683 5865 21692 5899
rect 21640 5856 21692 5865
rect 22376 5856 22428 5908
rect 19248 5788 19300 5840
rect 21180 5788 21232 5840
rect 17684 5720 17736 5772
rect 18328 5720 18380 5772
rect 18512 5720 18564 5772
rect 12256 5584 12308 5636
rect 11980 5516 12032 5568
rect 12992 5584 13044 5636
rect 13084 5516 13136 5568
rect 14188 5584 14240 5636
rect 14648 5584 14700 5636
rect 14832 5652 14884 5704
rect 15752 5652 15804 5704
rect 16028 5695 16080 5704
rect 16028 5661 16037 5695
rect 16037 5661 16071 5695
rect 16071 5661 16080 5695
rect 16028 5652 16080 5661
rect 16212 5695 16264 5704
rect 16212 5661 16221 5695
rect 16221 5661 16255 5695
rect 16255 5661 16264 5695
rect 16212 5652 16264 5661
rect 17316 5695 17368 5704
rect 15292 5584 15344 5636
rect 17316 5661 17325 5695
rect 17325 5661 17359 5695
rect 17359 5661 17368 5695
rect 17316 5652 17368 5661
rect 17868 5652 17920 5704
rect 20628 5720 20680 5772
rect 20444 5652 20496 5704
rect 22192 5720 22244 5772
rect 21272 5695 21324 5704
rect 21272 5661 21281 5695
rect 21281 5661 21315 5695
rect 21315 5661 21324 5695
rect 21272 5652 21324 5661
rect 21456 5652 21508 5704
rect 22928 5763 22980 5772
rect 22928 5729 22937 5763
rect 22937 5729 22971 5763
rect 22971 5729 22980 5763
rect 22928 5720 22980 5729
rect 23112 5652 23164 5704
rect 17408 5584 17460 5636
rect 17592 5516 17644 5568
rect 18788 5627 18840 5636
rect 18788 5593 18797 5627
rect 18797 5593 18831 5627
rect 18831 5593 18840 5627
rect 18788 5584 18840 5593
rect 19432 5516 19484 5568
rect 20352 5516 20404 5568
rect 22376 5516 22428 5568
rect 6630 5414 6682 5466
rect 6694 5414 6746 5466
rect 6758 5414 6810 5466
rect 6822 5414 6874 5466
rect 6886 5414 6938 5466
rect 12311 5414 12363 5466
rect 12375 5414 12427 5466
rect 12439 5414 12491 5466
rect 12503 5414 12555 5466
rect 12567 5414 12619 5466
rect 17992 5414 18044 5466
rect 18056 5414 18108 5466
rect 18120 5414 18172 5466
rect 18184 5414 18236 5466
rect 18248 5414 18300 5466
rect 23673 5414 23725 5466
rect 23737 5414 23789 5466
rect 23801 5414 23853 5466
rect 23865 5414 23917 5466
rect 23929 5414 23981 5466
rect 2964 5312 3016 5364
rect 3240 5312 3292 5364
rect 5816 5355 5868 5364
rect 4252 5244 4304 5296
rect 5816 5321 5825 5355
rect 5825 5321 5859 5355
rect 5859 5321 5868 5355
rect 5816 5312 5868 5321
rect 7380 5312 7432 5364
rect 11612 5312 11664 5364
rect 12532 5312 12584 5364
rect 13176 5312 13228 5364
rect 14372 5312 14424 5364
rect 6368 5244 6420 5296
rect 1768 5108 1820 5160
rect 2136 5176 2188 5228
rect 2320 5219 2372 5228
rect 2320 5185 2329 5219
rect 2329 5185 2363 5219
rect 2363 5185 2372 5219
rect 2320 5176 2372 5185
rect 3608 5176 3660 5228
rect 3148 5151 3200 5160
rect 3148 5117 3157 5151
rect 3157 5117 3191 5151
rect 3191 5117 3200 5151
rect 3148 5108 3200 5117
rect 4252 5108 4304 5160
rect 5264 5108 5316 5160
rect 6644 5176 6696 5228
rect 6736 5219 6788 5228
rect 6736 5185 6745 5219
rect 6745 5185 6779 5219
rect 6779 5185 6788 5219
rect 6736 5176 6788 5185
rect 7012 5176 7064 5228
rect 7748 5176 7800 5228
rect 8576 5219 8628 5228
rect 8576 5185 8585 5219
rect 8585 5185 8619 5219
rect 8619 5185 8628 5219
rect 8576 5176 8628 5185
rect 11060 5176 11112 5228
rect 13360 5176 13412 5228
rect 14096 5244 14148 5296
rect 14648 5287 14700 5296
rect 14648 5253 14657 5287
rect 14657 5253 14691 5287
rect 14691 5253 14700 5287
rect 14648 5244 14700 5253
rect 14832 5244 14884 5296
rect 14280 5176 14332 5228
rect 15292 5244 15344 5296
rect 16120 5312 16172 5364
rect 16212 5312 16264 5364
rect 17684 5312 17736 5364
rect 18788 5312 18840 5364
rect 21364 5355 21416 5364
rect 21364 5321 21373 5355
rect 21373 5321 21407 5355
rect 21407 5321 21416 5355
rect 21364 5312 21416 5321
rect 22100 5355 22152 5364
rect 22100 5321 22109 5355
rect 22109 5321 22143 5355
rect 22143 5321 22152 5355
rect 22100 5312 22152 5321
rect 18512 5244 18564 5296
rect 19524 5287 19576 5296
rect 19524 5253 19533 5287
rect 19533 5253 19567 5287
rect 19567 5253 19576 5287
rect 19524 5244 19576 5253
rect 19616 5244 19668 5296
rect 22560 5287 22612 5296
rect 22560 5253 22569 5287
rect 22569 5253 22603 5287
rect 22603 5253 22612 5287
rect 22560 5244 22612 5253
rect 6460 5108 6512 5160
rect 9680 5151 9732 5160
rect 4988 5040 5040 5092
rect 8576 5083 8628 5092
rect 8576 5049 8585 5083
rect 8585 5049 8619 5083
rect 8619 5049 8628 5083
rect 8576 5040 8628 5049
rect 9680 5117 9689 5151
rect 9689 5117 9723 5151
rect 9723 5117 9732 5151
rect 9680 5108 9732 5117
rect 12072 5108 12124 5160
rect 15752 5108 15804 5160
rect 16856 5176 16908 5228
rect 17408 5219 17460 5228
rect 17408 5185 17417 5219
rect 17417 5185 17451 5219
rect 17451 5185 17460 5219
rect 17408 5176 17460 5185
rect 17868 5176 17920 5228
rect 19432 5219 19484 5228
rect 19432 5185 19441 5219
rect 19441 5185 19475 5219
rect 19475 5185 19484 5219
rect 19432 5176 19484 5185
rect 22928 5244 22980 5296
rect 13728 5040 13780 5092
rect 17592 5108 17644 5160
rect 17684 5151 17736 5160
rect 17684 5117 17693 5151
rect 17693 5117 17727 5151
rect 17727 5117 17736 5151
rect 18328 5151 18380 5160
rect 17684 5108 17736 5117
rect 18328 5117 18337 5151
rect 18337 5117 18371 5151
rect 18371 5117 18380 5151
rect 18328 5108 18380 5117
rect 18420 5108 18472 5160
rect 3516 4972 3568 5024
rect 9128 5015 9180 5024
rect 9128 4981 9137 5015
rect 9137 4981 9171 5015
rect 9171 4981 9180 5015
rect 9128 4972 9180 4981
rect 14464 4972 14516 5024
rect 18880 5040 18932 5092
rect 23112 5176 23164 5228
rect 18696 4972 18748 5024
rect 19432 4972 19484 5024
rect 20168 4972 20220 5024
rect 3790 4870 3842 4922
rect 3854 4870 3906 4922
rect 3918 4870 3970 4922
rect 3982 4870 4034 4922
rect 4046 4870 4098 4922
rect 9471 4870 9523 4922
rect 9535 4870 9587 4922
rect 9599 4870 9651 4922
rect 9663 4870 9715 4922
rect 9727 4870 9779 4922
rect 15152 4870 15204 4922
rect 15216 4870 15268 4922
rect 15280 4870 15332 4922
rect 15344 4870 15396 4922
rect 15408 4870 15460 4922
rect 20833 4870 20885 4922
rect 20897 4870 20949 4922
rect 20961 4870 21013 4922
rect 21025 4870 21077 4922
rect 21089 4870 21141 4922
rect 2228 4768 2280 4820
rect 2780 4768 2832 4820
rect 7196 4768 7248 4820
rect 9128 4768 9180 4820
rect 10140 4768 10192 4820
rect 10784 4768 10836 4820
rect 11152 4768 11204 4820
rect 12900 4768 12952 4820
rect 13084 4768 13136 4820
rect 16212 4768 16264 4820
rect 16764 4768 16816 4820
rect 18696 4768 18748 4820
rect 20536 4811 20588 4820
rect 4344 4700 4396 4752
rect 5264 4700 5316 4752
rect 1768 4564 1820 4616
rect 2320 4607 2372 4616
rect 2320 4573 2329 4607
rect 2329 4573 2363 4607
rect 2363 4573 2372 4607
rect 2320 4564 2372 4573
rect 2412 4564 2464 4616
rect 4160 4564 4212 4616
rect 5816 4632 5868 4684
rect 5540 4564 5592 4616
rect 5724 4607 5776 4616
rect 5724 4573 5733 4607
rect 5733 4573 5767 4607
rect 5767 4573 5776 4607
rect 5724 4564 5776 4573
rect 6552 4700 6604 4752
rect 6736 4700 6788 4752
rect 10048 4743 10100 4752
rect 6092 4632 6144 4684
rect 6644 4632 6696 4684
rect 10048 4709 10057 4743
rect 10057 4709 10091 4743
rect 10091 4709 10100 4743
rect 10048 4700 10100 4709
rect 7380 4632 7432 4684
rect 3424 4471 3476 4480
rect 3424 4437 3433 4471
rect 3433 4437 3467 4471
rect 3467 4437 3476 4471
rect 3424 4428 3476 4437
rect 4160 4428 4212 4480
rect 4344 4496 4396 4548
rect 5080 4496 5132 4548
rect 5356 4496 5408 4548
rect 7932 4564 7984 4616
rect 8484 4632 8536 4684
rect 9864 4632 9916 4684
rect 10416 4632 10468 4684
rect 7564 4539 7616 4548
rect 7564 4505 7573 4539
rect 7573 4505 7607 4539
rect 7607 4505 7616 4539
rect 7564 4496 7616 4505
rect 10324 4607 10376 4616
rect 10324 4573 10333 4607
rect 10333 4573 10367 4607
rect 10367 4573 10376 4607
rect 10324 4564 10376 4573
rect 11704 4564 11756 4616
rect 12532 4700 12584 4752
rect 20536 4777 20545 4811
rect 20545 4777 20579 4811
rect 20579 4777 20588 4811
rect 20536 4768 20588 4777
rect 13452 4632 13504 4684
rect 12532 4607 12584 4616
rect 12532 4573 12541 4607
rect 12541 4573 12575 4607
rect 12575 4573 12584 4607
rect 13360 4607 13412 4616
rect 12532 4564 12584 4573
rect 13360 4573 13369 4607
rect 13369 4573 13403 4607
rect 13403 4573 13412 4607
rect 13360 4564 13412 4573
rect 13728 4607 13780 4616
rect 12072 4496 12124 4548
rect 12808 4496 12860 4548
rect 13728 4573 13737 4607
rect 13737 4573 13771 4607
rect 13771 4573 13780 4607
rect 13728 4564 13780 4573
rect 14372 4607 14424 4616
rect 14372 4573 14381 4607
rect 14381 4573 14415 4607
rect 14415 4573 14424 4607
rect 14372 4564 14424 4573
rect 16028 4564 16080 4616
rect 16212 4607 16264 4616
rect 16212 4573 16221 4607
rect 16221 4573 16255 4607
rect 16255 4573 16264 4607
rect 16212 4564 16264 4573
rect 13544 4539 13596 4548
rect 13544 4505 13553 4539
rect 13553 4505 13587 4539
rect 13587 4505 13596 4539
rect 13544 4496 13596 4505
rect 15844 4496 15896 4548
rect 16488 4607 16540 4616
rect 16488 4573 16497 4607
rect 16497 4573 16531 4607
rect 16531 4573 16540 4607
rect 16488 4564 16540 4573
rect 17316 4564 17368 4616
rect 19432 4607 19484 4616
rect 19432 4573 19441 4607
rect 19441 4573 19475 4607
rect 19475 4573 19484 4607
rect 19432 4564 19484 4573
rect 21456 4700 21508 4752
rect 22100 4675 22152 4684
rect 22100 4641 22109 4675
rect 22109 4641 22143 4675
rect 22143 4641 22152 4675
rect 22100 4632 22152 4641
rect 22376 4632 22428 4684
rect 20444 4607 20496 4616
rect 16580 4539 16632 4548
rect 16580 4505 16589 4539
rect 16589 4505 16623 4539
rect 16623 4505 16632 4539
rect 16580 4496 16632 4505
rect 16948 4496 17000 4548
rect 4436 4428 4488 4480
rect 9312 4428 9364 4480
rect 11980 4428 12032 4480
rect 15752 4428 15804 4480
rect 18604 4428 18656 4480
rect 20444 4573 20453 4607
rect 20453 4573 20487 4607
rect 20487 4573 20496 4607
rect 20444 4564 20496 4573
rect 23112 4564 23164 4616
rect 20812 4496 20864 4548
rect 6630 4326 6682 4378
rect 6694 4326 6746 4378
rect 6758 4326 6810 4378
rect 6822 4326 6874 4378
rect 6886 4326 6938 4378
rect 12311 4326 12363 4378
rect 12375 4326 12427 4378
rect 12439 4326 12491 4378
rect 12503 4326 12555 4378
rect 12567 4326 12619 4378
rect 17992 4326 18044 4378
rect 18056 4326 18108 4378
rect 18120 4326 18172 4378
rect 18184 4326 18236 4378
rect 18248 4326 18300 4378
rect 23673 4326 23725 4378
rect 23737 4326 23789 4378
rect 23801 4326 23853 4378
rect 23865 4326 23917 4378
rect 23929 4326 23981 4378
rect 7012 4224 7064 4276
rect 8484 4267 8536 4276
rect 8484 4233 8493 4267
rect 8493 4233 8527 4267
rect 8527 4233 8536 4267
rect 8484 4224 8536 4233
rect 10324 4224 10376 4276
rect 12072 4267 12124 4276
rect 12072 4233 12081 4267
rect 12081 4233 12115 4267
rect 12115 4233 12124 4267
rect 12072 4224 12124 4233
rect 14372 4224 14424 4276
rect 14556 4267 14608 4276
rect 14556 4233 14565 4267
rect 14565 4233 14599 4267
rect 14599 4233 14608 4267
rect 14556 4224 14608 4233
rect 16028 4224 16080 4276
rect 18328 4224 18380 4276
rect 18512 4267 18564 4276
rect 18512 4233 18521 4267
rect 18521 4233 18555 4267
rect 18555 4233 18564 4267
rect 18512 4224 18564 4233
rect 2320 4156 2372 4208
rect 4436 4156 4488 4208
rect 6368 4156 6420 4208
rect 6552 4156 6604 4208
rect 1860 4131 1912 4140
rect 1860 4097 1869 4131
rect 1869 4097 1903 4131
rect 1903 4097 1912 4131
rect 1860 4088 1912 4097
rect 2044 4088 2096 4140
rect 2596 4131 2648 4140
rect 2596 4097 2605 4131
rect 2605 4097 2639 4131
rect 2639 4097 2648 4131
rect 2596 4088 2648 4097
rect 4252 4088 4304 4140
rect 1952 3952 2004 4004
rect 3700 4020 3752 4072
rect 4896 4088 4948 4140
rect 5356 4131 5408 4140
rect 5356 4097 5365 4131
rect 5365 4097 5399 4131
rect 5399 4097 5408 4131
rect 7564 4156 7616 4208
rect 9036 4156 9088 4208
rect 5356 4088 5408 4097
rect 5448 4020 5500 4072
rect 1676 3927 1728 3936
rect 1676 3893 1685 3927
rect 1685 3893 1719 3927
rect 1719 3893 1728 3927
rect 1676 3884 1728 3893
rect 1860 3884 1912 3936
rect 4160 3952 4212 4004
rect 4988 3952 5040 4004
rect 8300 4088 8352 4140
rect 8668 4088 8720 4140
rect 10692 4131 10744 4140
rect 7196 4063 7248 4072
rect 7196 4029 7205 4063
rect 7205 4029 7239 4063
rect 7239 4029 7248 4063
rect 7196 4020 7248 4029
rect 8208 4020 8260 4072
rect 10692 4097 10701 4131
rect 10701 4097 10735 4131
rect 10735 4097 10744 4131
rect 10692 4088 10744 4097
rect 10784 4131 10836 4140
rect 10784 4097 10793 4131
rect 10793 4097 10827 4131
rect 10827 4097 10836 4131
rect 11704 4131 11756 4140
rect 10784 4088 10836 4097
rect 11704 4097 11713 4131
rect 11713 4097 11747 4131
rect 11747 4097 11756 4131
rect 11704 4088 11756 4097
rect 13820 4156 13872 4208
rect 14096 4088 14148 4140
rect 15752 4131 15804 4140
rect 8944 4020 8996 4072
rect 10968 4020 11020 4072
rect 7288 3952 7340 4004
rect 9220 3952 9272 4004
rect 12072 4020 12124 4072
rect 2872 3927 2924 3936
rect 2872 3893 2881 3927
rect 2881 3893 2915 3927
rect 2915 3893 2924 3927
rect 2872 3884 2924 3893
rect 3424 3884 3476 3936
rect 4344 3884 4396 3936
rect 7012 3884 7064 3936
rect 9128 3884 9180 3936
rect 12164 3952 12216 4004
rect 14740 4020 14792 4072
rect 14924 4020 14976 4072
rect 15752 4097 15761 4131
rect 15761 4097 15795 4131
rect 15795 4097 15804 4131
rect 15752 4088 15804 4097
rect 15936 4131 15988 4140
rect 15936 4097 15945 4131
rect 15945 4097 15979 4131
rect 15979 4097 15988 4131
rect 15936 4088 15988 4097
rect 16120 4131 16172 4140
rect 16120 4097 16129 4131
rect 16129 4097 16163 4131
rect 16163 4097 16172 4131
rect 16120 4088 16172 4097
rect 17500 4088 17552 4140
rect 18052 4088 18104 4140
rect 18880 4199 18932 4208
rect 18880 4165 18889 4199
rect 18889 4165 18923 4199
rect 18923 4165 18932 4199
rect 18880 4156 18932 4165
rect 19064 4131 19116 4140
rect 19064 4097 19073 4131
rect 19073 4097 19107 4131
rect 19107 4097 19116 4131
rect 19064 4088 19116 4097
rect 19984 4131 20036 4140
rect 19984 4097 19993 4131
rect 19993 4097 20027 4131
rect 20027 4097 20036 4131
rect 19984 4088 20036 4097
rect 20168 4131 20220 4140
rect 20168 4097 20177 4131
rect 20177 4097 20211 4131
rect 20211 4097 20220 4131
rect 20168 4088 20220 4097
rect 20352 4131 20404 4140
rect 20352 4097 20361 4131
rect 20361 4097 20395 4131
rect 20395 4097 20404 4131
rect 20352 4088 20404 4097
rect 20536 4131 20588 4140
rect 20536 4097 20545 4131
rect 20545 4097 20579 4131
rect 20579 4097 20588 4131
rect 20536 4088 20588 4097
rect 20812 4131 20864 4140
rect 20812 4097 20821 4131
rect 20821 4097 20855 4131
rect 20855 4097 20864 4131
rect 20812 4088 20864 4097
rect 21180 4088 21232 4140
rect 22468 4088 22520 4140
rect 18512 4020 18564 4072
rect 16948 3952 17000 4004
rect 17868 3952 17920 4004
rect 12808 3884 12860 3936
rect 13636 3884 13688 3936
rect 16580 3884 16632 3936
rect 18696 3884 18748 3936
rect 22376 3884 22428 3936
rect 3790 3782 3842 3834
rect 3854 3782 3906 3834
rect 3918 3782 3970 3834
rect 3982 3782 4034 3834
rect 4046 3782 4098 3834
rect 9471 3782 9523 3834
rect 9535 3782 9587 3834
rect 9599 3782 9651 3834
rect 9663 3782 9715 3834
rect 9727 3782 9779 3834
rect 15152 3782 15204 3834
rect 15216 3782 15268 3834
rect 15280 3782 15332 3834
rect 15344 3782 15396 3834
rect 15408 3782 15460 3834
rect 20833 3782 20885 3834
rect 20897 3782 20949 3834
rect 20961 3782 21013 3834
rect 21025 3782 21077 3834
rect 21089 3782 21141 3834
rect 2596 3680 2648 3732
rect 2780 3612 2832 3664
rect 1676 3476 1728 3528
rect 2596 3476 2648 3528
rect 2688 3519 2740 3528
rect 2688 3485 2697 3519
rect 2697 3485 2731 3519
rect 2731 3485 2740 3519
rect 2688 3476 2740 3485
rect 3424 3476 3476 3528
rect 4344 3680 4396 3732
rect 9220 3680 9272 3732
rect 9312 3680 9364 3732
rect 9588 3680 9640 3732
rect 13360 3680 13412 3732
rect 13544 3680 13596 3732
rect 14556 3680 14608 3732
rect 6460 3612 6512 3664
rect 8484 3612 8536 3664
rect 15936 3680 15988 3732
rect 18144 3680 18196 3732
rect 21824 3723 21876 3732
rect 18788 3612 18840 3664
rect 4988 3587 5040 3596
rect 4988 3553 4997 3587
rect 4997 3553 5031 3587
rect 5031 3553 5040 3587
rect 4988 3544 5040 3553
rect 5356 3544 5408 3596
rect 3976 3476 4028 3528
rect 5172 3476 5224 3528
rect 6552 3544 6604 3596
rect 10600 3544 10652 3596
rect 12072 3587 12124 3596
rect 7380 3476 7432 3528
rect 8300 3519 8352 3528
rect 8300 3485 8309 3519
rect 8309 3485 8343 3519
rect 8343 3485 8352 3519
rect 8300 3476 8352 3485
rect 8484 3519 8536 3528
rect 8484 3485 8493 3519
rect 8493 3485 8527 3519
rect 8527 3485 8536 3519
rect 8484 3476 8536 3485
rect 8944 3476 8996 3528
rect 9128 3519 9180 3528
rect 9128 3485 9137 3519
rect 9137 3485 9171 3519
rect 9171 3485 9180 3519
rect 9128 3476 9180 3485
rect 9312 3519 9364 3528
rect 9312 3485 9321 3519
rect 9321 3485 9355 3519
rect 9355 3485 9364 3519
rect 9312 3476 9364 3485
rect 9496 3476 9548 3528
rect 11704 3519 11756 3528
rect 11704 3485 11713 3519
rect 11713 3485 11747 3519
rect 11747 3485 11756 3519
rect 11704 3476 11756 3485
rect 12072 3553 12081 3587
rect 12081 3553 12115 3587
rect 12115 3553 12124 3587
rect 12072 3544 12124 3553
rect 12256 3587 12308 3596
rect 12256 3553 12265 3587
rect 12265 3553 12299 3587
rect 12299 3553 12308 3587
rect 12256 3544 12308 3553
rect 13452 3519 13504 3528
rect 13452 3485 13461 3519
rect 13461 3485 13495 3519
rect 13495 3485 13504 3519
rect 13452 3476 13504 3485
rect 13544 3519 13596 3528
rect 13544 3485 13553 3519
rect 13553 3485 13587 3519
rect 13587 3485 13596 3519
rect 15752 3544 15804 3596
rect 13544 3476 13596 3485
rect 15844 3519 15896 3528
rect 3332 3451 3384 3460
rect 3332 3417 3341 3451
rect 3341 3417 3375 3451
rect 3375 3417 3384 3451
rect 3332 3408 3384 3417
rect 4896 3451 4948 3460
rect 4896 3417 4905 3451
rect 4905 3417 4939 3451
rect 4939 3417 4948 3451
rect 4896 3408 4948 3417
rect 5816 3408 5868 3460
rect 13360 3408 13412 3460
rect 15844 3485 15853 3519
rect 15853 3485 15887 3519
rect 15887 3485 15896 3519
rect 15844 3476 15896 3485
rect 16120 3519 16172 3528
rect 16120 3485 16129 3519
rect 16129 3485 16163 3519
rect 16163 3485 16172 3519
rect 16120 3476 16172 3485
rect 16580 3519 16632 3528
rect 16580 3485 16589 3519
rect 16589 3485 16623 3519
rect 16623 3485 16632 3519
rect 16580 3476 16632 3485
rect 16948 3519 17000 3528
rect 16948 3485 16957 3519
rect 16957 3485 16991 3519
rect 16991 3485 17000 3519
rect 16948 3476 17000 3485
rect 18144 3544 18196 3596
rect 18696 3587 18748 3596
rect 18696 3553 18705 3587
rect 18705 3553 18739 3587
rect 18739 3553 18748 3587
rect 18696 3544 18748 3553
rect 21824 3689 21833 3723
rect 21833 3689 21867 3723
rect 21867 3689 21876 3723
rect 21824 3680 21876 3689
rect 22376 3723 22428 3732
rect 22376 3689 22385 3723
rect 22385 3689 22419 3723
rect 22419 3689 22428 3723
rect 22376 3680 22428 3689
rect 19340 3612 19392 3664
rect 20536 3544 20588 3596
rect 7564 3340 7616 3392
rect 7656 3340 7708 3392
rect 11152 3383 11204 3392
rect 11152 3349 11161 3383
rect 11161 3349 11195 3383
rect 11195 3349 11204 3383
rect 11152 3340 11204 3349
rect 11244 3340 11296 3392
rect 12256 3340 12308 3392
rect 13452 3340 13504 3392
rect 14648 3340 14700 3392
rect 18052 3476 18104 3528
rect 18236 3519 18288 3528
rect 18236 3485 18245 3519
rect 18245 3485 18279 3519
rect 18279 3485 18288 3519
rect 18236 3476 18288 3485
rect 18512 3519 18564 3528
rect 18512 3485 18547 3519
rect 18547 3485 18564 3519
rect 18512 3476 18564 3485
rect 18788 3476 18840 3528
rect 19984 3476 20036 3528
rect 20168 3519 20220 3528
rect 20168 3485 20177 3519
rect 20177 3485 20211 3519
rect 20211 3485 20220 3519
rect 20168 3476 20220 3485
rect 20352 3519 20404 3528
rect 20352 3485 20361 3519
rect 20361 3485 20395 3519
rect 20395 3485 20404 3519
rect 20352 3476 20404 3485
rect 21180 3519 21232 3528
rect 21180 3485 21189 3519
rect 21189 3485 21223 3519
rect 21223 3485 21232 3519
rect 21180 3476 21232 3485
rect 23388 3476 23440 3528
rect 17868 3408 17920 3460
rect 18880 3408 18932 3460
rect 6630 3238 6682 3290
rect 6694 3238 6746 3290
rect 6758 3238 6810 3290
rect 6822 3238 6874 3290
rect 6886 3238 6938 3290
rect 12311 3238 12363 3290
rect 12375 3238 12427 3290
rect 12439 3238 12491 3290
rect 12503 3238 12555 3290
rect 12567 3238 12619 3290
rect 17992 3238 18044 3290
rect 18056 3238 18108 3290
rect 18120 3238 18172 3290
rect 18184 3238 18236 3290
rect 18248 3238 18300 3290
rect 23673 3238 23725 3290
rect 23737 3238 23789 3290
rect 23801 3238 23853 3290
rect 23865 3238 23917 3290
rect 23929 3238 23981 3290
rect 1860 3136 1912 3188
rect 2596 3179 2648 3188
rect 1952 3000 2004 3052
rect 2596 3145 2605 3179
rect 2605 3145 2639 3179
rect 2639 3145 2648 3179
rect 2596 3136 2648 3145
rect 5540 3136 5592 3188
rect 8208 3136 8260 3188
rect 5356 3068 5408 3120
rect 2504 3000 2556 3052
rect 3516 3043 3568 3052
rect 3516 3009 3525 3043
rect 3525 3009 3559 3043
rect 3559 3009 3568 3043
rect 3516 3000 3568 3009
rect 3976 3043 4028 3052
rect 3976 3009 3985 3043
rect 3985 3009 4019 3043
rect 4019 3009 4028 3043
rect 3976 3000 4028 3009
rect 4252 3000 4304 3052
rect 4436 3043 4488 3052
rect 4436 3009 4445 3043
rect 4445 3009 4479 3043
rect 4479 3009 4488 3043
rect 4436 3000 4488 3009
rect 5724 3000 5776 3052
rect 5816 3043 5868 3052
rect 5816 3009 5825 3043
rect 5825 3009 5859 3043
rect 5859 3009 5868 3043
rect 7012 3043 7064 3052
rect 5816 3000 5868 3009
rect 7012 3009 7021 3043
rect 7021 3009 7055 3043
rect 7055 3009 7064 3043
rect 7012 3000 7064 3009
rect 9312 3136 9364 3188
rect 9588 3136 9640 3188
rect 9864 3179 9916 3188
rect 9864 3145 9873 3179
rect 9873 3145 9907 3179
rect 9907 3145 9916 3179
rect 9864 3136 9916 3145
rect 8576 3068 8628 3120
rect 11244 3136 11296 3188
rect 11428 3136 11480 3188
rect 12348 3136 12400 3188
rect 13544 3136 13596 3188
rect 13636 3179 13688 3188
rect 13636 3145 13645 3179
rect 13645 3145 13679 3179
rect 13679 3145 13688 3179
rect 13636 3136 13688 3145
rect 14556 3136 14608 3188
rect 14740 3179 14792 3188
rect 14740 3145 14749 3179
rect 14749 3145 14783 3179
rect 14783 3145 14792 3179
rect 14740 3136 14792 3145
rect 16856 3179 16908 3188
rect 16856 3145 16865 3179
rect 16865 3145 16899 3179
rect 16899 3145 16908 3179
rect 16856 3136 16908 3145
rect 18328 3136 18380 3188
rect 19524 3136 19576 3188
rect 10692 3068 10744 3120
rect 10600 3043 10652 3052
rect 3424 2932 3476 2984
rect 5448 2932 5500 2984
rect 5632 2975 5684 2984
rect 5632 2941 5641 2975
rect 5641 2941 5675 2975
rect 5675 2941 5684 2975
rect 5632 2932 5684 2941
rect 10600 3009 10609 3043
rect 10609 3009 10643 3043
rect 10643 3009 10652 3043
rect 10600 3000 10652 3009
rect 11060 3000 11112 3052
rect 12164 3000 12216 3052
rect 13268 3000 13320 3052
rect 14648 3043 14700 3052
rect 14648 3009 14657 3043
rect 14657 3009 14691 3043
rect 14691 3009 14700 3043
rect 14648 3000 14700 3009
rect 14832 3043 14884 3052
rect 14832 3009 14841 3043
rect 14841 3009 14875 3043
rect 14875 3009 14884 3043
rect 14832 3000 14884 3009
rect 17040 3043 17092 3052
rect 2136 2864 2188 2916
rect 3148 2864 3200 2916
rect 4160 2796 4212 2848
rect 4896 2864 4948 2916
rect 8576 2864 8628 2916
rect 11428 2932 11480 2984
rect 12072 2932 12124 2984
rect 17040 3009 17049 3043
rect 17049 3009 17083 3043
rect 17083 3009 17092 3043
rect 17868 3068 17920 3120
rect 18604 3111 18656 3120
rect 18604 3077 18613 3111
rect 18613 3077 18647 3111
rect 18647 3077 18656 3111
rect 18604 3068 18656 3077
rect 17316 3043 17368 3052
rect 17040 3000 17092 3009
rect 17316 3009 17325 3043
rect 17325 3009 17359 3043
rect 17359 3009 17368 3043
rect 17316 3000 17368 3009
rect 18696 3043 18748 3052
rect 18696 3009 18705 3043
rect 18705 3009 18739 3043
rect 18739 3009 18748 3043
rect 20628 3068 20680 3120
rect 18696 3000 18748 3009
rect 19064 2932 19116 2984
rect 11244 2864 11296 2916
rect 17592 2864 17644 2916
rect 19432 2864 19484 2916
rect 20168 2864 20220 2916
rect 4988 2796 5040 2848
rect 6092 2796 6144 2848
rect 10416 2796 10468 2848
rect 15752 2796 15804 2848
rect 18328 2796 18380 2848
rect 21456 2796 21508 2848
rect 22744 2796 22796 2848
rect 3790 2694 3842 2746
rect 3854 2694 3906 2746
rect 3918 2694 3970 2746
rect 3982 2694 4034 2746
rect 4046 2694 4098 2746
rect 9471 2694 9523 2746
rect 9535 2694 9587 2746
rect 9599 2694 9651 2746
rect 9663 2694 9715 2746
rect 9727 2694 9779 2746
rect 15152 2694 15204 2746
rect 15216 2694 15268 2746
rect 15280 2694 15332 2746
rect 15344 2694 15396 2746
rect 15408 2694 15460 2746
rect 20833 2694 20885 2746
rect 20897 2694 20949 2746
rect 20961 2694 21013 2746
rect 21025 2694 21077 2746
rect 21089 2694 21141 2746
rect 4436 2592 4488 2644
rect 4896 2524 4948 2576
rect 5816 2592 5868 2644
rect 6184 2592 6236 2644
rect 2780 2320 2832 2372
rect 4160 2388 4212 2440
rect 4344 2388 4396 2440
rect 5172 2431 5224 2440
rect 5172 2397 5181 2431
rect 5181 2397 5215 2431
rect 5215 2397 5224 2431
rect 5172 2388 5224 2397
rect 6460 2388 6512 2440
rect 7380 2388 7432 2440
rect 12348 2592 12400 2644
rect 14464 2592 14516 2644
rect 17316 2592 17368 2644
rect 18604 2592 18656 2644
rect 19432 2635 19484 2644
rect 19432 2601 19441 2635
rect 19441 2601 19475 2635
rect 19475 2601 19484 2635
rect 19432 2592 19484 2601
rect 20628 2592 20680 2644
rect 7656 2499 7708 2508
rect 7656 2465 7665 2499
rect 7665 2465 7699 2499
rect 7699 2465 7708 2499
rect 7656 2456 7708 2465
rect 16304 2456 16356 2508
rect 18880 2456 18932 2508
rect 9220 2388 9272 2440
rect 9864 2431 9916 2440
rect 9864 2397 9873 2431
rect 9873 2397 9907 2431
rect 9907 2397 9916 2431
rect 9864 2388 9916 2397
rect 10508 2431 10560 2440
rect 10508 2397 10517 2431
rect 10517 2397 10551 2431
rect 10551 2397 10560 2431
rect 10508 2388 10560 2397
rect 11152 2431 11204 2440
rect 11152 2397 11161 2431
rect 11161 2397 11195 2431
rect 11195 2397 11204 2431
rect 11152 2388 11204 2397
rect 11796 2388 11848 2440
rect 12716 2388 12768 2440
rect 13084 2388 13136 2440
rect 13728 2388 13780 2440
rect 14372 2388 14424 2440
rect 15016 2388 15068 2440
rect 15660 2388 15712 2440
rect 16948 2388 17000 2440
rect 19524 2388 19576 2440
rect 20812 2388 20864 2440
rect 22100 2388 22152 2440
rect 6000 2320 6052 2372
rect 4712 2252 4764 2304
rect 6630 2150 6682 2202
rect 6694 2150 6746 2202
rect 6758 2150 6810 2202
rect 6822 2150 6874 2202
rect 6886 2150 6938 2202
rect 12311 2150 12363 2202
rect 12375 2150 12427 2202
rect 12439 2150 12491 2202
rect 12503 2150 12555 2202
rect 12567 2150 12619 2202
rect 17992 2150 18044 2202
rect 18056 2150 18108 2202
rect 18120 2150 18172 2202
rect 18184 2150 18236 2202
rect 18248 2150 18300 2202
rect 23673 2150 23725 2202
rect 23737 2150 23789 2202
rect 23801 2150 23853 2202
rect 23865 2150 23917 2202
rect 23929 2150 23981 2202
rect 1492 1164 1544 1216
rect 7656 1164 7708 1216
<< metal2 >>
rect 2502 24200 2558 25000
rect 7470 24200 7526 25000
rect 12438 24200 12494 25000
rect 17406 24200 17462 25000
rect 22374 24200 22430 25000
rect 2516 21690 2544 24200
rect 3790 22332 4098 22341
rect 3790 22330 3796 22332
rect 3852 22330 3876 22332
rect 3932 22330 3956 22332
rect 4012 22330 4036 22332
rect 4092 22330 4098 22332
rect 3852 22278 3854 22330
rect 4034 22278 4036 22330
rect 3790 22276 3796 22278
rect 3852 22276 3876 22278
rect 3932 22276 3956 22278
rect 4012 22276 4036 22278
rect 4092 22276 4098 22278
rect 3790 22267 4098 22276
rect 7484 21962 7512 24200
rect 9471 22332 9779 22341
rect 9471 22330 9477 22332
rect 9533 22330 9557 22332
rect 9613 22330 9637 22332
rect 9693 22330 9717 22332
rect 9773 22330 9779 22332
rect 9533 22278 9535 22330
rect 9715 22278 9717 22330
rect 9471 22276 9477 22278
rect 9533 22276 9557 22278
rect 9613 22276 9637 22278
rect 9693 22276 9717 22278
rect 9773 22276 9779 22278
rect 9471 22267 9779 22276
rect 10508 22024 10560 22030
rect 10508 21966 10560 21972
rect 7472 21956 7524 21962
rect 7472 21898 7524 21904
rect 6276 21888 6328 21894
rect 6276 21830 6328 21836
rect 8944 21888 8996 21894
rect 8944 21830 8996 21836
rect 2504 21684 2556 21690
rect 2504 21626 2556 21632
rect 5816 21684 5868 21690
rect 5816 21626 5868 21632
rect 5356 21616 5408 21622
rect 5356 21558 5408 21564
rect 5446 21584 5502 21593
rect 2780 21548 2832 21554
rect 2780 21490 2832 21496
rect 2044 21480 2096 21486
rect 2044 21422 2096 21428
rect 1860 21344 1912 21350
rect 1860 21286 1912 21292
rect 1676 20868 1728 20874
rect 1676 20810 1728 20816
rect 1584 19780 1636 19786
rect 1584 19722 1636 19728
rect 1596 12442 1624 19722
rect 1688 14618 1716 20810
rect 1872 15094 1900 21286
rect 2056 20942 2084 21422
rect 2044 20936 2096 20942
rect 2044 20878 2096 20884
rect 2056 20398 2084 20878
rect 2044 20392 2096 20398
rect 2044 20334 2096 20340
rect 2056 19922 2084 20334
rect 2044 19916 2096 19922
rect 2044 19858 2096 19864
rect 2792 19394 2820 21490
rect 3790 21244 4098 21253
rect 3790 21242 3796 21244
rect 3852 21242 3876 21244
rect 3932 21242 3956 21244
rect 4012 21242 4036 21244
rect 4092 21242 4098 21244
rect 3852 21190 3854 21242
rect 4034 21190 4036 21242
rect 3790 21188 3796 21190
rect 3852 21188 3876 21190
rect 3932 21188 3956 21190
rect 4012 21188 4036 21190
rect 4092 21188 4098 21190
rect 3790 21179 4098 21188
rect 5368 21010 5396 21558
rect 5446 21519 5448 21528
rect 5500 21519 5502 21528
rect 5448 21490 5500 21496
rect 5356 21004 5408 21010
rect 5356 20946 5408 20952
rect 4712 20868 4764 20874
rect 4712 20810 4764 20816
rect 3148 20800 3200 20806
rect 3148 20742 3200 20748
rect 3516 20800 3568 20806
rect 3516 20742 3568 20748
rect 2792 19366 2912 19394
rect 2780 19304 2832 19310
rect 2780 19246 2832 19252
rect 2792 18766 2820 19246
rect 2780 18760 2832 18766
rect 2780 18702 2832 18708
rect 2596 18624 2648 18630
rect 2596 18566 2648 18572
rect 2320 18284 2372 18290
rect 2320 18226 2372 18232
rect 2228 15360 2280 15366
rect 2228 15302 2280 15308
rect 1860 15088 1912 15094
rect 1860 15030 1912 15036
rect 2136 15088 2188 15094
rect 2136 15030 2188 15036
rect 1768 15020 1820 15026
rect 1768 14962 1820 14968
rect 1676 14612 1728 14618
rect 1676 14554 1728 14560
rect 1584 12436 1636 12442
rect 1584 12378 1636 12384
rect 1676 12096 1728 12102
rect 1676 12038 1728 12044
rect 1688 11762 1716 12038
rect 1780 11898 1808 14962
rect 1952 14340 2004 14346
rect 1952 14282 2004 14288
rect 1860 13864 1912 13870
rect 1860 13806 1912 13812
rect 1768 11892 1820 11898
rect 1768 11834 1820 11840
rect 1676 11756 1728 11762
rect 1676 11698 1728 11704
rect 1872 11694 1900 13806
rect 1964 12866 1992 14282
rect 2044 13728 2096 13734
rect 2044 13670 2096 13676
rect 2056 12986 2084 13670
rect 2044 12980 2096 12986
rect 2044 12922 2096 12928
rect 1964 12838 2084 12866
rect 1952 12640 2004 12646
rect 1952 12582 2004 12588
rect 1964 12170 1992 12582
rect 2056 12374 2084 12838
rect 2044 12368 2096 12374
rect 2044 12310 2096 12316
rect 1952 12164 2004 12170
rect 1952 12106 2004 12112
rect 1964 11694 1992 12106
rect 1860 11688 1912 11694
rect 1860 11630 1912 11636
rect 1952 11688 2004 11694
rect 1952 11630 2004 11636
rect 1872 11286 1900 11630
rect 1860 11280 1912 11286
rect 1860 11222 1912 11228
rect 1584 11144 1636 11150
rect 1584 11086 1636 11092
rect 1596 10810 1624 11086
rect 1584 10804 1636 10810
rect 1584 10746 1636 10752
rect 1676 9920 1728 9926
rect 1676 9862 1728 9868
rect 1688 9178 1716 9862
rect 1964 9518 1992 11630
rect 2056 10742 2084 12310
rect 2148 12238 2176 15030
rect 2240 14414 2268 15302
rect 2332 15065 2360 18226
rect 2412 17604 2464 17610
rect 2412 17546 2464 17552
rect 2318 15056 2374 15065
rect 2318 14991 2320 15000
rect 2372 14991 2374 15000
rect 2320 14962 2372 14968
rect 2332 14414 2360 14962
rect 2228 14408 2280 14414
rect 2228 14350 2280 14356
rect 2320 14408 2372 14414
rect 2320 14350 2372 14356
rect 2320 13796 2372 13802
rect 2320 13738 2372 13744
rect 2332 13326 2360 13738
rect 2320 13320 2372 13326
rect 2320 13262 2372 13268
rect 2136 12232 2188 12238
rect 2136 12174 2188 12180
rect 2320 12232 2372 12238
rect 2320 12174 2372 12180
rect 2228 12096 2280 12102
rect 2228 12038 2280 12044
rect 2136 11552 2188 11558
rect 2136 11494 2188 11500
rect 2044 10736 2096 10742
rect 2044 10678 2096 10684
rect 2148 10470 2176 11494
rect 2136 10464 2188 10470
rect 2136 10406 2188 10412
rect 2240 9586 2268 12038
rect 2332 10606 2360 12174
rect 2424 11234 2452 17546
rect 2504 15496 2556 15502
rect 2504 15438 2556 15444
rect 2516 13938 2544 15438
rect 2504 13932 2556 13938
rect 2504 13874 2556 13880
rect 2516 13530 2544 13874
rect 2504 13524 2556 13530
rect 2504 13466 2556 13472
rect 2516 11898 2544 13466
rect 2608 12918 2636 18566
rect 2792 18222 2820 18702
rect 2780 18216 2832 18222
rect 2700 18176 2780 18204
rect 2700 17678 2728 18176
rect 2780 18158 2832 18164
rect 2688 17672 2740 17678
rect 2688 17614 2740 17620
rect 2700 17134 2728 17614
rect 2688 17128 2740 17134
rect 2688 17070 2740 17076
rect 2700 16590 2728 17070
rect 2688 16584 2740 16590
rect 2688 16526 2740 16532
rect 2780 16516 2832 16522
rect 2780 16458 2832 16464
rect 2688 15972 2740 15978
rect 2688 15914 2740 15920
rect 2700 15434 2728 15914
rect 2688 15428 2740 15434
rect 2688 15370 2740 15376
rect 2688 14408 2740 14414
rect 2688 14350 2740 14356
rect 2700 13326 2728 14350
rect 2792 13818 2820 16458
rect 2884 14822 2912 19366
rect 2964 17536 3016 17542
rect 2964 17478 3016 17484
rect 2872 14816 2924 14822
rect 2872 14758 2924 14764
rect 2872 14272 2924 14278
rect 2872 14214 2924 14220
rect 2884 14006 2912 14214
rect 2872 14000 2924 14006
rect 2872 13942 2924 13948
rect 2976 13954 3004 17478
rect 3056 16584 3108 16590
rect 3056 16526 3108 16532
rect 3068 15910 3096 16526
rect 3160 15978 3188 20742
rect 3424 19372 3476 19378
rect 3424 19314 3476 19320
rect 3332 18080 3384 18086
rect 3332 18022 3384 18028
rect 3148 15972 3200 15978
rect 3148 15914 3200 15920
rect 3056 15904 3108 15910
rect 3056 15846 3108 15852
rect 3068 15570 3096 15846
rect 3056 15564 3108 15570
rect 3056 15506 3108 15512
rect 3068 15026 3096 15506
rect 3344 15434 3372 18022
rect 3332 15428 3384 15434
rect 3332 15370 3384 15376
rect 3148 15360 3200 15366
rect 3148 15302 3200 15308
rect 3160 15144 3188 15302
rect 3240 15156 3292 15162
rect 3160 15116 3240 15144
rect 3056 15020 3108 15026
rect 3056 14962 3108 14968
rect 3068 14074 3096 14962
rect 3160 14822 3188 15116
rect 3240 15098 3292 15104
rect 3148 14816 3200 14822
rect 3148 14758 3200 14764
rect 3240 14476 3292 14482
rect 3160 14436 3240 14464
rect 3056 14068 3108 14074
rect 3056 14010 3108 14016
rect 2976 13926 3096 13954
rect 2792 13790 3004 13818
rect 2688 13320 2740 13326
rect 2688 13262 2740 13268
rect 2780 13252 2832 13258
rect 2780 13194 2832 13200
rect 2792 12918 2820 13194
rect 2596 12912 2648 12918
rect 2596 12854 2648 12860
rect 2780 12912 2832 12918
rect 2780 12854 2832 12860
rect 2688 12844 2740 12850
rect 2688 12786 2740 12792
rect 2596 12640 2648 12646
rect 2596 12582 2648 12588
rect 2608 12306 2636 12582
rect 2596 12300 2648 12306
rect 2596 12242 2648 12248
rect 2700 11898 2728 12786
rect 2792 12628 2820 12854
rect 2792 12600 2912 12628
rect 2778 12472 2834 12481
rect 2778 12407 2834 12416
rect 2504 11892 2556 11898
rect 2504 11834 2556 11840
rect 2688 11892 2740 11898
rect 2688 11834 2740 11840
rect 2424 11206 2544 11234
rect 2412 11144 2464 11150
rect 2412 11086 2464 11092
rect 2320 10600 2372 10606
rect 2320 10542 2372 10548
rect 2228 9580 2280 9586
rect 2228 9522 2280 9528
rect 1952 9512 2004 9518
rect 1952 9454 2004 9460
rect 2228 9444 2280 9450
rect 2228 9386 2280 9392
rect 1676 9172 1728 9178
rect 1676 9114 1728 9120
rect 2136 8968 2188 8974
rect 2136 8910 2188 8916
rect 1952 8560 2004 8566
rect 1952 8502 2004 8508
rect 1964 7886 1992 8502
rect 2148 8430 2176 8910
rect 2136 8424 2188 8430
rect 2136 8366 2188 8372
rect 1952 7880 2004 7886
rect 1952 7822 2004 7828
rect 1964 7410 1992 7822
rect 2148 7750 2176 8366
rect 2240 7886 2268 9386
rect 2332 9110 2360 10542
rect 2320 9104 2372 9110
rect 2320 9046 2372 9052
rect 2424 8430 2452 11086
rect 2516 10266 2544 11206
rect 2700 10656 2728 11834
rect 2792 11558 2820 12407
rect 2884 11778 2912 12600
rect 2976 11898 3004 13790
rect 2964 11892 3016 11898
rect 2964 11834 3016 11840
rect 2884 11762 3004 11778
rect 2884 11756 3016 11762
rect 2884 11750 2964 11756
rect 2964 11698 3016 11704
rect 2780 11552 2832 11558
rect 2780 11494 2832 11500
rect 2872 11144 2924 11150
rect 2872 11086 2924 11092
rect 2780 10668 2832 10674
rect 2700 10628 2780 10656
rect 2596 10532 2648 10538
rect 2596 10474 2648 10480
rect 2504 10260 2556 10266
rect 2504 10202 2556 10208
rect 2608 9042 2636 10474
rect 2700 10198 2728 10628
rect 2780 10610 2832 10616
rect 2884 10554 2912 11086
rect 2976 10810 3004 11698
rect 2964 10804 3016 10810
rect 2964 10746 3016 10752
rect 2792 10526 2912 10554
rect 2688 10192 2740 10198
rect 2688 10134 2740 10140
rect 2792 9654 2820 10526
rect 3068 10198 3096 13926
rect 3056 10192 3108 10198
rect 3056 10134 3108 10140
rect 3056 10056 3108 10062
rect 3056 9998 3108 10004
rect 2780 9648 2832 9654
rect 2780 9590 2832 9596
rect 2872 9444 2924 9450
rect 2872 9386 2924 9392
rect 2596 9036 2648 9042
rect 2596 8978 2648 8984
rect 2608 8838 2636 8978
rect 2596 8832 2648 8838
rect 2596 8774 2648 8780
rect 2780 8492 2832 8498
rect 2780 8434 2832 8440
rect 2412 8424 2464 8430
rect 2412 8366 2464 8372
rect 2688 8424 2740 8430
rect 2688 8366 2740 8372
rect 2228 7880 2280 7886
rect 2228 7822 2280 7828
rect 2136 7744 2188 7750
rect 2136 7686 2188 7692
rect 1768 7404 1820 7410
rect 1768 7346 1820 7352
rect 1952 7404 2004 7410
rect 1952 7346 2004 7352
rect 1780 5710 1808 7346
rect 2044 6792 2096 6798
rect 2044 6734 2096 6740
rect 2056 5914 2084 6734
rect 2044 5908 2096 5914
rect 2044 5850 2096 5856
rect 1768 5704 1820 5710
rect 1768 5646 1820 5652
rect 1952 5704 2004 5710
rect 1952 5646 2004 5652
rect 1780 5166 1808 5646
rect 1860 5568 1912 5574
rect 1860 5510 1912 5516
rect 1768 5160 1820 5166
rect 1768 5102 1820 5108
rect 1780 4622 1808 5102
rect 1768 4616 1820 4622
rect 1768 4558 1820 4564
rect 1872 4146 1900 5510
rect 1860 4140 1912 4146
rect 1860 4082 1912 4088
rect 1872 3942 1900 4082
rect 1964 4010 1992 5646
rect 2056 4146 2084 5850
rect 2148 5234 2176 7686
rect 2136 5228 2188 5234
rect 2136 5170 2188 5176
rect 2240 4826 2268 7822
rect 2320 7404 2372 7410
rect 2320 7346 2372 7352
rect 2332 5234 2360 7346
rect 2412 7268 2464 7274
rect 2412 7210 2464 7216
rect 2424 6322 2452 7210
rect 2596 6656 2648 6662
rect 2596 6598 2648 6604
rect 2608 6322 2636 6598
rect 2412 6316 2464 6322
rect 2412 6258 2464 6264
rect 2596 6316 2648 6322
rect 2596 6258 2648 6264
rect 2320 5228 2372 5234
rect 2372 5188 2452 5216
rect 2320 5170 2372 5176
rect 2228 4820 2280 4826
rect 2228 4762 2280 4768
rect 2424 4622 2452 5188
rect 2320 4616 2372 4622
rect 2320 4558 2372 4564
rect 2412 4616 2464 4622
rect 2412 4558 2464 4564
rect 2332 4214 2360 4558
rect 2320 4208 2372 4214
rect 2320 4150 2372 4156
rect 2044 4140 2096 4146
rect 2044 4082 2096 4088
rect 2596 4140 2648 4146
rect 2596 4082 2648 4088
rect 1952 4004 2004 4010
rect 1952 3946 2004 3952
rect 1676 3936 1728 3942
rect 1676 3878 1728 3884
rect 1860 3936 1912 3942
rect 1860 3878 1912 3884
rect 1688 3534 1716 3878
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 1872 3194 1900 3878
rect 1860 3188 1912 3194
rect 1860 3130 1912 3136
rect 1964 3058 1992 3946
rect 2608 3738 2636 4082
rect 2596 3732 2648 3738
rect 2516 3692 2596 3720
rect 2516 3058 2544 3692
rect 2596 3674 2648 3680
rect 2700 3534 2728 8366
rect 2792 8022 2820 8434
rect 2780 8016 2832 8022
rect 2780 7958 2832 7964
rect 2884 7546 2912 9386
rect 3068 8906 3096 9998
rect 3160 9654 3188 14436
rect 3240 14418 3292 14424
rect 3240 14340 3292 14346
rect 3240 14282 3292 14288
rect 3252 11354 3280 14282
rect 3344 13190 3372 15370
rect 3436 15162 3464 19314
rect 3424 15156 3476 15162
rect 3424 15098 3476 15104
rect 3424 14816 3476 14822
rect 3424 14758 3476 14764
rect 3436 14328 3464 14758
rect 3528 14482 3556 20742
rect 4344 20460 4396 20466
rect 4344 20402 4396 20408
rect 3790 20156 4098 20165
rect 3790 20154 3796 20156
rect 3852 20154 3876 20156
rect 3932 20154 3956 20156
rect 4012 20154 4036 20156
rect 4092 20154 4098 20156
rect 3852 20102 3854 20154
rect 4034 20102 4036 20154
rect 3790 20100 3796 20102
rect 3852 20100 3876 20102
rect 3932 20100 3956 20102
rect 4012 20100 4036 20102
rect 4092 20100 4098 20102
rect 3790 20091 4098 20100
rect 3608 19712 3660 19718
rect 3608 19654 3660 19660
rect 3516 14476 3568 14482
rect 3516 14418 3568 14424
rect 3516 14340 3568 14346
rect 3436 14300 3516 14328
rect 3516 14282 3568 14288
rect 3528 13394 3556 14282
rect 3516 13388 3568 13394
rect 3516 13330 3568 13336
rect 3528 13258 3556 13330
rect 3516 13252 3568 13258
rect 3516 13194 3568 13200
rect 3332 13184 3384 13190
rect 3332 13126 3384 13132
rect 3332 12844 3384 12850
rect 3332 12786 3384 12792
rect 3344 12481 3372 12786
rect 3424 12708 3476 12714
rect 3424 12650 3476 12656
rect 3330 12472 3386 12481
rect 3330 12407 3386 12416
rect 3332 12164 3384 12170
rect 3332 12106 3384 12112
rect 3344 11830 3372 12106
rect 3332 11824 3384 11830
rect 3332 11766 3384 11772
rect 3240 11348 3292 11354
rect 3240 11290 3292 11296
rect 3344 10606 3372 11766
rect 3332 10600 3384 10606
rect 3332 10542 3384 10548
rect 3344 10130 3372 10542
rect 3332 10124 3384 10130
rect 3332 10066 3384 10072
rect 3436 10062 3464 12650
rect 3516 11756 3568 11762
rect 3516 11698 3568 11704
rect 3528 11150 3556 11698
rect 3516 11144 3568 11150
rect 3516 11086 3568 11092
rect 3516 10464 3568 10470
rect 3516 10406 3568 10412
rect 3424 10056 3476 10062
rect 3424 9998 3476 10004
rect 3240 9988 3292 9994
rect 3240 9930 3292 9936
rect 3148 9648 3200 9654
rect 3148 9590 3200 9596
rect 3252 9450 3280 9930
rect 3528 9674 3556 10406
rect 3344 9646 3556 9674
rect 3344 9518 3372 9646
rect 3424 9580 3476 9586
rect 3476 9540 3556 9568
rect 3424 9522 3476 9528
rect 3332 9512 3384 9518
rect 3528 9489 3556 9540
rect 3332 9454 3384 9460
rect 3514 9480 3570 9489
rect 3240 9444 3292 9450
rect 3514 9415 3570 9424
rect 3240 9386 3292 9392
rect 3056 8900 3108 8906
rect 3056 8842 3108 8848
rect 2964 8424 3016 8430
rect 2964 8366 3016 8372
rect 2872 7540 2924 7546
rect 2872 7482 2924 7488
rect 2884 7410 2912 7482
rect 2872 7404 2924 7410
rect 2872 7346 2924 7352
rect 2976 7206 3004 8366
rect 2964 7200 3016 7206
rect 2964 7142 3016 7148
rect 2976 6798 3004 7142
rect 2964 6792 3016 6798
rect 2964 6734 3016 6740
rect 3068 6322 3096 8842
rect 3252 8566 3280 9386
rect 3424 9172 3476 9178
rect 3424 9114 3476 9120
rect 3240 8560 3292 8566
rect 3240 8502 3292 8508
rect 3252 8362 3280 8502
rect 3332 8492 3384 8498
rect 3332 8434 3384 8440
rect 3240 8356 3292 8362
rect 3240 8298 3292 8304
rect 3344 8090 3372 8434
rect 3332 8084 3384 8090
rect 3332 8026 3384 8032
rect 3240 8016 3292 8022
rect 3240 7958 3292 7964
rect 3252 7002 3280 7958
rect 3240 6996 3292 7002
rect 3240 6938 3292 6944
rect 3252 6798 3280 6938
rect 3240 6792 3292 6798
rect 3240 6734 3292 6740
rect 2780 6316 2832 6322
rect 2780 6258 2832 6264
rect 3056 6316 3108 6322
rect 3056 6258 3108 6264
rect 2792 4826 2820 6258
rect 2964 6180 3016 6186
rect 2964 6122 3016 6128
rect 2872 5636 2924 5642
rect 2872 5578 2924 5584
rect 2780 4820 2832 4826
rect 2780 4762 2832 4768
rect 2792 3670 2820 4762
rect 2884 3942 2912 5578
rect 2976 5574 3004 6122
rect 2964 5568 3016 5574
rect 2964 5510 3016 5516
rect 2976 5370 3004 5510
rect 3252 5370 3280 6734
rect 2964 5364 3016 5370
rect 2964 5306 3016 5312
rect 3240 5364 3292 5370
rect 3240 5306 3292 5312
rect 3148 5160 3200 5166
rect 3148 5102 3200 5108
rect 2872 3936 2924 3942
rect 2872 3878 2924 3884
rect 2780 3664 2832 3670
rect 2780 3606 2832 3612
rect 2596 3528 2648 3534
rect 2596 3470 2648 3476
rect 2688 3528 2740 3534
rect 2688 3470 2740 3476
rect 2608 3194 2636 3470
rect 2596 3188 2648 3194
rect 2596 3130 2648 3136
rect 1952 3052 2004 3058
rect 1952 2994 2004 3000
rect 2504 3052 2556 3058
rect 2504 2994 2556 3000
rect 3160 2922 3188 5102
rect 3436 4486 3464 9114
rect 3516 8424 3568 8430
rect 3516 8366 3568 8372
rect 3528 5846 3556 8366
rect 3516 5840 3568 5846
rect 3516 5782 3568 5788
rect 3620 5234 3648 19654
rect 4356 19378 4384 20402
rect 4436 19712 4488 19718
rect 4436 19654 4488 19660
rect 4344 19372 4396 19378
rect 4344 19314 4396 19320
rect 3790 19068 4098 19077
rect 3790 19066 3796 19068
rect 3852 19066 3876 19068
rect 3932 19066 3956 19068
rect 4012 19066 4036 19068
rect 4092 19066 4098 19068
rect 3852 19014 3854 19066
rect 4034 19014 4036 19066
rect 3790 19012 3796 19014
rect 3852 19012 3876 19014
rect 3932 19012 3956 19014
rect 4012 19012 4036 19014
rect 4092 19012 4098 19014
rect 3790 19003 4098 19012
rect 3790 17980 4098 17989
rect 3790 17978 3796 17980
rect 3852 17978 3876 17980
rect 3932 17978 3956 17980
rect 4012 17978 4036 17980
rect 4092 17978 4098 17980
rect 3852 17926 3854 17978
rect 4034 17926 4036 17978
rect 3790 17924 3796 17926
rect 3852 17924 3876 17926
rect 3932 17924 3956 17926
rect 4012 17924 4036 17926
rect 4092 17924 4098 17926
rect 3790 17915 4098 17924
rect 3790 16892 4098 16901
rect 3790 16890 3796 16892
rect 3852 16890 3876 16892
rect 3932 16890 3956 16892
rect 4012 16890 4036 16892
rect 4092 16890 4098 16892
rect 3852 16838 3854 16890
rect 4034 16838 4036 16890
rect 3790 16836 3796 16838
rect 3852 16836 3876 16838
rect 3932 16836 3956 16838
rect 4012 16836 4036 16838
rect 4092 16836 4098 16838
rect 3790 16827 4098 16836
rect 4356 16182 4384 19314
rect 4344 16176 4396 16182
rect 4344 16118 4396 16124
rect 3790 15804 4098 15813
rect 3790 15802 3796 15804
rect 3852 15802 3876 15804
rect 3932 15802 3956 15804
rect 4012 15802 4036 15804
rect 4092 15802 4098 15804
rect 3852 15750 3854 15802
rect 4034 15750 4036 15802
rect 3790 15748 3796 15750
rect 3852 15748 3876 15750
rect 3932 15748 3956 15750
rect 4012 15748 4036 15750
rect 4092 15748 4098 15750
rect 3790 15739 4098 15748
rect 3700 15496 3752 15502
rect 3700 15438 3752 15444
rect 3712 14074 3740 15438
rect 4252 15428 4304 15434
rect 4252 15370 4304 15376
rect 4160 15088 4212 15094
rect 4160 15030 4212 15036
rect 3790 14716 4098 14725
rect 3790 14714 3796 14716
rect 3852 14714 3876 14716
rect 3932 14714 3956 14716
rect 4012 14714 4036 14716
rect 4092 14714 4098 14716
rect 3852 14662 3854 14714
rect 4034 14662 4036 14714
rect 3790 14660 3796 14662
rect 3852 14660 3876 14662
rect 3932 14660 3956 14662
rect 4012 14660 4036 14662
rect 4092 14660 4098 14662
rect 3790 14651 4098 14660
rect 3700 14068 3752 14074
rect 3700 14010 3752 14016
rect 3700 13728 3752 13734
rect 3700 13670 3752 13676
rect 3712 13462 3740 13670
rect 3790 13628 4098 13637
rect 3790 13626 3796 13628
rect 3852 13626 3876 13628
rect 3932 13626 3956 13628
rect 4012 13626 4036 13628
rect 4092 13626 4098 13628
rect 3852 13574 3854 13626
rect 4034 13574 4036 13626
rect 3790 13572 3796 13574
rect 3852 13572 3876 13574
rect 3932 13572 3956 13574
rect 4012 13572 4036 13574
rect 4092 13572 4098 13574
rect 3790 13563 4098 13572
rect 3700 13456 3752 13462
rect 3700 13398 3752 13404
rect 3976 13252 4028 13258
rect 3976 13194 4028 13200
rect 3988 12918 4016 13194
rect 3976 12912 4028 12918
rect 3976 12854 4028 12860
rect 3790 12540 4098 12549
rect 3790 12538 3796 12540
rect 3852 12538 3876 12540
rect 3932 12538 3956 12540
rect 4012 12538 4036 12540
rect 4092 12538 4098 12540
rect 3852 12486 3854 12538
rect 4034 12486 4036 12538
rect 3790 12484 3796 12486
rect 3852 12484 3876 12486
rect 3932 12484 3956 12486
rect 4012 12484 4036 12486
rect 4092 12484 4098 12486
rect 3790 12475 4098 12484
rect 4172 12442 4200 15030
rect 4264 14550 4292 15370
rect 4252 14544 4304 14550
rect 4252 14486 4304 14492
rect 4448 13410 4476 19654
rect 4528 15360 4580 15366
rect 4528 15302 4580 15308
rect 4540 13462 4568 15302
rect 4620 14952 4672 14958
rect 4620 14894 4672 14900
rect 4632 14550 4660 14894
rect 4724 14618 4752 20810
rect 5724 19780 5776 19786
rect 5724 19722 5776 19728
rect 5172 19508 5224 19514
rect 5172 19450 5224 19456
rect 5080 17128 5132 17134
rect 5080 17070 5132 17076
rect 4896 16448 4948 16454
rect 4896 16390 4948 16396
rect 4712 14612 4764 14618
rect 4712 14554 4764 14560
rect 4620 14544 4672 14550
rect 4620 14486 4672 14492
rect 4620 14408 4672 14414
rect 4620 14350 4672 14356
rect 4632 13530 4660 14350
rect 4620 13524 4672 13530
rect 4620 13466 4672 13472
rect 4264 13394 4476 13410
rect 4528 13456 4580 13462
rect 4528 13398 4580 13404
rect 4252 13388 4476 13394
rect 4304 13382 4476 13388
rect 4252 13330 4304 13336
rect 4252 13252 4304 13258
rect 4252 13194 4304 13200
rect 4344 13252 4396 13258
rect 4344 13194 4396 13200
rect 4264 12850 4292 13194
rect 4356 12986 4384 13194
rect 4344 12980 4396 12986
rect 4344 12922 4396 12928
rect 4252 12844 4304 12850
rect 4252 12786 4304 12792
rect 4252 12640 4304 12646
rect 4252 12582 4304 12588
rect 4160 12436 4212 12442
rect 4160 12378 4212 12384
rect 3700 12232 3752 12238
rect 3700 12174 3752 12180
rect 4160 12232 4212 12238
rect 4160 12174 4212 12180
rect 3712 9364 3740 12174
rect 3790 11452 4098 11461
rect 3790 11450 3796 11452
rect 3852 11450 3876 11452
rect 3932 11450 3956 11452
rect 4012 11450 4036 11452
rect 4092 11450 4098 11452
rect 3852 11398 3854 11450
rect 4034 11398 4036 11450
rect 3790 11396 3796 11398
rect 3852 11396 3876 11398
rect 3932 11396 3956 11398
rect 4012 11396 4036 11398
rect 4092 11396 4098 11398
rect 3790 11387 4098 11396
rect 4172 11336 4200 12174
rect 3988 11308 4200 11336
rect 3884 11280 3936 11286
rect 3988 11268 4016 11308
rect 3936 11240 4016 11268
rect 3884 11222 3936 11228
rect 4068 11212 4120 11218
rect 4068 11154 4120 11160
rect 4160 11212 4212 11218
rect 4160 11154 4212 11160
rect 4080 10742 4108 11154
rect 4068 10736 4120 10742
rect 4068 10678 4120 10684
rect 4172 10538 4200 11154
rect 4264 11082 4292 12582
rect 4344 12096 4396 12102
rect 4344 12038 4396 12044
rect 4356 11286 4384 12038
rect 4344 11280 4396 11286
rect 4344 11222 4396 11228
rect 4344 11144 4396 11150
rect 4344 11086 4396 11092
rect 4252 11076 4304 11082
rect 4252 11018 4304 11024
rect 4356 10810 4384 11086
rect 4252 10804 4304 10810
rect 4252 10746 4304 10752
rect 4344 10804 4396 10810
rect 4344 10746 4396 10752
rect 4160 10532 4212 10538
rect 4160 10474 4212 10480
rect 3790 10364 4098 10373
rect 3790 10362 3796 10364
rect 3852 10362 3876 10364
rect 3932 10362 3956 10364
rect 4012 10362 4036 10364
rect 4092 10362 4098 10364
rect 3852 10310 3854 10362
rect 4034 10310 4036 10362
rect 3790 10308 3796 10310
rect 3852 10308 3876 10310
rect 3932 10308 3956 10310
rect 4012 10308 4036 10310
rect 4092 10308 4098 10310
rect 3790 10299 4098 10308
rect 4172 10130 4200 10474
rect 4160 10124 4212 10130
rect 4160 10066 4212 10072
rect 4264 9654 4292 10746
rect 4252 9648 4304 9654
rect 4252 9590 4304 9596
rect 4160 9580 4212 9586
rect 4160 9522 4212 9528
rect 3792 9376 3844 9382
rect 3712 9336 3792 9364
rect 3792 9318 3844 9324
rect 3790 9276 4098 9285
rect 3790 9274 3796 9276
rect 3852 9274 3876 9276
rect 3932 9274 3956 9276
rect 4012 9274 4036 9276
rect 4092 9274 4098 9276
rect 3852 9222 3854 9274
rect 4034 9222 4036 9274
rect 3790 9220 3796 9222
rect 3852 9220 3876 9222
rect 3932 9220 3956 9222
rect 4012 9220 4036 9222
rect 4092 9220 4098 9222
rect 3790 9211 4098 9220
rect 4172 9178 4200 9522
rect 4160 9172 4212 9178
rect 4160 9114 4212 9120
rect 3884 8968 3936 8974
rect 3936 8916 4200 8922
rect 3884 8910 4200 8916
rect 3896 8894 4200 8910
rect 3790 8188 4098 8197
rect 3790 8186 3796 8188
rect 3852 8186 3876 8188
rect 3932 8186 3956 8188
rect 4012 8186 4036 8188
rect 4092 8186 4098 8188
rect 3852 8134 3854 8186
rect 4034 8134 4036 8186
rect 3790 8132 3796 8134
rect 3852 8132 3876 8134
rect 3932 8132 3956 8134
rect 4012 8132 4036 8134
rect 4092 8132 4098 8134
rect 3790 8123 4098 8132
rect 4172 8090 4200 8894
rect 4252 8900 4304 8906
rect 4252 8842 4304 8848
rect 4264 8498 4292 8842
rect 4252 8492 4304 8498
rect 4252 8434 4304 8440
rect 4160 8084 4212 8090
rect 4160 8026 4212 8032
rect 4264 7206 4292 8434
rect 4436 8424 4488 8430
rect 4436 8366 4488 8372
rect 4344 8356 4396 8362
rect 4344 8298 4396 8304
rect 4356 7886 4384 8298
rect 4448 7886 4476 8366
rect 4540 7954 4568 13398
rect 4908 11898 4936 16390
rect 4986 15056 5042 15065
rect 4986 14991 4988 15000
rect 5040 14991 5042 15000
rect 4988 14962 5040 14968
rect 4988 14884 5040 14890
rect 4988 14826 5040 14832
rect 5000 13530 5028 14826
rect 5092 14074 5120 17070
rect 5080 14068 5132 14074
rect 5080 14010 5132 14016
rect 4988 13524 5040 13530
rect 4988 13466 5040 13472
rect 5000 12918 5028 13466
rect 5184 13326 5212 19450
rect 5540 17536 5592 17542
rect 5540 17478 5592 17484
rect 5356 16992 5408 16998
rect 5356 16934 5408 16940
rect 5264 16448 5316 16454
rect 5264 16390 5316 16396
rect 5276 15337 5304 16390
rect 5262 15328 5318 15337
rect 5262 15263 5318 15272
rect 5264 15088 5316 15094
rect 5264 15030 5316 15036
rect 5276 14414 5304 15030
rect 5264 14408 5316 14414
rect 5264 14350 5316 14356
rect 5368 13870 5396 16934
rect 5448 14408 5500 14414
rect 5448 14350 5500 14356
rect 5460 13938 5488 14350
rect 5448 13932 5500 13938
rect 5448 13874 5500 13880
rect 5356 13864 5408 13870
rect 5356 13806 5408 13812
rect 5460 13394 5488 13874
rect 5448 13388 5500 13394
rect 5448 13330 5500 13336
rect 5172 13320 5224 13326
rect 5172 13262 5224 13268
rect 5264 13320 5316 13326
rect 5264 13262 5316 13268
rect 5276 13190 5304 13262
rect 5264 13184 5316 13190
rect 5264 13126 5316 13132
rect 4988 12912 5040 12918
rect 4988 12854 5040 12860
rect 5276 12850 5304 13126
rect 5264 12844 5316 12850
rect 5264 12786 5316 12792
rect 5460 12714 5488 13330
rect 5448 12708 5500 12714
rect 5448 12650 5500 12656
rect 4896 11892 4948 11898
rect 4896 11834 4948 11840
rect 5172 11824 5224 11830
rect 5172 11766 5224 11772
rect 4988 11756 5040 11762
rect 4988 11698 5040 11704
rect 4620 11688 4672 11694
rect 4620 11630 4672 11636
rect 4896 11688 4948 11694
rect 4896 11630 4948 11636
rect 4632 11218 4660 11630
rect 4620 11212 4672 11218
rect 4620 11154 4672 11160
rect 4632 10742 4660 11154
rect 4712 10804 4764 10810
rect 4712 10746 4764 10752
rect 4620 10736 4672 10742
rect 4620 10678 4672 10684
rect 4620 10600 4672 10606
rect 4620 10542 4672 10548
rect 4632 9518 4660 10542
rect 4620 9512 4672 9518
rect 4620 9454 4672 9460
rect 4632 8974 4660 9454
rect 4724 9382 4752 10746
rect 4804 10464 4856 10470
rect 4804 10406 4856 10412
rect 4712 9376 4764 9382
rect 4712 9318 4764 9324
rect 4620 8968 4672 8974
rect 4620 8910 4672 8916
rect 4528 7948 4580 7954
rect 4528 7890 4580 7896
rect 4344 7880 4396 7886
rect 4344 7822 4396 7828
rect 4436 7880 4488 7886
rect 4436 7822 4488 7828
rect 4448 7478 4476 7822
rect 4528 7812 4580 7818
rect 4528 7754 4580 7760
rect 4436 7472 4488 7478
rect 4436 7414 4488 7420
rect 4540 7274 4568 7754
rect 4816 7478 4844 10406
rect 4908 9110 4936 11630
rect 5000 10266 5028 11698
rect 4988 10260 5040 10266
rect 4988 10202 5040 10208
rect 5080 10056 5132 10062
rect 5184 10044 5212 11766
rect 5448 11756 5500 11762
rect 5448 11698 5500 11704
rect 5356 10600 5408 10606
rect 5356 10542 5408 10548
rect 5368 10062 5396 10542
rect 5132 10033 5212 10044
rect 5356 10056 5408 10062
rect 5132 10024 5226 10033
rect 5132 10016 5170 10024
rect 5080 9998 5132 10004
rect 5356 9998 5408 10004
rect 5170 9959 5226 9968
rect 5080 9920 5132 9926
rect 5132 9880 5212 9908
rect 5080 9862 5132 9868
rect 5080 9648 5132 9654
rect 5080 9590 5132 9596
rect 4896 9104 4948 9110
rect 4896 9046 4948 9052
rect 4988 8900 5040 8906
rect 4988 8842 5040 8848
rect 4896 8832 4948 8838
rect 4896 8774 4948 8780
rect 4908 8498 4936 8774
rect 4896 8492 4948 8498
rect 4896 8434 4948 8440
rect 4804 7472 4856 7478
rect 4804 7414 4856 7420
rect 4528 7268 4580 7274
rect 4528 7210 4580 7216
rect 4160 7200 4212 7206
rect 4160 7142 4212 7148
rect 4252 7200 4304 7206
rect 4252 7142 4304 7148
rect 3790 7100 4098 7109
rect 3790 7098 3796 7100
rect 3852 7098 3876 7100
rect 3932 7098 3956 7100
rect 4012 7098 4036 7100
rect 4092 7098 4098 7100
rect 3852 7046 3854 7098
rect 4034 7046 4036 7098
rect 3790 7044 3796 7046
rect 3852 7044 3876 7046
rect 3932 7044 3956 7046
rect 4012 7044 4036 7046
rect 4092 7044 4098 7046
rect 3790 7035 4098 7044
rect 4172 6390 4200 7142
rect 4160 6384 4212 6390
rect 4160 6326 4212 6332
rect 3700 6248 3752 6254
rect 3700 6190 3752 6196
rect 3712 5914 3740 6190
rect 3790 6012 4098 6021
rect 3790 6010 3796 6012
rect 3852 6010 3876 6012
rect 3932 6010 3956 6012
rect 4012 6010 4036 6012
rect 4092 6010 4098 6012
rect 3852 5958 3854 6010
rect 4034 5958 4036 6010
rect 3790 5956 3796 5958
rect 3852 5956 3876 5958
rect 3932 5956 3956 5958
rect 4012 5956 4036 5958
rect 4092 5956 4098 5958
rect 3790 5947 4098 5956
rect 3700 5908 3752 5914
rect 3700 5850 3752 5856
rect 3608 5228 3660 5234
rect 3608 5170 3660 5176
rect 3516 5024 3568 5030
rect 3516 4966 3568 4972
rect 3424 4480 3476 4486
rect 3424 4422 3476 4428
rect 3436 3942 3464 4422
rect 3424 3936 3476 3942
rect 3424 3878 3476 3884
rect 3436 3534 3464 3878
rect 3424 3528 3476 3534
rect 3330 3496 3386 3505
rect 3424 3470 3476 3476
rect 3330 3431 3332 3440
rect 3384 3431 3386 3440
rect 3332 3402 3384 3408
rect 3528 3058 3556 4966
rect 3790 4924 4098 4933
rect 3790 4922 3796 4924
rect 3852 4922 3876 4924
rect 3932 4922 3956 4924
rect 4012 4922 4036 4924
rect 4092 4922 4098 4924
rect 3852 4870 3854 4922
rect 4034 4870 4036 4922
rect 3790 4868 3796 4870
rect 3852 4868 3876 4870
rect 3932 4868 3956 4870
rect 4012 4868 4036 4870
rect 4092 4868 4098 4870
rect 3790 4859 4098 4868
rect 4172 4622 4200 6326
rect 4264 5574 4292 7142
rect 4816 6866 4844 7414
rect 4908 7410 4936 8434
rect 5000 8090 5028 8842
rect 4988 8084 5040 8090
rect 4988 8026 5040 8032
rect 4896 7404 4948 7410
rect 4896 7346 4948 7352
rect 4804 6860 4856 6866
rect 4804 6802 4856 6808
rect 4344 6724 4396 6730
rect 4344 6666 4396 6672
rect 4252 5568 4304 5574
rect 4252 5510 4304 5516
rect 4264 5302 4292 5510
rect 4252 5296 4304 5302
rect 4252 5238 4304 5244
rect 4252 5160 4304 5166
rect 4252 5102 4304 5108
rect 4160 4616 4212 4622
rect 4160 4558 4212 4564
rect 4160 4480 4212 4486
rect 4160 4422 4212 4428
rect 3700 4072 3752 4078
rect 3700 4014 3752 4020
rect 3516 3052 3568 3058
rect 3516 2994 3568 3000
rect 3424 2984 3476 2990
rect 3424 2926 3476 2932
rect 2136 2916 2188 2922
rect 2136 2858 2188 2864
rect 3148 2916 3200 2922
rect 3148 2858 3200 2864
rect 1492 1216 1544 1222
rect 1492 1158 1544 1164
rect 1504 800 1532 1158
rect 2148 800 2176 2858
rect 2780 2372 2832 2378
rect 2780 2314 2832 2320
rect 2792 800 2820 2314
rect 3436 800 3464 2926
rect 1490 0 1546 800
rect 2134 0 2190 800
rect 2778 0 2834 800
rect 3422 0 3478 800
rect 3712 762 3740 4014
rect 4172 4010 4200 4422
rect 4264 4146 4292 5102
rect 4356 4758 4384 6666
rect 4816 6322 4844 6802
rect 4804 6316 4856 6322
rect 4804 6258 4856 6264
rect 4804 6112 4856 6118
rect 4804 6054 4856 6060
rect 4816 5710 4844 6054
rect 4804 5704 4856 5710
rect 4804 5646 4856 5652
rect 5000 5642 5028 8026
rect 5092 7410 5120 9590
rect 5080 7404 5132 7410
rect 5080 7346 5132 7352
rect 5080 6792 5132 6798
rect 5080 6734 5132 6740
rect 5092 6390 5120 6734
rect 5080 6384 5132 6390
rect 5080 6326 5132 6332
rect 5184 6225 5212 9880
rect 5356 9648 5408 9654
rect 5356 9590 5408 9596
rect 5368 9489 5396 9590
rect 5354 9480 5410 9489
rect 5354 9415 5410 9424
rect 5356 6860 5408 6866
rect 5356 6802 5408 6808
rect 5368 6769 5396 6802
rect 5354 6760 5410 6769
rect 5354 6695 5410 6704
rect 5170 6216 5226 6225
rect 5170 6151 5226 6160
rect 5080 5704 5132 5710
rect 5080 5646 5132 5652
rect 5264 5704 5316 5710
rect 5264 5646 5316 5652
rect 4988 5636 5040 5642
rect 4988 5578 5040 5584
rect 4896 5568 4948 5574
rect 4896 5510 4948 5516
rect 4344 4752 4396 4758
rect 4344 4694 4396 4700
rect 4356 4554 4384 4694
rect 4344 4548 4396 4554
rect 4344 4490 4396 4496
rect 4436 4480 4488 4486
rect 4356 4428 4436 4434
rect 4356 4422 4488 4428
rect 4356 4406 4476 4422
rect 4252 4140 4304 4146
rect 4252 4082 4304 4088
rect 4160 4004 4212 4010
rect 4160 3946 4212 3952
rect 3790 3836 4098 3845
rect 3790 3834 3796 3836
rect 3852 3834 3876 3836
rect 3932 3834 3956 3836
rect 4012 3834 4036 3836
rect 4092 3834 4098 3836
rect 3852 3782 3854 3834
rect 4034 3782 4036 3834
rect 3790 3780 3796 3782
rect 3852 3780 3876 3782
rect 3932 3780 3956 3782
rect 4012 3780 4036 3782
rect 4092 3780 4098 3782
rect 3790 3771 4098 3780
rect 3976 3528 4028 3534
rect 3976 3470 4028 3476
rect 3988 3058 4016 3470
rect 4264 3058 4292 4082
rect 4356 3942 4384 4406
rect 4436 4208 4488 4214
rect 4436 4150 4488 4156
rect 4344 3936 4396 3942
rect 4344 3878 4396 3884
rect 4356 3777 4384 3878
rect 4342 3768 4398 3777
rect 4342 3703 4344 3712
rect 4396 3703 4398 3712
rect 4344 3674 4396 3680
rect 4448 3058 4476 4150
rect 4908 4146 4936 5510
rect 5000 5098 5028 5578
rect 4988 5092 5040 5098
rect 4988 5034 5040 5040
rect 4896 4140 4948 4146
rect 4896 4082 4948 4088
rect 4908 3466 4936 4082
rect 5000 4010 5028 5034
rect 5092 4554 5120 5646
rect 5276 5166 5304 5646
rect 5264 5160 5316 5166
rect 5264 5102 5316 5108
rect 5264 4752 5316 4758
rect 5264 4694 5316 4700
rect 5080 4548 5132 4554
rect 5080 4490 5132 4496
rect 4988 4004 5040 4010
rect 4988 3946 5040 3952
rect 5000 3602 5028 3946
rect 4988 3596 5040 3602
rect 4988 3538 5040 3544
rect 4896 3460 4948 3466
rect 4896 3402 4948 3408
rect 3976 3052 4028 3058
rect 3976 2994 4028 3000
rect 4252 3052 4304 3058
rect 4436 3052 4488 3058
rect 4304 3012 4384 3040
rect 4252 2994 4304 3000
rect 4160 2848 4212 2854
rect 4160 2790 4212 2796
rect 3790 2748 4098 2757
rect 3790 2746 3796 2748
rect 3852 2746 3876 2748
rect 3932 2746 3956 2748
rect 4012 2746 4036 2748
rect 4092 2746 4098 2748
rect 3852 2694 3854 2746
rect 4034 2694 4036 2746
rect 3790 2692 3796 2694
rect 3852 2692 3876 2694
rect 3932 2692 3956 2694
rect 4012 2692 4036 2694
rect 4092 2692 4098 2694
rect 3790 2683 4098 2692
rect 4172 2446 4200 2790
rect 4356 2446 4384 3012
rect 4436 2994 4488 3000
rect 4448 2650 4476 2994
rect 4908 2922 4936 3402
rect 4896 2916 4948 2922
rect 4896 2858 4948 2864
rect 4436 2644 4488 2650
rect 4436 2586 4488 2592
rect 4908 2582 4936 2858
rect 5000 2854 5028 3538
rect 5172 3528 5224 3534
rect 5172 3470 5224 3476
rect 4988 2848 5040 2854
rect 4988 2790 5040 2796
rect 4896 2576 4948 2582
rect 4896 2518 4948 2524
rect 5184 2446 5212 3470
rect 5276 3210 5304 4694
rect 5356 4548 5408 4554
rect 5356 4490 5408 4496
rect 5368 4146 5396 4490
rect 5356 4140 5408 4146
rect 5356 4082 5408 4088
rect 5368 3602 5396 4082
rect 5460 4078 5488 11698
rect 5552 10538 5580 17478
rect 5632 15020 5684 15026
rect 5632 14962 5684 14968
rect 5644 12850 5672 14962
rect 5736 13734 5764 19722
rect 5828 18970 5856 21626
rect 6184 21344 6236 21350
rect 6184 21286 6236 21292
rect 5908 19508 5960 19514
rect 5908 19450 5960 19456
rect 5816 18964 5868 18970
rect 5816 18906 5868 18912
rect 5828 18766 5856 18906
rect 5816 18760 5868 18766
rect 5816 18702 5868 18708
rect 5920 14498 5948 19450
rect 6196 14890 6224 21286
rect 6288 15162 6316 21830
rect 6630 21788 6938 21797
rect 6630 21786 6636 21788
rect 6692 21786 6716 21788
rect 6772 21786 6796 21788
rect 6852 21786 6876 21788
rect 6932 21786 6938 21788
rect 6692 21734 6694 21786
rect 6874 21734 6876 21786
rect 6630 21732 6636 21734
rect 6692 21732 6716 21734
rect 6772 21732 6796 21734
rect 6852 21732 6876 21734
rect 6932 21732 6938 21734
rect 6630 21723 6938 21732
rect 8852 21344 8904 21350
rect 8852 21286 8904 21292
rect 6630 20700 6938 20709
rect 6630 20698 6636 20700
rect 6692 20698 6716 20700
rect 6772 20698 6796 20700
rect 6852 20698 6876 20700
rect 6932 20698 6938 20700
rect 6692 20646 6694 20698
rect 6874 20646 6876 20698
rect 6630 20644 6636 20646
rect 6692 20644 6716 20646
rect 6772 20644 6796 20646
rect 6852 20644 6876 20646
rect 6932 20644 6938 20646
rect 6630 20635 6938 20644
rect 6630 19612 6938 19621
rect 6630 19610 6636 19612
rect 6692 19610 6716 19612
rect 6772 19610 6796 19612
rect 6852 19610 6876 19612
rect 6932 19610 6938 19612
rect 6692 19558 6694 19610
rect 6874 19558 6876 19610
rect 6630 19556 6636 19558
rect 6692 19556 6716 19558
rect 6772 19556 6796 19558
rect 6852 19556 6876 19558
rect 6932 19556 6938 19558
rect 6630 19547 6938 19556
rect 7564 19440 7616 19446
rect 7564 19382 7616 19388
rect 7472 19372 7524 19378
rect 7472 19314 7524 19320
rect 7484 18970 7512 19314
rect 7472 18964 7524 18970
rect 7472 18906 7524 18912
rect 6630 18524 6938 18533
rect 6630 18522 6636 18524
rect 6692 18522 6716 18524
rect 6772 18522 6796 18524
rect 6852 18522 6876 18524
rect 6932 18522 6938 18524
rect 6692 18470 6694 18522
rect 6874 18470 6876 18522
rect 6630 18468 6636 18470
rect 6692 18468 6716 18470
rect 6772 18468 6796 18470
rect 6852 18468 6876 18470
rect 6932 18468 6938 18470
rect 6630 18459 6938 18468
rect 7484 18358 7512 18906
rect 7472 18352 7524 18358
rect 7472 18294 7524 18300
rect 7104 17740 7156 17746
rect 7104 17682 7156 17688
rect 6368 17604 6420 17610
rect 6368 17546 6420 17552
rect 6276 15156 6328 15162
rect 6276 15098 6328 15104
rect 6184 14884 6236 14890
rect 6184 14826 6236 14832
rect 6000 14816 6052 14822
rect 6000 14758 6052 14764
rect 6092 14816 6144 14822
rect 6092 14758 6144 14764
rect 6012 14550 6040 14758
rect 5828 14470 5948 14498
rect 6000 14544 6052 14550
rect 6000 14486 6052 14492
rect 6104 14482 6132 14758
rect 6092 14476 6144 14482
rect 5724 13728 5776 13734
rect 5724 13670 5776 13676
rect 5632 12844 5684 12850
rect 5632 12786 5684 12792
rect 5644 12442 5672 12786
rect 5724 12640 5776 12646
rect 5724 12582 5776 12588
rect 5632 12436 5684 12442
rect 5632 12378 5684 12384
rect 5644 11898 5672 12378
rect 5632 11892 5684 11898
rect 5632 11834 5684 11840
rect 5632 11688 5684 11694
rect 5632 11630 5684 11636
rect 5644 10606 5672 11630
rect 5736 11218 5764 12582
rect 5724 11212 5776 11218
rect 5724 11154 5776 11160
rect 5828 11014 5856 14470
rect 6092 14418 6144 14424
rect 6092 14340 6144 14346
rect 6092 14282 6144 14288
rect 6184 14340 6236 14346
rect 6184 14282 6236 14288
rect 5908 13864 5960 13870
rect 5908 13806 5960 13812
rect 5920 12102 5948 13806
rect 6000 12844 6052 12850
rect 6000 12786 6052 12792
rect 5908 12096 5960 12102
rect 5908 12038 5960 12044
rect 5920 11150 5948 12038
rect 5908 11144 5960 11150
rect 5908 11086 5960 11092
rect 5816 11008 5868 11014
rect 5816 10950 5868 10956
rect 5724 10668 5776 10674
rect 5724 10610 5776 10616
rect 5632 10600 5684 10606
rect 5632 10542 5684 10548
rect 5540 10532 5592 10538
rect 5540 10474 5592 10480
rect 5540 10192 5592 10198
rect 5540 10134 5592 10140
rect 5552 10062 5580 10134
rect 5540 10056 5592 10062
rect 5540 9998 5592 10004
rect 5736 9518 5764 10610
rect 5816 10464 5868 10470
rect 5816 10406 5868 10412
rect 5828 9926 5856 10406
rect 5816 9920 5868 9926
rect 5816 9862 5868 9868
rect 5724 9512 5776 9518
rect 5722 9480 5724 9489
rect 5776 9480 5778 9489
rect 5722 9415 5778 9424
rect 5828 9353 5856 9862
rect 5920 9654 5948 11086
rect 6012 9994 6040 12786
rect 6104 11082 6132 14282
rect 6196 13938 6224 14282
rect 6184 13932 6236 13938
rect 6184 13874 6236 13880
rect 6196 13530 6224 13874
rect 6184 13524 6236 13530
rect 6184 13466 6236 13472
rect 6288 13394 6316 15098
rect 6276 13388 6328 13394
rect 6276 13330 6328 13336
rect 6288 12306 6316 13330
rect 6276 12300 6328 12306
rect 6276 12242 6328 12248
rect 6276 11756 6328 11762
rect 6276 11698 6328 11704
rect 6092 11076 6144 11082
rect 6092 11018 6144 11024
rect 6000 9988 6052 9994
rect 6000 9930 6052 9936
rect 5908 9648 5960 9654
rect 5908 9590 5960 9596
rect 5920 9450 5948 9590
rect 5908 9444 5960 9450
rect 5908 9386 5960 9392
rect 5814 9344 5870 9353
rect 5814 9279 5870 9288
rect 5920 8498 5948 9386
rect 6012 8974 6040 9930
rect 6000 8968 6052 8974
rect 6000 8910 6052 8916
rect 5908 8492 5960 8498
rect 5908 8434 5960 8440
rect 5816 8016 5868 8022
rect 5816 7958 5868 7964
rect 5828 7886 5856 7958
rect 5816 7880 5868 7886
rect 5736 7840 5816 7868
rect 5540 7268 5592 7274
rect 5540 7210 5592 7216
rect 5552 6934 5580 7210
rect 5540 6928 5592 6934
rect 5540 6870 5592 6876
rect 5552 6322 5580 6870
rect 5540 6316 5592 6322
rect 5540 6258 5592 6264
rect 5736 6254 5764 7840
rect 5816 7822 5868 7828
rect 5816 7744 5868 7750
rect 5816 7686 5868 7692
rect 5828 6866 5856 7686
rect 5908 7404 5960 7410
rect 5908 7346 5960 7352
rect 5920 7274 5948 7346
rect 5908 7268 5960 7274
rect 5908 7210 5960 7216
rect 5816 6860 5868 6866
rect 5816 6802 5868 6808
rect 5816 6724 5868 6730
rect 5816 6666 5868 6672
rect 5724 6248 5776 6254
rect 5724 6190 5776 6196
rect 5828 5370 5856 6666
rect 5920 6236 5948 7210
rect 6012 6866 6040 8910
rect 6104 8090 6132 11018
rect 6288 10198 6316 11698
rect 6380 10810 6408 17546
rect 6630 17436 6938 17445
rect 6630 17434 6636 17436
rect 6692 17434 6716 17436
rect 6772 17434 6796 17436
rect 6852 17434 6876 17436
rect 6932 17434 6938 17436
rect 6692 17382 6694 17434
rect 6874 17382 6876 17434
rect 6630 17380 6636 17382
rect 6692 17380 6716 17382
rect 6772 17380 6796 17382
rect 6852 17380 6876 17382
rect 6932 17380 6938 17382
rect 6630 17371 6938 17380
rect 7116 16658 7144 17682
rect 7104 16652 7156 16658
rect 7104 16594 7156 16600
rect 6460 16448 6512 16454
rect 6460 16390 6512 16396
rect 6368 10804 6420 10810
rect 6368 10746 6420 10752
rect 6472 10266 6500 16390
rect 6630 16348 6938 16357
rect 6630 16346 6636 16348
rect 6692 16346 6716 16348
rect 6772 16346 6796 16348
rect 6852 16346 6876 16348
rect 6932 16346 6938 16348
rect 6692 16294 6694 16346
rect 6874 16294 6876 16346
rect 6630 16292 6636 16294
rect 6692 16292 6716 16294
rect 6772 16292 6796 16294
rect 6852 16292 6876 16294
rect 6932 16292 6938 16294
rect 6630 16283 6938 16292
rect 7576 15858 7604 19382
rect 8024 19372 8076 19378
rect 8024 19314 8076 19320
rect 8036 17746 8064 19314
rect 8300 18692 8352 18698
rect 8300 18634 8352 18640
rect 8024 17740 8076 17746
rect 8024 17682 8076 17688
rect 8036 17202 8064 17682
rect 8024 17196 8076 17202
rect 8024 17138 8076 17144
rect 8208 17196 8260 17202
rect 8208 17138 8260 17144
rect 8220 16658 8248 17138
rect 8208 16652 8260 16658
rect 8208 16594 8260 16600
rect 8220 16250 8248 16594
rect 8208 16244 8260 16250
rect 8208 16186 8260 16192
rect 7484 15830 7604 15858
rect 6552 15428 6604 15434
rect 6552 15370 6604 15376
rect 6564 14618 6592 15370
rect 6630 15260 6938 15269
rect 6630 15258 6636 15260
rect 6692 15258 6716 15260
rect 6772 15258 6796 15260
rect 6852 15258 6876 15260
rect 6932 15258 6938 15260
rect 6692 15206 6694 15258
rect 6874 15206 6876 15258
rect 6630 15204 6636 15206
rect 6692 15204 6716 15206
rect 6772 15204 6796 15206
rect 6852 15204 6876 15206
rect 6932 15204 6938 15206
rect 6630 15195 6938 15204
rect 7010 15056 7066 15065
rect 7010 14991 7066 15000
rect 6644 14884 6696 14890
rect 6644 14826 6696 14832
rect 6552 14612 6604 14618
rect 6552 14554 6604 14560
rect 6656 14362 6684 14826
rect 7024 14414 7052 14991
rect 7196 14544 7248 14550
rect 7196 14486 7248 14492
rect 6564 14334 6684 14362
rect 7012 14408 7064 14414
rect 7208 14396 7236 14486
rect 7288 14476 7340 14482
rect 7288 14418 7340 14424
rect 7064 14368 7236 14396
rect 7012 14350 7064 14356
rect 6564 13258 6592 14334
rect 7012 14272 7064 14278
rect 7012 14214 7064 14220
rect 6630 14172 6938 14181
rect 6630 14170 6636 14172
rect 6692 14170 6716 14172
rect 6772 14170 6796 14172
rect 6852 14170 6876 14172
rect 6932 14170 6938 14172
rect 6692 14118 6694 14170
rect 6874 14118 6876 14170
rect 6630 14116 6636 14118
rect 6692 14116 6716 14118
rect 6772 14116 6796 14118
rect 6852 14116 6876 14118
rect 6932 14116 6938 14118
rect 6630 14107 6938 14116
rect 7024 13734 7052 14214
rect 7012 13728 7064 13734
rect 7012 13670 7064 13676
rect 6552 13252 6604 13258
rect 6552 13194 6604 13200
rect 6630 13084 6938 13093
rect 6630 13082 6636 13084
rect 6692 13082 6716 13084
rect 6772 13082 6796 13084
rect 6852 13082 6876 13084
rect 6932 13082 6938 13084
rect 6692 13030 6694 13082
rect 6874 13030 6876 13082
rect 6630 13028 6636 13030
rect 6692 13028 6716 13030
rect 6772 13028 6796 13030
rect 6852 13028 6876 13030
rect 6932 13028 6938 13030
rect 6630 13019 6938 13028
rect 6552 12980 6604 12986
rect 6552 12922 6604 12928
rect 6564 12238 6592 12922
rect 7024 12646 7052 13670
rect 7104 13456 7156 13462
rect 7104 13398 7156 13404
rect 7116 12714 7144 13398
rect 7208 13190 7236 14368
rect 7196 13184 7248 13190
rect 7196 13126 7248 13132
rect 7104 12708 7156 12714
rect 7104 12650 7156 12656
rect 7012 12640 7064 12646
rect 7012 12582 7064 12588
rect 6552 12232 6604 12238
rect 6552 12174 6604 12180
rect 7024 12170 7052 12582
rect 7196 12436 7248 12442
rect 7196 12378 7248 12384
rect 7208 12238 7236 12378
rect 7300 12374 7328 14418
rect 7380 14408 7432 14414
rect 7380 14350 7432 14356
rect 7392 12442 7420 14350
rect 7380 12436 7432 12442
rect 7380 12378 7432 12384
rect 7288 12368 7340 12374
rect 7288 12310 7340 12316
rect 7196 12232 7248 12238
rect 7196 12174 7248 12180
rect 7012 12164 7064 12170
rect 7012 12106 7064 12112
rect 6630 11996 6938 12005
rect 6630 11994 6636 11996
rect 6692 11994 6716 11996
rect 6772 11994 6796 11996
rect 6852 11994 6876 11996
rect 6932 11994 6938 11996
rect 6692 11942 6694 11994
rect 6874 11942 6876 11994
rect 6630 11940 6636 11942
rect 6692 11940 6716 11942
rect 6772 11940 6796 11942
rect 6852 11940 6876 11942
rect 6932 11940 6938 11942
rect 6630 11931 6938 11940
rect 7012 11892 7064 11898
rect 7012 11834 7064 11840
rect 6552 11552 6604 11558
rect 6552 11494 6604 11500
rect 6564 10674 6592 11494
rect 6630 10908 6938 10917
rect 6630 10906 6636 10908
rect 6692 10906 6716 10908
rect 6772 10906 6796 10908
rect 6852 10906 6876 10908
rect 6932 10906 6938 10908
rect 6692 10854 6694 10906
rect 6874 10854 6876 10906
rect 6630 10852 6636 10854
rect 6692 10852 6716 10854
rect 6772 10852 6796 10854
rect 6852 10852 6876 10854
rect 6932 10852 6938 10854
rect 6630 10843 6938 10852
rect 7024 10742 7052 11834
rect 7208 11830 7236 12174
rect 7196 11824 7248 11830
rect 7196 11766 7248 11772
rect 7196 11688 7248 11694
rect 7196 11630 7248 11636
rect 7012 10736 7064 10742
rect 7012 10678 7064 10684
rect 6552 10668 6604 10674
rect 6552 10610 6604 10616
rect 6828 10532 6880 10538
rect 6828 10474 6880 10480
rect 6460 10260 6512 10266
rect 6460 10202 6512 10208
rect 6276 10192 6328 10198
rect 6276 10134 6328 10140
rect 6184 10056 6236 10062
rect 6184 9998 6236 10004
rect 6092 8084 6144 8090
rect 6092 8026 6144 8032
rect 6000 6860 6052 6866
rect 6000 6802 6052 6808
rect 6012 6390 6040 6802
rect 6104 6798 6132 8026
rect 6092 6792 6144 6798
rect 6092 6734 6144 6740
rect 6000 6384 6052 6390
rect 6000 6326 6052 6332
rect 5920 6208 6132 6236
rect 5816 5364 5868 5370
rect 5816 5306 5868 5312
rect 5828 4690 5856 5306
rect 6104 4690 6132 6208
rect 5816 4684 5868 4690
rect 5816 4626 5868 4632
rect 6092 4684 6144 4690
rect 6092 4626 6144 4632
rect 5540 4616 5592 4622
rect 5540 4558 5592 4564
rect 5724 4616 5776 4622
rect 5724 4558 5776 4564
rect 5448 4072 5500 4078
rect 5448 4014 5500 4020
rect 5356 3596 5408 3602
rect 5356 3538 5408 3544
rect 5276 3182 5488 3210
rect 5552 3194 5580 4558
rect 5356 3120 5408 3126
rect 5356 3062 5408 3068
rect 4160 2440 4212 2446
rect 4160 2382 4212 2388
rect 4344 2440 4396 2446
rect 4344 2382 4396 2388
rect 5172 2440 5224 2446
rect 5172 2382 5224 2388
rect 4712 2304 4764 2310
rect 4712 2246 4764 2252
rect 3988 870 4108 898
rect 3988 762 4016 870
rect 4080 800 4108 870
rect 4724 800 4752 2246
rect 5368 800 5396 3062
rect 5460 2990 5488 3182
rect 5540 3188 5592 3194
rect 5540 3130 5592 3136
rect 5736 3058 5764 4558
rect 5816 3460 5868 3466
rect 5816 3402 5868 3408
rect 5828 3058 5856 3402
rect 5724 3052 5776 3058
rect 5724 2994 5776 3000
rect 5816 3052 5868 3058
rect 5816 2994 5868 3000
rect 5448 2984 5500 2990
rect 5632 2984 5684 2990
rect 5448 2926 5500 2932
rect 5630 2952 5632 2961
rect 5684 2952 5686 2961
rect 5630 2887 5686 2896
rect 5828 2650 5856 2994
rect 6104 2854 6132 4626
rect 6092 2848 6144 2854
rect 6092 2790 6144 2796
rect 6196 2650 6224 9998
rect 6288 9178 6316 10134
rect 6840 10130 6868 10474
rect 6828 10124 6880 10130
rect 6828 10066 6880 10072
rect 6840 9926 6868 10066
rect 7024 10033 7052 10678
rect 7104 10192 7156 10198
rect 7104 10134 7156 10140
rect 7010 10024 7066 10033
rect 7010 9959 7066 9968
rect 6828 9920 6880 9926
rect 6828 9862 6880 9868
rect 6630 9820 6938 9829
rect 6630 9818 6636 9820
rect 6692 9818 6716 9820
rect 6772 9818 6796 9820
rect 6852 9818 6876 9820
rect 6932 9818 6938 9820
rect 6692 9766 6694 9818
rect 6874 9766 6876 9818
rect 6630 9764 6636 9766
rect 6692 9764 6716 9766
rect 6772 9764 6796 9766
rect 6852 9764 6876 9766
rect 6932 9764 6938 9766
rect 6630 9755 6938 9764
rect 7024 9654 7052 9959
rect 7012 9648 7064 9654
rect 7012 9590 7064 9596
rect 6368 9376 6420 9382
rect 6368 9318 6420 9324
rect 6642 9344 6698 9353
rect 6276 9172 6328 9178
rect 6276 9114 6328 9120
rect 6276 9036 6328 9042
rect 6276 8978 6328 8984
rect 6288 8362 6316 8978
rect 6380 8430 6408 9318
rect 6642 9279 6698 9288
rect 6656 8974 6684 9279
rect 7116 9178 7144 10134
rect 7208 10062 7236 11630
rect 7300 11150 7328 12310
rect 7484 11354 7512 15830
rect 8220 15570 8248 16186
rect 8208 15564 8260 15570
rect 8208 15506 8260 15512
rect 7932 15360 7984 15366
rect 7932 15302 7984 15308
rect 7840 14952 7892 14958
rect 7840 14894 7892 14900
rect 7656 14816 7708 14822
rect 7656 14758 7708 14764
rect 7564 12844 7616 12850
rect 7564 12786 7616 12792
rect 7576 12442 7604 12786
rect 7564 12436 7616 12442
rect 7564 12378 7616 12384
rect 7668 11778 7696 14758
rect 7852 13870 7880 14894
rect 7944 14414 7972 15302
rect 8220 15026 8248 15506
rect 8208 15020 8260 15026
rect 8208 14962 8260 14968
rect 7932 14408 7984 14414
rect 7932 14350 7984 14356
rect 7840 13864 7892 13870
rect 7840 13806 7892 13812
rect 7748 13184 7800 13190
rect 7748 13126 7800 13132
rect 7760 12918 7788 13126
rect 7852 12986 7880 13806
rect 7840 12980 7892 12986
rect 7840 12922 7892 12928
rect 7748 12912 7800 12918
rect 7748 12854 7800 12860
rect 7852 12714 7880 12922
rect 7840 12708 7892 12714
rect 7840 12650 7892 12656
rect 7840 12164 7892 12170
rect 7840 12106 7892 12112
rect 7576 11750 7696 11778
rect 7852 11762 7880 12106
rect 7840 11756 7892 11762
rect 7472 11348 7524 11354
rect 7472 11290 7524 11296
rect 7288 11144 7340 11150
rect 7288 11086 7340 11092
rect 7472 11144 7524 11150
rect 7472 11086 7524 11092
rect 7380 11008 7432 11014
rect 7380 10950 7432 10956
rect 7288 10600 7340 10606
rect 7286 10568 7288 10577
rect 7340 10568 7342 10577
rect 7286 10503 7342 10512
rect 7300 10470 7328 10503
rect 7288 10464 7340 10470
rect 7288 10406 7340 10412
rect 7196 10056 7248 10062
rect 7196 9998 7248 10004
rect 7392 9926 7420 10950
rect 7380 9920 7432 9926
rect 7380 9862 7432 9868
rect 7288 9716 7340 9722
rect 7288 9658 7340 9664
rect 7196 9376 7248 9382
rect 7300 9364 7328 9658
rect 7248 9336 7328 9364
rect 7196 9318 7248 9324
rect 7104 9172 7156 9178
rect 7104 9114 7156 9120
rect 6644 8968 6696 8974
rect 6644 8910 6696 8916
rect 7012 8900 7064 8906
rect 7012 8842 7064 8848
rect 6630 8732 6938 8741
rect 6630 8730 6636 8732
rect 6692 8730 6716 8732
rect 6772 8730 6796 8732
rect 6852 8730 6876 8732
rect 6932 8730 6938 8732
rect 6692 8678 6694 8730
rect 6874 8678 6876 8730
rect 6630 8676 6636 8678
rect 6692 8676 6716 8678
rect 6772 8676 6796 8678
rect 6852 8676 6876 8678
rect 6932 8676 6938 8678
rect 6630 8667 6938 8676
rect 7024 8566 7052 8842
rect 7012 8560 7064 8566
rect 7012 8502 7064 8508
rect 6368 8424 6420 8430
rect 6368 8366 6420 8372
rect 6276 8356 6328 8362
rect 6276 8298 6328 8304
rect 6380 7750 6408 8366
rect 6552 7880 6604 7886
rect 6552 7822 6604 7828
rect 6460 7812 6512 7818
rect 6460 7754 6512 7760
rect 6368 7744 6420 7750
rect 6368 7686 6420 7692
rect 6276 6792 6328 6798
rect 6276 6734 6328 6740
rect 6288 6186 6316 6734
rect 6380 6458 6408 7686
rect 6368 6452 6420 6458
rect 6368 6394 6420 6400
rect 6276 6180 6328 6186
rect 6276 6122 6328 6128
rect 6288 5846 6316 6122
rect 6276 5840 6328 5846
rect 6276 5782 6328 5788
rect 6380 5302 6408 6394
rect 6472 6390 6500 7754
rect 6564 7274 6592 7822
rect 6630 7644 6938 7653
rect 6630 7642 6636 7644
rect 6692 7642 6716 7644
rect 6772 7642 6796 7644
rect 6852 7642 6876 7644
rect 6932 7642 6938 7644
rect 6692 7590 6694 7642
rect 6874 7590 6876 7642
rect 6630 7588 6636 7590
rect 6692 7588 6716 7590
rect 6772 7588 6796 7590
rect 6852 7588 6876 7590
rect 6932 7588 6938 7590
rect 6630 7579 6938 7588
rect 6552 7268 6604 7274
rect 6552 7210 6604 7216
rect 6552 6656 6604 6662
rect 6552 6598 6604 6604
rect 6460 6384 6512 6390
rect 6460 6326 6512 6332
rect 6564 6322 6592 6598
rect 6630 6556 6938 6565
rect 6630 6554 6636 6556
rect 6692 6554 6716 6556
rect 6772 6554 6796 6556
rect 6852 6554 6876 6556
rect 6932 6554 6938 6556
rect 6692 6502 6694 6554
rect 6874 6502 6876 6554
rect 6630 6500 6636 6502
rect 6692 6500 6716 6502
rect 6772 6500 6796 6502
rect 6852 6500 6876 6502
rect 6932 6500 6938 6502
rect 6630 6491 6938 6500
rect 7012 6452 7064 6458
rect 7012 6394 7064 6400
rect 6552 6316 6604 6322
rect 6552 6258 6604 6264
rect 6564 5710 6592 6258
rect 6920 6248 6972 6254
rect 6920 6190 6972 6196
rect 6932 5914 6960 6190
rect 6920 5908 6972 5914
rect 6920 5850 6972 5856
rect 6552 5704 6604 5710
rect 6552 5646 6604 5652
rect 7024 5574 7052 6394
rect 7012 5568 7064 5574
rect 7012 5510 7064 5516
rect 6630 5468 6938 5477
rect 6630 5466 6636 5468
rect 6692 5466 6716 5468
rect 6772 5466 6796 5468
rect 6852 5466 6876 5468
rect 6932 5466 6938 5468
rect 6692 5414 6694 5466
rect 6874 5414 6876 5466
rect 6630 5412 6636 5414
rect 6692 5412 6716 5414
rect 6772 5412 6796 5414
rect 6852 5412 6876 5414
rect 6932 5412 6938 5414
rect 6630 5403 6938 5412
rect 6368 5296 6420 5302
rect 6368 5238 6420 5244
rect 6274 5128 6330 5137
rect 6274 5063 6330 5072
rect 6288 2774 6316 5063
rect 6380 4214 6408 5238
rect 7024 5234 7052 5510
rect 6644 5228 6696 5234
rect 6644 5170 6696 5176
rect 6736 5228 6788 5234
rect 6736 5170 6788 5176
rect 7012 5228 7064 5234
rect 7012 5170 7064 5176
rect 6460 5160 6512 5166
rect 6460 5102 6512 5108
rect 6368 4208 6420 4214
rect 6368 4150 6420 4156
rect 6472 3670 6500 5102
rect 6552 4752 6604 4758
rect 6552 4694 6604 4700
rect 6564 4214 6592 4694
rect 6656 4690 6684 5170
rect 6748 4758 6776 5170
rect 6736 4752 6788 4758
rect 6736 4694 6788 4700
rect 6644 4684 6696 4690
rect 6644 4626 6696 4632
rect 6630 4380 6938 4389
rect 6630 4378 6636 4380
rect 6692 4378 6716 4380
rect 6772 4378 6796 4380
rect 6852 4378 6876 4380
rect 6932 4378 6938 4380
rect 6692 4326 6694 4378
rect 6874 4326 6876 4378
rect 6630 4324 6636 4326
rect 6692 4324 6716 4326
rect 6772 4324 6796 4326
rect 6852 4324 6876 4326
rect 6932 4324 6938 4326
rect 6630 4315 6938 4324
rect 7024 4282 7052 5170
rect 7012 4276 7064 4282
rect 7012 4218 7064 4224
rect 6552 4208 6604 4214
rect 7116 4162 7144 9114
rect 7208 4826 7236 9318
rect 7392 8378 7420 9862
rect 7484 9586 7512 11086
rect 7576 10198 7604 11750
rect 7840 11698 7892 11704
rect 7656 11620 7708 11626
rect 7656 11562 7708 11568
rect 7668 10470 7696 11562
rect 7852 11218 7880 11698
rect 7944 11286 7972 14350
rect 8220 13938 8248 14962
rect 8312 14618 8340 18634
rect 8392 16992 8444 16998
rect 8392 16934 8444 16940
rect 8404 16590 8432 16934
rect 8392 16584 8444 16590
rect 8392 16526 8444 16532
rect 8484 16448 8536 16454
rect 8484 16390 8536 16396
rect 8300 14612 8352 14618
rect 8300 14554 8352 14560
rect 8300 14340 8352 14346
rect 8300 14282 8352 14288
rect 8208 13932 8260 13938
rect 8208 13874 8260 13880
rect 8312 12850 8340 14282
rect 8116 12844 8168 12850
rect 8116 12786 8168 12792
rect 8300 12844 8352 12850
rect 8300 12786 8352 12792
rect 8024 12640 8076 12646
rect 8024 12582 8076 12588
rect 7932 11280 7984 11286
rect 7932 11222 7984 11228
rect 7840 11212 7892 11218
rect 7840 11154 7892 11160
rect 7932 10668 7984 10674
rect 7932 10610 7984 10616
rect 7748 10600 7800 10606
rect 7748 10542 7800 10548
rect 7656 10464 7708 10470
rect 7656 10406 7708 10412
rect 7564 10192 7616 10198
rect 7564 10134 7616 10140
rect 7668 9994 7696 10406
rect 7656 9988 7708 9994
rect 7656 9930 7708 9936
rect 7564 9920 7616 9926
rect 7616 9868 7696 9874
rect 7564 9862 7696 9868
rect 7576 9846 7696 9862
rect 7564 9716 7616 9722
rect 7564 9658 7616 9664
rect 7472 9580 7524 9586
rect 7472 9522 7524 9528
rect 7484 9382 7512 9522
rect 7472 9376 7524 9382
rect 7472 9318 7524 9324
rect 7484 8498 7512 9318
rect 7472 8492 7524 8498
rect 7472 8434 7524 8440
rect 7392 8350 7512 8378
rect 7380 8016 7432 8022
rect 7380 7958 7432 7964
rect 7288 7812 7340 7818
rect 7288 7754 7340 7760
rect 7300 7002 7328 7754
rect 7288 6996 7340 7002
rect 7288 6938 7340 6944
rect 7300 6798 7328 6938
rect 7392 6798 7420 7958
rect 7288 6792 7340 6798
rect 7288 6734 7340 6740
rect 7380 6792 7432 6798
rect 7380 6734 7432 6740
rect 7392 5370 7420 6734
rect 7380 5364 7432 5370
rect 7380 5306 7432 5312
rect 7196 4820 7248 4826
rect 7196 4762 7248 4768
rect 7392 4690 7420 5306
rect 7380 4684 7432 4690
rect 7380 4626 7432 4632
rect 6552 4150 6604 4156
rect 7024 4134 7144 4162
rect 7024 3942 7052 4134
rect 7196 4072 7248 4078
rect 7196 4014 7248 4020
rect 7012 3936 7064 3942
rect 7012 3878 7064 3884
rect 6460 3664 6512 3670
rect 6460 3606 6512 3612
rect 6552 3596 6604 3602
rect 6552 3538 6604 3544
rect 6288 2746 6500 2774
rect 5816 2644 5868 2650
rect 5816 2586 5868 2592
rect 6184 2644 6236 2650
rect 6184 2586 6236 2592
rect 6472 2446 6500 2746
rect 6460 2440 6512 2446
rect 6460 2382 6512 2388
rect 6000 2372 6052 2378
rect 6000 2314 6052 2320
rect 6012 800 6040 2314
rect 6564 1986 6592 3538
rect 6630 3292 6938 3301
rect 6630 3290 6636 3292
rect 6692 3290 6716 3292
rect 6772 3290 6796 3292
rect 6852 3290 6876 3292
rect 6932 3290 6938 3292
rect 6692 3238 6694 3290
rect 6874 3238 6876 3290
rect 6630 3236 6636 3238
rect 6692 3236 6716 3238
rect 6772 3236 6796 3238
rect 6852 3236 6876 3238
rect 6932 3236 6938 3238
rect 6630 3227 6938 3236
rect 7024 3058 7052 3878
rect 7208 3641 7236 4014
rect 7288 4004 7340 4010
rect 7288 3946 7340 3952
rect 7194 3632 7250 3641
rect 7194 3567 7250 3576
rect 7012 3052 7064 3058
rect 7012 2994 7064 3000
rect 6630 2204 6938 2213
rect 6630 2202 6636 2204
rect 6692 2202 6716 2204
rect 6772 2202 6796 2204
rect 6852 2202 6876 2204
rect 6932 2202 6938 2204
rect 6692 2150 6694 2202
rect 6874 2150 6876 2202
rect 6630 2148 6636 2150
rect 6692 2148 6716 2150
rect 6772 2148 6796 2150
rect 6852 2148 6876 2150
rect 6932 2148 6938 2150
rect 6630 2139 6938 2148
rect 6564 1958 6684 1986
rect 6656 800 6684 1958
rect 7300 800 7328 3946
rect 7392 3534 7420 4626
rect 7380 3528 7432 3534
rect 7380 3470 7432 3476
rect 7484 2774 7512 8350
rect 7576 7274 7604 9658
rect 7668 9586 7696 9846
rect 7656 9580 7708 9586
rect 7656 9522 7708 9528
rect 7668 8634 7696 9522
rect 7760 9518 7788 10542
rect 7840 10056 7892 10062
rect 7840 9998 7892 10004
rect 7852 9722 7880 9998
rect 7944 9926 7972 10610
rect 8036 10130 8064 12582
rect 8128 11558 8156 12786
rect 8208 12368 8260 12374
rect 8208 12310 8260 12316
rect 8220 12238 8248 12310
rect 8312 12306 8340 12786
rect 8300 12300 8352 12306
rect 8300 12242 8352 12248
rect 8208 12232 8260 12238
rect 8208 12174 8260 12180
rect 8116 11552 8168 11558
rect 8116 11494 8168 11500
rect 8024 10124 8076 10130
rect 8024 10066 8076 10072
rect 7932 9920 7984 9926
rect 7932 9862 7984 9868
rect 7840 9716 7892 9722
rect 7840 9658 7892 9664
rect 7748 9512 7800 9518
rect 7748 9454 7800 9460
rect 7656 8628 7708 8634
rect 7656 8570 7708 8576
rect 7760 8090 7788 9454
rect 8300 8560 8352 8566
rect 8300 8502 8352 8508
rect 7840 8492 7892 8498
rect 7840 8434 7892 8440
rect 7748 8084 7800 8090
rect 7748 8026 7800 8032
rect 7852 7342 7880 8434
rect 7932 8288 7984 8294
rect 7932 8230 7984 8236
rect 8116 8288 8168 8294
rect 8116 8230 8168 8236
rect 7944 7954 7972 8230
rect 7932 7948 7984 7954
rect 7932 7890 7984 7896
rect 8024 7880 8076 7886
rect 8024 7822 8076 7828
rect 7932 7404 7984 7410
rect 8036 7392 8064 7822
rect 7984 7364 8064 7392
rect 7932 7346 7984 7352
rect 7840 7336 7892 7342
rect 7840 7278 7892 7284
rect 7564 7268 7616 7274
rect 7564 7210 7616 7216
rect 7944 7206 7972 7346
rect 7840 7200 7892 7206
rect 7840 7142 7892 7148
rect 7932 7200 7984 7206
rect 7932 7142 7984 7148
rect 7748 6792 7800 6798
rect 7748 6734 7800 6740
rect 7760 6662 7788 6734
rect 7748 6656 7800 6662
rect 7748 6598 7800 6604
rect 7654 6352 7710 6361
rect 7654 6287 7710 6296
rect 7668 6186 7696 6287
rect 7656 6180 7708 6186
rect 7656 6122 7708 6128
rect 7760 6118 7788 6598
rect 7748 6112 7800 6118
rect 7748 6054 7800 6060
rect 7852 5778 7880 7142
rect 7840 5772 7892 5778
rect 7840 5714 7892 5720
rect 7748 5704 7800 5710
rect 7748 5646 7800 5652
rect 7760 5234 7788 5646
rect 7852 5556 7880 5714
rect 7944 5710 7972 7142
rect 8024 6316 8076 6322
rect 8024 6258 8076 6264
rect 7932 5704 7984 5710
rect 7932 5646 7984 5652
rect 8036 5556 8064 6258
rect 8128 5710 8156 8230
rect 8208 7404 8260 7410
rect 8208 7346 8260 7352
rect 8220 6322 8248 7346
rect 8312 6798 8340 8502
rect 8496 7993 8524 16390
rect 8668 12912 8720 12918
rect 8668 12854 8720 12860
rect 8680 11762 8708 12854
rect 8864 12782 8892 21286
rect 8956 12850 8984 21830
rect 9128 21616 9180 21622
rect 9128 21558 9180 21564
rect 9140 21010 9168 21558
rect 10520 21554 10548 21966
rect 12452 21894 12480 24200
rect 15152 22332 15460 22341
rect 15152 22330 15158 22332
rect 15214 22330 15238 22332
rect 15294 22330 15318 22332
rect 15374 22330 15398 22332
rect 15454 22330 15460 22332
rect 15214 22278 15216 22330
rect 15396 22278 15398 22330
rect 15152 22276 15158 22278
rect 15214 22276 15238 22278
rect 15294 22276 15318 22278
rect 15374 22276 15398 22278
rect 15454 22276 15460 22278
rect 15152 22267 15460 22276
rect 17420 21962 17448 24200
rect 20833 22332 21141 22341
rect 20833 22330 20839 22332
rect 20895 22330 20919 22332
rect 20975 22330 20999 22332
rect 21055 22330 21079 22332
rect 21135 22330 21141 22332
rect 20895 22278 20897 22330
rect 21077 22278 21079 22330
rect 20833 22276 20839 22278
rect 20895 22276 20919 22278
rect 20975 22276 20999 22278
rect 21055 22276 21079 22278
rect 21135 22276 21141 22278
rect 20833 22267 21141 22276
rect 21180 22092 21232 22098
rect 21180 22034 21232 22040
rect 19984 22024 20036 22030
rect 19984 21966 20036 21972
rect 17408 21956 17460 21962
rect 17408 21898 17460 21904
rect 11336 21888 11388 21894
rect 11336 21830 11388 21836
rect 12440 21888 12492 21894
rect 12440 21830 12492 21836
rect 14004 21888 14056 21894
rect 14004 21830 14056 21836
rect 15108 21888 15160 21894
rect 15108 21830 15160 21836
rect 15660 21888 15712 21894
rect 15660 21830 15712 21836
rect 17684 21888 17736 21894
rect 17684 21830 17736 21836
rect 10508 21548 10560 21554
rect 10508 21490 10560 21496
rect 11348 21350 11376 21830
rect 12311 21788 12619 21797
rect 12311 21786 12317 21788
rect 12373 21786 12397 21788
rect 12453 21786 12477 21788
rect 12533 21786 12557 21788
rect 12613 21786 12619 21788
rect 12373 21734 12375 21786
rect 12555 21734 12557 21786
rect 12311 21732 12317 21734
rect 12373 21732 12397 21734
rect 12453 21732 12477 21734
rect 12533 21732 12557 21734
rect 12613 21732 12619 21734
rect 12311 21723 12619 21732
rect 13820 21616 13872 21622
rect 13872 21564 13952 21570
rect 13820 21558 13952 21564
rect 13084 21548 13136 21554
rect 13832 21542 13952 21558
rect 14016 21554 14044 21830
rect 14556 21616 14608 21622
rect 14556 21558 14608 21564
rect 13084 21490 13136 21496
rect 12900 21412 12952 21418
rect 12900 21354 12952 21360
rect 11336 21344 11388 21350
rect 11336 21286 11388 21292
rect 11796 21344 11848 21350
rect 11796 21286 11848 21292
rect 9471 21244 9779 21253
rect 9471 21242 9477 21244
rect 9533 21242 9557 21244
rect 9613 21242 9637 21244
rect 9693 21242 9717 21244
rect 9773 21242 9779 21244
rect 9533 21190 9535 21242
rect 9715 21190 9717 21242
rect 9471 21188 9477 21190
rect 9533 21188 9557 21190
rect 9613 21188 9637 21190
rect 9693 21188 9717 21190
rect 9773 21188 9779 21190
rect 9471 21179 9779 21188
rect 11348 21146 11376 21286
rect 9404 21140 9456 21146
rect 9404 21082 9456 21088
rect 11336 21140 11388 21146
rect 11336 21082 11388 21088
rect 9128 21004 9180 21010
rect 9128 20946 9180 20952
rect 9036 20460 9088 20466
rect 9140 20448 9168 20946
rect 9416 20874 9444 21082
rect 11348 20874 11376 21082
rect 11808 20942 11836 21286
rect 11796 20936 11848 20942
rect 11796 20878 11848 20884
rect 12716 20936 12768 20942
rect 12768 20896 12848 20924
rect 12716 20878 12768 20884
rect 9404 20868 9456 20874
rect 9404 20810 9456 20816
rect 11244 20868 11296 20874
rect 11244 20810 11296 20816
rect 11336 20868 11388 20874
rect 11336 20810 11388 20816
rect 10048 20800 10100 20806
rect 10048 20742 10100 20748
rect 9088 20420 9168 20448
rect 9036 20402 9088 20408
rect 9140 19922 9168 20420
rect 9471 20156 9779 20165
rect 9471 20154 9477 20156
rect 9533 20154 9557 20156
rect 9613 20154 9637 20156
rect 9693 20154 9717 20156
rect 9773 20154 9779 20156
rect 9533 20102 9535 20154
rect 9715 20102 9717 20154
rect 9471 20100 9477 20102
rect 9533 20100 9557 20102
rect 9613 20100 9637 20102
rect 9693 20100 9717 20102
rect 9773 20100 9779 20102
rect 9471 20091 9779 20100
rect 9128 19916 9180 19922
rect 9128 19858 9180 19864
rect 9140 19394 9168 19858
rect 9048 19378 9168 19394
rect 9036 19372 9168 19378
rect 9088 19366 9168 19372
rect 9036 19314 9088 19320
rect 9140 18834 9168 19366
rect 9471 19068 9779 19077
rect 9471 19066 9477 19068
rect 9533 19066 9557 19068
rect 9613 19066 9637 19068
rect 9693 19066 9717 19068
rect 9773 19066 9779 19068
rect 9533 19014 9535 19066
rect 9715 19014 9717 19066
rect 9471 19012 9477 19014
rect 9533 19012 9557 19014
rect 9613 19012 9637 19014
rect 9693 19012 9717 19014
rect 9773 19012 9779 19014
rect 9471 19003 9779 19012
rect 9128 18828 9180 18834
rect 9128 18770 9180 18776
rect 9140 18426 9168 18770
rect 9128 18420 9180 18426
rect 9128 18362 9180 18368
rect 9140 17746 9168 18362
rect 9471 17980 9779 17989
rect 9471 17978 9477 17980
rect 9533 17978 9557 17980
rect 9613 17978 9637 17980
rect 9693 17978 9717 17980
rect 9773 17978 9779 17980
rect 9533 17926 9535 17978
rect 9715 17926 9717 17978
rect 9471 17924 9477 17926
rect 9533 17924 9557 17926
rect 9613 17924 9637 17926
rect 9693 17924 9717 17926
rect 9773 17924 9779 17926
rect 9471 17915 9779 17924
rect 9128 17740 9180 17746
rect 9128 17682 9180 17688
rect 9220 16992 9272 16998
rect 9220 16934 9272 16940
rect 9232 16250 9260 16934
rect 9471 16892 9779 16901
rect 9471 16890 9477 16892
rect 9533 16890 9557 16892
rect 9613 16890 9637 16892
rect 9693 16890 9717 16892
rect 9773 16890 9779 16892
rect 9533 16838 9535 16890
rect 9715 16838 9717 16890
rect 9471 16836 9477 16838
rect 9533 16836 9557 16838
rect 9613 16836 9637 16838
rect 9693 16836 9717 16838
rect 9773 16836 9779 16838
rect 9471 16827 9779 16836
rect 9220 16244 9272 16250
rect 9220 16186 9272 16192
rect 9471 15804 9779 15813
rect 9471 15802 9477 15804
rect 9533 15802 9557 15804
rect 9613 15802 9637 15804
rect 9693 15802 9717 15804
rect 9773 15802 9779 15804
rect 9533 15750 9535 15802
rect 9715 15750 9717 15802
rect 9471 15748 9477 15750
rect 9533 15748 9557 15750
rect 9613 15748 9637 15750
rect 9693 15748 9717 15750
rect 9773 15748 9779 15750
rect 9471 15739 9779 15748
rect 9471 14716 9779 14725
rect 9471 14714 9477 14716
rect 9533 14714 9557 14716
rect 9613 14714 9637 14716
rect 9693 14714 9717 14716
rect 9773 14714 9779 14716
rect 9533 14662 9535 14714
rect 9715 14662 9717 14714
rect 9471 14660 9477 14662
rect 9533 14660 9557 14662
rect 9613 14660 9637 14662
rect 9693 14660 9717 14662
rect 9773 14660 9779 14662
rect 9471 14651 9779 14660
rect 9312 14544 9364 14550
rect 9312 14486 9364 14492
rect 9324 14414 9352 14486
rect 9312 14408 9364 14414
rect 9312 14350 9364 14356
rect 9680 14408 9732 14414
rect 9680 14350 9732 14356
rect 9404 14340 9456 14346
rect 9404 14282 9456 14288
rect 9220 14272 9272 14278
rect 9220 14214 9272 14220
rect 9232 12986 9260 14214
rect 9416 13682 9444 14282
rect 9692 13938 9720 14350
rect 10060 13938 10088 20742
rect 11060 20596 11112 20602
rect 11060 20538 11112 20544
rect 10784 19712 10836 19718
rect 10784 19654 10836 19660
rect 10600 18624 10652 18630
rect 10600 18566 10652 18572
rect 10416 17536 10468 17542
rect 10416 17478 10468 17484
rect 10140 15564 10192 15570
rect 10140 15506 10192 15512
rect 10152 14074 10180 15506
rect 10140 14068 10192 14074
rect 10140 14010 10192 14016
rect 9680 13932 9732 13938
rect 9680 13874 9732 13880
rect 10048 13932 10100 13938
rect 10048 13874 10100 13880
rect 9324 13654 9444 13682
rect 9220 12980 9272 12986
rect 9220 12922 9272 12928
rect 9324 12850 9352 13654
rect 9471 13628 9779 13637
rect 9471 13626 9477 13628
rect 9533 13626 9557 13628
rect 9613 13626 9637 13628
rect 9693 13626 9717 13628
rect 9773 13626 9779 13628
rect 9533 13574 9535 13626
rect 9715 13574 9717 13626
rect 9471 13572 9477 13574
rect 9533 13572 9557 13574
rect 9613 13572 9637 13574
rect 9693 13572 9717 13574
rect 9773 13572 9779 13574
rect 9471 13563 9779 13572
rect 10060 13462 10088 13874
rect 10324 13728 10376 13734
rect 10324 13670 10376 13676
rect 10048 13456 10100 13462
rect 10048 13398 10100 13404
rect 10336 13394 10364 13670
rect 10324 13388 10376 13394
rect 10324 13330 10376 13336
rect 10140 13252 10192 13258
rect 10140 13194 10192 13200
rect 10152 12918 10180 13194
rect 10140 12912 10192 12918
rect 10140 12854 10192 12860
rect 10428 12850 10456 17478
rect 10508 14544 10560 14550
rect 10508 14486 10560 14492
rect 8944 12844 8996 12850
rect 8944 12786 8996 12792
rect 9036 12844 9088 12850
rect 9036 12786 9088 12792
rect 9312 12844 9364 12850
rect 9312 12786 9364 12792
rect 10416 12844 10468 12850
rect 10416 12786 10468 12792
rect 8852 12776 8904 12782
rect 8852 12718 8904 12724
rect 8760 12640 8812 12646
rect 8760 12582 8812 12588
rect 8668 11756 8720 11762
rect 8668 11698 8720 11704
rect 8576 11076 8628 11082
rect 8576 11018 8628 11024
rect 8588 10266 8616 11018
rect 8576 10260 8628 10266
rect 8576 10202 8628 10208
rect 8668 8832 8720 8838
rect 8668 8774 8720 8780
rect 8680 8498 8708 8774
rect 8668 8492 8720 8498
rect 8668 8434 8720 8440
rect 8482 7984 8538 7993
rect 8482 7919 8538 7928
rect 8576 7540 8628 7546
rect 8576 7482 8628 7488
rect 8392 7268 8444 7274
rect 8392 7210 8444 7216
rect 8404 7002 8432 7210
rect 8392 6996 8444 7002
rect 8392 6938 8444 6944
rect 8300 6792 8352 6798
rect 8300 6734 8352 6740
rect 8404 6610 8432 6938
rect 8404 6582 8524 6610
rect 8298 6488 8354 6497
rect 8496 6458 8524 6582
rect 8298 6423 8354 6432
rect 8392 6452 8444 6458
rect 8312 6390 8340 6423
rect 8392 6394 8444 6400
rect 8484 6452 8536 6458
rect 8484 6394 8536 6400
rect 8300 6384 8352 6390
rect 8300 6326 8352 6332
rect 8208 6316 8260 6322
rect 8208 6258 8260 6264
rect 8404 6118 8432 6394
rect 8392 6112 8444 6118
rect 8392 6054 8444 6060
rect 8116 5704 8168 5710
rect 8116 5646 8168 5652
rect 7852 5528 8064 5556
rect 7748 5228 7800 5234
rect 7748 5170 7800 5176
rect 7932 4616 7984 4622
rect 7932 4558 7984 4564
rect 7564 4548 7616 4554
rect 7564 4490 7616 4496
rect 7576 4214 7604 4490
rect 7564 4208 7616 4214
rect 7564 4150 7616 4156
rect 7576 3398 7604 4150
rect 7654 3768 7710 3777
rect 7654 3703 7710 3712
rect 7668 3398 7696 3703
rect 7564 3392 7616 3398
rect 7564 3334 7616 3340
rect 7656 3392 7708 3398
rect 7656 3334 7708 3340
rect 7392 2746 7512 2774
rect 7392 2446 7420 2746
rect 7656 2508 7708 2514
rect 7656 2450 7708 2456
rect 7380 2440 7432 2446
rect 7380 2382 7432 2388
rect 7668 1222 7696 2450
rect 7656 1216 7708 1222
rect 7656 1158 7708 1164
rect 7944 800 7972 4558
rect 8036 4185 8064 5528
rect 8484 5568 8536 5574
rect 8484 5510 8536 5516
rect 8496 4690 8524 5510
rect 8588 5234 8616 7482
rect 8680 5710 8708 8434
rect 8772 5778 8800 12582
rect 9048 8566 9076 12786
rect 9471 12540 9779 12549
rect 9471 12538 9477 12540
rect 9533 12538 9557 12540
rect 9613 12538 9637 12540
rect 9693 12538 9717 12540
rect 9773 12538 9779 12540
rect 9533 12486 9535 12538
rect 9715 12486 9717 12538
rect 9471 12484 9477 12486
rect 9533 12484 9557 12486
rect 9613 12484 9637 12486
rect 9693 12484 9717 12486
rect 9773 12484 9779 12486
rect 9471 12475 9779 12484
rect 10520 12434 10548 14486
rect 10428 12406 10548 12434
rect 9312 12096 9364 12102
rect 9312 12038 9364 12044
rect 9220 11892 9272 11898
rect 9220 11834 9272 11840
rect 9128 11756 9180 11762
rect 9128 11698 9180 11704
rect 9140 10742 9168 11698
rect 9232 11150 9260 11834
rect 9324 11762 9352 12038
rect 9312 11756 9364 11762
rect 9312 11698 9364 11704
rect 10232 11756 10284 11762
rect 10232 11698 10284 11704
rect 9220 11144 9272 11150
rect 9220 11086 9272 11092
rect 9128 10736 9180 10742
rect 9128 10678 9180 10684
rect 9324 10674 9352 11698
rect 10048 11688 10100 11694
rect 10048 11630 10100 11636
rect 9864 11552 9916 11558
rect 9864 11494 9916 11500
rect 9471 11452 9779 11461
rect 9471 11450 9477 11452
rect 9533 11450 9557 11452
rect 9613 11450 9637 11452
rect 9693 11450 9717 11452
rect 9773 11450 9779 11452
rect 9533 11398 9535 11450
rect 9715 11398 9717 11450
rect 9471 11396 9477 11398
rect 9533 11396 9557 11398
rect 9613 11396 9637 11398
rect 9693 11396 9717 11398
rect 9773 11396 9779 11398
rect 9471 11387 9779 11396
rect 9876 11218 9904 11494
rect 9864 11212 9916 11218
rect 9864 11154 9916 11160
rect 9772 11144 9824 11150
rect 9772 11086 9824 11092
rect 9784 11014 9812 11086
rect 10060 11082 10088 11630
rect 10048 11076 10100 11082
rect 10048 11018 10100 11024
rect 9772 11008 9824 11014
rect 9772 10950 9824 10956
rect 9312 10668 9364 10674
rect 9312 10610 9364 10616
rect 10060 10606 10088 11018
rect 10048 10600 10100 10606
rect 10048 10542 10100 10548
rect 9471 10364 9779 10373
rect 9471 10362 9477 10364
rect 9533 10362 9557 10364
rect 9613 10362 9637 10364
rect 9693 10362 9717 10364
rect 9773 10362 9779 10364
rect 9533 10310 9535 10362
rect 9715 10310 9717 10362
rect 9471 10308 9477 10310
rect 9533 10308 9557 10310
rect 9613 10308 9637 10310
rect 9693 10308 9717 10310
rect 9773 10308 9779 10310
rect 9471 10299 9779 10308
rect 9680 10124 9732 10130
rect 9680 10066 9732 10072
rect 9128 10056 9180 10062
rect 9128 9998 9180 10004
rect 9312 10056 9364 10062
rect 9312 9998 9364 10004
rect 9140 9586 9168 9998
rect 9128 9580 9180 9586
rect 9128 9522 9180 9528
rect 9324 9518 9352 9998
rect 9692 9654 9720 10066
rect 10060 10062 10088 10542
rect 10244 10538 10272 11698
rect 10232 10532 10284 10538
rect 10232 10474 10284 10480
rect 10048 10056 10100 10062
rect 10048 9998 10100 10004
rect 9680 9648 9732 9654
rect 9680 9590 9732 9596
rect 9956 9580 10008 9586
rect 9956 9522 10008 9528
rect 9312 9512 9364 9518
rect 9126 9480 9182 9489
rect 9496 9512 9548 9518
rect 9312 9454 9364 9460
rect 9494 9480 9496 9489
rect 9548 9480 9550 9489
rect 9126 9415 9182 9424
rect 9494 9415 9550 9424
rect 9140 8634 9168 9415
rect 9312 9376 9364 9382
rect 9312 9318 9364 9324
rect 9864 9376 9916 9382
rect 9864 9318 9916 9324
rect 9324 9178 9352 9318
rect 9471 9276 9779 9285
rect 9471 9274 9477 9276
rect 9533 9274 9557 9276
rect 9613 9274 9637 9276
rect 9693 9274 9717 9276
rect 9773 9274 9779 9276
rect 9533 9222 9535 9274
rect 9715 9222 9717 9274
rect 9471 9220 9477 9222
rect 9533 9220 9557 9222
rect 9613 9220 9637 9222
rect 9693 9220 9717 9222
rect 9773 9220 9779 9222
rect 9471 9211 9779 9220
rect 9876 9178 9904 9318
rect 9312 9172 9364 9178
rect 9312 9114 9364 9120
rect 9864 9172 9916 9178
rect 9864 9114 9916 9120
rect 9772 8968 9824 8974
rect 9772 8910 9824 8916
rect 9128 8628 9180 8634
rect 9128 8570 9180 8576
rect 9036 8560 9088 8566
rect 9036 8502 9088 8508
rect 8944 8492 8996 8498
rect 8944 8434 8996 8440
rect 8956 8090 8984 8434
rect 9312 8424 9364 8430
rect 9312 8366 9364 8372
rect 9220 8288 9272 8294
rect 9220 8230 9272 8236
rect 8944 8084 8996 8090
rect 8944 8026 8996 8032
rect 8956 7410 8984 8026
rect 9036 7812 9088 7818
rect 9036 7754 9088 7760
rect 9048 7546 9076 7754
rect 9036 7540 9088 7546
rect 9036 7482 9088 7488
rect 8944 7404 8996 7410
rect 8944 7346 8996 7352
rect 9232 6866 9260 8230
rect 9324 7954 9352 8366
rect 9784 8294 9812 8910
rect 9864 8356 9916 8362
rect 9864 8298 9916 8304
rect 9772 8288 9824 8294
rect 9772 8230 9824 8236
rect 9471 8188 9779 8197
rect 9471 8186 9477 8188
rect 9533 8186 9557 8188
rect 9613 8186 9637 8188
rect 9693 8186 9717 8188
rect 9773 8186 9779 8188
rect 9533 8134 9535 8186
rect 9715 8134 9717 8186
rect 9471 8132 9477 8134
rect 9533 8132 9557 8134
rect 9613 8132 9637 8134
rect 9693 8132 9717 8134
rect 9773 8132 9779 8134
rect 9471 8123 9779 8132
rect 9312 7948 9364 7954
rect 9312 7890 9364 7896
rect 9680 7948 9732 7954
rect 9680 7890 9732 7896
rect 9324 7274 9352 7890
rect 9692 7274 9720 7890
rect 9876 7834 9904 8298
rect 9784 7806 9904 7834
rect 9784 7478 9812 7806
rect 9864 7744 9916 7750
rect 9864 7686 9916 7692
rect 9772 7472 9824 7478
rect 9772 7414 9824 7420
rect 9312 7268 9364 7274
rect 9312 7210 9364 7216
rect 9680 7268 9732 7274
rect 9680 7210 9732 7216
rect 9471 7100 9779 7109
rect 9471 7098 9477 7100
rect 9533 7098 9557 7100
rect 9613 7098 9637 7100
rect 9693 7098 9717 7100
rect 9773 7098 9779 7100
rect 9533 7046 9535 7098
rect 9715 7046 9717 7098
rect 9471 7044 9477 7046
rect 9533 7044 9557 7046
rect 9613 7044 9637 7046
rect 9693 7044 9717 7046
rect 9773 7044 9779 7046
rect 9471 7035 9779 7044
rect 9876 6934 9904 7686
rect 9864 6928 9916 6934
rect 9864 6870 9916 6876
rect 9968 6866 9996 9522
rect 10048 8968 10100 8974
rect 10048 8910 10100 8916
rect 9220 6860 9272 6866
rect 9220 6802 9272 6808
rect 9956 6860 10008 6866
rect 9956 6802 10008 6808
rect 9312 6792 9364 6798
rect 9772 6792 9824 6798
rect 9364 6752 9536 6780
rect 9312 6734 9364 6740
rect 9220 6724 9272 6730
rect 9220 6666 9272 6672
rect 8942 6488 8998 6497
rect 8942 6423 8944 6432
rect 8996 6423 8998 6432
rect 8944 6394 8996 6400
rect 8852 6384 8904 6390
rect 8850 6352 8852 6361
rect 8904 6352 8906 6361
rect 8850 6287 8906 6296
rect 9128 6316 9180 6322
rect 9128 6258 9180 6264
rect 9140 6186 9168 6258
rect 9128 6180 9180 6186
rect 9128 6122 9180 6128
rect 9232 5914 9260 6666
rect 9508 6322 9536 6752
rect 9772 6734 9824 6740
rect 9680 6452 9732 6458
rect 9784 6440 9812 6734
rect 9954 6624 10010 6633
rect 9954 6559 10010 6568
rect 9732 6412 9812 6440
rect 9680 6394 9732 6400
rect 9968 6390 9996 6559
rect 10060 6458 10088 8910
rect 10244 8566 10272 10474
rect 10232 8560 10284 8566
rect 10232 8502 10284 8508
rect 10324 7404 10376 7410
rect 10244 7364 10324 7392
rect 10140 7336 10192 7342
rect 10140 7278 10192 7284
rect 10048 6452 10100 6458
rect 10152 6440 10180 7278
rect 10244 6662 10272 7364
rect 10324 7346 10376 7352
rect 10324 7200 10376 7206
rect 10324 7142 10376 7148
rect 10232 6656 10284 6662
rect 10336 6633 10364 7142
rect 10428 6798 10456 12406
rect 10508 12232 10560 12238
rect 10508 12174 10560 12180
rect 10520 11762 10548 12174
rect 10508 11756 10560 11762
rect 10508 11698 10560 11704
rect 10612 11150 10640 18566
rect 10692 16448 10744 16454
rect 10692 16390 10744 16396
rect 10704 15638 10732 16390
rect 10692 15632 10744 15638
rect 10692 15574 10744 15580
rect 10796 13938 10824 19654
rect 10876 18692 10928 18698
rect 10876 18634 10928 18640
rect 10888 17270 10916 18634
rect 10876 17264 10928 17270
rect 10876 17206 10928 17212
rect 11072 14482 11100 20538
rect 11256 15502 11284 20810
rect 11348 20262 11376 20810
rect 12716 20800 12768 20806
rect 12716 20742 12768 20748
rect 12311 20700 12619 20709
rect 12311 20698 12317 20700
rect 12373 20698 12397 20700
rect 12453 20698 12477 20700
rect 12533 20698 12557 20700
rect 12613 20698 12619 20700
rect 12373 20646 12375 20698
rect 12555 20646 12557 20698
rect 12311 20644 12317 20646
rect 12373 20644 12397 20646
rect 12453 20644 12477 20646
rect 12533 20644 12557 20646
rect 12613 20644 12619 20646
rect 12311 20635 12619 20644
rect 12728 20466 12756 20742
rect 12072 20460 12124 20466
rect 12072 20402 12124 20408
rect 12164 20460 12216 20466
rect 12164 20402 12216 20408
rect 12716 20460 12768 20466
rect 12716 20402 12768 20408
rect 11336 20256 11388 20262
rect 11336 20198 11388 20204
rect 11348 19718 11376 20198
rect 12084 20058 12112 20402
rect 12072 20052 12124 20058
rect 12072 19994 12124 20000
rect 12176 19922 12204 20402
rect 12164 19916 12216 19922
rect 12164 19858 12216 19864
rect 11336 19712 11388 19718
rect 11336 19654 11388 19660
rect 11244 15496 11296 15502
rect 11244 15438 11296 15444
rect 11152 15360 11204 15366
rect 11152 15302 11204 15308
rect 11060 14476 11112 14482
rect 11060 14418 11112 14424
rect 11164 14346 11192 15302
rect 11152 14340 11204 14346
rect 11152 14282 11204 14288
rect 11348 14278 11376 19654
rect 12311 19612 12619 19621
rect 12311 19610 12317 19612
rect 12373 19610 12397 19612
rect 12453 19610 12477 19612
rect 12533 19610 12557 19612
rect 12613 19610 12619 19612
rect 12373 19558 12375 19610
rect 12555 19558 12557 19610
rect 12311 19556 12317 19558
rect 12373 19556 12397 19558
rect 12453 19556 12477 19558
rect 12533 19556 12557 19558
rect 12613 19556 12619 19558
rect 12311 19547 12619 19556
rect 11980 19508 12032 19514
rect 11980 19450 12032 19456
rect 11796 17536 11848 17542
rect 11796 17478 11848 17484
rect 11704 16992 11756 16998
rect 11704 16934 11756 16940
rect 11716 16114 11744 16934
rect 11808 16658 11836 17478
rect 11888 17060 11940 17066
rect 11888 17002 11940 17008
rect 11796 16652 11848 16658
rect 11796 16594 11848 16600
rect 11900 16590 11928 17002
rect 11888 16584 11940 16590
rect 11888 16526 11940 16532
rect 11992 16114 12020 19450
rect 12072 18692 12124 18698
rect 12072 18634 12124 18640
rect 12084 17678 12112 18634
rect 12311 18524 12619 18533
rect 12311 18522 12317 18524
rect 12373 18522 12397 18524
rect 12453 18522 12477 18524
rect 12533 18522 12557 18524
rect 12613 18522 12619 18524
rect 12373 18470 12375 18522
rect 12555 18470 12557 18522
rect 12311 18468 12317 18470
rect 12373 18468 12397 18470
rect 12453 18468 12477 18470
rect 12533 18468 12557 18470
rect 12613 18468 12619 18470
rect 12311 18459 12619 18468
rect 12164 17808 12216 17814
rect 12164 17750 12216 17756
rect 12072 17672 12124 17678
rect 12072 17614 12124 17620
rect 12176 17338 12204 17750
rect 12311 17436 12619 17445
rect 12311 17434 12317 17436
rect 12373 17434 12397 17436
rect 12453 17434 12477 17436
rect 12533 17434 12557 17436
rect 12613 17434 12619 17436
rect 12373 17382 12375 17434
rect 12555 17382 12557 17434
rect 12311 17380 12317 17382
rect 12373 17380 12397 17382
rect 12453 17380 12477 17382
rect 12533 17380 12557 17382
rect 12613 17380 12619 17382
rect 12311 17371 12619 17380
rect 12164 17332 12216 17338
rect 12164 17274 12216 17280
rect 12176 16590 12204 17274
rect 12716 16652 12768 16658
rect 12716 16594 12768 16600
rect 12164 16584 12216 16590
rect 12164 16526 12216 16532
rect 12072 16448 12124 16454
rect 12072 16390 12124 16396
rect 11704 16108 11756 16114
rect 11704 16050 11756 16056
rect 11980 16108 12032 16114
rect 11980 16050 12032 16056
rect 11428 15564 11480 15570
rect 11428 15506 11480 15512
rect 11336 14272 11388 14278
rect 11336 14214 11388 14220
rect 10692 13932 10744 13938
rect 10692 13874 10744 13880
rect 10784 13932 10836 13938
rect 10784 13874 10836 13880
rect 10704 13326 10732 13874
rect 10692 13320 10744 13326
rect 10692 13262 10744 13268
rect 10704 12442 10732 13262
rect 10692 12436 10744 12442
rect 10692 12378 10744 12384
rect 10796 12306 10824 13874
rect 11348 13530 11376 14214
rect 11336 13524 11388 13530
rect 11336 13466 11388 13472
rect 11152 12776 11204 12782
rect 11152 12718 11204 12724
rect 10968 12436 11020 12442
rect 10968 12378 11020 12384
rect 10784 12300 10836 12306
rect 10784 12242 10836 12248
rect 10692 12232 10744 12238
rect 10692 12174 10744 12180
rect 10600 11144 10652 11150
rect 10600 11086 10652 11092
rect 10506 10704 10562 10713
rect 10506 10639 10562 10648
rect 10520 10470 10548 10639
rect 10508 10464 10560 10470
rect 10508 10406 10560 10412
rect 10520 9926 10548 10406
rect 10600 9988 10652 9994
rect 10600 9930 10652 9936
rect 10508 9920 10560 9926
rect 10506 9888 10508 9897
rect 10560 9888 10562 9897
rect 10506 9823 10562 9832
rect 10508 8356 10560 8362
rect 10508 8298 10560 8304
rect 10416 6792 10468 6798
rect 10416 6734 10468 6740
rect 10232 6598 10284 6604
rect 10322 6624 10378 6633
rect 10322 6559 10378 6568
rect 10152 6412 10272 6440
rect 10048 6394 10100 6400
rect 9956 6384 10008 6390
rect 9956 6326 10008 6332
rect 10244 6322 10272 6412
rect 9496 6316 9548 6322
rect 9496 6258 9548 6264
rect 10140 6316 10192 6322
rect 10140 6258 10192 6264
rect 10232 6316 10284 6322
rect 10232 6258 10284 6264
rect 10048 6248 10100 6254
rect 10048 6190 10100 6196
rect 9471 6012 9779 6021
rect 9471 6010 9477 6012
rect 9533 6010 9557 6012
rect 9613 6010 9637 6012
rect 9693 6010 9717 6012
rect 9773 6010 9779 6012
rect 9533 5958 9535 6010
rect 9715 5958 9717 6010
rect 9471 5956 9477 5958
rect 9533 5956 9557 5958
rect 9613 5956 9637 5958
rect 9693 5956 9717 5958
rect 9773 5956 9779 5958
rect 9471 5947 9779 5956
rect 9220 5908 9272 5914
rect 9220 5850 9272 5856
rect 8760 5772 8812 5778
rect 8760 5714 8812 5720
rect 8668 5704 8720 5710
rect 8668 5646 8720 5652
rect 9126 5536 9182 5545
rect 9126 5471 9182 5480
rect 8576 5228 8628 5234
rect 8628 5188 8708 5216
rect 8576 5170 8628 5176
rect 8576 5092 8628 5098
rect 8576 5034 8628 5040
rect 8484 4684 8536 4690
rect 8484 4626 8536 4632
rect 8484 4276 8536 4282
rect 8484 4218 8536 4224
rect 8022 4176 8078 4185
rect 8022 4111 8078 4120
rect 8300 4140 8352 4146
rect 8300 4082 8352 4088
rect 8208 4072 8260 4078
rect 8208 4014 8260 4020
rect 8220 3194 8248 4014
rect 8312 3534 8340 4082
rect 8496 3670 8524 4218
rect 8484 3664 8536 3670
rect 8484 3606 8536 3612
rect 8300 3528 8352 3534
rect 8300 3470 8352 3476
rect 8484 3528 8536 3534
rect 8588 3516 8616 5034
rect 8680 4146 8708 5188
rect 9140 5030 9168 5471
rect 9680 5160 9732 5166
rect 9678 5128 9680 5137
rect 9732 5128 9734 5137
rect 9678 5063 9734 5072
rect 9128 5024 9180 5030
rect 9128 4966 9180 4972
rect 9471 4924 9779 4933
rect 9471 4922 9477 4924
rect 9533 4922 9557 4924
rect 9613 4922 9637 4924
rect 9693 4922 9717 4924
rect 9773 4922 9779 4924
rect 9533 4870 9535 4922
rect 9715 4870 9717 4922
rect 9471 4868 9477 4870
rect 9533 4868 9557 4870
rect 9613 4868 9637 4870
rect 9693 4868 9717 4870
rect 9773 4868 9779 4870
rect 9471 4859 9779 4868
rect 9128 4820 9180 4826
rect 9128 4762 9180 4768
rect 9036 4208 9088 4214
rect 9036 4150 9088 4156
rect 8668 4140 8720 4146
rect 8668 4082 8720 4088
rect 8680 4049 8708 4082
rect 8944 4072 8996 4078
rect 8666 4040 8722 4049
rect 8944 4014 8996 4020
rect 8666 3975 8722 3984
rect 8956 3534 8984 4014
rect 8536 3488 8616 3516
rect 8484 3470 8536 3476
rect 8208 3188 8260 3194
rect 8208 3130 8260 3136
rect 8588 3126 8616 3488
rect 8944 3528 8996 3534
rect 8944 3470 8996 3476
rect 9048 3380 9076 4150
rect 9140 3942 9168 4762
rect 10060 4758 10088 6190
rect 10152 5817 10180 6258
rect 10138 5808 10194 5817
rect 10138 5743 10194 5752
rect 10244 5710 10272 6258
rect 10140 5704 10192 5710
rect 10140 5646 10192 5652
rect 10232 5704 10284 5710
rect 10232 5646 10284 5652
rect 10152 4826 10180 5646
rect 10140 4820 10192 4826
rect 10140 4762 10192 4768
rect 10048 4752 10100 4758
rect 10048 4694 10100 4700
rect 10428 4690 10456 6734
rect 10520 6254 10548 8298
rect 10612 7886 10640 9930
rect 10704 8498 10732 12174
rect 10784 11756 10836 11762
rect 10784 11698 10836 11704
rect 10692 8492 10744 8498
rect 10692 8434 10744 8440
rect 10796 8294 10824 11698
rect 10980 11558 11008 12378
rect 11060 11824 11112 11830
rect 11060 11766 11112 11772
rect 10968 11552 11020 11558
rect 10968 11494 11020 11500
rect 10968 11076 11020 11082
rect 10968 11018 11020 11024
rect 10876 10804 10928 10810
rect 10876 10746 10928 10752
rect 10888 8634 10916 10746
rect 10980 9586 11008 11018
rect 11072 9586 11100 11766
rect 10968 9580 11020 9586
rect 10968 9522 11020 9528
rect 11060 9580 11112 9586
rect 11060 9522 11112 9528
rect 11060 9376 11112 9382
rect 11060 9318 11112 9324
rect 10968 8832 11020 8838
rect 10968 8774 11020 8780
rect 10876 8628 10928 8634
rect 10876 8570 10928 8576
rect 10784 8288 10836 8294
rect 10784 8230 10836 8236
rect 10600 7880 10652 7886
rect 10600 7822 10652 7828
rect 10784 7880 10836 7886
rect 10784 7822 10836 7828
rect 10600 7268 10652 7274
rect 10600 7210 10652 7216
rect 10612 6866 10640 7210
rect 10600 6860 10652 6866
rect 10600 6802 10652 6808
rect 10600 6656 10652 6662
rect 10600 6598 10652 6604
rect 10508 6248 10560 6254
rect 10508 6190 10560 6196
rect 10520 5710 10548 6190
rect 10612 6118 10640 6598
rect 10796 6186 10824 7822
rect 10980 7818 11008 8774
rect 10968 7812 11020 7818
rect 10968 7754 11020 7760
rect 10876 7744 10928 7750
rect 10876 7686 10928 7692
rect 10784 6180 10836 6186
rect 10784 6122 10836 6128
rect 10600 6112 10652 6118
rect 10600 6054 10652 6060
rect 10692 6112 10744 6118
rect 10692 6054 10744 6060
rect 10508 5704 10560 5710
rect 10508 5646 10560 5652
rect 10704 5574 10732 6054
rect 10796 5710 10824 6122
rect 10888 5817 10916 7686
rect 10980 7478 11008 7754
rect 10968 7472 11020 7478
rect 10968 7414 11020 7420
rect 11072 7342 11100 9318
rect 11164 8090 11192 12718
rect 11244 11756 11296 11762
rect 11244 11698 11296 11704
rect 11256 8922 11284 11698
rect 11256 8894 11376 8922
rect 11152 8084 11204 8090
rect 11152 8026 11204 8032
rect 11164 7834 11192 8026
rect 11164 7806 11284 7834
rect 11152 7744 11204 7750
rect 11152 7686 11204 7692
rect 11060 7336 11112 7342
rect 11164 7313 11192 7686
rect 11256 7546 11284 7806
rect 11244 7540 11296 7546
rect 11244 7482 11296 7488
rect 11060 7278 11112 7284
rect 11150 7304 11206 7313
rect 10968 6724 11020 6730
rect 10968 6666 11020 6672
rect 10980 6186 11008 6666
rect 11072 6458 11100 7278
rect 11150 7239 11206 7248
rect 11256 7154 11284 7482
rect 11164 7126 11284 7154
rect 11164 6934 11192 7126
rect 11244 6996 11296 7002
rect 11244 6938 11296 6944
rect 11152 6928 11204 6934
rect 11152 6870 11204 6876
rect 11152 6792 11204 6798
rect 11152 6734 11204 6740
rect 11060 6452 11112 6458
rect 11060 6394 11112 6400
rect 10968 6180 11020 6186
rect 10968 6122 11020 6128
rect 10874 5808 10930 5817
rect 10874 5743 10930 5752
rect 10784 5704 10836 5710
rect 10784 5646 10836 5652
rect 10692 5568 10744 5574
rect 10692 5510 10744 5516
rect 11072 5234 11100 6394
rect 11060 5228 11112 5234
rect 11060 5170 11112 5176
rect 11164 4826 11192 6734
rect 11256 6390 11284 6938
rect 11348 6662 11376 8894
rect 11336 6656 11388 6662
rect 11336 6598 11388 6604
rect 11244 6384 11296 6390
rect 11244 6326 11296 6332
rect 11440 5846 11468 15506
rect 11612 13728 11664 13734
rect 11612 13670 11664 13676
rect 11624 11898 11652 13670
rect 11716 13326 11744 16050
rect 11796 15496 11848 15502
rect 11796 15438 11848 15444
rect 11888 15496 11940 15502
rect 11888 15438 11940 15444
rect 11808 15094 11836 15438
rect 11900 15162 11928 15438
rect 11888 15156 11940 15162
rect 11888 15098 11940 15104
rect 11796 15088 11848 15094
rect 11796 15030 11848 15036
rect 11808 14890 11836 15030
rect 11796 14884 11848 14890
rect 11796 14826 11848 14832
rect 11808 14346 11836 14826
rect 11900 14550 11928 15098
rect 11888 14544 11940 14550
rect 11888 14486 11940 14492
rect 11796 14340 11848 14346
rect 11796 14282 11848 14288
rect 11808 13870 11836 14282
rect 11796 13864 11848 13870
rect 11796 13806 11848 13812
rect 11704 13320 11756 13326
rect 11704 13262 11756 13268
rect 11716 12918 11744 13262
rect 11704 12912 11756 12918
rect 11704 12854 11756 12860
rect 11808 12850 11836 13806
rect 11888 13184 11940 13190
rect 11888 13126 11940 13132
rect 11900 12986 11928 13126
rect 11888 12980 11940 12986
rect 11888 12922 11940 12928
rect 11796 12844 11848 12850
rect 11796 12786 11848 12792
rect 11808 12646 11836 12786
rect 11796 12640 11848 12646
rect 11796 12582 11848 12588
rect 11900 12170 11928 12922
rect 11992 12850 12020 16050
rect 12084 15978 12112 16390
rect 12311 16348 12619 16357
rect 12311 16346 12317 16348
rect 12373 16346 12397 16348
rect 12453 16346 12477 16348
rect 12533 16346 12557 16348
rect 12613 16346 12619 16348
rect 12373 16294 12375 16346
rect 12555 16294 12557 16346
rect 12311 16292 12317 16294
rect 12373 16292 12397 16294
rect 12453 16292 12477 16294
rect 12533 16292 12557 16294
rect 12613 16292 12619 16294
rect 12311 16283 12619 16292
rect 12164 16040 12216 16046
rect 12164 15982 12216 15988
rect 12072 15972 12124 15978
rect 12072 15914 12124 15920
rect 12176 14532 12204 15982
rect 12311 15260 12619 15269
rect 12311 15258 12317 15260
rect 12373 15258 12397 15260
rect 12453 15258 12477 15260
rect 12533 15258 12557 15260
rect 12613 15258 12619 15260
rect 12373 15206 12375 15258
rect 12555 15206 12557 15258
rect 12311 15204 12317 15206
rect 12373 15204 12397 15206
rect 12453 15204 12477 15206
rect 12533 15204 12557 15206
rect 12613 15204 12619 15206
rect 12311 15195 12619 15204
rect 12624 15020 12676 15026
rect 12624 14962 12676 14968
rect 12084 14504 12204 14532
rect 12084 13326 12112 14504
rect 12348 14476 12400 14482
rect 12176 14436 12348 14464
rect 12072 13320 12124 13326
rect 12072 13262 12124 13268
rect 12072 12912 12124 12918
rect 12072 12854 12124 12860
rect 11980 12844 12032 12850
rect 11980 12786 12032 12792
rect 11992 12442 12020 12786
rect 11980 12436 12032 12442
rect 11980 12378 12032 12384
rect 12084 12306 12112 12854
rect 12176 12442 12204 14436
rect 12348 14418 12400 14424
rect 12636 14362 12664 14962
rect 12728 14482 12756 16594
rect 12820 14618 12848 20896
rect 12912 19922 12940 21354
rect 13096 20777 13124 21490
rect 13268 21480 13320 21486
rect 13268 21422 13320 21428
rect 13924 21434 13952 21542
rect 14004 21548 14056 21554
rect 14004 21490 14056 21496
rect 14096 21548 14148 21554
rect 14096 21490 14148 21496
rect 14108 21434 14136 21490
rect 13280 20806 13308 21422
rect 13924 21406 14136 21434
rect 14372 21412 14424 21418
rect 13452 21072 13504 21078
rect 13452 21014 13504 21020
rect 13636 21072 13688 21078
rect 13636 21014 13688 21020
rect 13360 20868 13412 20874
rect 13360 20810 13412 20816
rect 13268 20800 13320 20806
rect 13082 20768 13138 20777
rect 13268 20742 13320 20748
rect 13082 20703 13138 20712
rect 13176 20460 13228 20466
rect 13176 20402 13228 20408
rect 12900 19916 12952 19922
rect 12900 19858 12952 19864
rect 13084 19780 13136 19786
rect 13084 19722 13136 19728
rect 12992 19304 13044 19310
rect 12992 19246 13044 19252
rect 12900 18828 12952 18834
rect 12900 18770 12952 18776
rect 12912 18222 12940 18770
rect 13004 18766 13032 19246
rect 12992 18760 13044 18766
rect 12992 18702 13044 18708
rect 12900 18216 12952 18222
rect 12900 18158 12952 18164
rect 12912 17542 12940 18158
rect 12900 17536 12952 17542
rect 12900 17478 12952 17484
rect 13004 16946 13032 18702
rect 13096 17066 13124 19722
rect 13188 17202 13216 20402
rect 13280 19990 13308 20742
rect 13372 20641 13400 20810
rect 13358 20632 13414 20641
rect 13358 20567 13414 20576
rect 13268 19984 13320 19990
rect 13266 19952 13268 19961
rect 13320 19952 13322 19961
rect 13266 19887 13322 19896
rect 13464 19854 13492 21014
rect 13648 20534 13676 21014
rect 13636 20528 13688 20534
rect 13636 20470 13688 20476
rect 13544 20460 13596 20466
rect 13544 20402 13596 20408
rect 13452 19848 13504 19854
rect 13452 19790 13504 19796
rect 13268 18828 13320 18834
rect 13268 18770 13320 18776
rect 13280 18086 13308 18770
rect 13360 18760 13412 18766
rect 13360 18702 13412 18708
rect 13268 18080 13320 18086
rect 13268 18022 13320 18028
rect 13372 17954 13400 18702
rect 13556 18426 13584 20402
rect 13634 20360 13690 20369
rect 13634 20295 13636 20304
rect 13688 20295 13690 20304
rect 13636 20266 13688 20272
rect 13544 18420 13596 18426
rect 13544 18362 13596 18368
rect 13280 17926 13400 17954
rect 13280 17610 13308 17926
rect 13820 17672 13872 17678
rect 13820 17614 13872 17620
rect 13268 17604 13320 17610
rect 13268 17546 13320 17552
rect 13176 17196 13228 17202
rect 13176 17138 13228 17144
rect 13084 17060 13136 17066
rect 13084 17002 13136 17008
rect 13004 16918 13124 16946
rect 13096 16590 13124 16918
rect 13280 16794 13308 17546
rect 13636 17128 13688 17134
rect 13636 17070 13688 17076
rect 13268 16788 13320 16794
rect 13268 16730 13320 16736
rect 12992 16584 13044 16590
rect 12992 16526 13044 16532
rect 13084 16584 13136 16590
rect 13084 16526 13136 16532
rect 12900 15428 12952 15434
rect 12900 15370 12952 15376
rect 12912 15094 12940 15370
rect 12900 15088 12952 15094
rect 12900 15030 12952 15036
rect 12900 14952 12952 14958
rect 12900 14894 12952 14900
rect 12808 14612 12860 14618
rect 12808 14554 12860 14560
rect 12716 14476 12768 14482
rect 12716 14418 12768 14424
rect 12808 14408 12860 14414
rect 12636 14334 12756 14362
rect 12808 14350 12860 14356
rect 12311 14172 12619 14181
rect 12311 14170 12317 14172
rect 12373 14170 12397 14172
rect 12453 14170 12477 14172
rect 12533 14170 12557 14172
rect 12613 14170 12619 14172
rect 12373 14118 12375 14170
rect 12555 14118 12557 14170
rect 12311 14116 12317 14118
rect 12373 14116 12397 14118
rect 12453 14116 12477 14118
rect 12533 14116 12557 14118
rect 12613 14116 12619 14118
rect 12311 14107 12619 14116
rect 12728 13938 12756 14334
rect 12820 14074 12848 14350
rect 12808 14068 12860 14074
rect 12808 14010 12860 14016
rect 12716 13932 12768 13938
rect 12716 13874 12768 13880
rect 12311 13084 12619 13093
rect 12311 13082 12317 13084
rect 12373 13082 12397 13084
rect 12453 13082 12477 13084
rect 12533 13082 12557 13084
rect 12613 13082 12619 13084
rect 12373 13030 12375 13082
rect 12555 13030 12557 13082
rect 12311 13028 12317 13030
rect 12373 13028 12397 13030
rect 12453 13028 12477 13030
rect 12533 13028 12557 13030
rect 12613 13028 12619 13030
rect 12311 13019 12619 13028
rect 12728 12918 12756 13874
rect 12716 12912 12768 12918
rect 12716 12854 12768 12860
rect 12912 12850 12940 14894
rect 13004 13258 13032 16526
rect 13084 15904 13136 15910
rect 13084 15846 13136 15852
rect 13096 15026 13124 15846
rect 13280 15706 13308 16730
rect 13268 15700 13320 15706
rect 13268 15642 13320 15648
rect 13544 15496 13596 15502
rect 13544 15438 13596 15444
rect 13084 15020 13136 15026
rect 13084 14962 13136 14968
rect 13268 15020 13320 15026
rect 13268 14962 13320 14968
rect 13280 14328 13308 14962
rect 13556 14890 13584 15438
rect 13544 14884 13596 14890
rect 13544 14826 13596 14832
rect 13360 14816 13412 14822
rect 13360 14758 13412 14764
rect 13372 14550 13400 14758
rect 13360 14544 13412 14550
rect 13360 14486 13412 14492
rect 13556 14414 13584 14826
rect 13544 14408 13596 14414
rect 13544 14350 13596 14356
rect 13360 14340 13412 14346
rect 13280 14300 13360 14328
rect 13360 14282 13412 14288
rect 13082 14104 13138 14113
rect 13082 14039 13138 14048
rect 13096 14006 13124 14039
rect 13084 14000 13136 14006
rect 13084 13942 13136 13948
rect 13372 13462 13400 14282
rect 13360 13456 13412 13462
rect 13360 13398 13412 13404
rect 12992 13252 13044 13258
rect 12992 13194 13044 13200
rect 12900 12844 12952 12850
rect 12900 12786 12952 12792
rect 12532 12640 12584 12646
rect 12532 12582 12584 12588
rect 12164 12436 12216 12442
rect 12164 12378 12216 12384
rect 12544 12374 12572 12582
rect 12532 12368 12584 12374
rect 12532 12310 12584 12316
rect 12072 12300 12124 12306
rect 12072 12242 12124 12248
rect 11888 12164 11940 12170
rect 11888 12106 11940 12112
rect 11612 11892 11664 11898
rect 11612 11834 11664 11840
rect 11704 11824 11756 11830
rect 11900 11812 11928 12106
rect 11980 11824 12032 11830
rect 11900 11784 11980 11812
rect 11704 11766 11756 11772
rect 11980 11766 12032 11772
rect 11716 10742 11744 11766
rect 12084 11762 12112 12242
rect 12311 11996 12619 12005
rect 12311 11994 12317 11996
rect 12373 11994 12397 11996
rect 12453 11994 12477 11996
rect 12533 11994 12557 11996
rect 12613 11994 12619 11996
rect 12373 11942 12375 11994
rect 12555 11942 12557 11994
rect 12311 11940 12317 11942
rect 12373 11940 12397 11942
rect 12453 11940 12477 11942
rect 12533 11940 12557 11942
rect 12613 11940 12619 11942
rect 12311 11931 12619 11940
rect 12716 11824 12768 11830
rect 12622 11792 12678 11801
rect 12072 11756 12124 11762
rect 12716 11766 12768 11772
rect 12622 11727 12678 11736
rect 12072 11698 12124 11704
rect 12636 11150 12664 11727
rect 11888 11144 11940 11150
rect 11888 11086 11940 11092
rect 12624 11144 12676 11150
rect 12624 11086 12676 11092
rect 11900 10810 11928 11086
rect 12164 11008 12216 11014
rect 12164 10950 12216 10956
rect 11888 10804 11940 10810
rect 11888 10746 11940 10752
rect 11704 10736 11756 10742
rect 11704 10678 11756 10684
rect 12176 10452 12204 10950
rect 12311 10908 12619 10917
rect 12311 10906 12317 10908
rect 12373 10906 12397 10908
rect 12453 10906 12477 10908
rect 12533 10906 12557 10908
rect 12613 10906 12619 10908
rect 12373 10854 12375 10906
rect 12555 10854 12557 10906
rect 12311 10852 12317 10854
rect 12373 10852 12397 10854
rect 12453 10852 12477 10854
rect 12533 10852 12557 10854
rect 12613 10852 12619 10854
rect 12311 10843 12619 10852
rect 12256 10464 12308 10470
rect 12176 10424 12256 10452
rect 12256 10406 12308 10412
rect 12268 10198 12296 10406
rect 12256 10192 12308 10198
rect 12256 10134 12308 10140
rect 12728 10062 12756 11766
rect 13004 11082 13032 13194
rect 13372 12918 13400 13398
rect 13360 12912 13412 12918
rect 13360 12854 13412 12860
rect 13176 12844 13228 12850
rect 13176 12786 13228 12792
rect 13188 12434 13216 12786
rect 13096 12406 13216 12434
rect 13096 11354 13124 12406
rect 13176 12368 13228 12374
rect 13174 12336 13176 12345
rect 13228 12336 13230 12345
rect 13174 12271 13230 12280
rect 13268 12300 13320 12306
rect 13188 11898 13216 12271
rect 13268 12242 13320 12248
rect 13176 11892 13228 11898
rect 13176 11834 13228 11840
rect 13280 11370 13308 12242
rect 13372 12102 13400 12854
rect 13360 12096 13412 12102
rect 13360 12038 13412 12044
rect 13084 11348 13136 11354
rect 13084 11290 13136 11296
rect 13188 11342 13308 11370
rect 13372 11676 13400 12038
rect 13452 11688 13504 11694
rect 13372 11648 13452 11676
rect 13084 11144 13136 11150
rect 13084 11086 13136 11092
rect 12992 11076 13044 11082
rect 12992 11018 13044 11024
rect 13096 10985 13124 11086
rect 13082 10976 13138 10985
rect 13082 10911 13138 10920
rect 13096 10792 13124 10911
rect 13004 10764 13124 10792
rect 12900 10736 12952 10742
rect 13004 10724 13032 10764
rect 12952 10696 13032 10724
rect 12900 10678 12952 10684
rect 13084 10668 13136 10674
rect 13084 10610 13136 10616
rect 12808 10600 12860 10606
rect 12808 10542 12860 10548
rect 12716 10056 12768 10062
rect 12716 9998 12768 10004
rect 12716 9920 12768 9926
rect 12716 9862 12768 9868
rect 12311 9820 12619 9829
rect 12311 9818 12317 9820
rect 12373 9818 12397 9820
rect 12453 9818 12477 9820
rect 12533 9818 12557 9820
rect 12613 9818 12619 9820
rect 12373 9766 12375 9818
rect 12555 9766 12557 9818
rect 12311 9764 12317 9766
rect 12373 9764 12397 9766
rect 12453 9764 12477 9766
rect 12533 9764 12557 9766
rect 12613 9764 12619 9766
rect 12311 9755 12619 9764
rect 11612 9512 11664 9518
rect 11612 9454 11664 9460
rect 11624 8974 11652 9454
rect 12072 9444 12124 9450
rect 12072 9386 12124 9392
rect 11520 8968 11572 8974
rect 11520 8910 11572 8916
rect 11612 8968 11664 8974
rect 11612 8910 11664 8916
rect 11532 6730 11560 8910
rect 11624 8430 11652 8910
rect 11704 8900 11756 8906
rect 11704 8842 11756 8848
rect 11716 8498 11744 8842
rect 12084 8634 12112 9386
rect 12624 9376 12676 9382
rect 12624 9318 12676 9324
rect 12636 9042 12664 9318
rect 12624 9036 12676 9042
rect 12624 8978 12676 8984
rect 12311 8732 12619 8741
rect 12311 8730 12317 8732
rect 12373 8730 12397 8732
rect 12453 8730 12477 8732
rect 12533 8730 12557 8732
rect 12613 8730 12619 8732
rect 12373 8678 12375 8730
rect 12555 8678 12557 8730
rect 12311 8676 12317 8678
rect 12373 8676 12397 8678
rect 12453 8676 12477 8678
rect 12533 8676 12557 8678
rect 12613 8676 12619 8678
rect 12311 8667 12619 8676
rect 12072 8628 12124 8634
rect 12072 8570 12124 8576
rect 11704 8492 11756 8498
rect 11704 8434 11756 8440
rect 11888 8492 11940 8498
rect 11888 8434 11940 8440
rect 12164 8492 12216 8498
rect 12164 8434 12216 8440
rect 11612 8424 11664 8430
rect 11612 8366 11664 8372
rect 11624 7478 11652 8366
rect 11704 8016 11756 8022
rect 11756 7976 11836 8004
rect 11704 7958 11756 7964
rect 11612 7472 11664 7478
rect 11612 7414 11664 7420
rect 11624 6934 11652 7414
rect 11704 7200 11756 7206
rect 11704 7142 11756 7148
rect 11612 6928 11664 6934
rect 11612 6870 11664 6876
rect 11520 6724 11572 6730
rect 11520 6666 11572 6672
rect 11716 6662 11744 7142
rect 11612 6656 11664 6662
rect 11612 6598 11664 6604
rect 11704 6656 11756 6662
rect 11704 6598 11756 6604
rect 11624 5846 11652 6598
rect 11716 5953 11744 6598
rect 11808 6304 11836 7976
rect 11900 7546 11928 8434
rect 11980 7880 12032 7886
rect 11980 7822 12032 7828
rect 11888 7540 11940 7546
rect 11888 7482 11940 7488
rect 11992 6633 12020 7822
rect 12072 7540 12124 7546
rect 12072 7482 12124 7488
rect 12084 7206 12112 7482
rect 12176 7426 12204 8434
rect 12311 7644 12619 7653
rect 12311 7642 12317 7644
rect 12373 7642 12397 7644
rect 12453 7642 12477 7644
rect 12533 7642 12557 7644
rect 12613 7642 12619 7644
rect 12373 7590 12375 7642
rect 12555 7590 12557 7642
rect 12311 7588 12317 7590
rect 12373 7588 12397 7590
rect 12453 7588 12477 7590
rect 12533 7588 12557 7590
rect 12613 7588 12619 7590
rect 12311 7579 12619 7588
rect 12728 7546 12756 9862
rect 12820 9450 12848 10542
rect 12900 10532 12952 10538
rect 12900 10474 12952 10480
rect 12808 9444 12860 9450
rect 12808 9386 12860 9392
rect 12912 9382 12940 10474
rect 12992 10056 13044 10062
rect 12992 9998 13044 10004
rect 13004 9654 13032 9998
rect 12992 9648 13044 9654
rect 12992 9590 13044 9596
rect 12900 9376 12952 9382
rect 12900 9318 12952 9324
rect 12912 8906 12940 9318
rect 13096 9110 13124 10610
rect 13188 9178 13216 11342
rect 13372 11268 13400 11648
rect 13452 11630 13504 11636
rect 13544 11552 13596 11558
rect 13544 11494 13596 11500
rect 13556 11354 13584 11494
rect 13544 11348 13596 11354
rect 13544 11290 13596 11296
rect 13280 11240 13400 11268
rect 13280 9994 13308 11240
rect 13452 11144 13504 11150
rect 13452 11086 13504 11092
rect 13360 11076 13412 11082
rect 13360 11018 13412 11024
rect 13372 10810 13400 11018
rect 13464 10849 13492 11086
rect 13450 10840 13506 10849
rect 13360 10804 13412 10810
rect 13450 10775 13506 10784
rect 13360 10746 13412 10752
rect 13372 10198 13400 10746
rect 13464 10470 13492 10775
rect 13452 10464 13504 10470
rect 13452 10406 13504 10412
rect 13556 10266 13584 11290
rect 13648 10810 13676 17070
rect 13832 16574 13860 17614
rect 13740 16546 13860 16574
rect 13740 12782 13768 16546
rect 13924 16436 13952 21406
rect 14372 21354 14424 21360
rect 14280 20936 14332 20942
rect 14280 20878 14332 20884
rect 14188 19236 14240 19242
rect 14188 19178 14240 19184
rect 14004 18352 14056 18358
rect 14004 18294 14056 18300
rect 14016 17338 14044 18294
rect 14004 17332 14056 17338
rect 14004 17274 14056 17280
rect 14096 17332 14148 17338
rect 14096 17274 14148 17280
rect 14108 17218 14136 17274
rect 13832 16408 13952 16436
rect 14016 17190 14136 17218
rect 13832 14618 13860 16408
rect 13912 15904 13964 15910
rect 13912 15846 13964 15852
rect 13924 15502 13952 15846
rect 13912 15496 13964 15502
rect 13912 15438 13964 15444
rect 13820 14612 13872 14618
rect 13820 14554 13872 14560
rect 13728 12776 13780 12782
rect 13728 12718 13780 12724
rect 13740 12434 13768 12718
rect 13740 12406 13860 12434
rect 13728 11688 13780 11694
rect 13728 11630 13780 11636
rect 13636 10804 13688 10810
rect 13636 10746 13688 10752
rect 13544 10260 13596 10266
rect 13544 10202 13596 10208
rect 13360 10192 13412 10198
rect 13360 10134 13412 10140
rect 13740 10130 13768 11630
rect 13832 11150 13860 12406
rect 13820 11144 13872 11150
rect 13820 11086 13872 11092
rect 13924 10849 13952 15438
rect 14016 14346 14044 17190
rect 14096 17128 14148 17134
rect 14096 17070 14148 17076
rect 14108 16726 14136 17070
rect 14096 16720 14148 16726
rect 14096 16662 14148 16668
rect 14200 16590 14228 19178
rect 14292 18970 14320 20878
rect 14280 18964 14332 18970
rect 14280 18906 14332 18912
rect 14384 18698 14412 21354
rect 14568 21078 14596 21558
rect 15120 21554 15148 21830
rect 15108 21548 15160 21554
rect 15108 21490 15160 21496
rect 14924 21480 14976 21486
rect 14924 21422 14976 21428
rect 15016 21480 15068 21486
rect 15016 21422 15068 21428
rect 14648 21344 14700 21350
rect 14648 21286 14700 21292
rect 14464 21072 14516 21078
rect 14464 21014 14516 21020
rect 14556 21072 14608 21078
rect 14556 21014 14608 21020
rect 14476 20777 14504 21014
rect 14462 20768 14518 20777
rect 14462 20703 14518 20712
rect 14660 20262 14688 21286
rect 14832 20868 14884 20874
rect 14832 20810 14884 20816
rect 14740 20460 14792 20466
rect 14740 20402 14792 20408
rect 14648 20256 14700 20262
rect 14648 20198 14700 20204
rect 14660 19854 14688 20198
rect 14648 19848 14700 19854
rect 14648 19790 14700 19796
rect 14752 19378 14780 20402
rect 14844 20398 14872 20810
rect 14936 20602 14964 21422
rect 14924 20596 14976 20602
rect 14924 20538 14976 20544
rect 14924 20460 14976 20466
rect 14924 20402 14976 20408
rect 14832 20392 14884 20398
rect 14832 20334 14884 20340
rect 14936 19904 14964 20402
rect 15028 20058 15056 21422
rect 15152 21244 15460 21253
rect 15152 21242 15158 21244
rect 15214 21242 15238 21244
rect 15294 21242 15318 21244
rect 15374 21242 15398 21244
rect 15454 21242 15460 21244
rect 15214 21190 15216 21242
rect 15396 21190 15398 21242
rect 15152 21188 15158 21190
rect 15214 21188 15238 21190
rect 15294 21188 15318 21190
rect 15374 21188 15398 21190
rect 15454 21188 15460 21190
rect 15152 21179 15460 21188
rect 15568 21072 15620 21078
rect 15568 21014 15620 21020
rect 15476 20936 15528 20942
rect 15476 20878 15528 20884
rect 15292 20868 15344 20874
rect 15292 20810 15344 20816
rect 15304 20312 15332 20810
rect 15488 20806 15516 20878
rect 15384 20800 15436 20806
rect 15384 20742 15436 20748
rect 15476 20800 15528 20806
rect 15476 20742 15528 20748
rect 15396 20534 15424 20742
rect 15384 20528 15436 20534
rect 15384 20470 15436 20476
rect 15580 20466 15608 21014
rect 15672 20942 15700 21830
rect 16210 21584 16266 21593
rect 17696 21554 17724 21830
rect 17992 21788 18300 21797
rect 17992 21786 17998 21788
rect 18054 21786 18078 21788
rect 18134 21786 18158 21788
rect 18214 21786 18238 21788
rect 18294 21786 18300 21788
rect 18054 21734 18056 21786
rect 18236 21734 18238 21786
rect 17992 21732 17998 21734
rect 18054 21732 18078 21734
rect 18134 21732 18158 21734
rect 18214 21732 18238 21734
rect 18294 21732 18300 21734
rect 17992 21723 18300 21732
rect 19996 21690 20024 21966
rect 21192 21690 21220 22034
rect 22388 22030 22416 24200
rect 22376 22024 22428 22030
rect 22376 21966 22428 21972
rect 22376 21888 22428 21894
rect 22376 21830 22428 21836
rect 19156 21684 19208 21690
rect 19156 21626 19208 21632
rect 19984 21684 20036 21690
rect 19984 21626 20036 21632
rect 21180 21684 21232 21690
rect 21180 21626 21232 21632
rect 16210 21519 16266 21528
rect 17040 21548 17092 21554
rect 15752 21412 15804 21418
rect 15752 21354 15804 21360
rect 15660 20936 15712 20942
rect 15660 20878 15712 20884
rect 15660 20800 15712 20806
rect 15660 20742 15712 20748
rect 15568 20460 15620 20466
rect 15568 20402 15620 20408
rect 15476 20324 15528 20330
rect 15304 20284 15476 20312
rect 15476 20266 15528 20272
rect 15152 20156 15460 20165
rect 15152 20154 15158 20156
rect 15214 20154 15238 20156
rect 15294 20154 15318 20156
rect 15374 20154 15398 20156
rect 15454 20154 15460 20156
rect 15214 20102 15216 20154
rect 15396 20102 15398 20154
rect 15152 20100 15158 20102
rect 15214 20100 15238 20102
rect 15294 20100 15318 20102
rect 15374 20100 15398 20102
rect 15454 20100 15460 20102
rect 15152 20091 15460 20100
rect 15016 20052 15068 20058
rect 15016 19994 15068 20000
rect 15292 19984 15344 19990
rect 15290 19952 15292 19961
rect 15344 19952 15346 19961
rect 15016 19916 15068 19922
rect 14936 19876 15016 19904
rect 15290 19887 15346 19896
rect 15384 19916 15436 19922
rect 15016 19858 15068 19864
rect 15384 19858 15436 19864
rect 15396 19825 15424 19858
rect 15382 19816 15438 19825
rect 15382 19751 15438 19760
rect 14924 19712 14976 19718
rect 14924 19654 14976 19660
rect 14556 19372 14608 19378
rect 14740 19372 14792 19378
rect 14556 19314 14608 19320
rect 14660 19332 14740 19360
rect 14464 19168 14516 19174
rect 14464 19110 14516 19116
rect 14476 18766 14504 19110
rect 14568 18970 14596 19314
rect 14556 18964 14608 18970
rect 14556 18906 14608 18912
rect 14464 18760 14516 18766
rect 14464 18702 14516 18708
rect 14372 18692 14424 18698
rect 14372 18634 14424 18640
rect 14556 18692 14608 18698
rect 14556 18634 14608 18640
rect 14464 18624 14516 18630
rect 14384 18572 14464 18578
rect 14384 18566 14516 18572
rect 14384 18550 14504 18566
rect 14280 17060 14332 17066
rect 14280 17002 14332 17008
rect 14292 16794 14320 17002
rect 14384 16998 14412 18550
rect 14464 18148 14516 18154
rect 14464 18090 14516 18096
rect 14476 17678 14504 18090
rect 14568 17882 14596 18634
rect 14556 17876 14608 17882
rect 14556 17818 14608 17824
rect 14464 17672 14516 17678
rect 14464 17614 14516 17620
rect 14556 17196 14608 17202
rect 14556 17138 14608 17144
rect 14464 17128 14516 17134
rect 14464 17070 14516 17076
rect 14372 16992 14424 16998
rect 14372 16934 14424 16940
rect 14280 16788 14332 16794
rect 14280 16730 14332 16736
rect 14188 16584 14240 16590
rect 14188 16526 14240 16532
rect 14292 16436 14320 16730
rect 14384 16590 14412 16934
rect 14372 16584 14424 16590
rect 14372 16526 14424 16532
rect 14372 16448 14424 16454
rect 14292 16408 14372 16436
rect 14372 16390 14424 16396
rect 14096 16040 14148 16046
rect 14096 15982 14148 15988
rect 14004 14340 14056 14346
rect 14004 14282 14056 14288
rect 14108 13734 14136 15982
rect 14188 14952 14240 14958
rect 14188 14894 14240 14900
rect 14200 14482 14228 14894
rect 14188 14476 14240 14482
rect 14188 14418 14240 14424
rect 14280 14408 14332 14414
rect 14280 14350 14332 14356
rect 14188 14340 14240 14346
rect 14188 14282 14240 14288
rect 14096 13728 14148 13734
rect 14096 13670 14148 13676
rect 14004 13184 14056 13190
rect 14004 13126 14056 13132
rect 14016 12238 14044 13126
rect 14108 12782 14136 13670
rect 14096 12776 14148 12782
rect 14096 12718 14148 12724
rect 14004 12232 14056 12238
rect 14004 12174 14056 12180
rect 14200 11830 14228 14282
rect 14292 13870 14320 14350
rect 14280 13864 14332 13870
rect 14280 13806 14332 13812
rect 14280 13320 14332 13326
rect 14280 13262 14332 13268
rect 14292 12866 14320 13262
rect 14384 13002 14412 16390
rect 14476 13938 14504 17070
rect 14568 14414 14596 17138
rect 14660 16658 14688 19332
rect 14740 19314 14792 19320
rect 14832 19168 14884 19174
rect 14832 19110 14884 19116
rect 14844 18902 14872 19110
rect 14832 18896 14884 18902
rect 14832 18838 14884 18844
rect 14740 18692 14792 18698
rect 14740 18634 14792 18640
rect 14752 18426 14780 18634
rect 14740 18420 14792 18426
rect 14740 18362 14792 18368
rect 14832 18284 14884 18290
rect 14832 18226 14884 18232
rect 14844 17610 14872 18226
rect 14832 17604 14884 17610
rect 14832 17546 14884 17552
rect 14740 17060 14792 17066
rect 14740 17002 14792 17008
rect 14752 16726 14780 17002
rect 14844 16794 14872 17546
rect 14936 16794 14964 19654
rect 15198 19408 15254 19417
rect 15198 19343 15200 19352
rect 15252 19343 15254 19352
rect 15200 19314 15252 19320
rect 15212 19242 15240 19314
rect 15200 19236 15252 19242
rect 15200 19178 15252 19184
rect 15488 19122 15516 20266
rect 15580 19242 15608 20402
rect 15672 19310 15700 20742
rect 15764 20602 15792 21354
rect 16224 21078 16252 21519
rect 17040 21490 17092 21496
rect 17684 21548 17736 21554
rect 17684 21490 17736 21496
rect 16488 21344 16540 21350
rect 16540 21292 16620 21298
rect 16488 21286 16620 21292
rect 16500 21270 16620 21286
rect 16500 21146 16528 21270
rect 16488 21140 16540 21146
rect 16488 21082 16540 21088
rect 16212 21072 16264 21078
rect 16212 21014 16264 21020
rect 16120 20936 16172 20942
rect 16120 20878 16172 20884
rect 15752 20596 15804 20602
rect 15752 20538 15804 20544
rect 15752 20460 15804 20466
rect 15752 20402 15804 20408
rect 15936 20460 15988 20466
rect 15936 20402 15988 20408
rect 15764 19938 15792 20402
rect 15764 19910 15884 19938
rect 15750 19544 15806 19553
rect 15750 19479 15806 19488
rect 15764 19446 15792 19479
rect 15752 19440 15804 19446
rect 15752 19382 15804 19388
rect 15660 19304 15712 19310
rect 15660 19246 15712 19252
rect 15568 19236 15620 19242
rect 15568 19178 15620 19184
rect 15488 19094 15608 19122
rect 15152 19068 15460 19077
rect 15152 19066 15158 19068
rect 15214 19066 15238 19068
rect 15294 19066 15318 19068
rect 15374 19066 15398 19068
rect 15454 19066 15460 19068
rect 15214 19014 15216 19066
rect 15396 19014 15398 19066
rect 15152 19012 15158 19014
rect 15214 19012 15238 19014
rect 15294 19012 15318 19014
rect 15374 19012 15398 19014
rect 15454 19012 15460 19014
rect 15152 19003 15460 19012
rect 15292 18964 15344 18970
rect 15292 18906 15344 18912
rect 15304 18698 15332 18906
rect 15292 18692 15344 18698
rect 15292 18634 15344 18640
rect 15304 18170 15332 18634
rect 15028 18142 15332 18170
rect 15476 18216 15528 18222
rect 15476 18158 15528 18164
rect 15028 17796 15056 18142
rect 15152 17980 15460 17989
rect 15152 17978 15158 17980
rect 15214 17978 15238 17980
rect 15294 17978 15318 17980
rect 15374 17978 15398 17980
rect 15454 17978 15460 17980
rect 15214 17926 15216 17978
rect 15396 17926 15398 17978
rect 15152 17924 15158 17926
rect 15214 17924 15238 17926
rect 15294 17924 15318 17926
rect 15374 17924 15398 17926
rect 15454 17924 15460 17926
rect 15152 17915 15460 17924
rect 15028 17768 15148 17796
rect 15016 17264 15068 17270
rect 15016 17206 15068 17212
rect 14832 16788 14884 16794
rect 14832 16730 14884 16736
rect 14924 16788 14976 16794
rect 14924 16730 14976 16736
rect 14740 16720 14792 16726
rect 14740 16662 14792 16668
rect 14648 16652 14700 16658
rect 14648 16594 14700 16600
rect 14660 14464 14688 16594
rect 14740 16244 14792 16250
rect 14740 16186 14792 16192
rect 14752 15502 14780 16186
rect 15028 15706 15056 17206
rect 15120 17134 15148 17768
rect 15108 17128 15160 17134
rect 15108 17070 15160 17076
rect 15292 17128 15344 17134
rect 15292 17070 15344 17076
rect 15304 16998 15332 17070
rect 15292 16992 15344 16998
rect 15292 16934 15344 16940
rect 15152 16892 15460 16901
rect 15152 16890 15158 16892
rect 15214 16890 15238 16892
rect 15294 16890 15318 16892
rect 15374 16890 15398 16892
rect 15454 16890 15460 16892
rect 15214 16838 15216 16890
rect 15396 16838 15398 16890
rect 15152 16836 15158 16838
rect 15214 16836 15238 16838
rect 15294 16836 15318 16838
rect 15374 16836 15398 16838
rect 15454 16836 15460 16838
rect 15152 16827 15460 16836
rect 15152 15804 15460 15813
rect 15152 15802 15158 15804
rect 15214 15802 15238 15804
rect 15294 15802 15318 15804
rect 15374 15802 15398 15804
rect 15454 15802 15460 15804
rect 15214 15750 15216 15802
rect 15396 15750 15398 15802
rect 15152 15748 15158 15750
rect 15214 15748 15238 15750
rect 15294 15748 15318 15750
rect 15374 15748 15398 15750
rect 15454 15748 15460 15750
rect 15152 15739 15460 15748
rect 15016 15700 15068 15706
rect 15016 15642 15068 15648
rect 15016 15564 15068 15570
rect 15016 15506 15068 15512
rect 14740 15496 14792 15502
rect 14740 15438 14792 15444
rect 14752 15366 14780 15438
rect 14740 15360 14792 15366
rect 14740 15302 14792 15308
rect 14924 15020 14976 15026
rect 14924 14962 14976 14968
rect 14832 14884 14884 14890
rect 14832 14826 14884 14832
rect 14660 14436 14780 14464
rect 14556 14408 14608 14414
rect 14556 14350 14608 14356
rect 14464 13932 14516 13938
rect 14464 13874 14516 13880
rect 14476 13326 14504 13874
rect 14464 13320 14516 13326
rect 14464 13262 14516 13268
rect 14568 13190 14596 14350
rect 14648 14340 14700 14346
rect 14648 14282 14700 14288
rect 14660 13326 14688 14282
rect 14752 13394 14780 14436
rect 14740 13388 14792 13394
rect 14740 13330 14792 13336
rect 14648 13320 14700 13326
rect 14648 13262 14700 13268
rect 14556 13184 14608 13190
rect 14556 13126 14608 13132
rect 14648 13184 14700 13190
rect 14648 13126 14700 13132
rect 14384 12974 14596 13002
rect 14292 12838 14504 12866
rect 14372 12300 14424 12306
rect 14476 12288 14504 12838
rect 14424 12260 14504 12288
rect 14372 12242 14424 12248
rect 14280 12232 14332 12238
rect 14278 12200 14280 12209
rect 14332 12200 14334 12209
rect 14278 12135 14334 12144
rect 14188 11824 14240 11830
rect 14188 11766 14240 11772
rect 14372 11552 14424 11558
rect 14372 11494 14424 11500
rect 14280 11144 14332 11150
rect 14278 11112 14280 11121
rect 14332 11112 14334 11121
rect 14188 11076 14240 11082
rect 14278 11047 14334 11056
rect 14188 11018 14240 11024
rect 14200 10985 14228 11018
rect 14186 10976 14242 10985
rect 14186 10911 14242 10920
rect 13910 10840 13966 10849
rect 13910 10775 13966 10784
rect 13912 10736 13964 10742
rect 13912 10678 13964 10684
rect 13924 10266 13952 10678
rect 13912 10260 13964 10266
rect 13912 10202 13964 10208
rect 13728 10124 13780 10130
rect 13728 10066 13780 10072
rect 13268 9988 13320 9994
rect 13268 9930 13320 9936
rect 13176 9172 13228 9178
rect 13176 9114 13228 9120
rect 13084 9104 13136 9110
rect 13084 9046 13136 9052
rect 13096 8974 13124 9046
rect 13084 8968 13136 8974
rect 13084 8910 13136 8916
rect 12900 8900 12952 8906
rect 12900 8842 12952 8848
rect 12808 8628 12860 8634
rect 12808 8570 12860 8576
rect 12820 7750 12848 8570
rect 12900 8288 12952 8294
rect 12900 8230 12952 8236
rect 12808 7744 12860 7750
rect 12808 7686 12860 7692
rect 12716 7540 12768 7546
rect 12716 7482 12768 7488
rect 12176 7398 12296 7426
rect 12164 7336 12216 7342
rect 12164 7278 12216 7284
rect 12072 7200 12124 7206
rect 12072 7142 12124 7148
rect 12176 6866 12204 7278
rect 12164 6860 12216 6866
rect 12164 6802 12216 6808
rect 12268 6712 12296 7398
rect 12716 7268 12768 7274
rect 12716 7210 12768 7216
rect 12348 6996 12400 7002
rect 12348 6938 12400 6944
rect 12084 6684 12296 6712
rect 11978 6624 12034 6633
rect 11978 6559 12034 6568
rect 11980 6316 12032 6322
rect 11808 6276 11980 6304
rect 11980 6258 12032 6264
rect 11702 5944 11758 5953
rect 11702 5879 11704 5888
rect 11756 5879 11758 5888
rect 11704 5850 11756 5856
rect 11428 5840 11480 5846
rect 11428 5782 11480 5788
rect 11612 5840 11664 5846
rect 11716 5819 11744 5850
rect 11612 5782 11664 5788
rect 10784 4820 10836 4826
rect 10784 4762 10836 4768
rect 11152 4820 11204 4826
rect 11152 4762 11204 4768
rect 9864 4684 9916 4690
rect 9864 4626 9916 4632
rect 10416 4684 10468 4690
rect 10416 4626 10468 4632
rect 9312 4480 9364 4486
rect 9312 4422 9364 4428
rect 9220 4004 9272 4010
rect 9220 3946 9272 3952
rect 9128 3936 9180 3942
rect 9128 3878 9180 3884
rect 9140 3534 9168 3878
rect 9232 3738 9260 3946
rect 9324 3738 9352 4422
rect 9471 3836 9779 3845
rect 9471 3834 9477 3836
rect 9533 3834 9557 3836
rect 9613 3834 9637 3836
rect 9693 3834 9717 3836
rect 9773 3834 9779 3836
rect 9533 3782 9535 3834
rect 9715 3782 9717 3834
rect 9471 3780 9477 3782
rect 9533 3780 9557 3782
rect 9613 3780 9637 3782
rect 9693 3780 9717 3782
rect 9773 3780 9779 3782
rect 9471 3771 9779 3780
rect 9220 3732 9272 3738
rect 9220 3674 9272 3680
rect 9312 3732 9364 3738
rect 9312 3674 9364 3680
rect 9588 3732 9640 3738
rect 9588 3674 9640 3680
rect 9232 3590 9536 3618
rect 9128 3528 9180 3534
rect 9128 3470 9180 3476
rect 9232 3380 9260 3590
rect 9508 3534 9536 3590
rect 9312 3528 9364 3534
rect 9312 3470 9364 3476
rect 9496 3528 9548 3534
rect 9496 3470 9548 3476
rect 9048 3352 9260 3380
rect 9324 3194 9352 3470
rect 9600 3194 9628 3674
rect 9876 3194 9904 4626
rect 10324 4616 10376 4622
rect 10324 4558 10376 4564
rect 10336 4282 10364 4558
rect 10324 4276 10376 4282
rect 10324 4218 10376 4224
rect 10796 4146 10824 4762
rect 10692 4140 10744 4146
rect 10692 4082 10744 4088
rect 10784 4140 10836 4146
rect 10784 4082 10836 4088
rect 10600 3596 10652 3602
rect 10600 3538 10652 3544
rect 9312 3188 9364 3194
rect 9312 3130 9364 3136
rect 9588 3188 9640 3194
rect 9588 3130 9640 3136
rect 9864 3188 9916 3194
rect 9864 3130 9916 3136
rect 8576 3120 8628 3126
rect 8576 3062 8628 3068
rect 10612 3058 10640 3538
rect 10704 3126 10732 4082
rect 10968 4072 11020 4078
rect 10968 4014 11020 4020
rect 10692 3120 10744 3126
rect 10980 3097 11008 4014
rect 11152 3392 11204 3398
rect 11152 3334 11204 3340
rect 11244 3392 11296 3398
rect 11244 3334 11296 3340
rect 10692 3062 10744 3068
rect 10966 3088 11022 3097
rect 10600 3052 10652 3058
rect 10966 3023 11022 3032
rect 11060 3052 11112 3058
rect 10600 2994 10652 3000
rect 11060 2994 11112 3000
rect 10612 2938 10640 2994
rect 11072 2961 11100 2994
rect 8576 2916 8628 2922
rect 8576 2858 8628 2864
rect 10428 2910 10640 2938
rect 11058 2952 11114 2961
rect 8588 800 8616 2858
rect 10428 2854 10456 2910
rect 11164 2938 11192 3334
rect 11256 3194 11284 3334
rect 11440 3194 11468 5782
rect 11992 5658 12020 6258
rect 12084 5914 12112 6684
rect 12360 6662 12388 6938
rect 12348 6656 12400 6662
rect 12162 6624 12218 6633
rect 12348 6598 12400 6604
rect 12162 6559 12218 6568
rect 12176 6322 12204 6559
rect 12311 6556 12619 6565
rect 12311 6554 12317 6556
rect 12373 6554 12397 6556
rect 12453 6554 12477 6556
rect 12533 6554 12557 6556
rect 12613 6554 12619 6556
rect 12373 6502 12375 6554
rect 12555 6502 12557 6554
rect 12311 6500 12317 6502
rect 12373 6500 12397 6502
rect 12453 6500 12477 6502
rect 12533 6500 12557 6502
rect 12613 6500 12619 6502
rect 12311 6491 12619 6500
rect 12164 6316 12216 6322
rect 12164 6258 12216 6264
rect 12728 6254 12756 7210
rect 12820 7002 12848 7686
rect 12912 7410 12940 8230
rect 13188 7886 13216 9114
rect 13280 8566 13308 9930
rect 13636 9580 13688 9586
rect 13636 9522 13688 9528
rect 13648 8974 13676 9522
rect 13636 8968 13688 8974
rect 13636 8910 13688 8916
rect 13268 8560 13320 8566
rect 13268 8502 13320 8508
rect 13648 8362 13676 8910
rect 13740 8906 13768 10066
rect 14384 9586 14412 11494
rect 14476 9994 14504 12260
rect 14568 11234 14596 12974
rect 14660 11354 14688 13126
rect 14752 12918 14780 13330
rect 14740 12912 14792 12918
rect 14740 12854 14792 12860
rect 14740 12232 14792 12238
rect 14740 12174 14792 12180
rect 14752 11558 14780 12174
rect 14740 11552 14792 11558
rect 14740 11494 14792 11500
rect 14648 11348 14700 11354
rect 14648 11290 14700 11296
rect 14738 11248 14794 11257
rect 14568 11206 14688 11234
rect 14660 10674 14688 11206
rect 14738 11183 14794 11192
rect 14648 10668 14700 10674
rect 14648 10610 14700 10616
rect 14464 9988 14516 9994
rect 14464 9930 14516 9936
rect 14660 9926 14688 10610
rect 14752 10062 14780 11183
rect 14844 10810 14872 14826
rect 14936 14618 14964 14962
rect 14924 14612 14976 14618
rect 14924 14554 14976 14560
rect 14924 13932 14976 13938
rect 14924 13874 14976 13880
rect 14936 11257 14964 13874
rect 15028 12306 15056 15506
rect 15200 15496 15252 15502
rect 15200 15438 15252 15444
rect 15212 14958 15240 15438
rect 15488 15162 15516 18158
rect 15580 15978 15608 19094
rect 15672 18970 15700 19246
rect 15660 18964 15712 18970
rect 15660 18906 15712 18912
rect 15752 18760 15804 18766
rect 15752 18702 15804 18708
rect 15660 18624 15712 18630
rect 15660 18566 15712 18572
rect 15672 16590 15700 18566
rect 15764 18057 15792 18702
rect 15750 18048 15806 18057
rect 15750 17983 15806 17992
rect 15856 17626 15884 19910
rect 15948 19718 15976 20402
rect 16028 19848 16080 19854
rect 16028 19790 16080 19796
rect 15936 19712 15988 19718
rect 15936 19654 15988 19660
rect 15948 19378 15976 19654
rect 15936 19372 15988 19378
rect 15936 19314 15988 19320
rect 16040 18970 16068 19790
rect 16028 18964 16080 18970
rect 16028 18906 16080 18912
rect 16132 18442 16160 20878
rect 16304 20460 16356 20466
rect 16304 20402 16356 20408
rect 16316 20262 16344 20402
rect 16304 20256 16356 20262
rect 16304 20198 16356 20204
rect 16304 19984 16356 19990
rect 16304 19926 16356 19932
rect 16488 19984 16540 19990
rect 16488 19926 16540 19932
rect 16040 18414 16160 18442
rect 16316 19836 16344 19926
rect 16396 19848 16448 19854
rect 16316 19808 16396 19836
rect 16040 18086 16068 18414
rect 16120 18352 16172 18358
rect 16120 18294 16172 18300
rect 16132 18086 16160 18294
rect 16028 18080 16080 18086
rect 16028 18022 16080 18028
rect 16120 18080 16172 18086
rect 16120 18022 16172 18028
rect 15764 17598 15884 17626
rect 15764 17134 15792 17598
rect 15844 17536 15896 17542
rect 15844 17478 15896 17484
rect 15752 17128 15804 17134
rect 15752 17070 15804 17076
rect 15752 16720 15804 16726
rect 15752 16662 15804 16668
rect 15660 16584 15712 16590
rect 15660 16526 15712 16532
rect 15568 15972 15620 15978
rect 15568 15914 15620 15920
rect 15660 15904 15712 15910
rect 15660 15846 15712 15852
rect 15672 15502 15700 15846
rect 15660 15496 15712 15502
rect 15660 15438 15712 15444
rect 15764 15178 15792 16662
rect 15856 16590 15884 17478
rect 15936 17196 15988 17202
rect 15936 17138 15988 17144
rect 15844 16584 15896 16590
rect 15844 16526 15896 16532
rect 15476 15156 15528 15162
rect 15764 15150 15884 15178
rect 15476 15098 15528 15104
rect 15200 14952 15252 14958
rect 15200 14894 15252 14900
rect 15152 14716 15460 14725
rect 15152 14714 15158 14716
rect 15214 14714 15238 14716
rect 15294 14714 15318 14716
rect 15374 14714 15398 14716
rect 15454 14714 15460 14716
rect 15214 14662 15216 14714
rect 15396 14662 15398 14714
rect 15152 14660 15158 14662
rect 15214 14660 15238 14662
rect 15294 14660 15318 14662
rect 15374 14660 15398 14662
rect 15454 14660 15460 14662
rect 15152 14651 15460 14660
rect 15200 14544 15252 14550
rect 15200 14486 15252 14492
rect 15212 14006 15240 14486
rect 15384 14476 15436 14482
rect 15384 14418 15436 14424
rect 15396 14278 15424 14418
rect 15488 14346 15516 15098
rect 15568 15020 15620 15026
rect 15568 14962 15620 14968
rect 15476 14340 15528 14346
rect 15476 14282 15528 14288
rect 15384 14272 15436 14278
rect 15384 14214 15436 14220
rect 15200 14000 15252 14006
rect 15200 13942 15252 13948
rect 15476 13728 15528 13734
rect 15476 13670 15528 13676
rect 15152 13628 15460 13637
rect 15152 13626 15158 13628
rect 15214 13626 15238 13628
rect 15294 13626 15318 13628
rect 15374 13626 15398 13628
rect 15454 13626 15460 13628
rect 15214 13574 15216 13626
rect 15396 13574 15398 13626
rect 15152 13572 15158 13574
rect 15214 13572 15238 13574
rect 15294 13572 15318 13574
rect 15374 13572 15398 13574
rect 15454 13572 15460 13574
rect 15152 13563 15460 13572
rect 15488 13326 15516 13670
rect 15292 13320 15344 13326
rect 15292 13262 15344 13268
rect 15476 13320 15528 13326
rect 15476 13262 15528 13268
rect 15304 13190 15332 13262
rect 15292 13184 15344 13190
rect 15292 13126 15344 13132
rect 15476 13184 15528 13190
rect 15476 13126 15528 13132
rect 15152 12540 15460 12549
rect 15152 12538 15158 12540
rect 15214 12538 15238 12540
rect 15294 12538 15318 12540
rect 15374 12538 15398 12540
rect 15454 12538 15460 12540
rect 15214 12486 15216 12538
rect 15396 12486 15398 12538
rect 15152 12484 15158 12486
rect 15214 12484 15238 12486
rect 15294 12484 15318 12486
rect 15374 12484 15398 12486
rect 15454 12484 15460 12486
rect 15152 12475 15460 12484
rect 15488 12442 15516 13126
rect 15476 12436 15528 12442
rect 15476 12378 15528 12384
rect 15016 12300 15068 12306
rect 15016 12242 15068 12248
rect 15108 11824 15160 11830
rect 15106 11792 15108 11801
rect 15160 11792 15162 11801
rect 15106 11727 15162 11736
rect 15152 11452 15460 11461
rect 15152 11450 15158 11452
rect 15214 11450 15238 11452
rect 15294 11450 15318 11452
rect 15374 11450 15398 11452
rect 15454 11450 15460 11452
rect 15214 11398 15216 11450
rect 15396 11398 15398 11450
rect 15152 11396 15158 11398
rect 15214 11396 15238 11398
rect 15294 11396 15318 11398
rect 15374 11396 15398 11398
rect 15454 11396 15460 11398
rect 15152 11387 15460 11396
rect 15016 11280 15068 11286
rect 14922 11248 14978 11257
rect 15016 11222 15068 11228
rect 14922 11183 14978 11192
rect 14924 11144 14976 11150
rect 14922 11112 14924 11121
rect 14976 11112 14978 11121
rect 14922 11047 14978 11056
rect 15028 10826 15056 11222
rect 15384 11212 15436 11218
rect 15384 11154 15436 11160
rect 15108 11076 15160 11082
rect 15108 11018 15160 11024
rect 15120 10849 15148 11018
rect 14832 10804 14884 10810
rect 14832 10746 14884 10752
rect 14936 10798 15056 10826
rect 15106 10840 15162 10849
rect 14936 10674 14964 10798
rect 15106 10775 15162 10784
rect 15396 10674 15424 11154
rect 15488 10742 15516 12378
rect 15580 12374 15608 14962
rect 15660 14272 15712 14278
rect 15660 14214 15712 14220
rect 15672 14113 15700 14214
rect 15658 14104 15714 14113
rect 15658 14039 15714 14048
rect 15856 14006 15884 15150
rect 15948 14414 15976 17138
rect 16040 16998 16068 18022
rect 16028 16992 16080 16998
rect 16028 16934 16080 16940
rect 16040 16833 16068 16934
rect 16026 16824 16082 16833
rect 16026 16759 16082 16768
rect 16040 16726 16068 16759
rect 16028 16720 16080 16726
rect 16028 16662 16080 16668
rect 16132 15366 16160 18022
rect 16316 17678 16344 19808
rect 16396 19790 16448 19796
rect 16500 19514 16528 19926
rect 16488 19508 16540 19514
rect 16488 19450 16540 19456
rect 16592 18834 16620 21270
rect 16672 20936 16724 20942
rect 16672 20878 16724 20884
rect 16948 20936 17000 20942
rect 16948 20878 17000 20884
rect 16684 20369 16712 20878
rect 16960 20466 16988 20878
rect 16948 20460 17000 20466
rect 16948 20402 17000 20408
rect 16670 20360 16726 20369
rect 16670 20295 16726 20304
rect 16764 19984 16816 19990
rect 16764 19926 16816 19932
rect 16672 19440 16724 19446
rect 16776 19417 16804 19926
rect 17052 19854 17080 21490
rect 18328 20936 18380 20942
rect 18328 20878 18380 20884
rect 17992 20700 18300 20709
rect 17992 20698 17998 20700
rect 18054 20698 18078 20700
rect 18134 20698 18158 20700
rect 18214 20698 18238 20700
rect 18294 20698 18300 20700
rect 18054 20646 18056 20698
rect 18236 20646 18238 20698
rect 17992 20644 17998 20646
rect 18054 20644 18078 20646
rect 18134 20644 18158 20646
rect 18214 20644 18238 20646
rect 18294 20644 18300 20646
rect 17866 20632 17922 20641
rect 17992 20635 18300 20644
rect 17316 20596 17368 20602
rect 17866 20567 17868 20576
rect 17316 20538 17368 20544
rect 17920 20567 17922 20576
rect 17868 20538 17920 20544
rect 17328 20448 17356 20538
rect 17684 20460 17736 20466
rect 17328 20420 17448 20448
rect 17040 19848 17092 19854
rect 16854 19816 16910 19825
rect 17040 19790 17092 19796
rect 16854 19751 16856 19760
rect 16908 19751 16910 19760
rect 16856 19722 16908 19728
rect 16672 19382 16724 19388
rect 16762 19408 16818 19417
rect 16580 18828 16632 18834
rect 16580 18770 16632 18776
rect 16684 18766 16712 19382
rect 16762 19343 16818 19352
rect 16488 18760 16540 18766
rect 16488 18702 16540 18708
rect 16672 18760 16724 18766
rect 16672 18702 16724 18708
rect 16948 18760 17000 18766
rect 16948 18702 17000 18708
rect 16500 18426 16528 18702
rect 16488 18420 16540 18426
rect 16488 18362 16540 18368
rect 16304 17672 16356 17678
rect 16304 17614 16356 17620
rect 16488 17672 16540 17678
rect 16488 17614 16540 17620
rect 16316 16726 16344 17614
rect 16396 17536 16448 17542
rect 16396 17478 16448 17484
rect 16408 17134 16436 17478
rect 16396 17128 16448 17134
rect 16396 17070 16448 17076
rect 16304 16720 16356 16726
rect 16304 16662 16356 16668
rect 16212 15496 16264 15502
rect 16212 15438 16264 15444
rect 16120 15360 16172 15366
rect 16120 15302 16172 15308
rect 16224 14822 16252 15438
rect 16316 14890 16344 16662
rect 16500 16046 16528 17614
rect 16580 17536 16632 17542
rect 16580 17478 16632 17484
rect 16488 16040 16540 16046
rect 16488 15982 16540 15988
rect 16592 15434 16620 17478
rect 16684 16454 16712 18702
rect 16856 18148 16908 18154
rect 16856 18090 16908 18096
rect 16672 16448 16724 16454
rect 16672 16390 16724 16396
rect 16684 15502 16712 16390
rect 16868 15638 16896 18090
rect 16960 18086 16988 18702
rect 16948 18080 17000 18086
rect 16948 18022 17000 18028
rect 16960 16522 16988 18022
rect 17052 17202 17080 19790
rect 17130 19544 17186 19553
rect 17130 19479 17186 19488
rect 17144 19378 17172 19479
rect 17314 19408 17370 19417
rect 17132 19372 17184 19378
rect 17314 19343 17316 19352
rect 17132 19314 17184 19320
rect 17368 19343 17370 19352
rect 17316 19314 17368 19320
rect 17132 18692 17184 18698
rect 17132 18634 17184 18640
rect 17040 17196 17092 17202
rect 17040 17138 17092 17144
rect 17052 16726 17080 17138
rect 17144 17066 17172 18634
rect 17420 18630 17448 20420
rect 17684 20402 17736 20408
rect 17696 20330 17724 20402
rect 17684 20324 17736 20330
rect 17684 20266 17736 20272
rect 17696 20040 17724 20266
rect 17512 20012 17724 20040
rect 17408 18624 17460 18630
rect 17408 18566 17460 18572
rect 17224 18420 17276 18426
rect 17224 18362 17276 18368
rect 17132 17060 17184 17066
rect 17132 17002 17184 17008
rect 17040 16720 17092 16726
rect 17040 16662 17092 16668
rect 17040 16584 17092 16590
rect 17040 16526 17092 16532
rect 16948 16516 17000 16522
rect 16948 16458 17000 16464
rect 17052 16096 17080 16526
rect 17144 16182 17172 17002
rect 17132 16176 17184 16182
rect 17132 16118 17184 16124
rect 16960 16068 17080 16096
rect 16856 15632 16908 15638
rect 16856 15574 16908 15580
rect 16672 15496 16724 15502
rect 16672 15438 16724 15444
rect 16580 15428 16632 15434
rect 16580 15370 16632 15376
rect 16396 15360 16448 15366
rect 16396 15302 16448 15308
rect 16488 15360 16540 15366
rect 16488 15302 16540 15308
rect 16408 15042 16436 15302
rect 16500 15162 16528 15302
rect 16488 15156 16540 15162
rect 16488 15098 16540 15104
rect 16408 15014 16528 15042
rect 16960 15026 16988 16068
rect 17040 15972 17092 15978
rect 17040 15914 17092 15920
rect 16304 14884 16356 14890
rect 16304 14826 16356 14832
rect 16212 14816 16264 14822
rect 16212 14758 16264 14764
rect 16224 14482 16252 14758
rect 16212 14476 16264 14482
rect 16212 14418 16264 14424
rect 15936 14408 15988 14414
rect 15936 14350 15988 14356
rect 16120 14272 16172 14278
rect 16120 14214 16172 14220
rect 16132 14074 16160 14214
rect 16120 14068 16172 14074
rect 16120 14010 16172 14016
rect 15844 14000 15896 14006
rect 15844 13942 15896 13948
rect 16028 14000 16080 14006
rect 16028 13942 16080 13948
rect 15752 13932 15804 13938
rect 15752 13874 15804 13880
rect 15936 13932 15988 13938
rect 15936 13874 15988 13880
rect 15660 13864 15712 13870
rect 15660 13806 15712 13812
rect 15672 13734 15700 13806
rect 15660 13728 15712 13734
rect 15660 13670 15712 13676
rect 15672 12918 15700 13670
rect 15764 13530 15792 13874
rect 15948 13841 15976 13874
rect 15934 13832 15990 13841
rect 15934 13767 15990 13776
rect 15752 13524 15804 13530
rect 15752 13466 15804 13472
rect 16040 13462 16068 13942
rect 16028 13456 16080 13462
rect 16028 13398 16080 13404
rect 16316 13274 16344 14826
rect 16396 14544 16448 14550
rect 16396 14486 16448 14492
rect 15844 13252 15896 13258
rect 15844 13194 15896 13200
rect 16132 13246 16344 13274
rect 15660 12912 15712 12918
rect 15660 12854 15712 12860
rect 15660 12776 15712 12782
rect 15660 12718 15712 12724
rect 15568 12368 15620 12374
rect 15568 12310 15620 12316
rect 15672 11694 15700 12718
rect 15856 12434 15884 13194
rect 16132 13190 16160 13246
rect 16120 13184 16172 13190
rect 16120 13126 16172 13132
rect 16304 13184 16356 13190
rect 16304 13126 16356 13132
rect 16118 13016 16174 13025
rect 16118 12951 16174 12960
rect 15934 12880 15990 12889
rect 15934 12815 15990 12824
rect 15948 12782 15976 12815
rect 16132 12782 16160 12951
rect 15936 12776 15988 12782
rect 15936 12718 15988 12724
rect 16120 12776 16172 12782
rect 16172 12736 16252 12764
rect 16120 12718 16172 12724
rect 15764 12406 15884 12434
rect 15764 12102 15792 12406
rect 16028 12164 16080 12170
rect 16028 12106 16080 12112
rect 16120 12164 16172 12170
rect 16120 12106 16172 12112
rect 15752 12096 15804 12102
rect 15752 12038 15804 12044
rect 15660 11688 15712 11694
rect 15660 11630 15712 11636
rect 15568 11552 15620 11558
rect 15568 11494 15620 11500
rect 15580 11286 15608 11494
rect 15568 11280 15620 11286
rect 15568 11222 15620 11228
rect 15764 11218 15792 12038
rect 15936 11552 15988 11558
rect 15936 11494 15988 11500
rect 15948 11218 15976 11494
rect 16040 11354 16068 12106
rect 16028 11348 16080 11354
rect 16028 11290 16080 11296
rect 16132 11234 16160 12106
rect 15752 11212 15804 11218
rect 15752 11154 15804 11160
rect 15936 11212 15988 11218
rect 15936 11154 15988 11160
rect 16040 11206 16160 11234
rect 15660 11008 15712 11014
rect 15566 10976 15622 10985
rect 15660 10950 15712 10956
rect 15752 11008 15804 11014
rect 15752 10950 15804 10956
rect 15566 10911 15622 10920
rect 15580 10742 15608 10911
rect 15476 10736 15528 10742
rect 15476 10678 15528 10684
rect 15568 10736 15620 10742
rect 15568 10678 15620 10684
rect 14924 10668 14976 10674
rect 14924 10610 14976 10616
rect 15384 10668 15436 10674
rect 15384 10610 15436 10616
rect 15016 10600 15068 10606
rect 15016 10542 15068 10548
rect 14740 10056 14792 10062
rect 14740 9998 14792 10004
rect 14648 9920 14700 9926
rect 14648 9862 14700 9868
rect 14372 9580 14424 9586
rect 14372 9522 14424 9528
rect 14648 9580 14700 9586
rect 14648 9522 14700 9528
rect 14660 9382 14688 9522
rect 14096 9376 14148 9382
rect 14096 9318 14148 9324
rect 14648 9376 14700 9382
rect 14648 9318 14700 9324
rect 14108 9178 14136 9318
rect 14096 9172 14148 9178
rect 14096 9114 14148 9120
rect 13728 8900 13780 8906
rect 13728 8842 13780 8848
rect 14108 8430 14136 9114
rect 14372 8968 14424 8974
rect 14372 8910 14424 8916
rect 14096 8424 14148 8430
rect 14096 8366 14148 8372
rect 13636 8356 13688 8362
rect 13636 8298 13688 8304
rect 13648 8090 13676 8298
rect 13636 8084 13688 8090
rect 13636 8026 13688 8032
rect 14108 8022 14136 8366
rect 14096 8016 14148 8022
rect 14096 7958 14148 7964
rect 14384 7954 14412 8910
rect 14556 8832 14608 8838
rect 14556 8774 14608 8780
rect 14372 7948 14424 7954
rect 14372 7890 14424 7896
rect 13176 7880 13228 7886
rect 13176 7822 13228 7828
rect 13544 7880 13596 7886
rect 13544 7822 13596 7828
rect 14464 7880 14516 7886
rect 14464 7822 14516 7828
rect 12900 7404 12952 7410
rect 12900 7346 12952 7352
rect 13176 7404 13228 7410
rect 13176 7346 13228 7352
rect 12898 7304 12954 7313
rect 12898 7239 12954 7248
rect 12912 7206 12940 7239
rect 12900 7200 12952 7206
rect 12900 7142 12952 7148
rect 12808 6996 12860 7002
rect 12808 6938 12860 6944
rect 13084 6928 13136 6934
rect 13084 6870 13136 6876
rect 12808 6860 12860 6866
rect 12808 6802 12860 6808
rect 12716 6248 12768 6254
rect 12622 6216 12678 6225
rect 12716 6190 12768 6196
rect 12622 6151 12624 6160
rect 12676 6151 12678 6160
rect 12624 6122 12676 6128
rect 12820 6118 12848 6802
rect 12912 6458 13032 6474
rect 12912 6452 13044 6458
rect 12912 6446 12992 6452
rect 12256 6112 12308 6118
rect 12256 6054 12308 6060
rect 12808 6112 12860 6118
rect 12808 6054 12860 6060
rect 12268 5930 12296 6054
rect 12072 5908 12124 5914
rect 12268 5902 12388 5930
rect 12072 5850 12124 5856
rect 12254 5808 12310 5817
rect 12254 5743 12310 5752
rect 11612 5636 11664 5642
rect 11992 5630 12204 5658
rect 12268 5642 12296 5743
rect 12360 5710 12388 5902
rect 12348 5704 12400 5710
rect 12348 5646 12400 5652
rect 11612 5578 11664 5584
rect 11624 5370 11652 5578
rect 11980 5568 12032 5574
rect 11980 5510 12032 5516
rect 11612 5364 11664 5370
rect 11612 5306 11664 5312
rect 11704 4616 11756 4622
rect 11704 4558 11756 4564
rect 11716 4146 11744 4558
rect 11992 4486 12020 5510
rect 12072 5160 12124 5166
rect 12072 5102 12124 5108
rect 12084 4554 12112 5102
rect 12072 4548 12124 4554
rect 12072 4490 12124 4496
rect 11980 4480 12032 4486
rect 11980 4422 12032 4428
rect 12084 4282 12112 4490
rect 12072 4276 12124 4282
rect 12176 4264 12204 5630
rect 12256 5636 12308 5642
rect 12256 5578 12308 5584
rect 12311 5468 12619 5477
rect 12311 5466 12317 5468
rect 12373 5466 12397 5468
rect 12453 5466 12477 5468
rect 12533 5466 12557 5468
rect 12613 5466 12619 5468
rect 12373 5414 12375 5466
rect 12555 5414 12557 5466
rect 12311 5412 12317 5414
rect 12373 5412 12397 5414
rect 12453 5412 12477 5414
rect 12533 5412 12557 5414
rect 12613 5412 12619 5414
rect 12311 5403 12619 5412
rect 12532 5364 12584 5370
rect 12532 5306 12584 5312
rect 12544 4758 12572 5306
rect 12912 4826 12940 6446
rect 12992 6394 13044 6400
rect 12992 6316 13044 6322
rect 12992 6258 13044 6264
rect 13004 5642 13032 6258
rect 13096 5658 13124 6870
rect 13188 6458 13216 7346
rect 13556 6934 13584 7822
rect 14476 7750 14504 7822
rect 14464 7744 14516 7750
rect 14464 7686 14516 7692
rect 13820 7200 13872 7206
rect 13820 7142 13872 7148
rect 13544 6928 13596 6934
rect 13544 6870 13596 6876
rect 13634 6760 13690 6769
rect 13634 6695 13690 6704
rect 13176 6452 13228 6458
rect 13176 6394 13228 6400
rect 12992 5636 13044 5642
rect 13096 5630 13216 5658
rect 12992 5578 13044 5584
rect 13084 5568 13136 5574
rect 13084 5510 13136 5516
rect 13096 4826 13124 5510
rect 13188 5370 13216 5630
rect 13176 5364 13228 5370
rect 13176 5306 13228 5312
rect 13360 5228 13412 5234
rect 13360 5170 13412 5176
rect 12900 4820 12952 4826
rect 12900 4762 12952 4768
rect 13084 4820 13136 4826
rect 13084 4762 13136 4768
rect 12532 4752 12584 4758
rect 12532 4694 12584 4700
rect 12544 4622 12572 4694
rect 13372 4622 13400 5170
rect 13452 4684 13504 4690
rect 13452 4626 13504 4632
rect 12532 4616 12584 4622
rect 13360 4616 13412 4622
rect 12532 4558 12584 4564
rect 13280 4576 13360 4604
rect 12808 4548 12860 4554
rect 12808 4490 12860 4496
rect 12311 4380 12619 4389
rect 12311 4378 12317 4380
rect 12373 4378 12397 4380
rect 12453 4378 12477 4380
rect 12533 4378 12557 4380
rect 12613 4378 12619 4380
rect 12373 4326 12375 4378
rect 12555 4326 12557 4378
rect 12311 4324 12317 4326
rect 12373 4324 12397 4326
rect 12453 4324 12477 4326
rect 12533 4324 12557 4326
rect 12613 4324 12619 4326
rect 12311 4315 12619 4324
rect 12176 4236 12296 4264
rect 12072 4218 12124 4224
rect 11704 4140 11756 4146
rect 11704 4082 11756 4088
rect 12072 4072 12124 4078
rect 11702 4040 11758 4049
rect 12072 4014 12124 4020
rect 11702 3975 11758 3984
rect 11716 3534 11744 3975
rect 12084 3602 12112 4014
rect 12164 4004 12216 4010
rect 12164 3946 12216 3952
rect 12072 3596 12124 3602
rect 12072 3538 12124 3544
rect 11704 3528 11756 3534
rect 11704 3470 11756 3476
rect 11244 3188 11296 3194
rect 11244 3130 11296 3136
rect 11428 3188 11480 3194
rect 11428 3130 11480 3136
rect 11440 2990 11468 3130
rect 12084 2990 12112 3538
rect 12176 3058 12204 3946
rect 12268 3602 12296 4236
rect 12820 3942 12848 4490
rect 12808 3936 12860 3942
rect 12808 3878 12860 3884
rect 12256 3596 12308 3602
rect 12256 3538 12308 3544
rect 12268 3398 12296 3538
rect 12256 3392 12308 3398
rect 12256 3334 12308 3340
rect 12311 3292 12619 3301
rect 12311 3290 12317 3292
rect 12373 3290 12397 3292
rect 12453 3290 12477 3292
rect 12533 3290 12557 3292
rect 12613 3290 12619 3292
rect 12373 3238 12375 3290
rect 12555 3238 12557 3290
rect 12311 3236 12317 3238
rect 12373 3236 12397 3238
rect 12453 3236 12477 3238
rect 12533 3236 12557 3238
rect 12613 3236 12619 3238
rect 12311 3227 12619 3236
rect 12348 3188 12400 3194
rect 12348 3130 12400 3136
rect 12164 3052 12216 3058
rect 12164 2994 12216 3000
rect 11428 2984 11480 2990
rect 11242 2952 11298 2961
rect 11164 2910 11242 2938
rect 11428 2926 11480 2932
rect 12072 2984 12124 2990
rect 12072 2926 12124 2932
rect 11058 2887 11114 2896
rect 11242 2887 11244 2896
rect 11296 2887 11298 2896
rect 11244 2858 11296 2864
rect 10416 2848 10468 2854
rect 10416 2790 10468 2796
rect 9471 2748 9779 2757
rect 9471 2746 9477 2748
rect 9533 2746 9557 2748
rect 9613 2746 9637 2748
rect 9693 2746 9717 2748
rect 9773 2746 9779 2748
rect 9533 2694 9535 2746
rect 9715 2694 9717 2746
rect 9471 2692 9477 2694
rect 9533 2692 9557 2694
rect 9613 2692 9637 2694
rect 9693 2692 9717 2694
rect 9773 2692 9779 2694
rect 9471 2683 9779 2692
rect 12360 2650 12388 3130
rect 13280 3058 13308 4576
rect 13360 4558 13412 4564
rect 13360 3732 13412 3738
rect 13360 3674 13412 3680
rect 13372 3466 13400 3674
rect 13464 3534 13492 4626
rect 13544 4548 13596 4554
rect 13544 4490 13596 4496
rect 13556 3738 13584 4490
rect 13648 3942 13676 6695
rect 13832 6118 13860 7142
rect 14476 6798 14504 7686
rect 14464 6792 14516 6798
rect 14464 6734 14516 6740
rect 14188 6724 14240 6730
rect 14188 6666 14240 6672
rect 14096 6656 14148 6662
rect 14096 6598 14148 6604
rect 13912 6316 13964 6322
rect 13912 6258 13964 6264
rect 13820 6112 13872 6118
rect 13820 6054 13872 6060
rect 13728 5092 13780 5098
rect 13728 5034 13780 5040
rect 13740 4622 13768 5034
rect 13728 4616 13780 4622
rect 13728 4558 13780 4564
rect 13832 4214 13860 6054
rect 13924 5778 13952 6258
rect 14108 6254 14136 6598
rect 14200 6322 14228 6666
rect 14188 6316 14240 6322
rect 14188 6258 14240 6264
rect 14096 6248 14148 6254
rect 14096 6190 14148 6196
rect 13912 5772 13964 5778
rect 13912 5714 13964 5720
rect 14108 5302 14136 6190
rect 14200 5642 14228 6258
rect 14464 5840 14516 5846
rect 14464 5782 14516 5788
rect 14188 5636 14240 5642
rect 14188 5578 14240 5584
rect 14372 5364 14424 5370
rect 14372 5306 14424 5312
rect 14096 5296 14148 5302
rect 14096 5238 14148 5244
rect 14278 5264 14334 5273
rect 13820 4208 13872 4214
rect 13820 4150 13872 4156
rect 14108 4146 14136 5238
rect 14278 5199 14280 5208
rect 14332 5199 14334 5208
rect 14280 5170 14332 5176
rect 14384 4622 14412 5306
rect 14476 5030 14504 5782
rect 14568 5137 14596 8774
rect 14660 8430 14688 9318
rect 14752 8537 14780 9998
rect 15028 9994 15056 10542
rect 15152 10364 15460 10373
rect 15152 10362 15158 10364
rect 15214 10362 15238 10364
rect 15294 10362 15318 10364
rect 15374 10362 15398 10364
rect 15454 10362 15460 10364
rect 15214 10310 15216 10362
rect 15396 10310 15398 10362
rect 15152 10308 15158 10310
rect 15214 10308 15238 10310
rect 15294 10308 15318 10310
rect 15374 10308 15398 10310
rect 15454 10308 15460 10310
rect 15152 10299 15460 10308
rect 15016 9988 15068 9994
rect 15016 9930 15068 9936
rect 15488 9722 15516 10678
rect 15672 10198 15700 10950
rect 15764 10810 15792 10950
rect 15752 10804 15804 10810
rect 15752 10746 15804 10752
rect 15764 10266 15792 10746
rect 15752 10260 15804 10266
rect 15752 10202 15804 10208
rect 15660 10192 15712 10198
rect 15660 10134 15712 10140
rect 16040 10062 16068 11206
rect 16120 11144 16172 11150
rect 16120 11086 16172 11092
rect 16028 10056 16080 10062
rect 16028 9998 16080 10004
rect 15568 9920 15620 9926
rect 15568 9862 15620 9868
rect 15580 9722 15608 9862
rect 15476 9716 15528 9722
rect 15476 9658 15528 9664
rect 15568 9716 15620 9722
rect 15568 9658 15620 9664
rect 15844 9512 15896 9518
rect 15844 9454 15896 9460
rect 15752 9444 15804 9450
rect 15752 9386 15804 9392
rect 15660 9376 15712 9382
rect 15660 9318 15712 9324
rect 15152 9276 15460 9285
rect 15152 9274 15158 9276
rect 15214 9274 15238 9276
rect 15294 9274 15318 9276
rect 15374 9274 15398 9276
rect 15454 9274 15460 9276
rect 15214 9222 15216 9274
rect 15396 9222 15398 9274
rect 15152 9220 15158 9222
rect 15214 9220 15238 9222
rect 15294 9220 15318 9222
rect 15374 9220 15398 9222
rect 15454 9220 15460 9222
rect 15152 9211 15460 9220
rect 15672 8906 15700 9318
rect 15660 8900 15712 8906
rect 15660 8842 15712 8848
rect 15384 8832 15436 8838
rect 15384 8774 15436 8780
rect 14738 8528 14794 8537
rect 14738 8463 14794 8472
rect 14648 8424 14700 8430
rect 14648 8366 14700 8372
rect 14660 7206 14688 8366
rect 15396 8294 15424 8774
rect 15016 8288 15068 8294
rect 15016 8230 15068 8236
rect 15384 8288 15436 8294
rect 15384 8230 15436 8236
rect 14830 7984 14886 7993
rect 14830 7919 14886 7928
rect 14844 7886 14872 7919
rect 14832 7880 14884 7886
rect 14832 7822 14884 7828
rect 14740 7744 14792 7750
rect 14740 7686 14792 7692
rect 14752 7478 14780 7686
rect 14740 7472 14792 7478
rect 14740 7414 14792 7420
rect 14648 7200 14700 7206
rect 14648 7142 14700 7148
rect 14844 6866 14872 7822
rect 15028 7410 15056 8230
rect 15152 8188 15460 8197
rect 15152 8186 15158 8188
rect 15214 8186 15238 8188
rect 15294 8186 15318 8188
rect 15374 8186 15398 8188
rect 15454 8186 15460 8188
rect 15214 8134 15216 8186
rect 15396 8134 15398 8186
rect 15152 8132 15158 8134
rect 15214 8132 15238 8134
rect 15294 8132 15318 8134
rect 15374 8132 15398 8134
rect 15454 8132 15460 8134
rect 15152 8123 15460 8132
rect 15476 7540 15528 7546
rect 15476 7482 15528 7488
rect 15016 7404 15068 7410
rect 15016 7346 15068 7352
rect 14924 7336 14976 7342
rect 14924 7278 14976 7284
rect 14832 6860 14884 6866
rect 14832 6802 14884 6808
rect 14740 6180 14792 6186
rect 14740 6122 14792 6128
rect 14752 5846 14780 6122
rect 14830 5944 14886 5953
rect 14830 5879 14886 5888
rect 14740 5840 14792 5846
rect 14740 5782 14792 5788
rect 14844 5710 14872 5879
rect 14832 5704 14884 5710
rect 14832 5646 14884 5652
rect 14648 5636 14700 5642
rect 14648 5578 14700 5584
rect 14660 5302 14688 5578
rect 14648 5296 14700 5302
rect 14648 5238 14700 5244
rect 14832 5296 14884 5302
rect 14832 5238 14884 5244
rect 14844 5137 14872 5238
rect 14554 5128 14610 5137
rect 14554 5063 14610 5072
rect 14830 5128 14886 5137
rect 14830 5063 14886 5072
rect 14464 5024 14516 5030
rect 14464 4966 14516 4972
rect 14372 4616 14424 4622
rect 14372 4558 14424 4564
rect 14384 4282 14412 4558
rect 14372 4276 14424 4282
rect 14372 4218 14424 4224
rect 14096 4140 14148 4146
rect 14096 4082 14148 4088
rect 13636 3936 13688 3942
rect 13636 3878 13688 3884
rect 13544 3732 13596 3738
rect 13544 3674 13596 3680
rect 13452 3528 13504 3534
rect 13452 3470 13504 3476
rect 13544 3528 13596 3534
rect 13544 3470 13596 3476
rect 13360 3460 13412 3466
rect 13360 3402 13412 3408
rect 13464 3398 13492 3470
rect 13452 3392 13504 3398
rect 13452 3334 13504 3340
rect 13556 3194 13584 3470
rect 13648 3369 13676 3878
rect 13634 3360 13690 3369
rect 13634 3295 13690 3304
rect 13648 3194 13676 3295
rect 13544 3188 13596 3194
rect 13544 3130 13596 3136
rect 13636 3188 13688 3194
rect 13636 3130 13688 3136
rect 13268 3052 13320 3058
rect 13268 2994 13320 3000
rect 14476 2650 14504 4966
rect 14568 4282 14596 5063
rect 14556 4276 14608 4282
rect 14556 4218 14608 4224
rect 14568 3738 14596 4218
rect 14936 4078 14964 7278
rect 15028 6390 15056 7346
rect 15152 7100 15460 7109
rect 15152 7098 15158 7100
rect 15214 7098 15238 7100
rect 15294 7098 15318 7100
rect 15374 7098 15398 7100
rect 15454 7098 15460 7100
rect 15214 7046 15216 7098
rect 15396 7046 15398 7098
rect 15152 7044 15158 7046
rect 15214 7044 15238 7046
rect 15294 7044 15318 7046
rect 15374 7044 15398 7046
rect 15454 7044 15460 7046
rect 15152 7035 15460 7044
rect 15016 6384 15068 6390
rect 15016 6326 15068 6332
rect 15016 6248 15068 6254
rect 15016 6190 15068 6196
rect 15028 5794 15056 6190
rect 15488 6186 15516 7482
rect 15672 7206 15700 8842
rect 15764 8838 15792 9386
rect 15856 9042 15884 9454
rect 16132 9382 16160 11086
rect 16224 10810 16252 12736
rect 16316 12442 16344 13126
rect 16304 12436 16356 12442
rect 16304 12378 16356 12384
rect 16212 10804 16264 10810
rect 16212 10746 16264 10752
rect 16408 10742 16436 14486
rect 16500 11014 16528 15014
rect 16948 15020 17000 15026
rect 16948 14962 17000 14968
rect 16580 14952 16632 14958
rect 16580 14894 16632 14900
rect 16592 13258 16620 14894
rect 16764 14408 16816 14414
rect 16764 14350 16816 14356
rect 16776 13258 16804 14350
rect 16960 14074 16988 14962
rect 16948 14068 17000 14074
rect 16948 14010 17000 14016
rect 16960 13938 16988 14010
rect 16948 13932 17000 13938
rect 16948 13874 17000 13880
rect 16948 13388 17000 13394
rect 16948 13330 17000 13336
rect 16856 13320 16908 13326
rect 16856 13262 16908 13268
rect 16580 13252 16632 13258
rect 16580 13194 16632 13200
rect 16764 13252 16816 13258
rect 16764 13194 16816 13200
rect 16672 12708 16724 12714
rect 16672 12650 16724 12656
rect 16488 11008 16540 11014
rect 16488 10950 16540 10956
rect 16396 10736 16448 10742
rect 16396 10678 16448 10684
rect 16408 10130 16436 10678
rect 16684 10538 16712 12650
rect 16672 10532 16724 10538
rect 16672 10474 16724 10480
rect 16488 10464 16540 10470
rect 16488 10406 16540 10412
rect 16396 10124 16448 10130
rect 16396 10066 16448 10072
rect 16500 9654 16528 10406
rect 16684 9994 16712 10474
rect 16776 10062 16804 13194
rect 16868 12646 16896 13262
rect 16960 13161 16988 13330
rect 16946 13152 17002 13161
rect 16946 13087 17002 13096
rect 16948 12844 17000 12850
rect 17052 12832 17080 15914
rect 17132 15904 17184 15910
rect 17132 15846 17184 15852
rect 17144 14482 17172 15846
rect 17132 14476 17184 14482
rect 17132 14418 17184 14424
rect 17236 14362 17264 18362
rect 17316 18080 17368 18086
rect 17316 18022 17368 18028
rect 17328 17610 17356 18022
rect 17512 17762 17540 20012
rect 17684 19916 17736 19922
rect 17684 19858 17736 19864
rect 17420 17734 17540 17762
rect 17316 17604 17368 17610
rect 17316 17546 17368 17552
rect 17316 17264 17368 17270
rect 17316 17206 17368 17212
rect 17328 16794 17356 17206
rect 17316 16788 17368 16794
rect 17316 16730 17368 16736
rect 17328 14958 17356 16730
rect 17420 16658 17448 17734
rect 17500 17672 17552 17678
rect 17500 17614 17552 17620
rect 17408 16652 17460 16658
rect 17408 16594 17460 16600
rect 17408 16516 17460 16522
rect 17408 16458 17460 16464
rect 17420 15434 17448 16458
rect 17408 15428 17460 15434
rect 17408 15370 17460 15376
rect 17316 14952 17368 14958
rect 17316 14894 17368 14900
rect 17408 14612 17460 14618
rect 17408 14554 17460 14560
rect 17420 14414 17448 14554
rect 17144 14334 17264 14362
rect 17316 14408 17368 14414
rect 17316 14350 17368 14356
rect 17408 14408 17460 14414
rect 17408 14350 17460 14356
rect 17144 13297 17172 14334
rect 17224 14272 17276 14278
rect 17224 14214 17276 14220
rect 17236 13977 17264 14214
rect 17222 13968 17278 13977
rect 17222 13903 17278 13912
rect 17328 13530 17356 14350
rect 17408 14068 17460 14074
rect 17408 14010 17460 14016
rect 17316 13524 17368 13530
rect 17316 13466 17368 13472
rect 17314 13424 17370 13433
rect 17314 13359 17370 13368
rect 17130 13288 17186 13297
rect 17130 13223 17186 13232
rect 17144 12850 17172 13223
rect 17224 12912 17276 12918
rect 17224 12854 17276 12860
rect 17000 12804 17080 12832
rect 17132 12844 17184 12850
rect 16948 12786 17000 12792
rect 17132 12786 17184 12792
rect 16856 12640 16908 12646
rect 16856 12582 16908 12588
rect 16868 12238 16896 12582
rect 16856 12232 16908 12238
rect 16856 12174 16908 12180
rect 16960 12170 16988 12786
rect 16948 12164 17000 12170
rect 16948 12106 17000 12112
rect 16960 11286 16988 12106
rect 16856 11280 16908 11286
rect 16856 11222 16908 11228
rect 16948 11280 17000 11286
rect 16948 11222 17000 11228
rect 16868 11150 16896 11222
rect 16856 11144 16908 11150
rect 16856 11086 16908 11092
rect 17144 10742 17172 12786
rect 17236 12209 17264 12854
rect 17222 12200 17278 12209
rect 17222 12135 17278 12144
rect 17132 10736 17184 10742
rect 17132 10678 17184 10684
rect 16764 10056 16816 10062
rect 16764 9998 16816 10004
rect 16672 9988 16724 9994
rect 16672 9930 16724 9936
rect 16948 9988 17000 9994
rect 16948 9930 17000 9936
rect 16488 9648 16540 9654
rect 16488 9590 16540 9596
rect 16684 9586 16712 9930
rect 16672 9580 16724 9586
rect 16672 9522 16724 9528
rect 16764 9580 16816 9586
rect 16764 9522 16816 9528
rect 16120 9376 16172 9382
rect 16120 9318 16172 9324
rect 16580 9376 16632 9382
rect 16580 9318 16632 9324
rect 16304 9104 16356 9110
rect 16304 9046 16356 9052
rect 15844 9036 15896 9042
rect 15844 8978 15896 8984
rect 15752 8832 15804 8838
rect 15752 8774 15804 8780
rect 15856 8566 15884 8978
rect 15844 8560 15896 8566
rect 16028 8560 16080 8566
rect 15844 8502 15896 8508
rect 15948 8508 16028 8514
rect 15948 8502 16080 8508
rect 15856 7546 15884 8502
rect 15948 8486 16068 8502
rect 15844 7540 15896 7546
rect 15844 7482 15896 7488
rect 15752 7404 15804 7410
rect 15752 7346 15804 7352
rect 15660 7200 15712 7206
rect 15660 7142 15712 7148
rect 15764 6934 15792 7346
rect 15752 6928 15804 6934
rect 15752 6870 15804 6876
rect 15476 6180 15528 6186
rect 15476 6122 15528 6128
rect 15152 6012 15460 6021
rect 15152 6010 15158 6012
rect 15214 6010 15238 6012
rect 15294 6010 15318 6012
rect 15374 6010 15398 6012
rect 15454 6010 15460 6012
rect 15214 5958 15216 6010
rect 15396 5958 15398 6010
rect 15152 5956 15158 5958
rect 15214 5956 15238 5958
rect 15294 5956 15318 5958
rect 15374 5956 15398 5958
rect 15454 5956 15460 5958
rect 15152 5947 15460 5956
rect 15488 5846 15516 6122
rect 15476 5840 15528 5846
rect 15028 5766 15332 5794
rect 15476 5782 15528 5788
rect 15304 5642 15332 5766
rect 15764 5710 15792 6870
rect 15948 6730 15976 8486
rect 16316 7954 16344 9046
rect 16592 9042 16620 9318
rect 16580 9036 16632 9042
rect 16580 8978 16632 8984
rect 16592 8566 16620 8978
rect 16580 8560 16632 8566
rect 16580 8502 16632 8508
rect 16304 7948 16356 7954
rect 16304 7890 16356 7896
rect 16592 7886 16620 8502
rect 16580 7880 16632 7886
rect 16580 7822 16632 7828
rect 16396 7404 16448 7410
rect 16396 7346 16448 7352
rect 16028 7200 16080 7206
rect 16028 7142 16080 7148
rect 15936 6724 15988 6730
rect 15936 6666 15988 6672
rect 15948 5778 15976 6666
rect 16040 6458 16068 7142
rect 16408 7002 16436 7346
rect 16396 6996 16448 7002
rect 16396 6938 16448 6944
rect 16028 6452 16080 6458
rect 16028 6394 16080 6400
rect 16592 6390 16620 7822
rect 16684 6866 16712 9522
rect 16776 8906 16804 9522
rect 16856 9444 16908 9450
rect 16856 9386 16908 9392
rect 16868 9110 16896 9386
rect 16856 9104 16908 9110
rect 16856 9046 16908 9052
rect 16764 8900 16816 8906
rect 16764 8842 16816 8848
rect 16776 7818 16804 8842
rect 16868 8634 16896 9046
rect 16960 9042 16988 9930
rect 17236 9926 17264 12135
rect 17328 11694 17356 13359
rect 17420 12753 17448 14010
rect 17406 12744 17462 12753
rect 17406 12679 17462 12688
rect 17408 12096 17460 12102
rect 17408 12038 17460 12044
rect 17420 11762 17448 12038
rect 17512 11898 17540 17614
rect 17592 17536 17644 17542
rect 17592 17478 17644 17484
rect 17604 16998 17632 17478
rect 17592 16992 17644 16998
rect 17592 16934 17644 16940
rect 17604 16046 17632 16934
rect 17592 16040 17644 16046
rect 17592 15982 17644 15988
rect 17604 13326 17632 15982
rect 17696 13802 17724 19858
rect 17868 19712 17920 19718
rect 17868 19654 17920 19660
rect 17776 18692 17828 18698
rect 17776 18634 17828 18640
rect 17788 17746 17816 18634
rect 17776 17740 17828 17746
rect 17776 17682 17828 17688
rect 17880 17678 17908 19654
rect 17992 19612 18300 19621
rect 17992 19610 17998 19612
rect 18054 19610 18078 19612
rect 18134 19610 18158 19612
rect 18214 19610 18238 19612
rect 18294 19610 18300 19612
rect 18054 19558 18056 19610
rect 18236 19558 18238 19610
rect 17992 19556 17998 19558
rect 18054 19556 18078 19558
rect 18134 19556 18158 19558
rect 18214 19556 18238 19558
rect 18294 19556 18300 19558
rect 17992 19547 18300 19556
rect 18340 18970 18368 20878
rect 18604 20460 18656 20466
rect 18604 20402 18656 20408
rect 18972 20460 19024 20466
rect 18972 20402 19024 20408
rect 18512 19372 18564 19378
rect 18512 19314 18564 19320
rect 18328 18964 18380 18970
rect 18328 18906 18380 18912
rect 18524 18766 18552 19314
rect 18512 18760 18564 18766
rect 18512 18702 18564 18708
rect 17992 18524 18300 18533
rect 17992 18522 17998 18524
rect 18054 18522 18078 18524
rect 18134 18522 18158 18524
rect 18214 18522 18238 18524
rect 18294 18522 18300 18524
rect 18054 18470 18056 18522
rect 18236 18470 18238 18522
rect 17992 18468 17998 18470
rect 18054 18468 18078 18470
rect 18134 18468 18158 18470
rect 18214 18468 18238 18470
rect 18294 18468 18300 18470
rect 17992 18459 18300 18468
rect 18420 18216 18472 18222
rect 18420 18158 18472 18164
rect 17868 17672 17920 17678
rect 17868 17614 17920 17620
rect 18328 17672 18380 17678
rect 18328 17614 18380 17620
rect 17992 17436 18300 17445
rect 17992 17434 17998 17436
rect 18054 17434 18078 17436
rect 18134 17434 18158 17436
rect 18214 17434 18238 17436
rect 18294 17434 18300 17436
rect 18054 17382 18056 17434
rect 18236 17382 18238 17434
rect 17992 17380 17998 17382
rect 18054 17380 18078 17382
rect 18134 17380 18158 17382
rect 18214 17380 18238 17382
rect 18294 17380 18300 17382
rect 17992 17371 18300 17380
rect 17868 17060 17920 17066
rect 17868 17002 17920 17008
rect 17776 16992 17828 16998
rect 17776 16934 17828 16940
rect 17788 16658 17816 16934
rect 17776 16652 17828 16658
rect 17776 16594 17828 16600
rect 17774 16552 17830 16561
rect 17774 16487 17830 16496
rect 17788 15978 17816 16487
rect 17880 16454 17908 17002
rect 18052 16992 18104 16998
rect 18052 16934 18104 16940
rect 18064 16561 18092 16934
rect 18340 16658 18368 17614
rect 18432 17202 18460 18158
rect 18524 17882 18552 18702
rect 18512 17876 18564 17882
rect 18512 17818 18564 17824
rect 18420 17196 18472 17202
rect 18420 17138 18472 17144
rect 18328 16652 18380 16658
rect 18328 16594 18380 16600
rect 18050 16552 18106 16561
rect 18050 16487 18106 16496
rect 18328 16516 18380 16522
rect 18328 16458 18380 16464
rect 17868 16448 17920 16454
rect 17868 16390 17920 16396
rect 17992 16348 18300 16357
rect 17992 16346 17998 16348
rect 18054 16346 18078 16348
rect 18134 16346 18158 16348
rect 18214 16346 18238 16348
rect 18294 16346 18300 16348
rect 18054 16294 18056 16346
rect 18236 16294 18238 16346
rect 17992 16292 17998 16294
rect 18054 16292 18078 16294
rect 18134 16292 18158 16294
rect 18214 16292 18238 16294
rect 18294 16292 18300 16294
rect 17992 16283 18300 16292
rect 18340 16250 18368 16458
rect 18328 16244 18380 16250
rect 18328 16186 18380 16192
rect 18432 16153 18460 17138
rect 18512 16788 18564 16794
rect 18512 16730 18564 16736
rect 18524 16658 18552 16730
rect 18512 16652 18564 16658
rect 18512 16594 18564 16600
rect 18418 16144 18474 16153
rect 18418 16079 18420 16088
rect 18472 16079 18474 16088
rect 18420 16050 18472 16056
rect 18432 16019 18460 16050
rect 18510 16008 18566 16017
rect 17776 15972 17828 15978
rect 18510 15943 18566 15952
rect 17776 15914 17828 15920
rect 17992 15260 18300 15269
rect 17992 15258 17998 15260
rect 18054 15258 18078 15260
rect 18134 15258 18158 15260
rect 18214 15258 18238 15260
rect 18294 15258 18300 15260
rect 18054 15206 18056 15258
rect 18236 15206 18238 15258
rect 17992 15204 17998 15206
rect 18054 15204 18078 15206
rect 18134 15204 18158 15206
rect 18214 15204 18238 15206
rect 18294 15204 18300 15206
rect 17992 15195 18300 15204
rect 18524 15094 18552 15943
rect 18512 15088 18564 15094
rect 18512 15030 18564 15036
rect 18328 14952 18380 14958
rect 18328 14894 18380 14900
rect 17992 14172 18300 14181
rect 17992 14170 17998 14172
rect 18054 14170 18078 14172
rect 18134 14170 18158 14172
rect 18214 14170 18238 14172
rect 18294 14170 18300 14172
rect 18054 14118 18056 14170
rect 18236 14118 18238 14170
rect 17992 14116 17998 14118
rect 18054 14116 18078 14118
rect 18134 14116 18158 14118
rect 18214 14116 18238 14118
rect 18294 14116 18300 14118
rect 17992 14107 18300 14116
rect 18234 13968 18290 13977
rect 17960 13932 18012 13938
rect 18234 13903 18236 13912
rect 17960 13874 18012 13880
rect 18288 13903 18290 13912
rect 18236 13874 18288 13880
rect 17684 13796 17736 13802
rect 17684 13738 17736 13744
rect 17972 13394 18000 13874
rect 17960 13388 18012 13394
rect 17880 13348 17960 13376
rect 17592 13320 17644 13326
rect 17592 13262 17644 13268
rect 17776 13184 17828 13190
rect 17682 13152 17738 13161
rect 17776 13126 17828 13132
rect 17682 13087 17738 13096
rect 17590 13016 17646 13025
rect 17696 12986 17724 13087
rect 17590 12951 17646 12960
rect 17684 12980 17736 12986
rect 17604 12918 17632 12951
rect 17684 12922 17736 12928
rect 17592 12912 17644 12918
rect 17592 12854 17644 12860
rect 17592 12640 17644 12646
rect 17592 12582 17644 12588
rect 17500 11892 17552 11898
rect 17500 11834 17552 11840
rect 17604 11762 17632 12582
rect 17684 12232 17736 12238
rect 17684 12174 17736 12180
rect 17408 11756 17460 11762
rect 17408 11698 17460 11704
rect 17592 11756 17644 11762
rect 17592 11698 17644 11704
rect 17316 11688 17368 11694
rect 17316 11630 17368 11636
rect 17592 10804 17644 10810
rect 17592 10746 17644 10752
rect 17604 10606 17632 10746
rect 17592 10600 17644 10606
rect 17592 10542 17644 10548
rect 17408 10464 17460 10470
rect 17408 10406 17460 10412
rect 17420 10062 17448 10406
rect 17696 10266 17724 12174
rect 17788 11762 17816 13126
rect 17880 12850 17908 13348
rect 17960 13330 18012 13336
rect 17992 13084 18300 13093
rect 17992 13082 17998 13084
rect 18054 13082 18078 13084
rect 18134 13082 18158 13084
rect 18214 13082 18238 13084
rect 18294 13082 18300 13084
rect 18054 13030 18056 13082
rect 18236 13030 18238 13082
rect 17992 13028 17998 13030
rect 18054 13028 18078 13030
rect 18134 13028 18158 13030
rect 18214 13028 18238 13030
rect 18294 13028 18300 13030
rect 17992 13019 18300 13028
rect 17868 12844 17920 12850
rect 17868 12786 17920 12792
rect 17866 12744 17922 12753
rect 17866 12679 17922 12688
rect 17880 12238 17908 12679
rect 17960 12300 18012 12306
rect 17960 12242 18012 12248
rect 17868 12232 17920 12238
rect 17868 12174 17920 12180
rect 17972 12084 18000 12242
rect 17880 12056 18000 12084
rect 17776 11756 17828 11762
rect 17776 11698 17828 11704
rect 17776 11144 17828 11150
rect 17776 11086 17828 11092
rect 17684 10260 17736 10266
rect 17684 10202 17736 10208
rect 17408 10056 17460 10062
rect 17500 10056 17552 10062
rect 17408 9998 17460 10004
rect 17498 10024 17500 10033
rect 17552 10024 17554 10033
rect 17498 9959 17554 9968
rect 17224 9920 17276 9926
rect 17224 9862 17276 9868
rect 17592 9920 17644 9926
rect 17592 9862 17644 9868
rect 17132 9648 17184 9654
rect 17132 9590 17184 9596
rect 17040 9172 17092 9178
rect 17144 9160 17172 9590
rect 17604 9586 17632 9862
rect 17592 9580 17644 9586
rect 17592 9522 17644 9528
rect 17592 9376 17644 9382
rect 17592 9318 17644 9324
rect 17092 9132 17172 9160
rect 17040 9114 17092 9120
rect 16948 9036 17000 9042
rect 16948 8978 17000 8984
rect 16856 8628 16908 8634
rect 16856 8570 16908 8576
rect 16764 7812 16816 7818
rect 16764 7754 16816 7760
rect 16776 7274 16804 7754
rect 16960 7410 16988 8978
rect 17052 7410 17080 9114
rect 17500 8832 17552 8838
rect 17500 8774 17552 8780
rect 17316 8628 17368 8634
rect 17316 8570 17368 8576
rect 17328 8430 17356 8570
rect 17316 8424 17368 8430
rect 17316 8366 17368 8372
rect 17132 8356 17184 8362
rect 17132 8298 17184 8304
rect 17144 7886 17172 8298
rect 17132 7880 17184 7886
rect 17132 7822 17184 7828
rect 17144 7546 17172 7822
rect 17132 7540 17184 7546
rect 17132 7482 17184 7488
rect 16948 7404 17000 7410
rect 16948 7346 17000 7352
rect 17040 7404 17092 7410
rect 17040 7346 17092 7352
rect 16764 7268 16816 7274
rect 16764 7210 16816 7216
rect 17328 6866 17356 8366
rect 17512 7290 17540 8774
rect 17604 7886 17632 9318
rect 17684 8424 17736 8430
rect 17684 8366 17736 8372
rect 17696 8090 17724 8366
rect 17684 8084 17736 8090
rect 17684 8026 17736 8032
rect 17592 7880 17644 7886
rect 17592 7822 17644 7828
rect 17604 7410 17632 7822
rect 17592 7404 17644 7410
rect 17592 7346 17644 7352
rect 17512 7262 17632 7290
rect 16672 6860 16724 6866
rect 16672 6802 16724 6808
rect 17316 6860 17368 6866
rect 17316 6802 17368 6808
rect 16672 6724 16724 6730
rect 16672 6666 16724 6672
rect 16580 6384 16632 6390
rect 16580 6326 16632 6332
rect 16028 6112 16080 6118
rect 16028 6054 16080 6060
rect 16212 6112 16264 6118
rect 16212 6054 16264 6060
rect 16040 5817 16068 6054
rect 16026 5808 16082 5817
rect 15936 5772 15988 5778
rect 16026 5743 16082 5752
rect 15936 5714 15988 5720
rect 16040 5710 16068 5743
rect 16224 5710 16252 6054
rect 15752 5704 15804 5710
rect 15752 5646 15804 5652
rect 16028 5704 16080 5710
rect 16028 5646 16080 5652
rect 16212 5704 16264 5710
rect 16212 5646 16264 5652
rect 15292 5636 15344 5642
rect 15292 5578 15344 5584
rect 15304 5302 15332 5578
rect 15292 5296 15344 5302
rect 15292 5238 15344 5244
rect 15764 5166 15792 5646
rect 15752 5160 15804 5166
rect 15752 5102 15804 5108
rect 15152 4924 15460 4933
rect 15152 4922 15158 4924
rect 15214 4922 15238 4924
rect 15294 4922 15318 4924
rect 15374 4922 15398 4924
rect 15454 4922 15460 4924
rect 15214 4870 15216 4922
rect 15396 4870 15398 4922
rect 15152 4868 15158 4870
rect 15214 4868 15238 4870
rect 15294 4868 15318 4870
rect 15374 4868 15398 4870
rect 15454 4868 15460 4870
rect 15152 4859 15460 4868
rect 15764 4486 15792 5102
rect 16040 4622 16068 5646
rect 16224 5370 16252 5646
rect 16120 5364 16172 5370
rect 16120 5306 16172 5312
rect 16212 5364 16264 5370
rect 16212 5306 16264 5312
rect 16132 5250 16160 5306
rect 16684 5273 16712 6666
rect 17500 6656 17552 6662
rect 17500 6598 17552 6604
rect 17316 6316 17368 6322
rect 17316 6258 17368 6264
rect 16764 5908 16816 5914
rect 16764 5850 16816 5856
rect 16670 5264 16726 5273
rect 16132 5222 16528 5250
rect 16212 4820 16264 4826
rect 16212 4762 16264 4768
rect 16224 4622 16252 4762
rect 16500 4622 16528 5222
rect 16670 5199 16726 5208
rect 16776 4826 16804 5850
rect 17328 5710 17356 6258
rect 17316 5704 17368 5710
rect 17316 5646 17368 5652
rect 17408 5636 17460 5642
rect 17408 5578 17460 5584
rect 17420 5234 17448 5578
rect 16856 5228 16908 5234
rect 16856 5170 16908 5176
rect 17408 5228 17460 5234
rect 17408 5170 17460 5176
rect 16764 4820 16816 4826
rect 16764 4762 16816 4768
rect 16028 4616 16080 4622
rect 16028 4558 16080 4564
rect 16212 4616 16264 4622
rect 16212 4558 16264 4564
rect 16488 4616 16540 4622
rect 16488 4558 16540 4564
rect 15844 4548 15896 4554
rect 15844 4490 15896 4496
rect 15752 4480 15804 4486
rect 15752 4422 15804 4428
rect 15752 4140 15804 4146
rect 15752 4082 15804 4088
rect 14740 4072 14792 4078
rect 14740 4014 14792 4020
rect 14924 4072 14976 4078
rect 14924 4014 14976 4020
rect 14556 3732 14608 3738
rect 14556 3674 14608 3680
rect 14568 3194 14596 3674
rect 14648 3392 14700 3398
rect 14648 3334 14700 3340
rect 14556 3188 14608 3194
rect 14556 3130 14608 3136
rect 14660 3058 14688 3334
rect 14752 3194 14780 4014
rect 15152 3836 15460 3845
rect 15152 3834 15158 3836
rect 15214 3834 15238 3836
rect 15294 3834 15318 3836
rect 15374 3834 15398 3836
rect 15454 3834 15460 3836
rect 15214 3782 15216 3834
rect 15396 3782 15398 3834
rect 15152 3780 15158 3782
rect 15214 3780 15238 3782
rect 15294 3780 15318 3782
rect 15374 3780 15398 3782
rect 15454 3780 15460 3782
rect 15152 3771 15460 3780
rect 15764 3602 15792 4082
rect 15752 3596 15804 3602
rect 15752 3538 15804 3544
rect 14830 3496 14886 3505
rect 14830 3431 14886 3440
rect 14740 3188 14792 3194
rect 14740 3130 14792 3136
rect 14844 3058 14872 3431
rect 14648 3052 14700 3058
rect 14648 2994 14700 3000
rect 14832 3052 14884 3058
rect 14832 2994 14884 3000
rect 15764 2854 15792 3538
rect 15856 3534 15884 4490
rect 16040 4282 16068 4558
rect 16580 4548 16632 4554
rect 16580 4490 16632 4496
rect 16028 4276 16080 4282
rect 16028 4218 16080 4224
rect 16118 4176 16174 4185
rect 15936 4140 15988 4146
rect 16118 4111 16120 4120
rect 15936 4082 15988 4088
rect 16172 4111 16174 4120
rect 16120 4082 16172 4088
rect 15948 3738 15976 4082
rect 15936 3732 15988 3738
rect 15936 3674 15988 3680
rect 16132 3534 16160 4082
rect 16592 3942 16620 4490
rect 16580 3936 16632 3942
rect 16580 3878 16632 3884
rect 16578 3632 16634 3641
rect 16578 3567 16634 3576
rect 16592 3534 16620 3567
rect 15844 3528 15896 3534
rect 15844 3470 15896 3476
rect 16120 3528 16172 3534
rect 16120 3470 16172 3476
rect 16580 3528 16632 3534
rect 16580 3470 16632 3476
rect 16868 3194 16896 5170
rect 17316 4616 17368 4622
rect 17316 4558 17368 4564
rect 16948 4548 17000 4554
rect 16948 4490 17000 4496
rect 16960 4010 16988 4490
rect 16948 4004 17000 4010
rect 16948 3946 17000 3952
rect 16948 3528 17000 3534
rect 16946 3496 16948 3505
rect 17000 3496 17002 3505
rect 16946 3431 17002 3440
rect 16856 3188 16908 3194
rect 16856 3130 16908 3136
rect 17038 3088 17094 3097
rect 17328 3058 17356 4558
rect 17512 4146 17540 6598
rect 17604 5574 17632 7262
rect 17788 6662 17816 11086
rect 17880 11082 17908 12056
rect 17992 11996 18300 12005
rect 17992 11994 17998 11996
rect 18054 11994 18078 11996
rect 18134 11994 18158 11996
rect 18214 11994 18238 11996
rect 18294 11994 18300 11996
rect 18054 11942 18056 11994
rect 18236 11942 18238 11994
rect 17992 11940 17998 11942
rect 18054 11940 18078 11942
rect 18134 11940 18158 11942
rect 18214 11940 18238 11942
rect 18294 11940 18300 11942
rect 17992 11931 18300 11940
rect 18236 11144 18288 11150
rect 18234 11112 18236 11121
rect 18288 11112 18290 11121
rect 17868 11076 17920 11082
rect 18234 11047 18290 11056
rect 17868 11018 17920 11024
rect 17992 10908 18300 10917
rect 17992 10906 17998 10908
rect 18054 10906 18078 10908
rect 18134 10906 18158 10908
rect 18214 10906 18238 10908
rect 18294 10906 18300 10908
rect 18054 10854 18056 10906
rect 18236 10854 18238 10906
rect 17992 10852 17998 10854
rect 18054 10852 18078 10854
rect 18134 10852 18158 10854
rect 18214 10852 18238 10854
rect 18294 10852 18300 10854
rect 17992 10843 18300 10852
rect 18052 10668 18104 10674
rect 18052 10610 18104 10616
rect 18064 10538 18092 10610
rect 18052 10532 18104 10538
rect 18052 10474 18104 10480
rect 17868 10192 17920 10198
rect 18340 10146 18368 14894
rect 18420 13456 18472 13462
rect 18616 13433 18644 20402
rect 18984 20058 19012 20402
rect 18972 20052 19024 20058
rect 18972 19994 19024 20000
rect 18696 19848 18748 19854
rect 18696 19790 18748 19796
rect 18708 19446 18736 19790
rect 18696 19440 18748 19446
rect 18696 19382 18748 19388
rect 18708 18290 18736 19382
rect 19168 19310 19196 21626
rect 20833 21244 21141 21253
rect 20833 21242 20839 21244
rect 20895 21242 20919 21244
rect 20975 21242 20999 21244
rect 21055 21242 21079 21244
rect 21135 21242 21141 21244
rect 20895 21190 20897 21242
rect 21077 21190 21079 21242
rect 20833 21188 20839 21190
rect 20895 21188 20919 21190
rect 20975 21188 20999 21190
rect 21055 21188 21079 21190
rect 21135 21188 21141 21190
rect 20833 21179 21141 21188
rect 21192 20942 21220 21626
rect 22388 21554 22416 21830
rect 23673 21788 23981 21797
rect 23673 21786 23679 21788
rect 23735 21786 23759 21788
rect 23815 21786 23839 21788
rect 23895 21786 23919 21788
rect 23975 21786 23981 21788
rect 23735 21734 23737 21786
rect 23917 21734 23919 21786
rect 23673 21732 23679 21734
rect 23735 21732 23759 21734
rect 23815 21732 23839 21734
rect 23895 21732 23919 21734
rect 23975 21732 23981 21734
rect 23673 21723 23981 21732
rect 21272 21548 21324 21554
rect 21272 21490 21324 21496
rect 22376 21548 22428 21554
rect 22376 21490 22428 21496
rect 21284 21146 21312 21490
rect 21272 21140 21324 21146
rect 21272 21082 21324 21088
rect 22100 21004 22152 21010
rect 22100 20946 22152 20952
rect 21180 20936 21232 20942
rect 21180 20878 21232 20884
rect 22112 20602 22140 20946
rect 22388 20942 22416 21490
rect 22376 20936 22428 20942
rect 22376 20878 22428 20884
rect 23673 20700 23981 20709
rect 23673 20698 23679 20700
rect 23735 20698 23759 20700
rect 23815 20698 23839 20700
rect 23895 20698 23919 20700
rect 23975 20698 23981 20700
rect 23735 20646 23737 20698
rect 23917 20646 23919 20698
rect 23673 20644 23679 20646
rect 23735 20644 23759 20646
rect 23815 20644 23839 20646
rect 23895 20644 23919 20646
rect 23975 20644 23981 20646
rect 23673 20635 23981 20644
rect 19432 20596 19484 20602
rect 19432 20538 19484 20544
rect 22100 20596 22152 20602
rect 22100 20538 22152 20544
rect 19444 20466 19472 20538
rect 19432 20460 19484 20466
rect 19432 20402 19484 20408
rect 20168 20460 20220 20466
rect 20168 20402 20220 20408
rect 22192 20460 22244 20466
rect 22192 20402 22244 20408
rect 19340 20324 19392 20330
rect 19340 20266 19392 20272
rect 19352 19378 19380 20266
rect 19444 19922 19472 20402
rect 20076 20392 20128 20398
rect 20076 20334 20128 20340
rect 19432 19916 19484 19922
rect 19432 19858 19484 19864
rect 19892 19712 19944 19718
rect 19892 19654 19944 19660
rect 19340 19372 19392 19378
rect 19340 19314 19392 19320
rect 19524 19372 19576 19378
rect 19524 19314 19576 19320
rect 19616 19372 19668 19378
rect 19616 19314 19668 19320
rect 18972 19304 19024 19310
rect 18972 19246 19024 19252
rect 19156 19304 19208 19310
rect 19156 19246 19208 19252
rect 18880 18964 18932 18970
rect 18880 18906 18932 18912
rect 18892 18834 18920 18906
rect 18880 18828 18932 18834
rect 18880 18770 18932 18776
rect 18984 18766 19012 19246
rect 18788 18760 18840 18766
rect 18788 18702 18840 18708
rect 18972 18760 19024 18766
rect 18972 18702 19024 18708
rect 18800 18426 18828 18702
rect 18788 18420 18840 18426
rect 18788 18362 18840 18368
rect 18696 18284 18748 18290
rect 18696 18226 18748 18232
rect 18708 14278 18736 18226
rect 18880 17332 18932 17338
rect 18880 17274 18932 17280
rect 18788 17128 18840 17134
rect 18788 17070 18840 17076
rect 18800 16522 18828 17070
rect 18788 16516 18840 16522
rect 18788 16458 18840 16464
rect 18892 16454 18920 17274
rect 18984 16998 19012 18702
rect 19248 18352 19300 18358
rect 19248 18294 19300 18300
rect 19260 17202 19288 18294
rect 19340 17604 19392 17610
rect 19340 17546 19392 17552
rect 19432 17604 19484 17610
rect 19432 17546 19484 17552
rect 19248 17196 19300 17202
rect 19248 17138 19300 17144
rect 18972 16992 19024 16998
rect 18972 16934 19024 16940
rect 19248 16992 19300 16998
rect 19248 16934 19300 16940
rect 18970 16824 19026 16833
rect 18970 16759 19026 16768
rect 18880 16448 18932 16454
rect 18880 16390 18932 16396
rect 18788 15564 18840 15570
rect 18788 15506 18840 15512
rect 18800 14822 18828 15506
rect 18788 14816 18840 14822
rect 18788 14758 18840 14764
rect 18696 14272 18748 14278
rect 18696 14214 18748 14220
rect 18420 13398 18472 13404
rect 18602 13424 18658 13433
rect 18432 12238 18460 13398
rect 18602 13359 18658 13368
rect 18512 12708 18564 12714
rect 18512 12650 18564 12656
rect 18420 12232 18472 12238
rect 18420 12174 18472 12180
rect 18420 11552 18472 11558
rect 18420 11494 18472 11500
rect 18432 11014 18460 11494
rect 18524 11234 18552 12650
rect 18604 12640 18656 12646
rect 18604 12582 18656 12588
rect 18616 12170 18644 12582
rect 18604 12164 18656 12170
rect 18604 12106 18656 12112
rect 18602 11248 18658 11257
rect 18524 11206 18602 11234
rect 18602 11183 18658 11192
rect 18616 11150 18644 11183
rect 18604 11144 18656 11150
rect 18510 11112 18566 11121
rect 18604 11086 18656 11092
rect 18510 11047 18566 11056
rect 18420 11008 18472 11014
rect 18420 10950 18472 10956
rect 18524 10266 18552 11047
rect 18708 10713 18736 14214
rect 18892 13734 18920 16390
rect 18984 15638 19012 16759
rect 19260 16726 19288 16934
rect 19248 16720 19300 16726
rect 19248 16662 19300 16668
rect 19156 16040 19208 16046
rect 19156 15982 19208 15988
rect 18972 15632 19024 15638
rect 18972 15574 19024 15580
rect 18880 13728 18932 13734
rect 18880 13670 18932 13676
rect 18788 13388 18840 13394
rect 18788 13330 18840 13336
rect 18800 11830 18828 13330
rect 18892 13190 18920 13670
rect 18880 13184 18932 13190
rect 18880 13126 18932 13132
rect 18788 11824 18840 11830
rect 18788 11766 18840 11772
rect 18892 11744 18920 13126
rect 18984 12442 19012 15574
rect 19064 15428 19116 15434
rect 19064 15370 19116 15376
rect 18972 12436 19024 12442
rect 18972 12378 19024 12384
rect 18972 11756 19024 11762
rect 18892 11716 18972 11744
rect 19076 11744 19104 15370
rect 19168 14346 19196 15982
rect 19248 15700 19300 15706
rect 19248 15642 19300 15648
rect 19260 15162 19288 15642
rect 19248 15156 19300 15162
rect 19248 15098 19300 15104
rect 19352 15094 19380 17546
rect 19444 16114 19472 17546
rect 19536 17338 19564 19314
rect 19628 18970 19656 19314
rect 19708 19168 19760 19174
rect 19708 19110 19760 19116
rect 19616 18964 19668 18970
rect 19616 18906 19668 18912
rect 19720 18766 19748 19110
rect 19904 18766 19932 19654
rect 20088 19310 20116 20334
rect 20076 19304 20128 19310
rect 20076 19246 20128 19252
rect 19708 18760 19760 18766
rect 19708 18702 19760 18708
rect 19892 18760 19944 18766
rect 19892 18702 19944 18708
rect 20076 18760 20128 18766
rect 20076 18702 20128 18708
rect 19904 18426 19932 18702
rect 19892 18420 19944 18426
rect 19892 18362 19944 18368
rect 19708 18284 19760 18290
rect 19708 18226 19760 18232
rect 19720 17746 19748 18226
rect 19892 18080 19944 18086
rect 19892 18022 19944 18028
rect 19800 17876 19852 17882
rect 19800 17818 19852 17824
rect 19708 17740 19760 17746
rect 19708 17682 19760 17688
rect 19524 17332 19576 17338
rect 19524 17274 19576 17280
rect 19720 17066 19748 17682
rect 19708 17060 19760 17066
rect 19708 17002 19760 17008
rect 19812 16114 19840 17818
rect 19432 16108 19484 16114
rect 19432 16050 19484 16056
rect 19616 16108 19668 16114
rect 19616 16050 19668 16056
rect 19800 16108 19852 16114
rect 19800 16050 19852 16056
rect 19444 15586 19472 16050
rect 19628 15706 19656 16050
rect 19708 15904 19760 15910
rect 19708 15846 19760 15852
rect 19616 15700 19668 15706
rect 19616 15642 19668 15648
rect 19444 15558 19656 15586
rect 19524 15496 19576 15502
rect 19524 15438 19576 15444
rect 19340 15088 19392 15094
rect 19340 15030 19392 15036
rect 19248 15020 19300 15026
rect 19248 14962 19300 14968
rect 19260 14498 19288 14962
rect 19338 14648 19394 14657
rect 19338 14583 19340 14592
rect 19392 14583 19394 14592
rect 19340 14554 19392 14560
rect 19260 14470 19472 14498
rect 19340 14408 19392 14414
rect 19340 14350 19392 14356
rect 19156 14340 19208 14346
rect 19156 14282 19208 14288
rect 19168 13870 19196 14282
rect 19156 13864 19208 13870
rect 19156 13806 19208 13812
rect 19168 13258 19196 13806
rect 19248 13320 19300 13326
rect 19248 13262 19300 13268
rect 19156 13252 19208 13258
rect 19156 13194 19208 13200
rect 19156 12436 19208 12442
rect 19156 12378 19208 12384
rect 19168 11898 19196 12378
rect 19156 11892 19208 11898
rect 19156 11834 19208 11840
rect 19076 11716 19196 11744
rect 18972 11698 19024 11704
rect 18788 11552 18840 11558
rect 18788 11494 18840 11500
rect 18800 11150 18828 11494
rect 18788 11144 18840 11150
rect 18788 11086 18840 11092
rect 18880 11076 18932 11082
rect 18880 11018 18932 11024
rect 18788 11008 18840 11014
rect 18788 10950 18840 10956
rect 18694 10704 18750 10713
rect 18694 10639 18750 10648
rect 18604 10600 18656 10606
rect 18604 10542 18656 10548
rect 18512 10260 18564 10266
rect 18512 10202 18564 10208
rect 17868 10134 17920 10140
rect 17880 9994 17908 10134
rect 18248 10118 18460 10146
rect 18144 10056 18196 10062
rect 18248 10044 18276 10118
rect 18196 10016 18276 10044
rect 18328 10056 18380 10062
rect 18144 9998 18196 10004
rect 18328 9998 18380 10004
rect 17868 9988 17920 9994
rect 17868 9930 17920 9936
rect 17992 9820 18300 9829
rect 17992 9818 17998 9820
rect 18054 9818 18078 9820
rect 18134 9818 18158 9820
rect 18214 9818 18238 9820
rect 18294 9818 18300 9820
rect 18054 9766 18056 9818
rect 18236 9766 18238 9818
rect 17992 9764 17998 9766
rect 18054 9764 18078 9766
rect 18134 9764 18158 9766
rect 18214 9764 18238 9766
rect 18294 9764 18300 9766
rect 17992 9755 18300 9764
rect 18340 9586 18368 9998
rect 18432 9586 18460 10118
rect 18328 9580 18380 9586
rect 18328 9522 18380 9528
rect 18420 9580 18472 9586
rect 18420 9522 18472 9528
rect 18328 8968 18380 8974
rect 18524 8956 18552 10202
rect 18380 8928 18552 8956
rect 18328 8910 18380 8916
rect 17992 8732 18300 8741
rect 17992 8730 17998 8732
rect 18054 8730 18078 8732
rect 18134 8730 18158 8732
rect 18214 8730 18238 8732
rect 18294 8730 18300 8732
rect 18054 8678 18056 8730
rect 18236 8678 18238 8730
rect 17992 8676 17998 8678
rect 18054 8676 18078 8678
rect 18134 8676 18158 8678
rect 18214 8676 18238 8678
rect 18294 8676 18300 8678
rect 17992 8667 18300 8676
rect 18234 8528 18290 8537
rect 18234 8463 18236 8472
rect 18288 8463 18290 8472
rect 18236 8434 18288 8440
rect 17992 7644 18300 7653
rect 17992 7642 17998 7644
rect 18054 7642 18078 7644
rect 18134 7642 18158 7644
rect 18214 7642 18238 7644
rect 18294 7642 18300 7644
rect 18054 7590 18056 7642
rect 18236 7590 18238 7642
rect 17992 7588 17998 7590
rect 18054 7588 18078 7590
rect 18134 7588 18158 7590
rect 18214 7588 18238 7590
rect 18294 7588 18300 7590
rect 17992 7579 18300 7588
rect 18340 7460 18368 8910
rect 18616 7886 18644 10542
rect 18708 9994 18736 10639
rect 18696 9988 18748 9994
rect 18696 9930 18748 9936
rect 18800 9674 18828 10950
rect 18892 10130 18920 11018
rect 18880 10124 18932 10130
rect 18880 10066 18932 10072
rect 18800 9646 18920 9674
rect 18892 8838 18920 9646
rect 18880 8832 18932 8838
rect 18880 8774 18932 8780
rect 18892 8498 18920 8774
rect 18880 8492 18932 8498
rect 18880 8434 18932 8440
rect 18604 7880 18656 7886
rect 18604 7822 18656 7828
rect 18420 7812 18472 7818
rect 18420 7754 18472 7760
rect 18248 7432 18368 7460
rect 17868 7404 17920 7410
rect 17868 7346 17920 7352
rect 17776 6656 17828 6662
rect 17776 6598 17828 6604
rect 17880 6304 17908 7346
rect 18248 6866 18276 7432
rect 18236 6860 18288 6866
rect 18236 6802 18288 6808
rect 18328 6792 18380 6798
rect 18328 6734 18380 6740
rect 17992 6556 18300 6565
rect 17992 6554 17998 6556
rect 18054 6554 18078 6556
rect 18134 6554 18158 6556
rect 18214 6554 18238 6556
rect 18294 6554 18300 6556
rect 18054 6502 18056 6554
rect 18236 6502 18238 6554
rect 17992 6500 17998 6502
rect 18054 6500 18078 6502
rect 18134 6500 18158 6502
rect 18214 6500 18238 6502
rect 18294 6500 18300 6502
rect 17992 6491 18300 6500
rect 18144 6452 18196 6458
rect 18144 6394 18196 6400
rect 17958 6352 18014 6361
rect 18156 6322 18184 6394
rect 17880 6296 17958 6304
rect 17880 6276 17960 6296
rect 18012 6287 18014 6296
rect 18144 6316 18196 6322
rect 17960 6258 18012 6264
rect 18144 6258 18196 6264
rect 18236 6248 18288 6254
rect 18236 6190 18288 6196
rect 17868 5840 17920 5846
rect 17868 5782 17920 5788
rect 17684 5772 17736 5778
rect 17684 5714 17736 5720
rect 17592 5568 17644 5574
rect 17592 5510 17644 5516
rect 17604 5166 17632 5510
rect 17696 5370 17724 5714
rect 17880 5710 17908 5782
rect 17868 5704 17920 5710
rect 17868 5646 17920 5652
rect 18248 5658 18276 6190
rect 18340 5778 18368 6734
rect 18432 5914 18460 7754
rect 18512 7404 18564 7410
rect 18512 7346 18564 7352
rect 18524 6730 18552 7346
rect 18512 6724 18564 6730
rect 18512 6666 18564 6672
rect 18524 6322 18552 6666
rect 18512 6316 18564 6322
rect 18512 6258 18564 6264
rect 18616 6186 18644 7822
rect 18984 7750 19012 11698
rect 19168 10810 19196 11716
rect 19156 10804 19208 10810
rect 19156 10746 19208 10752
rect 19062 10704 19118 10713
rect 19062 10639 19118 10648
rect 19156 10702 19208 10708
rect 19156 10644 19208 10650
rect 19076 10538 19104 10639
rect 19064 10532 19116 10538
rect 19064 10474 19116 10480
rect 18696 7744 18748 7750
rect 18696 7686 18748 7692
rect 18972 7744 19024 7750
rect 18972 7686 19024 7692
rect 18708 7206 18736 7686
rect 18696 7200 18748 7206
rect 18696 7142 18748 7148
rect 18512 6180 18564 6186
rect 18512 6122 18564 6128
rect 18604 6180 18656 6186
rect 18604 6122 18656 6128
rect 18420 5908 18472 5914
rect 18420 5850 18472 5856
rect 18524 5778 18552 6122
rect 18328 5772 18380 5778
rect 18328 5714 18380 5720
rect 18512 5772 18564 5778
rect 18512 5714 18564 5720
rect 17684 5364 17736 5370
rect 17684 5306 17736 5312
rect 17696 5166 17724 5306
rect 17880 5234 17908 5646
rect 18248 5630 18368 5658
rect 17992 5468 18300 5477
rect 17992 5466 17998 5468
rect 18054 5466 18078 5468
rect 18134 5466 18158 5468
rect 18214 5466 18238 5468
rect 18294 5466 18300 5468
rect 18054 5414 18056 5466
rect 18236 5414 18238 5466
rect 17992 5412 17998 5414
rect 18054 5412 18078 5414
rect 18134 5412 18158 5414
rect 18214 5412 18238 5414
rect 18294 5412 18300 5414
rect 17992 5403 18300 5412
rect 17868 5228 17920 5234
rect 17868 5170 17920 5176
rect 17592 5160 17644 5166
rect 17592 5102 17644 5108
rect 17684 5160 17736 5166
rect 17684 5102 17736 5108
rect 17500 4140 17552 4146
rect 17500 4082 17552 4088
rect 17880 4010 17908 5170
rect 18340 5166 18368 5630
rect 18512 5296 18564 5302
rect 18512 5238 18564 5244
rect 18328 5160 18380 5166
rect 18328 5102 18380 5108
rect 18420 5160 18472 5166
rect 18420 5102 18472 5108
rect 17992 4380 18300 4389
rect 17992 4378 17998 4380
rect 18054 4378 18078 4380
rect 18134 4378 18158 4380
rect 18214 4378 18238 4380
rect 18294 4378 18300 4380
rect 18054 4326 18056 4378
rect 18236 4326 18238 4378
rect 17992 4324 17998 4326
rect 18054 4324 18078 4326
rect 18134 4324 18158 4326
rect 18214 4324 18238 4326
rect 18294 4324 18300 4326
rect 17992 4315 18300 4324
rect 18328 4276 18380 4282
rect 18432 4264 18460 5102
rect 18524 4282 18552 5238
rect 18708 5030 18736 7142
rect 19076 6934 19104 10474
rect 19168 10062 19196 10644
rect 19260 10538 19288 13262
rect 19352 12986 19380 14350
rect 19340 12980 19392 12986
rect 19340 12922 19392 12928
rect 19340 12844 19392 12850
rect 19340 12786 19392 12792
rect 19352 12646 19380 12786
rect 19340 12640 19392 12646
rect 19340 12582 19392 12588
rect 19340 11688 19392 11694
rect 19340 11630 19392 11636
rect 19248 10532 19300 10538
rect 19248 10474 19300 10480
rect 19156 10056 19208 10062
rect 19156 9998 19208 10004
rect 19352 8362 19380 11630
rect 19444 8838 19472 14470
rect 19536 13870 19564 15438
rect 19628 14414 19656 15558
rect 19720 14550 19748 15846
rect 19812 15434 19840 16050
rect 19904 15570 19932 18022
rect 20088 17678 20116 18702
rect 20180 18352 20208 20402
rect 20833 20156 21141 20165
rect 20833 20154 20839 20156
rect 20895 20154 20919 20156
rect 20975 20154 20999 20156
rect 21055 20154 21079 20156
rect 21135 20154 21141 20156
rect 20895 20102 20897 20154
rect 21077 20102 21079 20154
rect 20833 20100 20839 20102
rect 20895 20100 20919 20102
rect 20975 20100 20999 20102
rect 21055 20100 21079 20102
rect 21135 20100 21141 20102
rect 20833 20091 21141 20100
rect 20444 19916 20496 19922
rect 20444 19858 20496 19864
rect 20260 19372 20312 19378
rect 20260 19314 20312 19320
rect 20272 18766 20300 19314
rect 20456 18766 20484 19858
rect 20996 19848 21048 19854
rect 20996 19790 21048 19796
rect 21008 19310 21036 19790
rect 21180 19372 21232 19378
rect 21180 19314 21232 19320
rect 22100 19372 22152 19378
rect 22100 19314 22152 19320
rect 20996 19304 21048 19310
rect 20996 19246 21048 19252
rect 20833 19068 21141 19077
rect 20833 19066 20839 19068
rect 20895 19066 20919 19068
rect 20975 19066 20999 19068
rect 21055 19066 21079 19068
rect 21135 19066 21141 19068
rect 20895 19014 20897 19066
rect 21077 19014 21079 19066
rect 20833 19012 20839 19014
rect 20895 19012 20919 19014
rect 20975 19012 20999 19014
rect 21055 19012 21079 19014
rect 21135 19012 21141 19014
rect 20833 19003 21141 19012
rect 20720 18896 20772 18902
rect 20720 18838 20772 18844
rect 20260 18760 20312 18766
rect 20444 18760 20496 18766
rect 20260 18702 20312 18708
rect 20364 18720 20444 18748
rect 20364 18358 20392 18720
rect 20444 18702 20496 18708
rect 20628 18692 20680 18698
rect 20628 18634 20680 18640
rect 20177 18290 20208 18352
rect 20352 18352 20404 18358
rect 20352 18294 20404 18300
rect 20165 18284 20217 18290
rect 20165 18226 20217 18232
rect 20260 18284 20312 18290
rect 20260 18226 20312 18232
rect 19984 17672 20036 17678
rect 19984 17614 20036 17620
rect 20076 17672 20128 17678
rect 20076 17614 20128 17620
rect 19996 16164 20024 17614
rect 20088 17270 20116 17614
rect 20076 17264 20128 17270
rect 20076 17206 20128 17212
rect 20180 16454 20208 18226
rect 20168 16448 20220 16454
rect 20168 16390 20220 16396
rect 20272 16250 20300 18226
rect 20352 17060 20404 17066
rect 20352 17002 20404 17008
rect 20364 16658 20392 17002
rect 20536 16720 20588 16726
rect 20536 16662 20588 16668
rect 20352 16652 20404 16658
rect 20352 16594 20404 16600
rect 20444 16584 20496 16590
rect 20444 16526 20496 16532
rect 20260 16244 20312 16250
rect 20260 16186 20312 16192
rect 20168 16176 20220 16182
rect 19996 16136 20168 16164
rect 20168 16118 20220 16124
rect 19892 15564 19944 15570
rect 19892 15506 19944 15512
rect 19800 15428 19852 15434
rect 19800 15370 19852 15376
rect 19904 15026 19932 15506
rect 19800 15020 19852 15026
rect 19800 14962 19852 14968
rect 19892 15020 19944 15026
rect 19892 14962 19944 14968
rect 19708 14544 19760 14550
rect 19708 14486 19760 14492
rect 19616 14408 19668 14414
rect 19616 14350 19668 14356
rect 19524 13864 19576 13870
rect 19524 13806 19576 13812
rect 19628 13818 19656 14350
rect 19812 14074 19840 14962
rect 20076 14340 20128 14346
rect 20076 14282 20128 14288
rect 19800 14068 19852 14074
rect 19800 14010 19852 14016
rect 19890 13968 19946 13977
rect 19890 13903 19946 13912
rect 19536 13410 19564 13806
rect 19628 13790 19840 13818
rect 19614 13560 19670 13569
rect 19812 13530 19840 13790
rect 19614 13495 19616 13504
rect 19668 13495 19670 13504
rect 19708 13524 19760 13530
rect 19616 13466 19668 13472
rect 19708 13466 19760 13472
rect 19800 13524 19852 13530
rect 19800 13466 19852 13472
rect 19720 13410 19748 13466
rect 19536 13394 19748 13410
rect 19524 13388 19748 13394
rect 19576 13382 19748 13388
rect 19524 13330 19576 13336
rect 19616 13252 19668 13258
rect 19616 13194 19668 13200
rect 19524 11824 19576 11830
rect 19524 11766 19576 11772
rect 19536 10470 19564 11766
rect 19628 11354 19656 13194
rect 19706 13152 19762 13161
rect 19706 13087 19762 13096
rect 19720 12306 19748 13087
rect 19904 12850 19932 13903
rect 19984 13728 20036 13734
rect 19984 13670 20036 13676
rect 19996 13258 20024 13670
rect 19984 13252 20036 13258
rect 19984 13194 20036 13200
rect 19996 12986 20024 13194
rect 19984 12980 20036 12986
rect 19984 12922 20036 12928
rect 19892 12844 19944 12850
rect 19892 12786 19944 12792
rect 19800 12708 19852 12714
rect 19800 12650 19852 12656
rect 19708 12300 19760 12306
rect 19708 12242 19760 12248
rect 19616 11348 19668 11354
rect 19616 11290 19668 11296
rect 19628 11082 19656 11290
rect 19720 11234 19748 12242
rect 19812 11898 19840 12650
rect 19800 11892 19852 11898
rect 19800 11834 19852 11840
rect 19996 11762 20024 12922
rect 19984 11756 20036 11762
rect 19984 11698 20036 11704
rect 19984 11552 20036 11558
rect 19984 11494 20036 11500
rect 19720 11206 19840 11234
rect 19708 11144 19760 11150
rect 19708 11086 19760 11092
rect 19616 11076 19668 11082
rect 19616 11018 19668 11024
rect 19720 10674 19748 11086
rect 19812 10674 19840 11206
rect 19996 10742 20024 11494
rect 20088 10826 20116 14282
rect 20180 12170 20208 16118
rect 20352 15700 20404 15706
rect 20352 15642 20404 15648
rect 20260 15020 20312 15026
rect 20260 14962 20312 14968
rect 20272 14278 20300 14962
rect 20364 14618 20392 15642
rect 20352 14612 20404 14618
rect 20352 14554 20404 14560
rect 20260 14272 20312 14278
rect 20260 14214 20312 14220
rect 20260 13932 20312 13938
rect 20260 13874 20312 13880
rect 20272 12986 20300 13874
rect 20364 13258 20392 14554
rect 20352 13252 20404 13258
rect 20352 13194 20404 13200
rect 20364 13161 20392 13194
rect 20350 13152 20406 13161
rect 20350 13087 20406 13096
rect 20260 12980 20312 12986
rect 20260 12922 20312 12928
rect 20260 12844 20312 12850
rect 20260 12786 20312 12792
rect 20352 12844 20404 12850
rect 20352 12786 20404 12792
rect 20272 12617 20300 12786
rect 20258 12608 20314 12617
rect 20258 12543 20314 12552
rect 20364 12442 20392 12786
rect 20352 12436 20404 12442
rect 20272 12406 20352 12434
rect 20168 12164 20220 12170
rect 20168 12106 20220 12112
rect 20088 10798 20208 10826
rect 19984 10736 20036 10742
rect 19984 10678 20036 10684
rect 19708 10668 19760 10674
rect 19708 10610 19760 10616
rect 19800 10668 19852 10674
rect 19800 10610 19852 10616
rect 19616 10600 19668 10606
rect 19616 10542 19668 10548
rect 19524 10464 19576 10470
rect 19524 10406 19576 10412
rect 19524 9580 19576 9586
rect 19524 9522 19576 9528
rect 19432 8832 19484 8838
rect 19432 8774 19484 8780
rect 19536 8430 19564 9522
rect 19628 9450 19656 10542
rect 19812 10470 19840 10610
rect 19800 10464 19852 10470
rect 19800 10406 19852 10412
rect 19996 9926 20024 10678
rect 20076 10668 20128 10674
rect 20076 10610 20128 10616
rect 20088 10062 20116 10610
rect 20076 10056 20128 10062
rect 20076 9998 20128 10004
rect 19984 9920 20036 9926
rect 19984 9862 20036 9868
rect 19800 9648 19852 9654
rect 19800 9590 19852 9596
rect 19616 9444 19668 9450
rect 19616 9386 19668 9392
rect 19628 8906 19656 9386
rect 19708 9376 19760 9382
rect 19708 9318 19760 9324
rect 19720 9110 19748 9318
rect 19708 9104 19760 9110
rect 19708 9046 19760 9052
rect 19616 8900 19668 8906
rect 19616 8842 19668 8848
rect 19616 8560 19668 8566
rect 19616 8502 19668 8508
rect 19524 8424 19576 8430
rect 19524 8366 19576 8372
rect 19340 8356 19392 8362
rect 19340 8298 19392 8304
rect 19248 7268 19300 7274
rect 19248 7210 19300 7216
rect 19064 6928 19116 6934
rect 19064 6870 19116 6876
rect 19260 6798 19288 7210
rect 19248 6792 19300 6798
rect 19248 6734 19300 6740
rect 18788 6656 18840 6662
rect 18788 6598 18840 6604
rect 19156 6656 19208 6662
rect 19156 6598 19208 6604
rect 18800 5914 18828 6598
rect 19168 6361 19196 6598
rect 19154 6352 19210 6361
rect 19154 6287 19156 6296
rect 19208 6287 19210 6296
rect 19156 6258 19208 6264
rect 18788 5908 18840 5914
rect 18788 5850 18840 5856
rect 19260 5846 19288 6734
rect 19352 6458 19380 8298
rect 19432 8016 19484 8022
rect 19432 7958 19484 7964
rect 19340 6452 19392 6458
rect 19340 6394 19392 6400
rect 19444 6338 19472 7958
rect 19524 7812 19576 7818
rect 19628 7800 19656 8502
rect 19576 7772 19656 7800
rect 19524 7754 19576 7760
rect 19812 7410 19840 9590
rect 19892 8968 19944 8974
rect 19892 8910 19944 8916
rect 19904 8634 19932 8910
rect 19892 8628 19944 8634
rect 19892 8570 19944 8576
rect 19996 8090 20024 9862
rect 19984 8084 20036 8090
rect 19984 8026 20036 8032
rect 19996 7750 20024 8026
rect 20088 7818 20116 9998
rect 20180 7954 20208 10798
rect 20272 9586 20300 12406
rect 20352 12378 20404 12384
rect 20456 10130 20484 16526
rect 20548 10606 20576 16662
rect 20640 12850 20668 18634
rect 20732 17338 20760 18838
rect 21192 18766 21220 19314
rect 21364 19304 21416 19310
rect 21364 19246 21416 19252
rect 21180 18760 21232 18766
rect 21180 18702 21232 18708
rect 20904 18624 20956 18630
rect 20904 18566 20956 18572
rect 20916 18193 20944 18566
rect 20902 18184 20958 18193
rect 20902 18119 20958 18128
rect 20833 17980 21141 17989
rect 20833 17978 20839 17980
rect 20895 17978 20919 17980
rect 20975 17978 20999 17980
rect 21055 17978 21079 17980
rect 21135 17978 21141 17980
rect 20895 17926 20897 17978
rect 21077 17926 21079 17978
rect 20833 17924 20839 17926
rect 20895 17924 20919 17926
rect 20975 17924 20999 17926
rect 21055 17924 21079 17926
rect 21135 17924 21141 17926
rect 20833 17915 21141 17924
rect 20812 17536 20864 17542
rect 20812 17478 20864 17484
rect 20904 17536 20956 17542
rect 20904 17478 20956 17484
rect 20720 17332 20772 17338
rect 20720 17274 20772 17280
rect 20824 17134 20852 17478
rect 20916 17202 20944 17478
rect 20904 17196 20956 17202
rect 20904 17138 20956 17144
rect 20720 17128 20772 17134
rect 20720 17070 20772 17076
rect 20812 17128 20864 17134
rect 20812 17070 20864 17076
rect 20732 14618 20760 17070
rect 20833 16892 21141 16901
rect 20833 16890 20839 16892
rect 20895 16890 20919 16892
rect 20975 16890 20999 16892
rect 21055 16890 21079 16892
rect 21135 16890 21141 16892
rect 20895 16838 20897 16890
rect 21077 16838 21079 16890
rect 20833 16836 20839 16838
rect 20895 16836 20919 16838
rect 20975 16836 20999 16838
rect 21055 16836 21079 16838
rect 21135 16836 21141 16838
rect 20833 16827 21141 16836
rect 20996 16448 21048 16454
rect 20996 16390 21048 16396
rect 21008 16250 21036 16390
rect 20996 16244 21048 16250
rect 20996 16186 21048 16192
rect 20812 16176 20864 16182
rect 20810 16144 20812 16153
rect 20864 16144 20866 16153
rect 20810 16079 20866 16088
rect 20996 16108 21048 16114
rect 20996 16050 21048 16056
rect 21008 15910 21036 16050
rect 21192 15978 21220 18702
rect 21180 15972 21232 15978
rect 21180 15914 21232 15920
rect 20996 15904 21048 15910
rect 20996 15846 21048 15852
rect 20833 15804 21141 15813
rect 20833 15802 20839 15804
rect 20895 15802 20919 15804
rect 20975 15802 20999 15804
rect 21055 15802 21079 15804
rect 21135 15802 21141 15804
rect 20895 15750 20897 15802
rect 21077 15750 21079 15802
rect 20833 15748 20839 15750
rect 20895 15748 20919 15750
rect 20975 15748 20999 15750
rect 21055 15748 21079 15750
rect 21135 15748 21141 15750
rect 20833 15739 21141 15748
rect 20812 15428 20864 15434
rect 20812 15370 20864 15376
rect 20824 14958 20852 15370
rect 21192 15026 21220 15914
rect 21272 15904 21324 15910
rect 21272 15846 21324 15852
rect 21180 15020 21232 15026
rect 21180 14962 21232 14968
rect 20812 14952 20864 14958
rect 20812 14894 20864 14900
rect 20833 14716 21141 14725
rect 20833 14714 20839 14716
rect 20895 14714 20919 14716
rect 20975 14714 20999 14716
rect 21055 14714 21079 14716
rect 21135 14714 21141 14716
rect 20895 14662 20897 14714
rect 21077 14662 21079 14714
rect 20833 14660 20839 14662
rect 20895 14660 20919 14662
rect 20975 14660 20999 14662
rect 21055 14660 21079 14662
rect 21135 14660 21141 14662
rect 20833 14651 21141 14660
rect 20720 14612 20772 14618
rect 20720 14554 20772 14560
rect 21284 14550 21312 15846
rect 21376 15502 21404 19246
rect 21732 19168 21784 19174
rect 21732 19110 21784 19116
rect 21456 18420 21508 18426
rect 21456 18362 21508 18368
rect 21364 15496 21416 15502
rect 21364 15438 21416 15444
rect 21364 14884 21416 14890
rect 21364 14826 21416 14832
rect 21272 14544 21324 14550
rect 21272 14486 21324 14492
rect 20994 13968 21050 13977
rect 20812 13898 20864 13904
rect 20994 13903 20996 13912
rect 21048 13903 21050 13912
rect 20996 13874 21048 13880
rect 20812 13840 20864 13846
rect 20824 13716 20852 13840
rect 20824 13688 21220 13716
rect 20833 13628 21141 13637
rect 20833 13626 20839 13628
rect 20895 13626 20919 13628
rect 20975 13626 20999 13628
rect 21055 13626 21079 13628
rect 21135 13626 21141 13628
rect 20895 13574 20897 13626
rect 21077 13574 21079 13626
rect 20833 13572 20839 13574
rect 20895 13572 20919 13574
rect 20975 13572 20999 13574
rect 21055 13572 21079 13574
rect 21135 13572 21141 13574
rect 20833 13563 21141 13572
rect 20904 13388 20956 13394
rect 20904 13330 20956 13336
rect 20628 12844 20680 12850
rect 20628 12786 20680 12792
rect 20720 12844 20772 12850
rect 20720 12786 20772 12792
rect 20628 12640 20680 12646
rect 20628 12582 20680 12588
rect 20640 12220 20668 12582
rect 20732 12434 20760 12786
rect 20916 12628 20944 13330
rect 21192 12696 21220 13688
rect 21376 12918 21404 14826
rect 21468 14414 21496 18362
rect 21744 14414 21772 19110
rect 22112 18630 22140 19314
rect 22100 18624 22152 18630
rect 22100 18566 22152 18572
rect 21824 17672 21876 17678
rect 21824 17614 21876 17620
rect 21836 16114 21864 17614
rect 22008 17536 22060 17542
rect 22008 17478 22060 17484
rect 22020 16153 22048 17478
rect 22006 16144 22062 16153
rect 21824 16108 21876 16114
rect 22006 16079 22062 16088
rect 21824 16050 21876 16056
rect 21916 16040 21968 16046
rect 21916 15982 21968 15988
rect 21824 14816 21876 14822
rect 21824 14758 21876 14764
rect 21456 14408 21508 14414
rect 21732 14408 21784 14414
rect 21508 14368 21588 14396
rect 21456 14350 21508 14356
rect 21456 14068 21508 14074
rect 21456 14010 21508 14016
rect 21468 13530 21496 14010
rect 21456 13524 21508 13530
rect 21456 13466 21508 13472
rect 21560 13394 21588 14368
rect 21732 14350 21784 14356
rect 21640 13932 21692 13938
rect 21640 13874 21692 13880
rect 21548 13388 21600 13394
rect 21548 13330 21600 13336
rect 21364 12912 21416 12918
rect 21270 12880 21326 12889
rect 21364 12854 21416 12860
rect 21270 12815 21272 12824
rect 21324 12815 21326 12824
rect 21272 12786 21324 12792
rect 21192 12668 21312 12696
rect 20916 12600 21220 12628
rect 20833 12540 21141 12549
rect 20833 12538 20839 12540
rect 20895 12538 20919 12540
rect 20975 12538 20999 12540
rect 21055 12538 21079 12540
rect 21135 12538 21141 12540
rect 20895 12486 20897 12538
rect 21077 12486 21079 12538
rect 20833 12484 20839 12486
rect 20895 12484 20919 12486
rect 20975 12484 20999 12486
rect 21055 12484 21079 12486
rect 21135 12484 21141 12486
rect 20833 12475 21141 12484
rect 20732 12406 21128 12434
rect 20812 12232 20864 12238
rect 20640 12192 20812 12220
rect 20732 10606 20760 12192
rect 20812 12174 20864 12180
rect 21100 11608 21128 12406
rect 21192 12102 21220 12600
rect 21284 12374 21312 12668
rect 21272 12368 21324 12374
rect 21272 12310 21324 12316
rect 21272 12164 21324 12170
rect 21272 12106 21324 12112
rect 21180 12096 21232 12102
rect 21180 12038 21232 12044
rect 21284 11744 21312 12106
rect 21376 11898 21404 12854
rect 21652 12374 21680 13874
rect 21744 12918 21772 14350
rect 21836 13802 21864 14758
rect 21824 13796 21876 13802
rect 21824 13738 21876 13744
rect 21732 12912 21784 12918
rect 21732 12854 21784 12860
rect 21640 12368 21692 12374
rect 21640 12310 21692 12316
rect 21640 12232 21692 12238
rect 21546 12200 21602 12209
rect 21640 12174 21692 12180
rect 21546 12135 21548 12144
rect 21600 12135 21602 12144
rect 21548 12106 21600 12112
rect 21456 12096 21508 12102
rect 21456 12038 21508 12044
rect 21364 11892 21416 11898
rect 21364 11834 21416 11840
rect 21364 11756 21416 11762
rect 21284 11716 21364 11744
rect 21364 11698 21416 11704
rect 21100 11580 21312 11608
rect 20833 11452 21141 11461
rect 20833 11450 20839 11452
rect 20895 11450 20919 11452
rect 20975 11450 20999 11452
rect 21055 11450 21079 11452
rect 21135 11450 21141 11452
rect 20895 11398 20897 11450
rect 21077 11398 21079 11450
rect 20833 11396 20839 11398
rect 20895 11396 20919 11398
rect 20975 11396 20999 11398
rect 21055 11396 21079 11398
rect 21135 11396 21141 11398
rect 20833 11387 21141 11396
rect 21180 11280 21232 11286
rect 21178 11248 21180 11257
rect 21232 11248 21234 11257
rect 21178 11183 21234 11192
rect 20536 10600 20588 10606
rect 20536 10542 20588 10548
rect 20720 10600 20772 10606
rect 20720 10542 20772 10548
rect 20444 10124 20496 10130
rect 20444 10066 20496 10072
rect 20352 10056 20404 10062
rect 20352 9998 20404 10004
rect 20260 9580 20312 9586
rect 20260 9522 20312 9528
rect 20260 8900 20312 8906
rect 20260 8842 20312 8848
rect 20168 7948 20220 7954
rect 20168 7890 20220 7896
rect 20076 7812 20128 7818
rect 20076 7754 20128 7760
rect 19984 7744 20036 7750
rect 19984 7686 20036 7692
rect 19524 7404 19576 7410
rect 19524 7346 19576 7352
rect 19800 7404 19852 7410
rect 19800 7346 19852 7352
rect 19536 6866 19564 7346
rect 19524 6860 19576 6866
rect 19524 6802 19576 6808
rect 19352 6310 19472 6338
rect 19248 5840 19300 5846
rect 19248 5782 19300 5788
rect 18788 5636 18840 5642
rect 18788 5578 18840 5584
rect 18800 5370 18828 5578
rect 18788 5364 18840 5370
rect 18788 5306 18840 5312
rect 18880 5092 18932 5098
rect 18880 5034 18932 5040
rect 18696 5024 18748 5030
rect 18696 4966 18748 4972
rect 18708 4826 18736 4966
rect 18696 4820 18748 4826
rect 18696 4762 18748 4768
rect 18604 4480 18656 4486
rect 18604 4422 18656 4428
rect 18380 4236 18460 4264
rect 18512 4276 18564 4282
rect 18328 4218 18380 4224
rect 18512 4218 18564 4224
rect 18052 4140 18104 4146
rect 18052 4082 18104 4088
rect 17868 4004 17920 4010
rect 17868 3946 17920 3952
rect 18064 3534 18092 4082
rect 18512 4072 18564 4078
rect 18512 4014 18564 4020
rect 18144 3732 18196 3738
rect 18144 3674 18196 3680
rect 18156 3602 18184 3674
rect 18144 3596 18196 3602
rect 18144 3538 18196 3544
rect 18524 3534 18552 4014
rect 18052 3528 18104 3534
rect 18052 3470 18104 3476
rect 18236 3528 18288 3534
rect 18236 3470 18288 3476
rect 18512 3528 18564 3534
rect 18512 3470 18564 3476
rect 17868 3460 17920 3466
rect 17868 3402 17920 3408
rect 17880 3126 17908 3402
rect 18248 3380 18276 3470
rect 18248 3352 18368 3380
rect 17992 3292 18300 3301
rect 17992 3290 17998 3292
rect 18054 3290 18078 3292
rect 18134 3290 18158 3292
rect 18214 3290 18238 3292
rect 18294 3290 18300 3292
rect 18054 3238 18056 3290
rect 18236 3238 18238 3290
rect 17992 3236 17998 3238
rect 18054 3236 18078 3238
rect 18134 3236 18158 3238
rect 18214 3236 18238 3238
rect 18294 3236 18300 3238
rect 17992 3227 18300 3236
rect 18340 3194 18368 3352
rect 18328 3188 18380 3194
rect 18328 3130 18380 3136
rect 18616 3126 18644 4422
rect 18892 4214 18920 5034
rect 18880 4208 18932 4214
rect 18880 4150 18932 4156
rect 18696 3936 18748 3942
rect 18696 3878 18748 3884
rect 18708 3602 18736 3878
rect 18788 3664 18840 3670
rect 18788 3606 18840 3612
rect 18696 3596 18748 3602
rect 18696 3538 18748 3544
rect 18800 3534 18828 3606
rect 18788 3528 18840 3534
rect 18788 3470 18840 3476
rect 18892 3466 18920 4150
rect 19064 4140 19116 4146
rect 19064 4082 19116 4088
rect 18880 3460 18932 3466
rect 18880 3402 18932 3408
rect 17868 3120 17920 3126
rect 17868 3062 17920 3068
rect 18604 3120 18656 3126
rect 18604 3062 18656 3068
rect 17038 3023 17040 3032
rect 17092 3023 17094 3032
rect 17316 3052 17368 3058
rect 17040 2994 17092 3000
rect 17316 2994 17368 3000
rect 15752 2848 15804 2854
rect 15752 2790 15804 2796
rect 15152 2748 15460 2757
rect 15152 2746 15158 2748
rect 15214 2746 15238 2748
rect 15294 2746 15318 2748
rect 15374 2746 15398 2748
rect 15454 2746 15460 2748
rect 15214 2694 15216 2746
rect 15396 2694 15398 2746
rect 15152 2692 15158 2694
rect 15214 2692 15238 2694
rect 15294 2692 15318 2694
rect 15374 2692 15398 2694
rect 15454 2692 15460 2694
rect 15152 2683 15460 2692
rect 17328 2650 17356 2994
rect 17592 2916 17644 2922
rect 17592 2858 17644 2864
rect 12348 2644 12400 2650
rect 12348 2586 12400 2592
rect 14464 2644 14516 2650
rect 14464 2586 14516 2592
rect 17316 2644 17368 2650
rect 17316 2586 17368 2592
rect 16304 2508 16356 2514
rect 16304 2450 16356 2456
rect 9220 2440 9272 2446
rect 9220 2382 9272 2388
rect 9864 2440 9916 2446
rect 9864 2382 9916 2388
rect 10508 2440 10560 2446
rect 10508 2382 10560 2388
rect 11152 2440 11204 2446
rect 11152 2382 11204 2388
rect 11796 2440 11848 2446
rect 11796 2382 11848 2388
rect 12716 2440 12768 2446
rect 12716 2382 12768 2388
rect 13084 2440 13136 2446
rect 13084 2382 13136 2388
rect 13728 2440 13780 2446
rect 13728 2382 13780 2388
rect 14372 2440 14424 2446
rect 14372 2382 14424 2388
rect 15016 2440 15068 2446
rect 15016 2382 15068 2388
rect 15660 2440 15712 2446
rect 15660 2382 15712 2388
rect 9232 800 9260 2382
rect 9876 800 9904 2382
rect 10520 800 10548 2382
rect 11164 800 11192 2382
rect 11808 800 11836 2382
rect 12311 2204 12619 2213
rect 12311 2202 12317 2204
rect 12373 2202 12397 2204
rect 12453 2202 12477 2204
rect 12533 2202 12557 2204
rect 12613 2202 12619 2204
rect 12373 2150 12375 2202
rect 12555 2150 12557 2202
rect 12311 2148 12317 2150
rect 12373 2148 12397 2150
rect 12453 2148 12477 2150
rect 12533 2148 12557 2150
rect 12613 2148 12619 2150
rect 12311 2139 12619 2148
rect 12452 870 12572 898
rect 12452 800 12480 870
rect 3712 734 4016 762
rect 4066 0 4122 800
rect 4710 0 4766 800
rect 5354 0 5410 800
rect 5998 0 6054 800
rect 6642 0 6698 800
rect 7286 0 7342 800
rect 7930 0 7986 800
rect 8574 0 8630 800
rect 9218 0 9274 800
rect 9862 0 9918 800
rect 10506 0 10562 800
rect 11150 0 11206 800
rect 11794 0 11850 800
rect 12438 0 12494 800
rect 12544 762 12572 870
rect 12728 762 12756 2382
rect 13096 800 13124 2382
rect 13740 800 13768 2382
rect 14384 800 14412 2382
rect 15028 800 15056 2382
rect 15672 800 15700 2382
rect 16316 800 16344 2450
rect 16948 2440 17000 2446
rect 16948 2382 17000 2388
rect 16960 800 16988 2382
rect 17604 800 17632 2858
rect 18328 2848 18380 2854
rect 18328 2790 18380 2796
rect 17992 2204 18300 2213
rect 17992 2202 17998 2204
rect 18054 2202 18078 2204
rect 18134 2202 18158 2204
rect 18214 2202 18238 2204
rect 18294 2202 18300 2204
rect 18054 2150 18056 2202
rect 18236 2150 18238 2202
rect 17992 2148 17998 2150
rect 18054 2148 18078 2150
rect 18134 2148 18158 2150
rect 18214 2148 18238 2150
rect 18294 2148 18300 2150
rect 17992 2139 18300 2148
rect 18340 1442 18368 2790
rect 18616 2650 18644 3062
rect 18696 3052 18748 3058
rect 18696 2994 18748 3000
rect 18708 2961 18736 2994
rect 19076 2990 19104 4082
rect 19352 3670 19380 6310
rect 19812 6304 19840 7346
rect 20272 7342 20300 8842
rect 20364 8566 20392 9998
rect 20732 9586 20760 10542
rect 20833 10364 21141 10373
rect 20833 10362 20839 10364
rect 20895 10362 20919 10364
rect 20975 10362 20999 10364
rect 21055 10362 21079 10364
rect 21135 10362 21141 10364
rect 20895 10310 20897 10362
rect 21077 10310 21079 10362
rect 20833 10308 20839 10310
rect 20895 10308 20919 10310
rect 20975 10308 20999 10310
rect 21055 10308 21079 10310
rect 21135 10308 21141 10310
rect 20833 10299 21141 10308
rect 21192 10062 21220 11183
rect 21180 10056 21232 10062
rect 21180 9998 21232 10004
rect 21192 9674 21220 9998
rect 21100 9646 21220 9674
rect 20628 9580 20680 9586
rect 20628 9522 20680 9528
rect 20720 9580 20772 9586
rect 20720 9522 20772 9528
rect 20352 8560 20404 8566
rect 20352 8502 20404 8508
rect 20640 8362 20668 9522
rect 20720 9444 20772 9450
rect 20720 9386 20772 9392
rect 20732 8566 20760 9386
rect 21100 9382 21128 9646
rect 21180 9580 21232 9586
rect 21180 9522 21232 9528
rect 21088 9376 21140 9382
rect 21088 9318 21140 9324
rect 20833 9276 21141 9285
rect 20833 9274 20839 9276
rect 20895 9274 20919 9276
rect 20975 9274 20999 9276
rect 21055 9274 21079 9276
rect 21135 9274 21141 9276
rect 20895 9222 20897 9274
rect 21077 9222 21079 9274
rect 20833 9220 20839 9222
rect 20895 9220 20919 9222
rect 20975 9220 20999 9222
rect 21055 9220 21079 9222
rect 21135 9220 21141 9222
rect 20833 9211 21141 9220
rect 21192 8974 21220 9522
rect 21180 8968 21232 8974
rect 21180 8910 21232 8916
rect 20720 8560 20772 8566
rect 20720 8502 20772 8508
rect 20720 8424 20772 8430
rect 20720 8366 20772 8372
rect 20628 8356 20680 8362
rect 20628 8298 20680 8304
rect 20628 7812 20680 7818
rect 20628 7754 20680 7760
rect 20640 7410 20668 7754
rect 20628 7404 20680 7410
rect 20628 7346 20680 7352
rect 20260 7336 20312 7342
rect 20260 7278 20312 7284
rect 19892 6316 19944 6322
rect 19812 6276 19892 6304
rect 19892 6258 19944 6264
rect 20536 6316 20588 6322
rect 20536 6258 20588 6264
rect 20352 6248 20404 6254
rect 20352 6190 20404 6196
rect 19616 6112 19668 6118
rect 19616 6054 19668 6060
rect 19432 5568 19484 5574
rect 19432 5510 19484 5516
rect 19444 5234 19472 5510
rect 19628 5302 19656 6054
rect 20364 5914 20392 6190
rect 20352 5908 20404 5914
rect 20352 5850 20404 5856
rect 20364 5574 20392 5850
rect 20444 5704 20496 5710
rect 20444 5646 20496 5652
rect 20352 5568 20404 5574
rect 20352 5510 20404 5516
rect 19524 5296 19576 5302
rect 19524 5238 19576 5244
rect 19616 5296 19668 5302
rect 19616 5238 19668 5244
rect 19432 5228 19484 5234
rect 19432 5170 19484 5176
rect 19432 5024 19484 5030
rect 19432 4966 19484 4972
rect 19444 4622 19472 4966
rect 19432 4616 19484 4622
rect 19432 4558 19484 4564
rect 19340 3664 19392 3670
rect 19340 3606 19392 3612
rect 19536 3194 19564 5238
rect 20168 5024 20220 5030
rect 20168 4966 20220 4972
rect 20180 4146 20208 4966
rect 20456 4622 20484 5646
rect 20548 4826 20576 6258
rect 20640 5778 20668 7346
rect 20732 6390 20760 8366
rect 20833 8188 21141 8197
rect 20833 8186 20839 8188
rect 20895 8186 20919 8188
rect 20975 8186 20999 8188
rect 21055 8186 21079 8188
rect 21135 8186 21141 8188
rect 20895 8134 20897 8186
rect 21077 8134 21079 8186
rect 20833 8132 20839 8134
rect 20895 8132 20919 8134
rect 20975 8132 20999 8134
rect 21055 8132 21079 8134
rect 21135 8132 21141 8134
rect 20833 8123 21141 8132
rect 21284 8022 21312 11580
rect 21376 11014 21404 11698
rect 21468 11150 21496 12038
rect 21456 11144 21508 11150
rect 21456 11086 21508 11092
rect 21364 11008 21416 11014
rect 21364 10950 21416 10956
rect 21652 10810 21680 12174
rect 21744 11762 21772 12854
rect 21732 11756 21784 11762
rect 21732 11698 21784 11704
rect 21732 11008 21784 11014
rect 21732 10950 21784 10956
rect 21640 10804 21692 10810
rect 21640 10746 21692 10752
rect 21548 10668 21600 10674
rect 21548 10610 21600 10616
rect 21560 10470 21588 10610
rect 21548 10464 21600 10470
rect 21548 10406 21600 10412
rect 21560 10062 21588 10406
rect 21548 10056 21600 10062
rect 21548 9998 21600 10004
rect 21456 9920 21508 9926
rect 21456 9862 21508 9868
rect 21364 9376 21416 9382
rect 21364 9318 21416 9324
rect 21376 9178 21404 9318
rect 21364 9172 21416 9178
rect 21364 9114 21416 9120
rect 21468 8974 21496 9862
rect 21548 9648 21600 9654
rect 21548 9590 21600 9596
rect 21364 8968 21416 8974
rect 21364 8910 21416 8916
rect 21456 8968 21508 8974
rect 21456 8910 21508 8916
rect 21272 8016 21324 8022
rect 21272 7958 21324 7964
rect 21180 7336 21232 7342
rect 21180 7278 21232 7284
rect 20833 7100 21141 7109
rect 20833 7098 20839 7100
rect 20895 7098 20919 7100
rect 20975 7098 20999 7100
rect 21055 7098 21079 7100
rect 21135 7098 21141 7100
rect 20895 7046 20897 7098
rect 21077 7046 21079 7098
rect 20833 7044 20839 7046
rect 20895 7044 20919 7046
rect 20975 7044 20999 7046
rect 21055 7044 21079 7046
rect 21135 7044 21141 7046
rect 20833 7035 21141 7044
rect 20720 6384 20772 6390
rect 20720 6326 20772 6332
rect 20833 6012 21141 6021
rect 20833 6010 20839 6012
rect 20895 6010 20919 6012
rect 20975 6010 20999 6012
rect 21055 6010 21079 6012
rect 21135 6010 21141 6012
rect 20895 5958 20897 6010
rect 21077 5958 21079 6010
rect 20833 5956 20839 5958
rect 20895 5956 20919 5958
rect 20975 5956 20999 5958
rect 21055 5956 21079 5958
rect 21135 5956 21141 5958
rect 20833 5947 21141 5956
rect 21192 5846 21220 7278
rect 21284 6798 21312 7958
rect 21272 6792 21324 6798
rect 21272 6734 21324 6740
rect 21376 6458 21404 8910
rect 21560 8498 21588 9590
rect 21652 9586 21680 10746
rect 21640 9580 21692 9586
rect 21640 9522 21692 9528
rect 21744 8566 21772 10950
rect 21732 8560 21784 8566
rect 21732 8502 21784 8508
rect 21548 8492 21600 8498
rect 21548 8434 21600 8440
rect 21640 8492 21692 8498
rect 21640 8434 21692 8440
rect 21560 8090 21588 8434
rect 21548 8084 21600 8090
rect 21548 8026 21600 8032
rect 21456 7880 21508 7886
rect 21456 7822 21508 7828
rect 21364 6452 21416 6458
rect 21364 6394 21416 6400
rect 21468 6338 21496 7822
rect 21546 6896 21602 6905
rect 21546 6831 21548 6840
rect 21600 6831 21602 6840
rect 21548 6802 21600 6808
rect 21560 6390 21588 6802
rect 21376 6310 21496 6338
rect 21548 6384 21600 6390
rect 21548 6326 21600 6332
rect 21180 5840 21232 5846
rect 21180 5782 21232 5788
rect 20628 5772 20680 5778
rect 20628 5714 20680 5720
rect 21192 5692 21220 5782
rect 21272 5704 21324 5710
rect 21192 5664 21272 5692
rect 21272 5646 21324 5652
rect 21376 5370 21404 6310
rect 21652 5914 21680 8434
rect 21836 8090 21864 13738
rect 21928 9654 21956 15982
rect 22020 15706 22048 16079
rect 22112 16017 22140 18566
rect 22204 18426 22232 20402
rect 23673 19612 23981 19621
rect 23673 19610 23679 19612
rect 23735 19610 23759 19612
rect 23815 19610 23839 19612
rect 23895 19610 23919 19612
rect 23975 19610 23981 19612
rect 23735 19558 23737 19610
rect 23917 19558 23919 19610
rect 23673 19556 23679 19558
rect 23735 19556 23759 19558
rect 23815 19556 23839 19558
rect 23895 19556 23919 19558
rect 23975 19556 23981 19558
rect 23673 19547 23981 19556
rect 22376 19236 22428 19242
rect 22376 19178 22428 19184
rect 22388 18970 22416 19178
rect 22376 18964 22428 18970
rect 22376 18906 22428 18912
rect 22388 18426 22416 18906
rect 23673 18524 23981 18533
rect 23673 18522 23679 18524
rect 23735 18522 23759 18524
rect 23815 18522 23839 18524
rect 23895 18522 23919 18524
rect 23975 18522 23981 18524
rect 23735 18470 23737 18522
rect 23917 18470 23919 18522
rect 23673 18468 23679 18470
rect 23735 18468 23759 18470
rect 23815 18468 23839 18470
rect 23895 18468 23919 18470
rect 23975 18468 23981 18470
rect 23673 18459 23981 18468
rect 22192 18420 22244 18426
rect 22192 18362 22244 18368
rect 22376 18420 22428 18426
rect 22376 18362 22428 18368
rect 22284 18284 22336 18290
rect 22284 18226 22336 18232
rect 22468 18284 22520 18290
rect 22468 18226 22520 18232
rect 22652 18284 22704 18290
rect 22652 18226 22704 18232
rect 22296 17202 22324 18226
rect 22284 17196 22336 17202
rect 22284 17138 22336 17144
rect 22296 16726 22324 17138
rect 22376 17128 22428 17134
rect 22376 17070 22428 17076
rect 22388 16794 22416 17070
rect 22376 16788 22428 16794
rect 22376 16730 22428 16736
rect 22284 16720 22336 16726
rect 22284 16662 22336 16668
rect 22284 16448 22336 16454
rect 22284 16390 22336 16396
rect 22098 16008 22154 16017
rect 22098 15943 22154 15952
rect 22008 15700 22060 15706
rect 22060 15660 22140 15688
rect 22008 15642 22060 15648
rect 22112 15026 22140 15660
rect 22296 15026 22324 16390
rect 22480 15162 22508 18226
rect 22664 17882 22692 18226
rect 22652 17876 22704 17882
rect 22652 17818 22704 17824
rect 23673 17436 23981 17445
rect 23673 17434 23679 17436
rect 23735 17434 23759 17436
rect 23815 17434 23839 17436
rect 23895 17434 23919 17436
rect 23975 17434 23981 17436
rect 23735 17382 23737 17434
rect 23917 17382 23919 17434
rect 23673 17380 23679 17382
rect 23735 17380 23759 17382
rect 23815 17380 23839 17382
rect 23895 17380 23919 17382
rect 23975 17380 23981 17382
rect 23673 17371 23981 17380
rect 22744 16992 22796 16998
rect 22744 16934 22796 16940
rect 22560 16040 22612 16046
rect 22560 15982 22612 15988
rect 22572 15638 22600 15982
rect 22652 15904 22704 15910
rect 22652 15846 22704 15852
rect 22560 15632 22612 15638
rect 22560 15574 22612 15580
rect 22468 15156 22520 15162
rect 22468 15098 22520 15104
rect 22008 15020 22060 15026
rect 22008 14962 22060 14968
rect 22100 15020 22152 15026
rect 22100 14962 22152 14968
rect 22284 15020 22336 15026
rect 22336 14980 22416 15008
rect 22284 14962 22336 14968
rect 22020 14396 22048 14962
rect 22284 14884 22336 14890
rect 22284 14826 22336 14832
rect 22100 14408 22152 14414
rect 22020 14368 22100 14396
rect 22100 14350 22152 14356
rect 22112 13394 22140 14350
rect 22296 13938 22324 14826
rect 22284 13932 22336 13938
rect 22284 13874 22336 13880
rect 22296 13734 22324 13874
rect 22284 13728 22336 13734
rect 22284 13670 22336 13676
rect 22282 13424 22338 13433
rect 22100 13388 22152 13394
rect 22282 13359 22338 13368
rect 22100 13330 22152 13336
rect 22112 12782 22140 13330
rect 22296 12986 22324 13359
rect 22284 12980 22336 12986
rect 22284 12922 22336 12928
rect 22100 12776 22152 12782
rect 22100 12718 22152 12724
rect 22008 12232 22060 12238
rect 22112 12220 22140 12718
rect 22388 12434 22416 14980
rect 22468 14272 22520 14278
rect 22468 14214 22520 14220
rect 22480 13326 22508 14214
rect 22572 13938 22600 15574
rect 22664 15502 22692 15846
rect 22756 15706 22784 16934
rect 23296 16516 23348 16522
rect 23296 16458 23348 16464
rect 22744 15700 22796 15706
rect 22744 15642 22796 15648
rect 22652 15496 22704 15502
rect 22652 15438 22704 15444
rect 22756 14006 22784 15642
rect 23020 15496 23072 15502
rect 23020 15438 23072 15444
rect 22836 15020 22888 15026
rect 22836 14962 22888 14968
rect 22848 14414 22876 14962
rect 22836 14408 22888 14414
rect 22836 14350 22888 14356
rect 22744 14000 22796 14006
rect 22664 13960 22744 13988
rect 22560 13932 22612 13938
rect 22560 13874 22612 13880
rect 22572 13841 22600 13874
rect 22558 13832 22614 13841
rect 22558 13767 22614 13776
rect 22664 13682 22692 13960
rect 22744 13942 22796 13948
rect 22572 13654 22692 13682
rect 22468 13320 22520 13326
rect 22468 13262 22520 13268
rect 22388 12406 22508 12434
rect 22284 12300 22336 12306
rect 22284 12242 22336 12248
rect 22192 12232 22244 12238
rect 22112 12192 22192 12220
rect 22008 12174 22060 12180
rect 22192 12174 22244 12180
rect 22020 10198 22048 12174
rect 22100 11756 22152 11762
rect 22100 11698 22152 11704
rect 22112 10266 22140 11698
rect 22100 10260 22152 10266
rect 22100 10202 22152 10208
rect 22008 10192 22060 10198
rect 22008 10134 22060 10140
rect 22204 10130 22232 12174
rect 22296 11354 22324 12242
rect 22376 12164 22428 12170
rect 22376 12106 22428 12112
rect 22284 11348 22336 11354
rect 22284 11290 22336 11296
rect 22388 10470 22416 12106
rect 22480 10606 22508 12406
rect 22572 10810 22600 13654
rect 22742 13288 22798 13297
rect 22742 13223 22798 13232
rect 22652 13184 22704 13190
rect 22652 13126 22704 13132
rect 22664 12850 22692 13126
rect 22756 12918 22784 13223
rect 22744 12912 22796 12918
rect 22744 12854 22796 12860
rect 22652 12844 22704 12850
rect 22652 12786 22704 12792
rect 22664 12170 22692 12786
rect 22744 12640 22796 12646
rect 22744 12582 22796 12588
rect 22652 12164 22704 12170
rect 22652 12106 22704 12112
rect 22652 11688 22704 11694
rect 22652 11630 22704 11636
rect 22664 11082 22692 11630
rect 22652 11076 22704 11082
rect 22652 11018 22704 11024
rect 22560 10804 22612 10810
rect 22560 10746 22612 10752
rect 22650 10704 22706 10713
rect 22650 10639 22652 10648
rect 22704 10639 22706 10648
rect 22652 10610 22704 10616
rect 22468 10600 22520 10606
rect 22468 10542 22520 10548
rect 22376 10464 22428 10470
rect 22376 10406 22428 10412
rect 22192 10124 22244 10130
rect 22192 10066 22244 10072
rect 22100 10056 22152 10062
rect 22100 9998 22152 10004
rect 21916 9648 21968 9654
rect 21916 9590 21968 9596
rect 22008 9172 22060 9178
rect 22008 9114 22060 9120
rect 21916 8968 21968 8974
rect 21916 8910 21968 8916
rect 21824 8084 21876 8090
rect 21824 8026 21876 8032
rect 21928 6662 21956 8910
rect 22020 7886 22048 9114
rect 22008 7880 22060 7886
rect 22008 7822 22060 7828
rect 22112 7274 22140 9998
rect 22204 9568 22232 10066
rect 22284 9580 22336 9586
rect 22204 9540 22284 9568
rect 22284 9522 22336 9528
rect 22388 9450 22416 10406
rect 22376 9444 22428 9450
rect 22376 9386 22428 9392
rect 22192 9376 22244 9382
rect 22192 9318 22244 9324
rect 22204 8838 22232 9318
rect 22376 9036 22428 9042
rect 22376 8978 22428 8984
rect 22192 8832 22244 8838
rect 22192 8774 22244 8780
rect 22100 7268 22152 7274
rect 22100 7210 22152 7216
rect 22204 7154 22232 8774
rect 22282 8392 22338 8401
rect 22282 8327 22284 8336
rect 22336 8327 22338 8336
rect 22284 8298 22336 8304
rect 22388 8242 22416 8978
rect 22480 8378 22508 10542
rect 22560 10464 22612 10470
rect 22560 10406 22612 10412
rect 22572 8498 22600 10406
rect 22664 9926 22692 10610
rect 22756 10198 22784 12582
rect 22848 12374 22876 14350
rect 22928 14272 22980 14278
rect 22928 14214 22980 14220
rect 22940 13258 22968 14214
rect 23032 13818 23060 15438
rect 23112 14816 23164 14822
rect 23112 14758 23164 14764
rect 23124 13938 23152 14758
rect 23112 13932 23164 13938
rect 23112 13874 23164 13880
rect 23032 13790 23152 13818
rect 23124 13258 23152 13790
rect 22928 13252 22980 13258
rect 22928 13194 22980 13200
rect 23112 13252 23164 13258
rect 23112 13194 23164 13200
rect 22940 12850 22968 13194
rect 22928 12844 22980 12850
rect 22928 12786 22980 12792
rect 22836 12368 22888 12374
rect 22836 12310 22888 12316
rect 22940 12306 22968 12786
rect 23020 12708 23072 12714
rect 23020 12650 23072 12656
rect 22928 12300 22980 12306
rect 22928 12242 22980 12248
rect 23032 11898 23060 12650
rect 23124 12434 23152 13194
rect 23124 12406 23244 12434
rect 23216 12238 23244 12406
rect 23204 12232 23256 12238
rect 23204 12174 23256 12180
rect 23020 11892 23072 11898
rect 23020 11834 23072 11840
rect 22928 11824 22980 11830
rect 22928 11766 22980 11772
rect 22836 10736 22888 10742
rect 22836 10678 22888 10684
rect 22744 10192 22796 10198
rect 22744 10134 22796 10140
rect 22652 9920 22704 9926
rect 22652 9862 22704 9868
rect 22664 9450 22692 9862
rect 22652 9444 22704 9450
rect 22652 9386 22704 9392
rect 22744 9376 22796 9382
rect 22744 9318 22796 9324
rect 22560 8492 22612 8498
rect 22560 8434 22612 8440
rect 22756 8430 22784 9318
rect 22848 9178 22876 10678
rect 22940 10044 22968 11766
rect 23020 11756 23072 11762
rect 23020 11698 23072 11704
rect 23112 11756 23164 11762
rect 23112 11698 23164 11704
rect 23032 11218 23060 11698
rect 23020 11212 23072 11218
rect 23020 11154 23072 11160
rect 23032 10690 23060 11154
rect 23124 10810 23152 11698
rect 23112 10804 23164 10810
rect 23112 10746 23164 10752
rect 23032 10662 23152 10690
rect 23020 10056 23072 10062
rect 22940 10016 23020 10044
rect 23020 9998 23072 10004
rect 22928 9512 22980 9518
rect 22928 9454 22980 9460
rect 22836 9172 22888 9178
rect 22836 9114 22888 9120
rect 22836 8492 22888 8498
rect 22836 8434 22888 8440
rect 22744 8424 22796 8430
rect 22480 8350 22600 8378
rect 22744 8366 22796 8372
rect 22296 8214 22416 8242
rect 22296 8022 22324 8214
rect 22284 8016 22336 8022
rect 22284 7958 22336 7964
rect 22296 7342 22324 7958
rect 22376 7948 22428 7954
rect 22376 7890 22428 7896
rect 22284 7336 22336 7342
rect 22284 7278 22336 7284
rect 22112 7126 22232 7154
rect 21916 6656 21968 6662
rect 21916 6598 21968 6604
rect 21824 6316 21876 6322
rect 21824 6258 21876 6264
rect 21640 5908 21692 5914
rect 21640 5850 21692 5856
rect 21456 5704 21508 5710
rect 21456 5646 21508 5652
rect 21364 5364 21416 5370
rect 21364 5306 21416 5312
rect 20833 4924 21141 4933
rect 20833 4922 20839 4924
rect 20895 4922 20919 4924
rect 20975 4922 20999 4924
rect 21055 4922 21079 4924
rect 21135 4922 21141 4924
rect 20895 4870 20897 4922
rect 21077 4870 21079 4922
rect 20833 4868 20839 4870
rect 20895 4868 20919 4870
rect 20975 4868 20999 4870
rect 21055 4868 21079 4870
rect 21135 4868 21141 4870
rect 20833 4859 21141 4868
rect 20536 4820 20588 4826
rect 20536 4762 20588 4768
rect 21468 4758 21496 5646
rect 21456 4752 21508 4758
rect 21456 4694 21508 4700
rect 20444 4616 20496 4622
rect 20444 4558 20496 4564
rect 20812 4548 20864 4554
rect 20812 4490 20864 4496
rect 20824 4146 20852 4490
rect 19984 4140 20036 4146
rect 19984 4082 20036 4088
rect 20168 4140 20220 4146
rect 20168 4082 20220 4088
rect 20352 4140 20404 4146
rect 20352 4082 20404 4088
rect 20536 4140 20588 4146
rect 20536 4082 20588 4088
rect 20812 4140 20864 4146
rect 20812 4082 20864 4088
rect 21180 4140 21232 4146
rect 21180 4082 21232 4088
rect 19996 3534 20024 4082
rect 20180 3534 20208 4082
rect 20364 3534 20392 4082
rect 20548 3602 20576 4082
rect 20833 3836 21141 3845
rect 20833 3834 20839 3836
rect 20895 3834 20919 3836
rect 20975 3834 20999 3836
rect 21055 3834 21079 3836
rect 21135 3834 21141 3836
rect 20895 3782 20897 3834
rect 21077 3782 21079 3834
rect 20833 3780 20839 3782
rect 20895 3780 20919 3782
rect 20975 3780 20999 3782
rect 21055 3780 21079 3782
rect 21135 3780 21141 3782
rect 20833 3771 21141 3780
rect 20536 3596 20588 3602
rect 20536 3538 20588 3544
rect 21192 3534 21220 4082
rect 21836 3738 21864 6258
rect 22112 5370 22140 7126
rect 22192 6724 22244 6730
rect 22192 6666 22244 6672
rect 22204 6322 22232 6666
rect 22192 6316 22244 6322
rect 22192 6258 22244 6264
rect 22204 5778 22232 6258
rect 22192 5772 22244 5778
rect 22192 5714 22244 5720
rect 22100 5364 22152 5370
rect 22100 5306 22152 5312
rect 22098 4720 22154 4729
rect 22098 4655 22100 4664
rect 22152 4655 22154 4664
rect 22100 4626 22152 4632
rect 22296 4570 22324 7278
rect 22388 7206 22416 7890
rect 22468 7744 22520 7750
rect 22468 7686 22520 7692
rect 22480 7410 22508 7686
rect 22468 7404 22520 7410
rect 22468 7346 22520 7352
rect 22376 7200 22428 7206
rect 22376 7142 22428 7148
rect 22388 6322 22416 7142
rect 22376 6316 22428 6322
rect 22376 6258 22428 6264
rect 22388 5914 22416 6258
rect 22376 5908 22428 5914
rect 22376 5850 22428 5856
rect 22376 5568 22428 5574
rect 22376 5510 22428 5516
rect 22388 4690 22416 5510
rect 22376 4684 22428 4690
rect 22376 4626 22428 4632
rect 22296 4542 22416 4570
rect 22388 3942 22416 4542
rect 22480 4146 22508 7346
rect 22572 5302 22600 8350
rect 22848 7546 22876 8434
rect 22940 7818 22968 9454
rect 23032 7886 23060 9998
rect 23124 9654 23152 10662
rect 23216 9926 23244 12174
rect 23308 11830 23336 16458
rect 23673 16348 23981 16357
rect 23673 16346 23679 16348
rect 23735 16346 23759 16348
rect 23815 16346 23839 16348
rect 23895 16346 23919 16348
rect 23975 16346 23981 16348
rect 23735 16294 23737 16346
rect 23917 16294 23919 16346
rect 23673 16292 23679 16294
rect 23735 16292 23759 16294
rect 23815 16292 23839 16294
rect 23895 16292 23919 16294
rect 23975 16292 23981 16294
rect 23673 16283 23981 16292
rect 23673 15260 23981 15269
rect 23673 15258 23679 15260
rect 23735 15258 23759 15260
rect 23815 15258 23839 15260
rect 23895 15258 23919 15260
rect 23975 15258 23981 15260
rect 23735 15206 23737 15258
rect 23917 15206 23919 15258
rect 23673 15204 23679 15206
rect 23735 15204 23759 15206
rect 23815 15204 23839 15206
rect 23895 15204 23919 15206
rect 23975 15204 23981 15206
rect 23673 15195 23981 15204
rect 23673 14172 23981 14181
rect 23673 14170 23679 14172
rect 23735 14170 23759 14172
rect 23815 14170 23839 14172
rect 23895 14170 23919 14172
rect 23975 14170 23981 14172
rect 23735 14118 23737 14170
rect 23917 14118 23919 14170
rect 23673 14116 23679 14118
rect 23735 14116 23759 14118
rect 23815 14116 23839 14118
rect 23895 14116 23919 14118
rect 23975 14116 23981 14118
rect 23673 14107 23981 14116
rect 23388 13796 23440 13802
rect 23388 13738 23440 13744
rect 23296 11824 23348 11830
rect 23296 11766 23348 11772
rect 23400 11286 23428 13738
rect 23673 13084 23981 13093
rect 23673 13082 23679 13084
rect 23735 13082 23759 13084
rect 23815 13082 23839 13084
rect 23895 13082 23919 13084
rect 23975 13082 23981 13084
rect 23735 13030 23737 13082
rect 23917 13030 23919 13082
rect 23673 13028 23679 13030
rect 23735 13028 23759 13030
rect 23815 13028 23839 13030
rect 23895 13028 23919 13030
rect 23975 13028 23981 13030
rect 23673 13019 23981 13028
rect 23673 11996 23981 12005
rect 23673 11994 23679 11996
rect 23735 11994 23759 11996
rect 23815 11994 23839 11996
rect 23895 11994 23919 11996
rect 23975 11994 23981 11996
rect 23735 11942 23737 11994
rect 23917 11942 23919 11994
rect 23673 11940 23679 11942
rect 23735 11940 23759 11942
rect 23815 11940 23839 11942
rect 23895 11940 23919 11942
rect 23975 11940 23981 11942
rect 23673 11931 23981 11940
rect 23388 11280 23440 11286
rect 23388 11222 23440 11228
rect 23296 11076 23348 11082
rect 23296 11018 23348 11024
rect 23204 9920 23256 9926
rect 23204 9862 23256 9868
rect 23216 9722 23244 9862
rect 23204 9716 23256 9722
rect 23204 9658 23256 9664
rect 23112 9648 23164 9654
rect 23308 9602 23336 11018
rect 23673 10908 23981 10917
rect 23673 10906 23679 10908
rect 23735 10906 23759 10908
rect 23815 10906 23839 10908
rect 23895 10906 23919 10908
rect 23975 10906 23981 10908
rect 23735 10854 23737 10906
rect 23917 10854 23919 10906
rect 23673 10852 23679 10854
rect 23735 10852 23759 10854
rect 23815 10852 23839 10854
rect 23895 10852 23919 10854
rect 23975 10852 23981 10854
rect 23673 10843 23981 10852
rect 23673 9820 23981 9829
rect 23673 9818 23679 9820
rect 23735 9818 23759 9820
rect 23815 9818 23839 9820
rect 23895 9818 23919 9820
rect 23975 9818 23981 9820
rect 23735 9766 23737 9818
rect 23917 9766 23919 9818
rect 23673 9764 23679 9766
rect 23735 9764 23759 9766
rect 23815 9764 23839 9766
rect 23895 9764 23919 9766
rect 23975 9764 23981 9766
rect 23673 9755 23981 9764
rect 23112 9590 23164 9596
rect 23124 9042 23152 9590
rect 23216 9574 23336 9602
rect 23112 9036 23164 9042
rect 23112 8978 23164 8984
rect 23216 8838 23244 9574
rect 23204 8832 23256 8838
rect 23204 8774 23256 8780
rect 23216 8634 23244 8774
rect 23673 8732 23981 8741
rect 23673 8730 23679 8732
rect 23735 8730 23759 8732
rect 23815 8730 23839 8732
rect 23895 8730 23919 8732
rect 23975 8730 23981 8732
rect 23735 8678 23737 8730
rect 23917 8678 23919 8730
rect 23673 8676 23679 8678
rect 23735 8676 23759 8678
rect 23815 8676 23839 8678
rect 23895 8676 23919 8678
rect 23975 8676 23981 8678
rect 23673 8667 23981 8676
rect 23204 8628 23256 8634
rect 23204 8570 23256 8576
rect 23020 7880 23072 7886
rect 23020 7822 23072 7828
rect 22928 7812 22980 7818
rect 22928 7754 22980 7760
rect 22836 7540 22888 7546
rect 22836 7482 22888 7488
rect 22940 7410 22968 7754
rect 22928 7404 22980 7410
rect 22928 7346 22980 7352
rect 22652 7200 22704 7206
rect 22652 7142 22704 7148
rect 22664 6798 22692 7142
rect 22940 7002 22968 7346
rect 22928 6996 22980 7002
rect 22928 6938 22980 6944
rect 22652 6792 22704 6798
rect 22652 6734 22704 6740
rect 22940 6458 22968 6938
rect 23032 6934 23060 7822
rect 23020 6928 23072 6934
rect 23020 6870 23072 6876
rect 23216 6866 23244 8570
rect 23673 7644 23981 7653
rect 23673 7642 23679 7644
rect 23735 7642 23759 7644
rect 23815 7642 23839 7644
rect 23895 7642 23919 7644
rect 23975 7642 23981 7644
rect 23735 7590 23737 7642
rect 23917 7590 23919 7642
rect 23673 7588 23679 7590
rect 23735 7588 23759 7590
rect 23815 7588 23839 7590
rect 23895 7588 23919 7590
rect 23975 7588 23981 7590
rect 23673 7579 23981 7588
rect 23204 6860 23256 6866
rect 23204 6802 23256 6808
rect 23673 6556 23981 6565
rect 23673 6554 23679 6556
rect 23735 6554 23759 6556
rect 23815 6554 23839 6556
rect 23895 6554 23919 6556
rect 23975 6554 23981 6556
rect 23735 6502 23737 6554
rect 23917 6502 23919 6554
rect 23673 6500 23679 6502
rect 23735 6500 23759 6502
rect 23815 6500 23839 6502
rect 23895 6500 23919 6502
rect 23975 6500 23981 6502
rect 23673 6491 23981 6500
rect 22928 6452 22980 6458
rect 22928 6394 22980 6400
rect 22928 6316 22980 6322
rect 22928 6258 22980 6264
rect 23112 6316 23164 6322
rect 23112 6258 23164 6264
rect 22940 5778 22968 6258
rect 22928 5772 22980 5778
rect 22928 5714 22980 5720
rect 22940 5302 22968 5714
rect 23124 5710 23152 6258
rect 23112 5704 23164 5710
rect 23112 5646 23164 5652
rect 22560 5296 22612 5302
rect 22560 5238 22612 5244
rect 22928 5296 22980 5302
rect 22928 5238 22980 5244
rect 23124 5234 23152 5646
rect 23673 5468 23981 5477
rect 23673 5466 23679 5468
rect 23735 5466 23759 5468
rect 23815 5466 23839 5468
rect 23895 5466 23919 5468
rect 23975 5466 23981 5468
rect 23735 5414 23737 5466
rect 23917 5414 23919 5466
rect 23673 5412 23679 5414
rect 23735 5412 23759 5414
rect 23815 5412 23839 5414
rect 23895 5412 23919 5414
rect 23975 5412 23981 5414
rect 23673 5403 23981 5412
rect 23112 5228 23164 5234
rect 23112 5170 23164 5176
rect 23124 4622 23152 5170
rect 23112 4616 23164 4622
rect 23112 4558 23164 4564
rect 23673 4380 23981 4389
rect 23673 4378 23679 4380
rect 23735 4378 23759 4380
rect 23815 4378 23839 4380
rect 23895 4378 23919 4380
rect 23975 4378 23981 4380
rect 23735 4326 23737 4378
rect 23917 4326 23919 4378
rect 23673 4324 23679 4326
rect 23735 4324 23759 4326
rect 23815 4324 23839 4326
rect 23895 4324 23919 4326
rect 23975 4324 23981 4326
rect 23673 4315 23981 4324
rect 22468 4140 22520 4146
rect 22468 4082 22520 4088
rect 22376 3936 22428 3942
rect 22376 3878 22428 3884
rect 22388 3738 22416 3878
rect 21824 3732 21876 3738
rect 21824 3674 21876 3680
rect 22376 3732 22428 3738
rect 22376 3674 22428 3680
rect 19984 3528 20036 3534
rect 19984 3470 20036 3476
rect 20168 3528 20220 3534
rect 20352 3528 20404 3534
rect 20168 3470 20220 3476
rect 20350 3496 20352 3505
rect 21180 3528 21232 3534
rect 20404 3496 20406 3505
rect 21180 3470 21232 3476
rect 23388 3528 23440 3534
rect 23388 3470 23440 3476
rect 20350 3431 20406 3440
rect 19524 3188 19576 3194
rect 19524 3130 19576 3136
rect 20628 3120 20680 3126
rect 20628 3062 20680 3068
rect 19064 2984 19116 2990
rect 18694 2952 18750 2961
rect 19064 2926 19116 2932
rect 18694 2887 18750 2896
rect 19432 2916 19484 2922
rect 19432 2858 19484 2864
rect 20168 2916 20220 2922
rect 20168 2858 20220 2864
rect 19444 2650 19472 2858
rect 18604 2644 18656 2650
rect 18604 2586 18656 2592
rect 19432 2644 19484 2650
rect 19432 2586 19484 2592
rect 18880 2508 18932 2514
rect 18880 2450 18932 2456
rect 18248 1414 18368 1442
rect 18248 800 18276 1414
rect 18892 800 18920 2450
rect 19524 2440 19576 2446
rect 19524 2382 19576 2388
rect 19536 800 19564 2382
rect 20180 800 20208 2858
rect 20640 2650 20668 3062
rect 21456 2848 21508 2854
rect 21456 2790 21508 2796
rect 22744 2848 22796 2854
rect 22744 2790 22796 2796
rect 20833 2748 21141 2757
rect 20833 2746 20839 2748
rect 20895 2746 20919 2748
rect 20975 2746 20999 2748
rect 21055 2746 21079 2748
rect 21135 2746 21141 2748
rect 20895 2694 20897 2746
rect 21077 2694 21079 2746
rect 20833 2692 20839 2694
rect 20895 2692 20919 2694
rect 20975 2692 20999 2694
rect 21055 2692 21079 2694
rect 21135 2692 21141 2694
rect 20833 2683 21141 2692
rect 20628 2644 20680 2650
rect 20628 2586 20680 2592
rect 20812 2440 20864 2446
rect 20812 2382 20864 2388
rect 20824 800 20852 2382
rect 21468 800 21496 2790
rect 22100 2440 22152 2446
rect 22100 2382 22152 2388
rect 22112 800 22140 2382
rect 22756 800 22784 2790
rect 23400 800 23428 3470
rect 23673 3292 23981 3301
rect 23673 3290 23679 3292
rect 23735 3290 23759 3292
rect 23815 3290 23839 3292
rect 23895 3290 23919 3292
rect 23975 3290 23981 3292
rect 23735 3238 23737 3290
rect 23917 3238 23919 3290
rect 23673 3236 23679 3238
rect 23735 3236 23759 3238
rect 23815 3236 23839 3238
rect 23895 3236 23919 3238
rect 23975 3236 23981 3238
rect 23673 3227 23981 3236
rect 23673 2204 23981 2213
rect 23673 2202 23679 2204
rect 23735 2202 23759 2204
rect 23815 2202 23839 2204
rect 23895 2202 23919 2204
rect 23975 2202 23981 2204
rect 23735 2150 23737 2202
rect 23917 2150 23919 2202
rect 23673 2148 23679 2150
rect 23735 2148 23759 2150
rect 23815 2148 23839 2150
rect 23895 2148 23919 2150
rect 23975 2148 23981 2150
rect 23673 2139 23981 2148
rect 12544 734 12756 762
rect 13082 0 13138 800
rect 13726 0 13782 800
rect 14370 0 14426 800
rect 15014 0 15070 800
rect 15658 0 15714 800
rect 16302 0 16358 800
rect 16946 0 17002 800
rect 17590 0 17646 800
rect 18234 0 18290 800
rect 18878 0 18934 800
rect 19522 0 19578 800
rect 20166 0 20222 800
rect 20810 0 20866 800
rect 21454 0 21510 800
rect 22098 0 22154 800
rect 22742 0 22798 800
rect 23386 0 23442 800
<< via2 >>
rect 3796 22330 3852 22332
rect 3876 22330 3932 22332
rect 3956 22330 4012 22332
rect 4036 22330 4092 22332
rect 3796 22278 3842 22330
rect 3842 22278 3852 22330
rect 3876 22278 3906 22330
rect 3906 22278 3918 22330
rect 3918 22278 3932 22330
rect 3956 22278 3970 22330
rect 3970 22278 3982 22330
rect 3982 22278 4012 22330
rect 4036 22278 4046 22330
rect 4046 22278 4092 22330
rect 3796 22276 3852 22278
rect 3876 22276 3932 22278
rect 3956 22276 4012 22278
rect 4036 22276 4092 22278
rect 9477 22330 9533 22332
rect 9557 22330 9613 22332
rect 9637 22330 9693 22332
rect 9717 22330 9773 22332
rect 9477 22278 9523 22330
rect 9523 22278 9533 22330
rect 9557 22278 9587 22330
rect 9587 22278 9599 22330
rect 9599 22278 9613 22330
rect 9637 22278 9651 22330
rect 9651 22278 9663 22330
rect 9663 22278 9693 22330
rect 9717 22278 9727 22330
rect 9727 22278 9773 22330
rect 9477 22276 9533 22278
rect 9557 22276 9613 22278
rect 9637 22276 9693 22278
rect 9717 22276 9773 22278
rect 3796 21242 3852 21244
rect 3876 21242 3932 21244
rect 3956 21242 4012 21244
rect 4036 21242 4092 21244
rect 3796 21190 3842 21242
rect 3842 21190 3852 21242
rect 3876 21190 3906 21242
rect 3906 21190 3918 21242
rect 3918 21190 3932 21242
rect 3956 21190 3970 21242
rect 3970 21190 3982 21242
rect 3982 21190 4012 21242
rect 4036 21190 4046 21242
rect 4046 21190 4092 21242
rect 3796 21188 3852 21190
rect 3876 21188 3932 21190
rect 3956 21188 4012 21190
rect 4036 21188 4092 21190
rect 5446 21548 5502 21584
rect 5446 21528 5448 21548
rect 5448 21528 5500 21548
rect 5500 21528 5502 21548
rect 2318 15020 2374 15056
rect 2318 15000 2320 15020
rect 2320 15000 2372 15020
rect 2372 15000 2374 15020
rect 2778 12416 2834 12472
rect 3796 20154 3852 20156
rect 3876 20154 3932 20156
rect 3956 20154 4012 20156
rect 4036 20154 4092 20156
rect 3796 20102 3842 20154
rect 3842 20102 3852 20154
rect 3876 20102 3906 20154
rect 3906 20102 3918 20154
rect 3918 20102 3932 20154
rect 3956 20102 3970 20154
rect 3970 20102 3982 20154
rect 3982 20102 4012 20154
rect 4036 20102 4046 20154
rect 4046 20102 4092 20154
rect 3796 20100 3852 20102
rect 3876 20100 3932 20102
rect 3956 20100 4012 20102
rect 4036 20100 4092 20102
rect 3330 12416 3386 12472
rect 3514 9424 3570 9480
rect 3796 19066 3852 19068
rect 3876 19066 3932 19068
rect 3956 19066 4012 19068
rect 4036 19066 4092 19068
rect 3796 19014 3842 19066
rect 3842 19014 3852 19066
rect 3876 19014 3906 19066
rect 3906 19014 3918 19066
rect 3918 19014 3932 19066
rect 3956 19014 3970 19066
rect 3970 19014 3982 19066
rect 3982 19014 4012 19066
rect 4036 19014 4046 19066
rect 4046 19014 4092 19066
rect 3796 19012 3852 19014
rect 3876 19012 3932 19014
rect 3956 19012 4012 19014
rect 4036 19012 4092 19014
rect 3796 17978 3852 17980
rect 3876 17978 3932 17980
rect 3956 17978 4012 17980
rect 4036 17978 4092 17980
rect 3796 17926 3842 17978
rect 3842 17926 3852 17978
rect 3876 17926 3906 17978
rect 3906 17926 3918 17978
rect 3918 17926 3932 17978
rect 3956 17926 3970 17978
rect 3970 17926 3982 17978
rect 3982 17926 4012 17978
rect 4036 17926 4046 17978
rect 4046 17926 4092 17978
rect 3796 17924 3852 17926
rect 3876 17924 3932 17926
rect 3956 17924 4012 17926
rect 4036 17924 4092 17926
rect 3796 16890 3852 16892
rect 3876 16890 3932 16892
rect 3956 16890 4012 16892
rect 4036 16890 4092 16892
rect 3796 16838 3842 16890
rect 3842 16838 3852 16890
rect 3876 16838 3906 16890
rect 3906 16838 3918 16890
rect 3918 16838 3932 16890
rect 3956 16838 3970 16890
rect 3970 16838 3982 16890
rect 3982 16838 4012 16890
rect 4036 16838 4046 16890
rect 4046 16838 4092 16890
rect 3796 16836 3852 16838
rect 3876 16836 3932 16838
rect 3956 16836 4012 16838
rect 4036 16836 4092 16838
rect 3796 15802 3852 15804
rect 3876 15802 3932 15804
rect 3956 15802 4012 15804
rect 4036 15802 4092 15804
rect 3796 15750 3842 15802
rect 3842 15750 3852 15802
rect 3876 15750 3906 15802
rect 3906 15750 3918 15802
rect 3918 15750 3932 15802
rect 3956 15750 3970 15802
rect 3970 15750 3982 15802
rect 3982 15750 4012 15802
rect 4036 15750 4046 15802
rect 4046 15750 4092 15802
rect 3796 15748 3852 15750
rect 3876 15748 3932 15750
rect 3956 15748 4012 15750
rect 4036 15748 4092 15750
rect 3796 14714 3852 14716
rect 3876 14714 3932 14716
rect 3956 14714 4012 14716
rect 4036 14714 4092 14716
rect 3796 14662 3842 14714
rect 3842 14662 3852 14714
rect 3876 14662 3906 14714
rect 3906 14662 3918 14714
rect 3918 14662 3932 14714
rect 3956 14662 3970 14714
rect 3970 14662 3982 14714
rect 3982 14662 4012 14714
rect 4036 14662 4046 14714
rect 4046 14662 4092 14714
rect 3796 14660 3852 14662
rect 3876 14660 3932 14662
rect 3956 14660 4012 14662
rect 4036 14660 4092 14662
rect 3796 13626 3852 13628
rect 3876 13626 3932 13628
rect 3956 13626 4012 13628
rect 4036 13626 4092 13628
rect 3796 13574 3842 13626
rect 3842 13574 3852 13626
rect 3876 13574 3906 13626
rect 3906 13574 3918 13626
rect 3918 13574 3932 13626
rect 3956 13574 3970 13626
rect 3970 13574 3982 13626
rect 3982 13574 4012 13626
rect 4036 13574 4046 13626
rect 4046 13574 4092 13626
rect 3796 13572 3852 13574
rect 3876 13572 3932 13574
rect 3956 13572 4012 13574
rect 4036 13572 4092 13574
rect 3796 12538 3852 12540
rect 3876 12538 3932 12540
rect 3956 12538 4012 12540
rect 4036 12538 4092 12540
rect 3796 12486 3842 12538
rect 3842 12486 3852 12538
rect 3876 12486 3906 12538
rect 3906 12486 3918 12538
rect 3918 12486 3932 12538
rect 3956 12486 3970 12538
rect 3970 12486 3982 12538
rect 3982 12486 4012 12538
rect 4036 12486 4046 12538
rect 4046 12486 4092 12538
rect 3796 12484 3852 12486
rect 3876 12484 3932 12486
rect 3956 12484 4012 12486
rect 4036 12484 4092 12486
rect 3796 11450 3852 11452
rect 3876 11450 3932 11452
rect 3956 11450 4012 11452
rect 4036 11450 4092 11452
rect 3796 11398 3842 11450
rect 3842 11398 3852 11450
rect 3876 11398 3906 11450
rect 3906 11398 3918 11450
rect 3918 11398 3932 11450
rect 3956 11398 3970 11450
rect 3970 11398 3982 11450
rect 3982 11398 4012 11450
rect 4036 11398 4046 11450
rect 4046 11398 4092 11450
rect 3796 11396 3852 11398
rect 3876 11396 3932 11398
rect 3956 11396 4012 11398
rect 4036 11396 4092 11398
rect 3796 10362 3852 10364
rect 3876 10362 3932 10364
rect 3956 10362 4012 10364
rect 4036 10362 4092 10364
rect 3796 10310 3842 10362
rect 3842 10310 3852 10362
rect 3876 10310 3906 10362
rect 3906 10310 3918 10362
rect 3918 10310 3932 10362
rect 3956 10310 3970 10362
rect 3970 10310 3982 10362
rect 3982 10310 4012 10362
rect 4036 10310 4046 10362
rect 4046 10310 4092 10362
rect 3796 10308 3852 10310
rect 3876 10308 3932 10310
rect 3956 10308 4012 10310
rect 4036 10308 4092 10310
rect 3796 9274 3852 9276
rect 3876 9274 3932 9276
rect 3956 9274 4012 9276
rect 4036 9274 4092 9276
rect 3796 9222 3842 9274
rect 3842 9222 3852 9274
rect 3876 9222 3906 9274
rect 3906 9222 3918 9274
rect 3918 9222 3932 9274
rect 3956 9222 3970 9274
rect 3970 9222 3982 9274
rect 3982 9222 4012 9274
rect 4036 9222 4046 9274
rect 4046 9222 4092 9274
rect 3796 9220 3852 9222
rect 3876 9220 3932 9222
rect 3956 9220 4012 9222
rect 4036 9220 4092 9222
rect 3796 8186 3852 8188
rect 3876 8186 3932 8188
rect 3956 8186 4012 8188
rect 4036 8186 4092 8188
rect 3796 8134 3842 8186
rect 3842 8134 3852 8186
rect 3876 8134 3906 8186
rect 3906 8134 3918 8186
rect 3918 8134 3932 8186
rect 3956 8134 3970 8186
rect 3970 8134 3982 8186
rect 3982 8134 4012 8186
rect 4036 8134 4046 8186
rect 4046 8134 4092 8186
rect 3796 8132 3852 8134
rect 3876 8132 3932 8134
rect 3956 8132 4012 8134
rect 4036 8132 4092 8134
rect 4986 15020 5042 15056
rect 4986 15000 4988 15020
rect 4988 15000 5040 15020
rect 5040 15000 5042 15020
rect 5262 15272 5318 15328
rect 5170 9968 5226 10024
rect 3796 7098 3852 7100
rect 3876 7098 3932 7100
rect 3956 7098 4012 7100
rect 4036 7098 4092 7100
rect 3796 7046 3842 7098
rect 3842 7046 3852 7098
rect 3876 7046 3906 7098
rect 3906 7046 3918 7098
rect 3918 7046 3932 7098
rect 3956 7046 3970 7098
rect 3970 7046 3982 7098
rect 3982 7046 4012 7098
rect 4036 7046 4046 7098
rect 4046 7046 4092 7098
rect 3796 7044 3852 7046
rect 3876 7044 3932 7046
rect 3956 7044 4012 7046
rect 4036 7044 4092 7046
rect 3796 6010 3852 6012
rect 3876 6010 3932 6012
rect 3956 6010 4012 6012
rect 4036 6010 4092 6012
rect 3796 5958 3842 6010
rect 3842 5958 3852 6010
rect 3876 5958 3906 6010
rect 3906 5958 3918 6010
rect 3918 5958 3932 6010
rect 3956 5958 3970 6010
rect 3970 5958 3982 6010
rect 3982 5958 4012 6010
rect 4036 5958 4046 6010
rect 4046 5958 4092 6010
rect 3796 5956 3852 5958
rect 3876 5956 3932 5958
rect 3956 5956 4012 5958
rect 4036 5956 4092 5958
rect 3330 3460 3386 3496
rect 3330 3440 3332 3460
rect 3332 3440 3384 3460
rect 3384 3440 3386 3460
rect 3796 4922 3852 4924
rect 3876 4922 3932 4924
rect 3956 4922 4012 4924
rect 4036 4922 4092 4924
rect 3796 4870 3842 4922
rect 3842 4870 3852 4922
rect 3876 4870 3906 4922
rect 3906 4870 3918 4922
rect 3918 4870 3932 4922
rect 3956 4870 3970 4922
rect 3970 4870 3982 4922
rect 3982 4870 4012 4922
rect 4036 4870 4046 4922
rect 4046 4870 4092 4922
rect 3796 4868 3852 4870
rect 3876 4868 3932 4870
rect 3956 4868 4012 4870
rect 4036 4868 4092 4870
rect 5354 9424 5410 9480
rect 5354 6704 5410 6760
rect 5170 6160 5226 6216
rect 3796 3834 3852 3836
rect 3876 3834 3932 3836
rect 3956 3834 4012 3836
rect 4036 3834 4092 3836
rect 3796 3782 3842 3834
rect 3842 3782 3852 3834
rect 3876 3782 3906 3834
rect 3906 3782 3918 3834
rect 3918 3782 3932 3834
rect 3956 3782 3970 3834
rect 3970 3782 3982 3834
rect 3982 3782 4012 3834
rect 4036 3782 4046 3834
rect 4046 3782 4092 3834
rect 3796 3780 3852 3782
rect 3876 3780 3932 3782
rect 3956 3780 4012 3782
rect 4036 3780 4092 3782
rect 4342 3732 4398 3768
rect 4342 3712 4344 3732
rect 4344 3712 4396 3732
rect 4396 3712 4398 3732
rect 3796 2746 3852 2748
rect 3876 2746 3932 2748
rect 3956 2746 4012 2748
rect 4036 2746 4092 2748
rect 3796 2694 3842 2746
rect 3842 2694 3852 2746
rect 3876 2694 3906 2746
rect 3906 2694 3918 2746
rect 3918 2694 3932 2746
rect 3956 2694 3970 2746
rect 3970 2694 3982 2746
rect 3982 2694 4012 2746
rect 4036 2694 4046 2746
rect 4046 2694 4092 2746
rect 3796 2692 3852 2694
rect 3876 2692 3932 2694
rect 3956 2692 4012 2694
rect 4036 2692 4092 2694
rect 6636 21786 6692 21788
rect 6716 21786 6772 21788
rect 6796 21786 6852 21788
rect 6876 21786 6932 21788
rect 6636 21734 6682 21786
rect 6682 21734 6692 21786
rect 6716 21734 6746 21786
rect 6746 21734 6758 21786
rect 6758 21734 6772 21786
rect 6796 21734 6810 21786
rect 6810 21734 6822 21786
rect 6822 21734 6852 21786
rect 6876 21734 6886 21786
rect 6886 21734 6932 21786
rect 6636 21732 6692 21734
rect 6716 21732 6772 21734
rect 6796 21732 6852 21734
rect 6876 21732 6932 21734
rect 6636 20698 6692 20700
rect 6716 20698 6772 20700
rect 6796 20698 6852 20700
rect 6876 20698 6932 20700
rect 6636 20646 6682 20698
rect 6682 20646 6692 20698
rect 6716 20646 6746 20698
rect 6746 20646 6758 20698
rect 6758 20646 6772 20698
rect 6796 20646 6810 20698
rect 6810 20646 6822 20698
rect 6822 20646 6852 20698
rect 6876 20646 6886 20698
rect 6886 20646 6932 20698
rect 6636 20644 6692 20646
rect 6716 20644 6772 20646
rect 6796 20644 6852 20646
rect 6876 20644 6932 20646
rect 6636 19610 6692 19612
rect 6716 19610 6772 19612
rect 6796 19610 6852 19612
rect 6876 19610 6932 19612
rect 6636 19558 6682 19610
rect 6682 19558 6692 19610
rect 6716 19558 6746 19610
rect 6746 19558 6758 19610
rect 6758 19558 6772 19610
rect 6796 19558 6810 19610
rect 6810 19558 6822 19610
rect 6822 19558 6852 19610
rect 6876 19558 6886 19610
rect 6886 19558 6932 19610
rect 6636 19556 6692 19558
rect 6716 19556 6772 19558
rect 6796 19556 6852 19558
rect 6876 19556 6932 19558
rect 6636 18522 6692 18524
rect 6716 18522 6772 18524
rect 6796 18522 6852 18524
rect 6876 18522 6932 18524
rect 6636 18470 6682 18522
rect 6682 18470 6692 18522
rect 6716 18470 6746 18522
rect 6746 18470 6758 18522
rect 6758 18470 6772 18522
rect 6796 18470 6810 18522
rect 6810 18470 6822 18522
rect 6822 18470 6852 18522
rect 6876 18470 6886 18522
rect 6886 18470 6932 18522
rect 6636 18468 6692 18470
rect 6716 18468 6772 18470
rect 6796 18468 6852 18470
rect 6876 18468 6932 18470
rect 5722 9460 5724 9480
rect 5724 9460 5776 9480
rect 5776 9460 5778 9480
rect 5722 9424 5778 9460
rect 5814 9288 5870 9344
rect 6636 17434 6692 17436
rect 6716 17434 6772 17436
rect 6796 17434 6852 17436
rect 6876 17434 6932 17436
rect 6636 17382 6682 17434
rect 6682 17382 6692 17434
rect 6716 17382 6746 17434
rect 6746 17382 6758 17434
rect 6758 17382 6772 17434
rect 6796 17382 6810 17434
rect 6810 17382 6822 17434
rect 6822 17382 6852 17434
rect 6876 17382 6886 17434
rect 6886 17382 6932 17434
rect 6636 17380 6692 17382
rect 6716 17380 6772 17382
rect 6796 17380 6852 17382
rect 6876 17380 6932 17382
rect 6636 16346 6692 16348
rect 6716 16346 6772 16348
rect 6796 16346 6852 16348
rect 6876 16346 6932 16348
rect 6636 16294 6682 16346
rect 6682 16294 6692 16346
rect 6716 16294 6746 16346
rect 6746 16294 6758 16346
rect 6758 16294 6772 16346
rect 6796 16294 6810 16346
rect 6810 16294 6822 16346
rect 6822 16294 6852 16346
rect 6876 16294 6886 16346
rect 6886 16294 6932 16346
rect 6636 16292 6692 16294
rect 6716 16292 6772 16294
rect 6796 16292 6852 16294
rect 6876 16292 6932 16294
rect 6636 15258 6692 15260
rect 6716 15258 6772 15260
rect 6796 15258 6852 15260
rect 6876 15258 6932 15260
rect 6636 15206 6682 15258
rect 6682 15206 6692 15258
rect 6716 15206 6746 15258
rect 6746 15206 6758 15258
rect 6758 15206 6772 15258
rect 6796 15206 6810 15258
rect 6810 15206 6822 15258
rect 6822 15206 6852 15258
rect 6876 15206 6886 15258
rect 6886 15206 6932 15258
rect 6636 15204 6692 15206
rect 6716 15204 6772 15206
rect 6796 15204 6852 15206
rect 6876 15204 6932 15206
rect 7010 15000 7066 15056
rect 6636 14170 6692 14172
rect 6716 14170 6772 14172
rect 6796 14170 6852 14172
rect 6876 14170 6932 14172
rect 6636 14118 6682 14170
rect 6682 14118 6692 14170
rect 6716 14118 6746 14170
rect 6746 14118 6758 14170
rect 6758 14118 6772 14170
rect 6796 14118 6810 14170
rect 6810 14118 6822 14170
rect 6822 14118 6852 14170
rect 6876 14118 6886 14170
rect 6886 14118 6932 14170
rect 6636 14116 6692 14118
rect 6716 14116 6772 14118
rect 6796 14116 6852 14118
rect 6876 14116 6932 14118
rect 6636 13082 6692 13084
rect 6716 13082 6772 13084
rect 6796 13082 6852 13084
rect 6876 13082 6932 13084
rect 6636 13030 6682 13082
rect 6682 13030 6692 13082
rect 6716 13030 6746 13082
rect 6746 13030 6758 13082
rect 6758 13030 6772 13082
rect 6796 13030 6810 13082
rect 6810 13030 6822 13082
rect 6822 13030 6852 13082
rect 6876 13030 6886 13082
rect 6886 13030 6932 13082
rect 6636 13028 6692 13030
rect 6716 13028 6772 13030
rect 6796 13028 6852 13030
rect 6876 13028 6932 13030
rect 6636 11994 6692 11996
rect 6716 11994 6772 11996
rect 6796 11994 6852 11996
rect 6876 11994 6932 11996
rect 6636 11942 6682 11994
rect 6682 11942 6692 11994
rect 6716 11942 6746 11994
rect 6746 11942 6758 11994
rect 6758 11942 6772 11994
rect 6796 11942 6810 11994
rect 6810 11942 6822 11994
rect 6822 11942 6852 11994
rect 6876 11942 6886 11994
rect 6886 11942 6932 11994
rect 6636 11940 6692 11942
rect 6716 11940 6772 11942
rect 6796 11940 6852 11942
rect 6876 11940 6932 11942
rect 6636 10906 6692 10908
rect 6716 10906 6772 10908
rect 6796 10906 6852 10908
rect 6876 10906 6932 10908
rect 6636 10854 6682 10906
rect 6682 10854 6692 10906
rect 6716 10854 6746 10906
rect 6746 10854 6758 10906
rect 6758 10854 6772 10906
rect 6796 10854 6810 10906
rect 6810 10854 6822 10906
rect 6822 10854 6852 10906
rect 6876 10854 6886 10906
rect 6886 10854 6932 10906
rect 6636 10852 6692 10854
rect 6716 10852 6772 10854
rect 6796 10852 6852 10854
rect 6876 10852 6932 10854
rect 5630 2932 5632 2952
rect 5632 2932 5684 2952
rect 5684 2932 5686 2952
rect 5630 2896 5686 2932
rect 7010 9968 7066 10024
rect 6636 9818 6692 9820
rect 6716 9818 6772 9820
rect 6796 9818 6852 9820
rect 6876 9818 6932 9820
rect 6636 9766 6682 9818
rect 6682 9766 6692 9818
rect 6716 9766 6746 9818
rect 6746 9766 6758 9818
rect 6758 9766 6772 9818
rect 6796 9766 6810 9818
rect 6810 9766 6822 9818
rect 6822 9766 6852 9818
rect 6876 9766 6886 9818
rect 6886 9766 6932 9818
rect 6636 9764 6692 9766
rect 6716 9764 6772 9766
rect 6796 9764 6852 9766
rect 6876 9764 6932 9766
rect 6642 9288 6698 9344
rect 7286 10548 7288 10568
rect 7288 10548 7340 10568
rect 7340 10548 7342 10568
rect 7286 10512 7342 10548
rect 6636 8730 6692 8732
rect 6716 8730 6772 8732
rect 6796 8730 6852 8732
rect 6876 8730 6932 8732
rect 6636 8678 6682 8730
rect 6682 8678 6692 8730
rect 6716 8678 6746 8730
rect 6746 8678 6758 8730
rect 6758 8678 6772 8730
rect 6796 8678 6810 8730
rect 6810 8678 6822 8730
rect 6822 8678 6852 8730
rect 6876 8678 6886 8730
rect 6886 8678 6932 8730
rect 6636 8676 6692 8678
rect 6716 8676 6772 8678
rect 6796 8676 6852 8678
rect 6876 8676 6932 8678
rect 6636 7642 6692 7644
rect 6716 7642 6772 7644
rect 6796 7642 6852 7644
rect 6876 7642 6932 7644
rect 6636 7590 6682 7642
rect 6682 7590 6692 7642
rect 6716 7590 6746 7642
rect 6746 7590 6758 7642
rect 6758 7590 6772 7642
rect 6796 7590 6810 7642
rect 6810 7590 6822 7642
rect 6822 7590 6852 7642
rect 6876 7590 6886 7642
rect 6886 7590 6932 7642
rect 6636 7588 6692 7590
rect 6716 7588 6772 7590
rect 6796 7588 6852 7590
rect 6876 7588 6932 7590
rect 6636 6554 6692 6556
rect 6716 6554 6772 6556
rect 6796 6554 6852 6556
rect 6876 6554 6932 6556
rect 6636 6502 6682 6554
rect 6682 6502 6692 6554
rect 6716 6502 6746 6554
rect 6746 6502 6758 6554
rect 6758 6502 6772 6554
rect 6796 6502 6810 6554
rect 6810 6502 6822 6554
rect 6822 6502 6852 6554
rect 6876 6502 6886 6554
rect 6886 6502 6932 6554
rect 6636 6500 6692 6502
rect 6716 6500 6772 6502
rect 6796 6500 6852 6502
rect 6876 6500 6932 6502
rect 6636 5466 6692 5468
rect 6716 5466 6772 5468
rect 6796 5466 6852 5468
rect 6876 5466 6932 5468
rect 6636 5414 6682 5466
rect 6682 5414 6692 5466
rect 6716 5414 6746 5466
rect 6746 5414 6758 5466
rect 6758 5414 6772 5466
rect 6796 5414 6810 5466
rect 6810 5414 6822 5466
rect 6822 5414 6852 5466
rect 6876 5414 6886 5466
rect 6886 5414 6932 5466
rect 6636 5412 6692 5414
rect 6716 5412 6772 5414
rect 6796 5412 6852 5414
rect 6876 5412 6932 5414
rect 6274 5072 6330 5128
rect 6636 4378 6692 4380
rect 6716 4378 6772 4380
rect 6796 4378 6852 4380
rect 6876 4378 6932 4380
rect 6636 4326 6682 4378
rect 6682 4326 6692 4378
rect 6716 4326 6746 4378
rect 6746 4326 6758 4378
rect 6758 4326 6772 4378
rect 6796 4326 6810 4378
rect 6810 4326 6822 4378
rect 6822 4326 6852 4378
rect 6876 4326 6886 4378
rect 6886 4326 6932 4378
rect 6636 4324 6692 4326
rect 6716 4324 6772 4326
rect 6796 4324 6852 4326
rect 6876 4324 6932 4326
rect 6636 3290 6692 3292
rect 6716 3290 6772 3292
rect 6796 3290 6852 3292
rect 6876 3290 6932 3292
rect 6636 3238 6682 3290
rect 6682 3238 6692 3290
rect 6716 3238 6746 3290
rect 6746 3238 6758 3290
rect 6758 3238 6772 3290
rect 6796 3238 6810 3290
rect 6810 3238 6822 3290
rect 6822 3238 6852 3290
rect 6876 3238 6886 3290
rect 6886 3238 6932 3290
rect 6636 3236 6692 3238
rect 6716 3236 6772 3238
rect 6796 3236 6852 3238
rect 6876 3236 6932 3238
rect 7194 3576 7250 3632
rect 6636 2202 6692 2204
rect 6716 2202 6772 2204
rect 6796 2202 6852 2204
rect 6876 2202 6932 2204
rect 6636 2150 6682 2202
rect 6682 2150 6692 2202
rect 6716 2150 6746 2202
rect 6746 2150 6758 2202
rect 6758 2150 6772 2202
rect 6796 2150 6810 2202
rect 6810 2150 6822 2202
rect 6822 2150 6852 2202
rect 6876 2150 6886 2202
rect 6886 2150 6932 2202
rect 6636 2148 6692 2150
rect 6716 2148 6772 2150
rect 6796 2148 6852 2150
rect 6876 2148 6932 2150
rect 7654 6296 7710 6352
rect 15158 22330 15214 22332
rect 15238 22330 15294 22332
rect 15318 22330 15374 22332
rect 15398 22330 15454 22332
rect 15158 22278 15204 22330
rect 15204 22278 15214 22330
rect 15238 22278 15268 22330
rect 15268 22278 15280 22330
rect 15280 22278 15294 22330
rect 15318 22278 15332 22330
rect 15332 22278 15344 22330
rect 15344 22278 15374 22330
rect 15398 22278 15408 22330
rect 15408 22278 15454 22330
rect 15158 22276 15214 22278
rect 15238 22276 15294 22278
rect 15318 22276 15374 22278
rect 15398 22276 15454 22278
rect 20839 22330 20895 22332
rect 20919 22330 20975 22332
rect 20999 22330 21055 22332
rect 21079 22330 21135 22332
rect 20839 22278 20885 22330
rect 20885 22278 20895 22330
rect 20919 22278 20949 22330
rect 20949 22278 20961 22330
rect 20961 22278 20975 22330
rect 20999 22278 21013 22330
rect 21013 22278 21025 22330
rect 21025 22278 21055 22330
rect 21079 22278 21089 22330
rect 21089 22278 21135 22330
rect 20839 22276 20895 22278
rect 20919 22276 20975 22278
rect 20999 22276 21055 22278
rect 21079 22276 21135 22278
rect 12317 21786 12373 21788
rect 12397 21786 12453 21788
rect 12477 21786 12533 21788
rect 12557 21786 12613 21788
rect 12317 21734 12363 21786
rect 12363 21734 12373 21786
rect 12397 21734 12427 21786
rect 12427 21734 12439 21786
rect 12439 21734 12453 21786
rect 12477 21734 12491 21786
rect 12491 21734 12503 21786
rect 12503 21734 12533 21786
rect 12557 21734 12567 21786
rect 12567 21734 12613 21786
rect 12317 21732 12373 21734
rect 12397 21732 12453 21734
rect 12477 21732 12533 21734
rect 12557 21732 12613 21734
rect 9477 21242 9533 21244
rect 9557 21242 9613 21244
rect 9637 21242 9693 21244
rect 9717 21242 9773 21244
rect 9477 21190 9523 21242
rect 9523 21190 9533 21242
rect 9557 21190 9587 21242
rect 9587 21190 9599 21242
rect 9599 21190 9613 21242
rect 9637 21190 9651 21242
rect 9651 21190 9663 21242
rect 9663 21190 9693 21242
rect 9717 21190 9727 21242
rect 9727 21190 9773 21242
rect 9477 21188 9533 21190
rect 9557 21188 9613 21190
rect 9637 21188 9693 21190
rect 9717 21188 9773 21190
rect 9477 20154 9533 20156
rect 9557 20154 9613 20156
rect 9637 20154 9693 20156
rect 9717 20154 9773 20156
rect 9477 20102 9523 20154
rect 9523 20102 9533 20154
rect 9557 20102 9587 20154
rect 9587 20102 9599 20154
rect 9599 20102 9613 20154
rect 9637 20102 9651 20154
rect 9651 20102 9663 20154
rect 9663 20102 9693 20154
rect 9717 20102 9727 20154
rect 9727 20102 9773 20154
rect 9477 20100 9533 20102
rect 9557 20100 9613 20102
rect 9637 20100 9693 20102
rect 9717 20100 9773 20102
rect 9477 19066 9533 19068
rect 9557 19066 9613 19068
rect 9637 19066 9693 19068
rect 9717 19066 9773 19068
rect 9477 19014 9523 19066
rect 9523 19014 9533 19066
rect 9557 19014 9587 19066
rect 9587 19014 9599 19066
rect 9599 19014 9613 19066
rect 9637 19014 9651 19066
rect 9651 19014 9663 19066
rect 9663 19014 9693 19066
rect 9717 19014 9727 19066
rect 9727 19014 9773 19066
rect 9477 19012 9533 19014
rect 9557 19012 9613 19014
rect 9637 19012 9693 19014
rect 9717 19012 9773 19014
rect 9477 17978 9533 17980
rect 9557 17978 9613 17980
rect 9637 17978 9693 17980
rect 9717 17978 9773 17980
rect 9477 17926 9523 17978
rect 9523 17926 9533 17978
rect 9557 17926 9587 17978
rect 9587 17926 9599 17978
rect 9599 17926 9613 17978
rect 9637 17926 9651 17978
rect 9651 17926 9663 17978
rect 9663 17926 9693 17978
rect 9717 17926 9727 17978
rect 9727 17926 9773 17978
rect 9477 17924 9533 17926
rect 9557 17924 9613 17926
rect 9637 17924 9693 17926
rect 9717 17924 9773 17926
rect 9477 16890 9533 16892
rect 9557 16890 9613 16892
rect 9637 16890 9693 16892
rect 9717 16890 9773 16892
rect 9477 16838 9523 16890
rect 9523 16838 9533 16890
rect 9557 16838 9587 16890
rect 9587 16838 9599 16890
rect 9599 16838 9613 16890
rect 9637 16838 9651 16890
rect 9651 16838 9663 16890
rect 9663 16838 9693 16890
rect 9717 16838 9727 16890
rect 9727 16838 9773 16890
rect 9477 16836 9533 16838
rect 9557 16836 9613 16838
rect 9637 16836 9693 16838
rect 9717 16836 9773 16838
rect 9477 15802 9533 15804
rect 9557 15802 9613 15804
rect 9637 15802 9693 15804
rect 9717 15802 9773 15804
rect 9477 15750 9523 15802
rect 9523 15750 9533 15802
rect 9557 15750 9587 15802
rect 9587 15750 9599 15802
rect 9599 15750 9613 15802
rect 9637 15750 9651 15802
rect 9651 15750 9663 15802
rect 9663 15750 9693 15802
rect 9717 15750 9727 15802
rect 9727 15750 9773 15802
rect 9477 15748 9533 15750
rect 9557 15748 9613 15750
rect 9637 15748 9693 15750
rect 9717 15748 9773 15750
rect 9477 14714 9533 14716
rect 9557 14714 9613 14716
rect 9637 14714 9693 14716
rect 9717 14714 9773 14716
rect 9477 14662 9523 14714
rect 9523 14662 9533 14714
rect 9557 14662 9587 14714
rect 9587 14662 9599 14714
rect 9599 14662 9613 14714
rect 9637 14662 9651 14714
rect 9651 14662 9663 14714
rect 9663 14662 9693 14714
rect 9717 14662 9727 14714
rect 9727 14662 9773 14714
rect 9477 14660 9533 14662
rect 9557 14660 9613 14662
rect 9637 14660 9693 14662
rect 9717 14660 9773 14662
rect 9477 13626 9533 13628
rect 9557 13626 9613 13628
rect 9637 13626 9693 13628
rect 9717 13626 9773 13628
rect 9477 13574 9523 13626
rect 9523 13574 9533 13626
rect 9557 13574 9587 13626
rect 9587 13574 9599 13626
rect 9599 13574 9613 13626
rect 9637 13574 9651 13626
rect 9651 13574 9663 13626
rect 9663 13574 9693 13626
rect 9717 13574 9727 13626
rect 9727 13574 9773 13626
rect 9477 13572 9533 13574
rect 9557 13572 9613 13574
rect 9637 13572 9693 13574
rect 9717 13572 9773 13574
rect 8482 7928 8538 7984
rect 8298 6432 8354 6488
rect 7654 3712 7710 3768
rect 9477 12538 9533 12540
rect 9557 12538 9613 12540
rect 9637 12538 9693 12540
rect 9717 12538 9773 12540
rect 9477 12486 9523 12538
rect 9523 12486 9533 12538
rect 9557 12486 9587 12538
rect 9587 12486 9599 12538
rect 9599 12486 9613 12538
rect 9637 12486 9651 12538
rect 9651 12486 9663 12538
rect 9663 12486 9693 12538
rect 9717 12486 9727 12538
rect 9727 12486 9773 12538
rect 9477 12484 9533 12486
rect 9557 12484 9613 12486
rect 9637 12484 9693 12486
rect 9717 12484 9773 12486
rect 9477 11450 9533 11452
rect 9557 11450 9613 11452
rect 9637 11450 9693 11452
rect 9717 11450 9773 11452
rect 9477 11398 9523 11450
rect 9523 11398 9533 11450
rect 9557 11398 9587 11450
rect 9587 11398 9599 11450
rect 9599 11398 9613 11450
rect 9637 11398 9651 11450
rect 9651 11398 9663 11450
rect 9663 11398 9693 11450
rect 9717 11398 9727 11450
rect 9727 11398 9773 11450
rect 9477 11396 9533 11398
rect 9557 11396 9613 11398
rect 9637 11396 9693 11398
rect 9717 11396 9773 11398
rect 9477 10362 9533 10364
rect 9557 10362 9613 10364
rect 9637 10362 9693 10364
rect 9717 10362 9773 10364
rect 9477 10310 9523 10362
rect 9523 10310 9533 10362
rect 9557 10310 9587 10362
rect 9587 10310 9599 10362
rect 9599 10310 9613 10362
rect 9637 10310 9651 10362
rect 9651 10310 9663 10362
rect 9663 10310 9693 10362
rect 9717 10310 9727 10362
rect 9727 10310 9773 10362
rect 9477 10308 9533 10310
rect 9557 10308 9613 10310
rect 9637 10308 9693 10310
rect 9717 10308 9773 10310
rect 9126 9424 9182 9480
rect 9494 9460 9496 9480
rect 9496 9460 9548 9480
rect 9548 9460 9550 9480
rect 9494 9424 9550 9460
rect 9477 9274 9533 9276
rect 9557 9274 9613 9276
rect 9637 9274 9693 9276
rect 9717 9274 9773 9276
rect 9477 9222 9523 9274
rect 9523 9222 9533 9274
rect 9557 9222 9587 9274
rect 9587 9222 9599 9274
rect 9599 9222 9613 9274
rect 9637 9222 9651 9274
rect 9651 9222 9663 9274
rect 9663 9222 9693 9274
rect 9717 9222 9727 9274
rect 9727 9222 9773 9274
rect 9477 9220 9533 9222
rect 9557 9220 9613 9222
rect 9637 9220 9693 9222
rect 9717 9220 9773 9222
rect 9477 8186 9533 8188
rect 9557 8186 9613 8188
rect 9637 8186 9693 8188
rect 9717 8186 9773 8188
rect 9477 8134 9523 8186
rect 9523 8134 9533 8186
rect 9557 8134 9587 8186
rect 9587 8134 9599 8186
rect 9599 8134 9613 8186
rect 9637 8134 9651 8186
rect 9651 8134 9663 8186
rect 9663 8134 9693 8186
rect 9717 8134 9727 8186
rect 9727 8134 9773 8186
rect 9477 8132 9533 8134
rect 9557 8132 9613 8134
rect 9637 8132 9693 8134
rect 9717 8132 9773 8134
rect 9477 7098 9533 7100
rect 9557 7098 9613 7100
rect 9637 7098 9693 7100
rect 9717 7098 9773 7100
rect 9477 7046 9523 7098
rect 9523 7046 9533 7098
rect 9557 7046 9587 7098
rect 9587 7046 9599 7098
rect 9599 7046 9613 7098
rect 9637 7046 9651 7098
rect 9651 7046 9663 7098
rect 9663 7046 9693 7098
rect 9717 7046 9727 7098
rect 9727 7046 9773 7098
rect 9477 7044 9533 7046
rect 9557 7044 9613 7046
rect 9637 7044 9693 7046
rect 9717 7044 9773 7046
rect 8942 6452 8998 6488
rect 8942 6432 8944 6452
rect 8944 6432 8996 6452
rect 8996 6432 8998 6452
rect 8850 6332 8852 6352
rect 8852 6332 8904 6352
rect 8904 6332 8906 6352
rect 8850 6296 8906 6332
rect 9954 6568 10010 6624
rect 12317 20698 12373 20700
rect 12397 20698 12453 20700
rect 12477 20698 12533 20700
rect 12557 20698 12613 20700
rect 12317 20646 12363 20698
rect 12363 20646 12373 20698
rect 12397 20646 12427 20698
rect 12427 20646 12439 20698
rect 12439 20646 12453 20698
rect 12477 20646 12491 20698
rect 12491 20646 12503 20698
rect 12503 20646 12533 20698
rect 12557 20646 12567 20698
rect 12567 20646 12613 20698
rect 12317 20644 12373 20646
rect 12397 20644 12453 20646
rect 12477 20644 12533 20646
rect 12557 20644 12613 20646
rect 12317 19610 12373 19612
rect 12397 19610 12453 19612
rect 12477 19610 12533 19612
rect 12557 19610 12613 19612
rect 12317 19558 12363 19610
rect 12363 19558 12373 19610
rect 12397 19558 12427 19610
rect 12427 19558 12439 19610
rect 12439 19558 12453 19610
rect 12477 19558 12491 19610
rect 12491 19558 12503 19610
rect 12503 19558 12533 19610
rect 12557 19558 12567 19610
rect 12567 19558 12613 19610
rect 12317 19556 12373 19558
rect 12397 19556 12453 19558
rect 12477 19556 12533 19558
rect 12557 19556 12613 19558
rect 12317 18522 12373 18524
rect 12397 18522 12453 18524
rect 12477 18522 12533 18524
rect 12557 18522 12613 18524
rect 12317 18470 12363 18522
rect 12363 18470 12373 18522
rect 12397 18470 12427 18522
rect 12427 18470 12439 18522
rect 12439 18470 12453 18522
rect 12477 18470 12491 18522
rect 12491 18470 12503 18522
rect 12503 18470 12533 18522
rect 12557 18470 12567 18522
rect 12567 18470 12613 18522
rect 12317 18468 12373 18470
rect 12397 18468 12453 18470
rect 12477 18468 12533 18470
rect 12557 18468 12613 18470
rect 12317 17434 12373 17436
rect 12397 17434 12453 17436
rect 12477 17434 12533 17436
rect 12557 17434 12613 17436
rect 12317 17382 12363 17434
rect 12363 17382 12373 17434
rect 12397 17382 12427 17434
rect 12427 17382 12439 17434
rect 12439 17382 12453 17434
rect 12477 17382 12491 17434
rect 12491 17382 12503 17434
rect 12503 17382 12533 17434
rect 12557 17382 12567 17434
rect 12567 17382 12613 17434
rect 12317 17380 12373 17382
rect 12397 17380 12453 17382
rect 12477 17380 12533 17382
rect 12557 17380 12613 17382
rect 10506 10648 10562 10704
rect 10506 9868 10508 9888
rect 10508 9868 10560 9888
rect 10560 9868 10562 9888
rect 10506 9832 10562 9868
rect 10322 6568 10378 6624
rect 9477 6010 9533 6012
rect 9557 6010 9613 6012
rect 9637 6010 9693 6012
rect 9717 6010 9773 6012
rect 9477 5958 9523 6010
rect 9523 5958 9533 6010
rect 9557 5958 9587 6010
rect 9587 5958 9599 6010
rect 9599 5958 9613 6010
rect 9637 5958 9651 6010
rect 9651 5958 9663 6010
rect 9663 5958 9693 6010
rect 9717 5958 9727 6010
rect 9727 5958 9773 6010
rect 9477 5956 9533 5958
rect 9557 5956 9613 5958
rect 9637 5956 9693 5958
rect 9717 5956 9773 5958
rect 9126 5480 9182 5536
rect 8022 4120 8078 4176
rect 9678 5108 9680 5128
rect 9680 5108 9732 5128
rect 9732 5108 9734 5128
rect 9678 5072 9734 5108
rect 9477 4922 9533 4924
rect 9557 4922 9613 4924
rect 9637 4922 9693 4924
rect 9717 4922 9773 4924
rect 9477 4870 9523 4922
rect 9523 4870 9533 4922
rect 9557 4870 9587 4922
rect 9587 4870 9599 4922
rect 9599 4870 9613 4922
rect 9637 4870 9651 4922
rect 9651 4870 9663 4922
rect 9663 4870 9693 4922
rect 9717 4870 9727 4922
rect 9727 4870 9773 4922
rect 9477 4868 9533 4870
rect 9557 4868 9613 4870
rect 9637 4868 9693 4870
rect 9717 4868 9773 4870
rect 8666 3984 8722 4040
rect 10138 5752 10194 5808
rect 11150 7248 11206 7304
rect 10874 5752 10930 5808
rect 12317 16346 12373 16348
rect 12397 16346 12453 16348
rect 12477 16346 12533 16348
rect 12557 16346 12613 16348
rect 12317 16294 12363 16346
rect 12363 16294 12373 16346
rect 12397 16294 12427 16346
rect 12427 16294 12439 16346
rect 12439 16294 12453 16346
rect 12477 16294 12491 16346
rect 12491 16294 12503 16346
rect 12503 16294 12533 16346
rect 12557 16294 12567 16346
rect 12567 16294 12613 16346
rect 12317 16292 12373 16294
rect 12397 16292 12453 16294
rect 12477 16292 12533 16294
rect 12557 16292 12613 16294
rect 12317 15258 12373 15260
rect 12397 15258 12453 15260
rect 12477 15258 12533 15260
rect 12557 15258 12613 15260
rect 12317 15206 12363 15258
rect 12363 15206 12373 15258
rect 12397 15206 12427 15258
rect 12427 15206 12439 15258
rect 12439 15206 12453 15258
rect 12477 15206 12491 15258
rect 12491 15206 12503 15258
rect 12503 15206 12533 15258
rect 12557 15206 12567 15258
rect 12567 15206 12613 15258
rect 12317 15204 12373 15206
rect 12397 15204 12453 15206
rect 12477 15204 12533 15206
rect 12557 15204 12613 15206
rect 13082 20712 13138 20768
rect 13358 20576 13414 20632
rect 13266 19932 13268 19952
rect 13268 19932 13320 19952
rect 13320 19932 13322 19952
rect 13266 19896 13322 19932
rect 13634 20324 13690 20360
rect 13634 20304 13636 20324
rect 13636 20304 13688 20324
rect 13688 20304 13690 20324
rect 12317 14170 12373 14172
rect 12397 14170 12453 14172
rect 12477 14170 12533 14172
rect 12557 14170 12613 14172
rect 12317 14118 12363 14170
rect 12363 14118 12373 14170
rect 12397 14118 12427 14170
rect 12427 14118 12439 14170
rect 12439 14118 12453 14170
rect 12477 14118 12491 14170
rect 12491 14118 12503 14170
rect 12503 14118 12533 14170
rect 12557 14118 12567 14170
rect 12567 14118 12613 14170
rect 12317 14116 12373 14118
rect 12397 14116 12453 14118
rect 12477 14116 12533 14118
rect 12557 14116 12613 14118
rect 12317 13082 12373 13084
rect 12397 13082 12453 13084
rect 12477 13082 12533 13084
rect 12557 13082 12613 13084
rect 12317 13030 12363 13082
rect 12363 13030 12373 13082
rect 12397 13030 12427 13082
rect 12427 13030 12439 13082
rect 12439 13030 12453 13082
rect 12477 13030 12491 13082
rect 12491 13030 12503 13082
rect 12503 13030 12533 13082
rect 12557 13030 12567 13082
rect 12567 13030 12613 13082
rect 12317 13028 12373 13030
rect 12397 13028 12453 13030
rect 12477 13028 12533 13030
rect 12557 13028 12613 13030
rect 13082 14048 13138 14104
rect 12317 11994 12373 11996
rect 12397 11994 12453 11996
rect 12477 11994 12533 11996
rect 12557 11994 12613 11996
rect 12317 11942 12363 11994
rect 12363 11942 12373 11994
rect 12397 11942 12427 11994
rect 12427 11942 12439 11994
rect 12439 11942 12453 11994
rect 12477 11942 12491 11994
rect 12491 11942 12503 11994
rect 12503 11942 12533 11994
rect 12557 11942 12567 11994
rect 12567 11942 12613 11994
rect 12317 11940 12373 11942
rect 12397 11940 12453 11942
rect 12477 11940 12533 11942
rect 12557 11940 12613 11942
rect 12622 11736 12678 11792
rect 12317 10906 12373 10908
rect 12397 10906 12453 10908
rect 12477 10906 12533 10908
rect 12557 10906 12613 10908
rect 12317 10854 12363 10906
rect 12363 10854 12373 10906
rect 12397 10854 12427 10906
rect 12427 10854 12439 10906
rect 12439 10854 12453 10906
rect 12477 10854 12491 10906
rect 12491 10854 12503 10906
rect 12503 10854 12533 10906
rect 12557 10854 12567 10906
rect 12567 10854 12613 10906
rect 12317 10852 12373 10854
rect 12397 10852 12453 10854
rect 12477 10852 12533 10854
rect 12557 10852 12613 10854
rect 13174 12316 13176 12336
rect 13176 12316 13228 12336
rect 13228 12316 13230 12336
rect 13174 12280 13230 12316
rect 13082 10920 13138 10976
rect 12317 9818 12373 9820
rect 12397 9818 12453 9820
rect 12477 9818 12533 9820
rect 12557 9818 12613 9820
rect 12317 9766 12363 9818
rect 12363 9766 12373 9818
rect 12397 9766 12427 9818
rect 12427 9766 12439 9818
rect 12439 9766 12453 9818
rect 12477 9766 12491 9818
rect 12491 9766 12503 9818
rect 12503 9766 12533 9818
rect 12557 9766 12567 9818
rect 12567 9766 12613 9818
rect 12317 9764 12373 9766
rect 12397 9764 12453 9766
rect 12477 9764 12533 9766
rect 12557 9764 12613 9766
rect 12317 8730 12373 8732
rect 12397 8730 12453 8732
rect 12477 8730 12533 8732
rect 12557 8730 12613 8732
rect 12317 8678 12363 8730
rect 12363 8678 12373 8730
rect 12397 8678 12427 8730
rect 12427 8678 12439 8730
rect 12439 8678 12453 8730
rect 12477 8678 12491 8730
rect 12491 8678 12503 8730
rect 12503 8678 12533 8730
rect 12557 8678 12567 8730
rect 12567 8678 12613 8730
rect 12317 8676 12373 8678
rect 12397 8676 12453 8678
rect 12477 8676 12533 8678
rect 12557 8676 12613 8678
rect 12317 7642 12373 7644
rect 12397 7642 12453 7644
rect 12477 7642 12533 7644
rect 12557 7642 12613 7644
rect 12317 7590 12363 7642
rect 12363 7590 12373 7642
rect 12397 7590 12427 7642
rect 12427 7590 12439 7642
rect 12439 7590 12453 7642
rect 12477 7590 12491 7642
rect 12491 7590 12503 7642
rect 12503 7590 12533 7642
rect 12557 7590 12567 7642
rect 12567 7590 12613 7642
rect 12317 7588 12373 7590
rect 12397 7588 12453 7590
rect 12477 7588 12533 7590
rect 12557 7588 12613 7590
rect 13450 10784 13506 10840
rect 14462 20712 14518 20768
rect 15158 21242 15214 21244
rect 15238 21242 15294 21244
rect 15318 21242 15374 21244
rect 15398 21242 15454 21244
rect 15158 21190 15204 21242
rect 15204 21190 15214 21242
rect 15238 21190 15268 21242
rect 15268 21190 15280 21242
rect 15280 21190 15294 21242
rect 15318 21190 15332 21242
rect 15332 21190 15344 21242
rect 15344 21190 15374 21242
rect 15398 21190 15408 21242
rect 15408 21190 15454 21242
rect 15158 21188 15214 21190
rect 15238 21188 15294 21190
rect 15318 21188 15374 21190
rect 15398 21188 15454 21190
rect 16210 21528 16266 21584
rect 17998 21786 18054 21788
rect 18078 21786 18134 21788
rect 18158 21786 18214 21788
rect 18238 21786 18294 21788
rect 17998 21734 18044 21786
rect 18044 21734 18054 21786
rect 18078 21734 18108 21786
rect 18108 21734 18120 21786
rect 18120 21734 18134 21786
rect 18158 21734 18172 21786
rect 18172 21734 18184 21786
rect 18184 21734 18214 21786
rect 18238 21734 18248 21786
rect 18248 21734 18294 21786
rect 17998 21732 18054 21734
rect 18078 21732 18134 21734
rect 18158 21732 18214 21734
rect 18238 21732 18294 21734
rect 15158 20154 15214 20156
rect 15238 20154 15294 20156
rect 15318 20154 15374 20156
rect 15398 20154 15454 20156
rect 15158 20102 15204 20154
rect 15204 20102 15214 20154
rect 15238 20102 15268 20154
rect 15268 20102 15280 20154
rect 15280 20102 15294 20154
rect 15318 20102 15332 20154
rect 15332 20102 15344 20154
rect 15344 20102 15374 20154
rect 15398 20102 15408 20154
rect 15408 20102 15454 20154
rect 15158 20100 15214 20102
rect 15238 20100 15294 20102
rect 15318 20100 15374 20102
rect 15398 20100 15454 20102
rect 15290 19932 15292 19952
rect 15292 19932 15344 19952
rect 15344 19932 15346 19952
rect 15290 19896 15346 19932
rect 15382 19760 15438 19816
rect 15198 19372 15254 19408
rect 15198 19352 15200 19372
rect 15200 19352 15252 19372
rect 15252 19352 15254 19372
rect 15750 19488 15806 19544
rect 15158 19066 15214 19068
rect 15238 19066 15294 19068
rect 15318 19066 15374 19068
rect 15398 19066 15454 19068
rect 15158 19014 15204 19066
rect 15204 19014 15214 19066
rect 15238 19014 15268 19066
rect 15268 19014 15280 19066
rect 15280 19014 15294 19066
rect 15318 19014 15332 19066
rect 15332 19014 15344 19066
rect 15344 19014 15374 19066
rect 15398 19014 15408 19066
rect 15408 19014 15454 19066
rect 15158 19012 15214 19014
rect 15238 19012 15294 19014
rect 15318 19012 15374 19014
rect 15398 19012 15454 19014
rect 15158 17978 15214 17980
rect 15238 17978 15294 17980
rect 15318 17978 15374 17980
rect 15398 17978 15454 17980
rect 15158 17926 15204 17978
rect 15204 17926 15214 17978
rect 15238 17926 15268 17978
rect 15268 17926 15280 17978
rect 15280 17926 15294 17978
rect 15318 17926 15332 17978
rect 15332 17926 15344 17978
rect 15344 17926 15374 17978
rect 15398 17926 15408 17978
rect 15408 17926 15454 17978
rect 15158 17924 15214 17926
rect 15238 17924 15294 17926
rect 15318 17924 15374 17926
rect 15398 17924 15454 17926
rect 15158 16890 15214 16892
rect 15238 16890 15294 16892
rect 15318 16890 15374 16892
rect 15398 16890 15454 16892
rect 15158 16838 15204 16890
rect 15204 16838 15214 16890
rect 15238 16838 15268 16890
rect 15268 16838 15280 16890
rect 15280 16838 15294 16890
rect 15318 16838 15332 16890
rect 15332 16838 15344 16890
rect 15344 16838 15374 16890
rect 15398 16838 15408 16890
rect 15408 16838 15454 16890
rect 15158 16836 15214 16838
rect 15238 16836 15294 16838
rect 15318 16836 15374 16838
rect 15398 16836 15454 16838
rect 15158 15802 15214 15804
rect 15238 15802 15294 15804
rect 15318 15802 15374 15804
rect 15398 15802 15454 15804
rect 15158 15750 15204 15802
rect 15204 15750 15214 15802
rect 15238 15750 15268 15802
rect 15268 15750 15280 15802
rect 15280 15750 15294 15802
rect 15318 15750 15332 15802
rect 15332 15750 15344 15802
rect 15344 15750 15374 15802
rect 15398 15750 15408 15802
rect 15408 15750 15454 15802
rect 15158 15748 15214 15750
rect 15238 15748 15294 15750
rect 15318 15748 15374 15750
rect 15398 15748 15454 15750
rect 14278 12180 14280 12200
rect 14280 12180 14332 12200
rect 14332 12180 14334 12200
rect 14278 12144 14334 12180
rect 14278 11092 14280 11112
rect 14280 11092 14332 11112
rect 14332 11092 14334 11112
rect 14278 11056 14334 11092
rect 14186 10920 14242 10976
rect 13910 10784 13966 10840
rect 11978 6568 12034 6624
rect 11702 5908 11758 5944
rect 11702 5888 11704 5908
rect 11704 5888 11756 5908
rect 11756 5888 11758 5908
rect 9477 3834 9533 3836
rect 9557 3834 9613 3836
rect 9637 3834 9693 3836
rect 9717 3834 9773 3836
rect 9477 3782 9523 3834
rect 9523 3782 9533 3834
rect 9557 3782 9587 3834
rect 9587 3782 9599 3834
rect 9599 3782 9613 3834
rect 9637 3782 9651 3834
rect 9651 3782 9663 3834
rect 9663 3782 9693 3834
rect 9717 3782 9727 3834
rect 9727 3782 9773 3834
rect 9477 3780 9533 3782
rect 9557 3780 9613 3782
rect 9637 3780 9693 3782
rect 9717 3780 9773 3782
rect 10966 3032 11022 3088
rect 11058 2896 11114 2952
rect 12162 6568 12218 6624
rect 12317 6554 12373 6556
rect 12397 6554 12453 6556
rect 12477 6554 12533 6556
rect 12557 6554 12613 6556
rect 12317 6502 12363 6554
rect 12363 6502 12373 6554
rect 12397 6502 12427 6554
rect 12427 6502 12439 6554
rect 12439 6502 12453 6554
rect 12477 6502 12491 6554
rect 12491 6502 12503 6554
rect 12503 6502 12533 6554
rect 12557 6502 12567 6554
rect 12567 6502 12613 6554
rect 12317 6500 12373 6502
rect 12397 6500 12453 6502
rect 12477 6500 12533 6502
rect 12557 6500 12613 6502
rect 14738 11192 14794 11248
rect 15750 17992 15806 18048
rect 15158 14714 15214 14716
rect 15238 14714 15294 14716
rect 15318 14714 15374 14716
rect 15398 14714 15454 14716
rect 15158 14662 15204 14714
rect 15204 14662 15214 14714
rect 15238 14662 15268 14714
rect 15268 14662 15280 14714
rect 15280 14662 15294 14714
rect 15318 14662 15332 14714
rect 15332 14662 15344 14714
rect 15344 14662 15374 14714
rect 15398 14662 15408 14714
rect 15408 14662 15454 14714
rect 15158 14660 15214 14662
rect 15238 14660 15294 14662
rect 15318 14660 15374 14662
rect 15398 14660 15454 14662
rect 15158 13626 15214 13628
rect 15238 13626 15294 13628
rect 15318 13626 15374 13628
rect 15398 13626 15454 13628
rect 15158 13574 15204 13626
rect 15204 13574 15214 13626
rect 15238 13574 15268 13626
rect 15268 13574 15280 13626
rect 15280 13574 15294 13626
rect 15318 13574 15332 13626
rect 15332 13574 15344 13626
rect 15344 13574 15374 13626
rect 15398 13574 15408 13626
rect 15408 13574 15454 13626
rect 15158 13572 15214 13574
rect 15238 13572 15294 13574
rect 15318 13572 15374 13574
rect 15398 13572 15454 13574
rect 15158 12538 15214 12540
rect 15238 12538 15294 12540
rect 15318 12538 15374 12540
rect 15398 12538 15454 12540
rect 15158 12486 15204 12538
rect 15204 12486 15214 12538
rect 15238 12486 15268 12538
rect 15268 12486 15280 12538
rect 15280 12486 15294 12538
rect 15318 12486 15332 12538
rect 15332 12486 15344 12538
rect 15344 12486 15374 12538
rect 15398 12486 15408 12538
rect 15408 12486 15454 12538
rect 15158 12484 15214 12486
rect 15238 12484 15294 12486
rect 15318 12484 15374 12486
rect 15398 12484 15454 12486
rect 15106 11772 15108 11792
rect 15108 11772 15160 11792
rect 15160 11772 15162 11792
rect 15106 11736 15162 11772
rect 15158 11450 15214 11452
rect 15238 11450 15294 11452
rect 15318 11450 15374 11452
rect 15398 11450 15454 11452
rect 15158 11398 15204 11450
rect 15204 11398 15214 11450
rect 15238 11398 15268 11450
rect 15268 11398 15280 11450
rect 15280 11398 15294 11450
rect 15318 11398 15332 11450
rect 15332 11398 15344 11450
rect 15344 11398 15374 11450
rect 15398 11398 15408 11450
rect 15408 11398 15454 11450
rect 15158 11396 15214 11398
rect 15238 11396 15294 11398
rect 15318 11396 15374 11398
rect 15398 11396 15454 11398
rect 14922 11192 14978 11248
rect 14922 11092 14924 11112
rect 14924 11092 14976 11112
rect 14976 11092 14978 11112
rect 14922 11056 14978 11092
rect 15106 10784 15162 10840
rect 15658 14048 15714 14104
rect 16026 16768 16082 16824
rect 16670 20304 16726 20360
rect 17998 20698 18054 20700
rect 18078 20698 18134 20700
rect 18158 20698 18214 20700
rect 18238 20698 18294 20700
rect 17998 20646 18044 20698
rect 18044 20646 18054 20698
rect 18078 20646 18108 20698
rect 18108 20646 18120 20698
rect 18120 20646 18134 20698
rect 18158 20646 18172 20698
rect 18172 20646 18184 20698
rect 18184 20646 18214 20698
rect 18238 20646 18248 20698
rect 18248 20646 18294 20698
rect 17998 20644 18054 20646
rect 18078 20644 18134 20646
rect 18158 20644 18214 20646
rect 18238 20644 18294 20646
rect 17866 20596 17922 20632
rect 17866 20576 17868 20596
rect 17868 20576 17920 20596
rect 17920 20576 17922 20596
rect 16854 19780 16910 19816
rect 16854 19760 16856 19780
rect 16856 19760 16908 19780
rect 16908 19760 16910 19780
rect 16762 19352 16818 19408
rect 17130 19488 17186 19544
rect 17314 19372 17370 19408
rect 17314 19352 17316 19372
rect 17316 19352 17368 19372
rect 17368 19352 17370 19372
rect 15934 13776 15990 13832
rect 16118 12960 16174 13016
rect 15934 12824 15990 12880
rect 15566 10920 15622 10976
rect 12898 7248 12954 7304
rect 12622 6180 12678 6216
rect 12622 6160 12624 6180
rect 12624 6160 12676 6180
rect 12676 6160 12678 6180
rect 12254 5752 12310 5808
rect 12317 5466 12373 5468
rect 12397 5466 12453 5468
rect 12477 5466 12533 5468
rect 12557 5466 12613 5468
rect 12317 5414 12363 5466
rect 12363 5414 12373 5466
rect 12397 5414 12427 5466
rect 12427 5414 12439 5466
rect 12439 5414 12453 5466
rect 12477 5414 12491 5466
rect 12491 5414 12503 5466
rect 12503 5414 12533 5466
rect 12557 5414 12567 5466
rect 12567 5414 12613 5466
rect 12317 5412 12373 5414
rect 12397 5412 12453 5414
rect 12477 5412 12533 5414
rect 12557 5412 12613 5414
rect 13634 6704 13690 6760
rect 12317 4378 12373 4380
rect 12397 4378 12453 4380
rect 12477 4378 12533 4380
rect 12557 4378 12613 4380
rect 12317 4326 12363 4378
rect 12363 4326 12373 4378
rect 12397 4326 12427 4378
rect 12427 4326 12439 4378
rect 12439 4326 12453 4378
rect 12477 4326 12491 4378
rect 12491 4326 12503 4378
rect 12503 4326 12533 4378
rect 12557 4326 12567 4378
rect 12567 4326 12613 4378
rect 12317 4324 12373 4326
rect 12397 4324 12453 4326
rect 12477 4324 12533 4326
rect 12557 4324 12613 4326
rect 11702 3984 11758 4040
rect 12317 3290 12373 3292
rect 12397 3290 12453 3292
rect 12477 3290 12533 3292
rect 12557 3290 12613 3292
rect 12317 3238 12363 3290
rect 12363 3238 12373 3290
rect 12397 3238 12427 3290
rect 12427 3238 12439 3290
rect 12439 3238 12453 3290
rect 12477 3238 12491 3290
rect 12491 3238 12503 3290
rect 12503 3238 12533 3290
rect 12557 3238 12567 3290
rect 12567 3238 12613 3290
rect 12317 3236 12373 3238
rect 12397 3236 12453 3238
rect 12477 3236 12533 3238
rect 12557 3236 12613 3238
rect 11242 2916 11298 2952
rect 11242 2896 11244 2916
rect 11244 2896 11296 2916
rect 11296 2896 11298 2916
rect 9477 2746 9533 2748
rect 9557 2746 9613 2748
rect 9637 2746 9693 2748
rect 9717 2746 9773 2748
rect 9477 2694 9523 2746
rect 9523 2694 9533 2746
rect 9557 2694 9587 2746
rect 9587 2694 9599 2746
rect 9599 2694 9613 2746
rect 9637 2694 9651 2746
rect 9651 2694 9663 2746
rect 9663 2694 9693 2746
rect 9717 2694 9727 2746
rect 9727 2694 9773 2746
rect 9477 2692 9533 2694
rect 9557 2692 9613 2694
rect 9637 2692 9693 2694
rect 9717 2692 9773 2694
rect 14278 5228 14334 5264
rect 14278 5208 14280 5228
rect 14280 5208 14332 5228
rect 14332 5208 14334 5228
rect 15158 10362 15214 10364
rect 15238 10362 15294 10364
rect 15318 10362 15374 10364
rect 15398 10362 15454 10364
rect 15158 10310 15204 10362
rect 15204 10310 15214 10362
rect 15238 10310 15268 10362
rect 15268 10310 15280 10362
rect 15280 10310 15294 10362
rect 15318 10310 15332 10362
rect 15332 10310 15344 10362
rect 15344 10310 15374 10362
rect 15398 10310 15408 10362
rect 15408 10310 15454 10362
rect 15158 10308 15214 10310
rect 15238 10308 15294 10310
rect 15318 10308 15374 10310
rect 15398 10308 15454 10310
rect 15158 9274 15214 9276
rect 15238 9274 15294 9276
rect 15318 9274 15374 9276
rect 15398 9274 15454 9276
rect 15158 9222 15204 9274
rect 15204 9222 15214 9274
rect 15238 9222 15268 9274
rect 15268 9222 15280 9274
rect 15280 9222 15294 9274
rect 15318 9222 15332 9274
rect 15332 9222 15344 9274
rect 15344 9222 15374 9274
rect 15398 9222 15408 9274
rect 15408 9222 15454 9274
rect 15158 9220 15214 9222
rect 15238 9220 15294 9222
rect 15318 9220 15374 9222
rect 15398 9220 15454 9222
rect 14738 8472 14794 8528
rect 14830 7928 14886 7984
rect 15158 8186 15214 8188
rect 15238 8186 15294 8188
rect 15318 8186 15374 8188
rect 15398 8186 15454 8188
rect 15158 8134 15204 8186
rect 15204 8134 15214 8186
rect 15238 8134 15268 8186
rect 15268 8134 15280 8186
rect 15280 8134 15294 8186
rect 15318 8134 15332 8186
rect 15332 8134 15344 8186
rect 15344 8134 15374 8186
rect 15398 8134 15408 8186
rect 15408 8134 15454 8186
rect 15158 8132 15214 8134
rect 15238 8132 15294 8134
rect 15318 8132 15374 8134
rect 15398 8132 15454 8134
rect 14830 5888 14886 5944
rect 14554 5072 14610 5128
rect 14830 5072 14886 5128
rect 13634 3304 13690 3360
rect 15158 7098 15214 7100
rect 15238 7098 15294 7100
rect 15318 7098 15374 7100
rect 15398 7098 15454 7100
rect 15158 7046 15204 7098
rect 15204 7046 15214 7098
rect 15238 7046 15268 7098
rect 15268 7046 15280 7098
rect 15280 7046 15294 7098
rect 15318 7046 15332 7098
rect 15332 7046 15344 7098
rect 15344 7046 15374 7098
rect 15398 7046 15408 7098
rect 15408 7046 15454 7098
rect 15158 7044 15214 7046
rect 15238 7044 15294 7046
rect 15318 7044 15374 7046
rect 15398 7044 15454 7046
rect 16946 13096 17002 13152
rect 17222 13912 17278 13968
rect 17314 13368 17370 13424
rect 17130 13232 17186 13288
rect 17222 12144 17278 12200
rect 15158 6010 15214 6012
rect 15238 6010 15294 6012
rect 15318 6010 15374 6012
rect 15398 6010 15454 6012
rect 15158 5958 15204 6010
rect 15204 5958 15214 6010
rect 15238 5958 15268 6010
rect 15268 5958 15280 6010
rect 15280 5958 15294 6010
rect 15318 5958 15332 6010
rect 15332 5958 15344 6010
rect 15344 5958 15374 6010
rect 15398 5958 15408 6010
rect 15408 5958 15454 6010
rect 15158 5956 15214 5958
rect 15238 5956 15294 5958
rect 15318 5956 15374 5958
rect 15398 5956 15454 5958
rect 17406 12688 17462 12744
rect 17998 19610 18054 19612
rect 18078 19610 18134 19612
rect 18158 19610 18214 19612
rect 18238 19610 18294 19612
rect 17998 19558 18044 19610
rect 18044 19558 18054 19610
rect 18078 19558 18108 19610
rect 18108 19558 18120 19610
rect 18120 19558 18134 19610
rect 18158 19558 18172 19610
rect 18172 19558 18184 19610
rect 18184 19558 18214 19610
rect 18238 19558 18248 19610
rect 18248 19558 18294 19610
rect 17998 19556 18054 19558
rect 18078 19556 18134 19558
rect 18158 19556 18214 19558
rect 18238 19556 18294 19558
rect 17998 18522 18054 18524
rect 18078 18522 18134 18524
rect 18158 18522 18214 18524
rect 18238 18522 18294 18524
rect 17998 18470 18044 18522
rect 18044 18470 18054 18522
rect 18078 18470 18108 18522
rect 18108 18470 18120 18522
rect 18120 18470 18134 18522
rect 18158 18470 18172 18522
rect 18172 18470 18184 18522
rect 18184 18470 18214 18522
rect 18238 18470 18248 18522
rect 18248 18470 18294 18522
rect 17998 18468 18054 18470
rect 18078 18468 18134 18470
rect 18158 18468 18214 18470
rect 18238 18468 18294 18470
rect 17998 17434 18054 17436
rect 18078 17434 18134 17436
rect 18158 17434 18214 17436
rect 18238 17434 18294 17436
rect 17998 17382 18044 17434
rect 18044 17382 18054 17434
rect 18078 17382 18108 17434
rect 18108 17382 18120 17434
rect 18120 17382 18134 17434
rect 18158 17382 18172 17434
rect 18172 17382 18184 17434
rect 18184 17382 18214 17434
rect 18238 17382 18248 17434
rect 18248 17382 18294 17434
rect 17998 17380 18054 17382
rect 18078 17380 18134 17382
rect 18158 17380 18214 17382
rect 18238 17380 18294 17382
rect 17774 16496 17830 16552
rect 18050 16496 18106 16552
rect 17998 16346 18054 16348
rect 18078 16346 18134 16348
rect 18158 16346 18214 16348
rect 18238 16346 18294 16348
rect 17998 16294 18044 16346
rect 18044 16294 18054 16346
rect 18078 16294 18108 16346
rect 18108 16294 18120 16346
rect 18120 16294 18134 16346
rect 18158 16294 18172 16346
rect 18172 16294 18184 16346
rect 18184 16294 18214 16346
rect 18238 16294 18248 16346
rect 18248 16294 18294 16346
rect 17998 16292 18054 16294
rect 18078 16292 18134 16294
rect 18158 16292 18214 16294
rect 18238 16292 18294 16294
rect 18418 16108 18474 16144
rect 18418 16088 18420 16108
rect 18420 16088 18472 16108
rect 18472 16088 18474 16108
rect 18510 15952 18566 16008
rect 17998 15258 18054 15260
rect 18078 15258 18134 15260
rect 18158 15258 18214 15260
rect 18238 15258 18294 15260
rect 17998 15206 18044 15258
rect 18044 15206 18054 15258
rect 18078 15206 18108 15258
rect 18108 15206 18120 15258
rect 18120 15206 18134 15258
rect 18158 15206 18172 15258
rect 18172 15206 18184 15258
rect 18184 15206 18214 15258
rect 18238 15206 18248 15258
rect 18248 15206 18294 15258
rect 17998 15204 18054 15206
rect 18078 15204 18134 15206
rect 18158 15204 18214 15206
rect 18238 15204 18294 15206
rect 17998 14170 18054 14172
rect 18078 14170 18134 14172
rect 18158 14170 18214 14172
rect 18238 14170 18294 14172
rect 17998 14118 18044 14170
rect 18044 14118 18054 14170
rect 18078 14118 18108 14170
rect 18108 14118 18120 14170
rect 18120 14118 18134 14170
rect 18158 14118 18172 14170
rect 18172 14118 18184 14170
rect 18184 14118 18214 14170
rect 18238 14118 18248 14170
rect 18248 14118 18294 14170
rect 17998 14116 18054 14118
rect 18078 14116 18134 14118
rect 18158 14116 18214 14118
rect 18238 14116 18294 14118
rect 18234 13932 18290 13968
rect 18234 13912 18236 13932
rect 18236 13912 18288 13932
rect 18288 13912 18290 13932
rect 17682 13096 17738 13152
rect 17590 12960 17646 13016
rect 17998 13082 18054 13084
rect 18078 13082 18134 13084
rect 18158 13082 18214 13084
rect 18238 13082 18294 13084
rect 17998 13030 18044 13082
rect 18044 13030 18054 13082
rect 18078 13030 18108 13082
rect 18108 13030 18120 13082
rect 18120 13030 18134 13082
rect 18158 13030 18172 13082
rect 18172 13030 18184 13082
rect 18184 13030 18214 13082
rect 18238 13030 18248 13082
rect 18248 13030 18294 13082
rect 17998 13028 18054 13030
rect 18078 13028 18134 13030
rect 18158 13028 18214 13030
rect 18238 13028 18294 13030
rect 17866 12688 17922 12744
rect 17498 10004 17500 10024
rect 17500 10004 17552 10024
rect 17552 10004 17554 10024
rect 17498 9968 17554 10004
rect 16026 5752 16082 5808
rect 15158 4922 15214 4924
rect 15238 4922 15294 4924
rect 15318 4922 15374 4924
rect 15398 4922 15454 4924
rect 15158 4870 15204 4922
rect 15204 4870 15214 4922
rect 15238 4870 15268 4922
rect 15268 4870 15280 4922
rect 15280 4870 15294 4922
rect 15318 4870 15332 4922
rect 15332 4870 15344 4922
rect 15344 4870 15374 4922
rect 15398 4870 15408 4922
rect 15408 4870 15454 4922
rect 15158 4868 15214 4870
rect 15238 4868 15294 4870
rect 15318 4868 15374 4870
rect 15398 4868 15454 4870
rect 16670 5208 16726 5264
rect 15158 3834 15214 3836
rect 15238 3834 15294 3836
rect 15318 3834 15374 3836
rect 15398 3834 15454 3836
rect 15158 3782 15204 3834
rect 15204 3782 15214 3834
rect 15238 3782 15268 3834
rect 15268 3782 15280 3834
rect 15280 3782 15294 3834
rect 15318 3782 15332 3834
rect 15332 3782 15344 3834
rect 15344 3782 15374 3834
rect 15398 3782 15408 3834
rect 15408 3782 15454 3834
rect 15158 3780 15214 3782
rect 15238 3780 15294 3782
rect 15318 3780 15374 3782
rect 15398 3780 15454 3782
rect 14830 3440 14886 3496
rect 16118 4140 16174 4176
rect 16118 4120 16120 4140
rect 16120 4120 16172 4140
rect 16172 4120 16174 4140
rect 16578 3576 16634 3632
rect 16946 3476 16948 3496
rect 16948 3476 17000 3496
rect 17000 3476 17002 3496
rect 16946 3440 17002 3476
rect 17038 3052 17094 3088
rect 17998 11994 18054 11996
rect 18078 11994 18134 11996
rect 18158 11994 18214 11996
rect 18238 11994 18294 11996
rect 17998 11942 18044 11994
rect 18044 11942 18054 11994
rect 18078 11942 18108 11994
rect 18108 11942 18120 11994
rect 18120 11942 18134 11994
rect 18158 11942 18172 11994
rect 18172 11942 18184 11994
rect 18184 11942 18214 11994
rect 18238 11942 18248 11994
rect 18248 11942 18294 11994
rect 17998 11940 18054 11942
rect 18078 11940 18134 11942
rect 18158 11940 18214 11942
rect 18238 11940 18294 11942
rect 18234 11092 18236 11112
rect 18236 11092 18288 11112
rect 18288 11092 18290 11112
rect 18234 11056 18290 11092
rect 17998 10906 18054 10908
rect 18078 10906 18134 10908
rect 18158 10906 18214 10908
rect 18238 10906 18294 10908
rect 17998 10854 18044 10906
rect 18044 10854 18054 10906
rect 18078 10854 18108 10906
rect 18108 10854 18120 10906
rect 18120 10854 18134 10906
rect 18158 10854 18172 10906
rect 18172 10854 18184 10906
rect 18184 10854 18214 10906
rect 18238 10854 18248 10906
rect 18248 10854 18294 10906
rect 17998 10852 18054 10854
rect 18078 10852 18134 10854
rect 18158 10852 18214 10854
rect 18238 10852 18294 10854
rect 20839 21242 20895 21244
rect 20919 21242 20975 21244
rect 20999 21242 21055 21244
rect 21079 21242 21135 21244
rect 20839 21190 20885 21242
rect 20885 21190 20895 21242
rect 20919 21190 20949 21242
rect 20949 21190 20961 21242
rect 20961 21190 20975 21242
rect 20999 21190 21013 21242
rect 21013 21190 21025 21242
rect 21025 21190 21055 21242
rect 21079 21190 21089 21242
rect 21089 21190 21135 21242
rect 20839 21188 20895 21190
rect 20919 21188 20975 21190
rect 20999 21188 21055 21190
rect 21079 21188 21135 21190
rect 23679 21786 23735 21788
rect 23759 21786 23815 21788
rect 23839 21786 23895 21788
rect 23919 21786 23975 21788
rect 23679 21734 23725 21786
rect 23725 21734 23735 21786
rect 23759 21734 23789 21786
rect 23789 21734 23801 21786
rect 23801 21734 23815 21786
rect 23839 21734 23853 21786
rect 23853 21734 23865 21786
rect 23865 21734 23895 21786
rect 23919 21734 23929 21786
rect 23929 21734 23975 21786
rect 23679 21732 23735 21734
rect 23759 21732 23815 21734
rect 23839 21732 23895 21734
rect 23919 21732 23975 21734
rect 23679 20698 23735 20700
rect 23759 20698 23815 20700
rect 23839 20698 23895 20700
rect 23919 20698 23975 20700
rect 23679 20646 23725 20698
rect 23725 20646 23735 20698
rect 23759 20646 23789 20698
rect 23789 20646 23801 20698
rect 23801 20646 23815 20698
rect 23839 20646 23853 20698
rect 23853 20646 23865 20698
rect 23865 20646 23895 20698
rect 23919 20646 23929 20698
rect 23929 20646 23975 20698
rect 23679 20644 23735 20646
rect 23759 20644 23815 20646
rect 23839 20644 23895 20646
rect 23919 20644 23975 20646
rect 18970 16768 19026 16824
rect 18602 13368 18658 13424
rect 18602 11192 18658 11248
rect 18510 11056 18566 11112
rect 19338 14612 19394 14648
rect 19338 14592 19340 14612
rect 19340 14592 19392 14612
rect 19392 14592 19394 14612
rect 18694 10648 18750 10704
rect 17998 9818 18054 9820
rect 18078 9818 18134 9820
rect 18158 9818 18214 9820
rect 18238 9818 18294 9820
rect 17998 9766 18044 9818
rect 18044 9766 18054 9818
rect 18078 9766 18108 9818
rect 18108 9766 18120 9818
rect 18120 9766 18134 9818
rect 18158 9766 18172 9818
rect 18172 9766 18184 9818
rect 18184 9766 18214 9818
rect 18238 9766 18248 9818
rect 18248 9766 18294 9818
rect 17998 9764 18054 9766
rect 18078 9764 18134 9766
rect 18158 9764 18214 9766
rect 18238 9764 18294 9766
rect 17998 8730 18054 8732
rect 18078 8730 18134 8732
rect 18158 8730 18214 8732
rect 18238 8730 18294 8732
rect 17998 8678 18044 8730
rect 18044 8678 18054 8730
rect 18078 8678 18108 8730
rect 18108 8678 18120 8730
rect 18120 8678 18134 8730
rect 18158 8678 18172 8730
rect 18172 8678 18184 8730
rect 18184 8678 18214 8730
rect 18238 8678 18248 8730
rect 18248 8678 18294 8730
rect 17998 8676 18054 8678
rect 18078 8676 18134 8678
rect 18158 8676 18214 8678
rect 18238 8676 18294 8678
rect 18234 8492 18290 8528
rect 18234 8472 18236 8492
rect 18236 8472 18288 8492
rect 18288 8472 18290 8492
rect 17998 7642 18054 7644
rect 18078 7642 18134 7644
rect 18158 7642 18214 7644
rect 18238 7642 18294 7644
rect 17998 7590 18044 7642
rect 18044 7590 18054 7642
rect 18078 7590 18108 7642
rect 18108 7590 18120 7642
rect 18120 7590 18134 7642
rect 18158 7590 18172 7642
rect 18172 7590 18184 7642
rect 18184 7590 18214 7642
rect 18238 7590 18248 7642
rect 18248 7590 18294 7642
rect 17998 7588 18054 7590
rect 18078 7588 18134 7590
rect 18158 7588 18214 7590
rect 18238 7588 18294 7590
rect 17998 6554 18054 6556
rect 18078 6554 18134 6556
rect 18158 6554 18214 6556
rect 18238 6554 18294 6556
rect 17998 6502 18044 6554
rect 18044 6502 18054 6554
rect 18078 6502 18108 6554
rect 18108 6502 18120 6554
rect 18120 6502 18134 6554
rect 18158 6502 18172 6554
rect 18172 6502 18184 6554
rect 18184 6502 18214 6554
rect 18238 6502 18248 6554
rect 18248 6502 18294 6554
rect 17998 6500 18054 6502
rect 18078 6500 18134 6502
rect 18158 6500 18214 6502
rect 18238 6500 18294 6502
rect 17958 6316 18014 6352
rect 17958 6296 17960 6316
rect 17960 6296 18012 6316
rect 18012 6296 18014 6316
rect 19062 10648 19118 10704
rect 17998 5466 18054 5468
rect 18078 5466 18134 5468
rect 18158 5466 18214 5468
rect 18238 5466 18294 5468
rect 17998 5414 18044 5466
rect 18044 5414 18054 5466
rect 18078 5414 18108 5466
rect 18108 5414 18120 5466
rect 18120 5414 18134 5466
rect 18158 5414 18172 5466
rect 18172 5414 18184 5466
rect 18184 5414 18214 5466
rect 18238 5414 18248 5466
rect 18248 5414 18294 5466
rect 17998 5412 18054 5414
rect 18078 5412 18134 5414
rect 18158 5412 18214 5414
rect 18238 5412 18294 5414
rect 17998 4378 18054 4380
rect 18078 4378 18134 4380
rect 18158 4378 18214 4380
rect 18238 4378 18294 4380
rect 17998 4326 18044 4378
rect 18044 4326 18054 4378
rect 18078 4326 18108 4378
rect 18108 4326 18120 4378
rect 18120 4326 18134 4378
rect 18158 4326 18172 4378
rect 18172 4326 18184 4378
rect 18184 4326 18214 4378
rect 18238 4326 18248 4378
rect 18248 4326 18294 4378
rect 17998 4324 18054 4326
rect 18078 4324 18134 4326
rect 18158 4324 18214 4326
rect 18238 4324 18294 4326
rect 20839 20154 20895 20156
rect 20919 20154 20975 20156
rect 20999 20154 21055 20156
rect 21079 20154 21135 20156
rect 20839 20102 20885 20154
rect 20885 20102 20895 20154
rect 20919 20102 20949 20154
rect 20949 20102 20961 20154
rect 20961 20102 20975 20154
rect 20999 20102 21013 20154
rect 21013 20102 21025 20154
rect 21025 20102 21055 20154
rect 21079 20102 21089 20154
rect 21089 20102 21135 20154
rect 20839 20100 20895 20102
rect 20919 20100 20975 20102
rect 20999 20100 21055 20102
rect 21079 20100 21135 20102
rect 20839 19066 20895 19068
rect 20919 19066 20975 19068
rect 20999 19066 21055 19068
rect 21079 19066 21135 19068
rect 20839 19014 20885 19066
rect 20885 19014 20895 19066
rect 20919 19014 20949 19066
rect 20949 19014 20961 19066
rect 20961 19014 20975 19066
rect 20999 19014 21013 19066
rect 21013 19014 21025 19066
rect 21025 19014 21055 19066
rect 21079 19014 21089 19066
rect 21089 19014 21135 19066
rect 20839 19012 20895 19014
rect 20919 19012 20975 19014
rect 20999 19012 21055 19014
rect 21079 19012 21135 19014
rect 19890 13912 19946 13968
rect 19614 13524 19670 13560
rect 19614 13504 19616 13524
rect 19616 13504 19668 13524
rect 19668 13504 19670 13524
rect 19706 13096 19762 13152
rect 20350 13096 20406 13152
rect 20258 12552 20314 12608
rect 19154 6316 19210 6352
rect 19154 6296 19156 6316
rect 19156 6296 19208 6316
rect 19208 6296 19210 6316
rect 20902 18128 20958 18184
rect 20839 17978 20895 17980
rect 20919 17978 20975 17980
rect 20999 17978 21055 17980
rect 21079 17978 21135 17980
rect 20839 17926 20885 17978
rect 20885 17926 20895 17978
rect 20919 17926 20949 17978
rect 20949 17926 20961 17978
rect 20961 17926 20975 17978
rect 20999 17926 21013 17978
rect 21013 17926 21025 17978
rect 21025 17926 21055 17978
rect 21079 17926 21089 17978
rect 21089 17926 21135 17978
rect 20839 17924 20895 17926
rect 20919 17924 20975 17926
rect 20999 17924 21055 17926
rect 21079 17924 21135 17926
rect 20839 16890 20895 16892
rect 20919 16890 20975 16892
rect 20999 16890 21055 16892
rect 21079 16890 21135 16892
rect 20839 16838 20885 16890
rect 20885 16838 20895 16890
rect 20919 16838 20949 16890
rect 20949 16838 20961 16890
rect 20961 16838 20975 16890
rect 20999 16838 21013 16890
rect 21013 16838 21025 16890
rect 21025 16838 21055 16890
rect 21079 16838 21089 16890
rect 21089 16838 21135 16890
rect 20839 16836 20895 16838
rect 20919 16836 20975 16838
rect 20999 16836 21055 16838
rect 21079 16836 21135 16838
rect 20810 16124 20812 16144
rect 20812 16124 20864 16144
rect 20864 16124 20866 16144
rect 20810 16088 20866 16124
rect 20839 15802 20895 15804
rect 20919 15802 20975 15804
rect 20999 15802 21055 15804
rect 21079 15802 21135 15804
rect 20839 15750 20885 15802
rect 20885 15750 20895 15802
rect 20919 15750 20949 15802
rect 20949 15750 20961 15802
rect 20961 15750 20975 15802
rect 20999 15750 21013 15802
rect 21013 15750 21025 15802
rect 21025 15750 21055 15802
rect 21079 15750 21089 15802
rect 21089 15750 21135 15802
rect 20839 15748 20895 15750
rect 20919 15748 20975 15750
rect 20999 15748 21055 15750
rect 21079 15748 21135 15750
rect 20839 14714 20895 14716
rect 20919 14714 20975 14716
rect 20999 14714 21055 14716
rect 21079 14714 21135 14716
rect 20839 14662 20885 14714
rect 20885 14662 20895 14714
rect 20919 14662 20949 14714
rect 20949 14662 20961 14714
rect 20961 14662 20975 14714
rect 20999 14662 21013 14714
rect 21013 14662 21025 14714
rect 21025 14662 21055 14714
rect 21079 14662 21089 14714
rect 21089 14662 21135 14714
rect 20839 14660 20895 14662
rect 20919 14660 20975 14662
rect 20999 14660 21055 14662
rect 21079 14660 21135 14662
rect 20994 13932 21050 13968
rect 20994 13912 20996 13932
rect 20996 13912 21048 13932
rect 21048 13912 21050 13932
rect 20839 13626 20895 13628
rect 20919 13626 20975 13628
rect 20999 13626 21055 13628
rect 21079 13626 21135 13628
rect 20839 13574 20885 13626
rect 20885 13574 20895 13626
rect 20919 13574 20949 13626
rect 20949 13574 20961 13626
rect 20961 13574 20975 13626
rect 20999 13574 21013 13626
rect 21013 13574 21025 13626
rect 21025 13574 21055 13626
rect 21079 13574 21089 13626
rect 21089 13574 21135 13626
rect 20839 13572 20895 13574
rect 20919 13572 20975 13574
rect 20999 13572 21055 13574
rect 21079 13572 21135 13574
rect 22006 16088 22062 16144
rect 21270 12844 21326 12880
rect 21270 12824 21272 12844
rect 21272 12824 21324 12844
rect 21324 12824 21326 12844
rect 20839 12538 20895 12540
rect 20919 12538 20975 12540
rect 20999 12538 21055 12540
rect 21079 12538 21135 12540
rect 20839 12486 20885 12538
rect 20885 12486 20895 12538
rect 20919 12486 20949 12538
rect 20949 12486 20961 12538
rect 20961 12486 20975 12538
rect 20999 12486 21013 12538
rect 21013 12486 21025 12538
rect 21025 12486 21055 12538
rect 21079 12486 21089 12538
rect 21089 12486 21135 12538
rect 20839 12484 20895 12486
rect 20919 12484 20975 12486
rect 20999 12484 21055 12486
rect 21079 12484 21135 12486
rect 21546 12164 21602 12200
rect 21546 12144 21548 12164
rect 21548 12144 21600 12164
rect 21600 12144 21602 12164
rect 20839 11450 20895 11452
rect 20919 11450 20975 11452
rect 20999 11450 21055 11452
rect 21079 11450 21135 11452
rect 20839 11398 20885 11450
rect 20885 11398 20895 11450
rect 20919 11398 20949 11450
rect 20949 11398 20961 11450
rect 20961 11398 20975 11450
rect 20999 11398 21013 11450
rect 21013 11398 21025 11450
rect 21025 11398 21055 11450
rect 21079 11398 21089 11450
rect 21089 11398 21135 11450
rect 20839 11396 20895 11398
rect 20919 11396 20975 11398
rect 20999 11396 21055 11398
rect 21079 11396 21135 11398
rect 21178 11228 21180 11248
rect 21180 11228 21232 11248
rect 21232 11228 21234 11248
rect 21178 11192 21234 11228
rect 17998 3290 18054 3292
rect 18078 3290 18134 3292
rect 18158 3290 18214 3292
rect 18238 3290 18294 3292
rect 17998 3238 18044 3290
rect 18044 3238 18054 3290
rect 18078 3238 18108 3290
rect 18108 3238 18120 3290
rect 18120 3238 18134 3290
rect 18158 3238 18172 3290
rect 18172 3238 18184 3290
rect 18184 3238 18214 3290
rect 18238 3238 18248 3290
rect 18248 3238 18294 3290
rect 17998 3236 18054 3238
rect 18078 3236 18134 3238
rect 18158 3236 18214 3238
rect 18238 3236 18294 3238
rect 17038 3032 17040 3052
rect 17040 3032 17092 3052
rect 17092 3032 17094 3052
rect 15158 2746 15214 2748
rect 15238 2746 15294 2748
rect 15318 2746 15374 2748
rect 15398 2746 15454 2748
rect 15158 2694 15204 2746
rect 15204 2694 15214 2746
rect 15238 2694 15268 2746
rect 15268 2694 15280 2746
rect 15280 2694 15294 2746
rect 15318 2694 15332 2746
rect 15332 2694 15344 2746
rect 15344 2694 15374 2746
rect 15398 2694 15408 2746
rect 15408 2694 15454 2746
rect 15158 2692 15214 2694
rect 15238 2692 15294 2694
rect 15318 2692 15374 2694
rect 15398 2692 15454 2694
rect 12317 2202 12373 2204
rect 12397 2202 12453 2204
rect 12477 2202 12533 2204
rect 12557 2202 12613 2204
rect 12317 2150 12363 2202
rect 12363 2150 12373 2202
rect 12397 2150 12427 2202
rect 12427 2150 12439 2202
rect 12439 2150 12453 2202
rect 12477 2150 12491 2202
rect 12491 2150 12503 2202
rect 12503 2150 12533 2202
rect 12557 2150 12567 2202
rect 12567 2150 12613 2202
rect 12317 2148 12373 2150
rect 12397 2148 12453 2150
rect 12477 2148 12533 2150
rect 12557 2148 12613 2150
rect 17998 2202 18054 2204
rect 18078 2202 18134 2204
rect 18158 2202 18214 2204
rect 18238 2202 18294 2204
rect 17998 2150 18044 2202
rect 18044 2150 18054 2202
rect 18078 2150 18108 2202
rect 18108 2150 18120 2202
rect 18120 2150 18134 2202
rect 18158 2150 18172 2202
rect 18172 2150 18184 2202
rect 18184 2150 18214 2202
rect 18238 2150 18248 2202
rect 18248 2150 18294 2202
rect 17998 2148 18054 2150
rect 18078 2148 18134 2150
rect 18158 2148 18214 2150
rect 18238 2148 18294 2150
rect 20839 10362 20895 10364
rect 20919 10362 20975 10364
rect 20999 10362 21055 10364
rect 21079 10362 21135 10364
rect 20839 10310 20885 10362
rect 20885 10310 20895 10362
rect 20919 10310 20949 10362
rect 20949 10310 20961 10362
rect 20961 10310 20975 10362
rect 20999 10310 21013 10362
rect 21013 10310 21025 10362
rect 21025 10310 21055 10362
rect 21079 10310 21089 10362
rect 21089 10310 21135 10362
rect 20839 10308 20895 10310
rect 20919 10308 20975 10310
rect 20999 10308 21055 10310
rect 21079 10308 21135 10310
rect 20839 9274 20895 9276
rect 20919 9274 20975 9276
rect 20999 9274 21055 9276
rect 21079 9274 21135 9276
rect 20839 9222 20885 9274
rect 20885 9222 20895 9274
rect 20919 9222 20949 9274
rect 20949 9222 20961 9274
rect 20961 9222 20975 9274
rect 20999 9222 21013 9274
rect 21013 9222 21025 9274
rect 21025 9222 21055 9274
rect 21079 9222 21089 9274
rect 21089 9222 21135 9274
rect 20839 9220 20895 9222
rect 20919 9220 20975 9222
rect 20999 9220 21055 9222
rect 21079 9220 21135 9222
rect 20839 8186 20895 8188
rect 20919 8186 20975 8188
rect 20999 8186 21055 8188
rect 21079 8186 21135 8188
rect 20839 8134 20885 8186
rect 20885 8134 20895 8186
rect 20919 8134 20949 8186
rect 20949 8134 20961 8186
rect 20961 8134 20975 8186
rect 20999 8134 21013 8186
rect 21013 8134 21025 8186
rect 21025 8134 21055 8186
rect 21079 8134 21089 8186
rect 21089 8134 21135 8186
rect 20839 8132 20895 8134
rect 20919 8132 20975 8134
rect 20999 8132 21055 8134
rect 21079 8132 21135 8134
rect 20839 7098 20895 7100
rect 20919 7098 20975 7100
rect 20999 7098 21055 7100
rect 21079 7098 21135 7100
rect 20839 7046 20885 7098
rect 20885 7046 20895 7098
rect 20919 7046 20949 7098
rect 20949 7046 20961 7098
rect 20961 7046 20975 7098
rect 20999 7046 21013 7098
rect 21013 7046 21025 7098
rect 21025 7046 21055 7098
rect 21079 7046 21089 7098
rect 21089 7046 21135 7098
rect 20839 7044 20895 7046
rect 20919 7044 20975 7046
rect 20999 7044 21055 7046
rect 21079 7044 21135 7046
rect 20839 6010 20895 6012
rect 20919 6010 20975 6012
rect 20999 6010 21055 6012
rect 21079 6010 21135 6012
rect 20839 5958 20885 6010
rect 20885 5958 20895 6010
rect 20919 5958 20949 6010
rect 20949 5958 20961 6010
rect 20961 5958 20975 6010
rect 20999 5958 21013 6010
rect 21013 5958 21025 6010
rect 21025 5958 21055 6010
rect 21079 5958 21089 6010
rect 21089 5958 21135 6010
rect 20839 5956 20895 5958
rect 20919 5956 20975 5958
rect 20999 5956 21055 5958
rect 21079 5956 21135 5958
rect 21546 6860 21602 6896
rect 21546 6840 21548 6860
rect 21548 6840 21600 6860
rect 21600 6840 21602 6860
rect 23679 19610 23735 19612
rect 23759 19610 23815 19612
rect 23839 19610 23895 19612
rect 23919 19610 23975 19612
rect 23679 19558 23725 19610
rect 23725 19558 23735 19610
rect 23759 19558 23789 19610
rect 23789 19558 23801 19610
rect 23801 19558 23815 19610
rect 23839 19558 23853 19610
rect 23853 19558 23865 19610
rect 23865 19558 23895 19610
rect 23919 19558 23929 19610
rect 23929 19558 23975 19610
rect 23679 19556 23735 19558
rect 23759 19556 23815 19558
rect 23839 19556 23895 19558
rect 23919 19556 23975 19558
rect 23679 18522 23735 18524
rect 23759 18522 23815 18524
rect 23839 18522 23895 18524
rect 23919 18522 23975 18524
rect 23679 18470 23725 18522
rect 23725 18470 23735 18522
rect 23759 18470 23789 18522
rect 23789 18470 23801 18522
rect 23801 18470 23815 18522
rect 23839 18470 23853 18522
rect 23853 18470 23865 18522
rect 23865 18470 23895 18522
rect 23919 18470 23929 18522
rect 23929 18470 23975 18522
rect 23679 18468 23735 18470
rect 23759 18468 23815 18470
rect 23839 18468 23895 18470
rect 23919 18468 23975 18470
rect 22098 15952 22154 16008
rect 23679 17434 23735 17436
rect 23759 17434 23815 17436
rect 23839 17434 23895 17436
rect 23919 17434 23975 17436
rect 23679 17382 23725 17434
rect 23725 17382 23735 17434
rect 23759 17382 23789 17434
rect 23789 17382 23801 17434
rect 23801 17382 23815 17434
rect 23839 17382 23853 17434
rect 23853 17382 23865 17434
rect 23865 17382 23895 17434
rect 23919 17382 23929 17434
rect 23929 17382 23975 17434
rect 23679 17380 23735 17382
rect 23759 17380 23815 17382
rect 23839 17380 23895 17382
rect 23919 17380 23975 17382
rect 22282 13368 22338 13424
rect 22558 13776 22614 13832
rect 22742 13232 22798 13288
rect 22650 10668 22706 10704
rect 22650 10648 22652 10668
rect 22652 10648 22704 10668
rect 22704 10648 22706 10668
rect 22282 8356 22338 8392
rect 22282 8336 22284 8356
rect 22284 8336 22336 8356
rect 22336 8336 22338 8356
rect 20839 4922 20895 4924
rect 20919 4922 20975 4924
rect 20999 4922 21055 4924
rect 21079 4922 21135 4924
rect 20839 4870 20885 4922
rect 20885 4870 20895 4922
rect 20919 4870 20949 4922
rect 20949 4870 20961 4922
rect 20961 4870 20975 4922
rect 20999 4870 21013 4922
rect 21013 4870 21025 4922
rect 21025 4870 21055 4922
rect 21079 4870 21089 4922
rect 21089 4870 21135 4922
rect 20839 4868 20895 4870
rect 20919 4868 20975 4870
rect 20999 4868 21055 4870
rect 21079 4868 21135 4870
rect 20839 3834 20895 3836
rect 20919 3834 20975 3836
rect 20999 3834 21055 3836
rect 21079 3834 21135 3836
rect 20839 3782 20885 3834
rect 20885 3782 20895 3834
rect 20919 3782 20949 3834
rect 20949 3782 20961 3834
rect 20961 3782 20975 3834
rect 20999 3782 21013 3834
rect 21013 3782 21025 3834
rect 21025 3782 21055 3834
rect 21079 3782 21089 3834
rect 21089 3782 21135 3834
rect 20839 3780 20895 3782
rect 20919 3780 20975 3782
rect 20999 3780 21055 3782
rect 21079 3780 21135 3782
rect 22098 4684 22154 4720
rect 22098 4664 22100 4684
rect 22100 4664 22152 4684
rect 22152 4664 22154 4684
rect 23679 16346 23735 16348
rect 23759 16346 23815 16348
rect 23839 16346 23895 16348
rect 23919 16346 23975 16348
rect 23679 16294 23725 16346
rect 23725 16294 23735 16346
rect 23759 16294 23789 16346
rect 23789 16294 23801 16346
rect 23801 16294 23815 16346
rect 23839 16294 23853 16346
rect 23853 16294 23865 16346
rect 23865 16294 23895 16346
rect 23919 16294 23929 16346
rect 23929 16294 23975 16346
rect 23679 16292 23735 16294
rect 23759 16292 23815 16294
rect 23839 16292 23895 16294
rect 23919 16292 23975 16294
rect 23679 15258 23735 15260
rect 23759 15258 23815 15260
rect 23839 15258 23895 15260
rect 23919 15258 23975 15260
rect 23679 15206 23725 15258
rect 23725 15206 23735 15258
rect 23759 15206 23789 15258
rect 23789 15206 23801 15258
rect 23801 15206 23815 15258
rect 23839 15206 23853 15258
rect 23853 15206 23865 15258
rect 23865 15206 23895 15258
rect 23919 15206 23929 15258
rect 23929 15206 23975 15258
rect 23679 15204 23735 15206
rect 23759 15204 23815 15206
rect 23839 15204 23895 15206
rect 23919 15204 23975 15206
rect 23679 14170 23735 14172
rect 23759 14170 23815 14172
rect 23839 14170 23895 14172
rect 23919 14170 23975 14172
rect 23679 14118 23725 14170
rect 23725 14118 23735 14170
rect 23759 14118 23789 14170
rect 23789 14118 23801 14170
rect 23801 14118 23815 14170
rect 23839 14118 23853 14170
rect 23853 14118 23865 14170
rect 23865 14118 23895 14170
rect 23919 14118 23929 14170
rect 23929 14118 23975 14170
rect 23679 14116 23735 14118
rect 23759 14116 23815 14118
rect 23839 14116 23895 14118
rect 23919 14116 23975 14118
rect 23679 13082 23735 13084
rect 23759 13082 23815 13084
rect 23839 13082 23895 13084
rect 23919 13082 23975 13084
rect 23679 13030 23725 13082
rect 23725 13030 23735 13082
rect 23759 13030 23789 13082
rect 23789 13030 23801 13082
rect 23801 13030 23815 13082
rect 23839 13030 23853 13082
rect 23853 13030 23865 13082
rect 23865 13030 23895 13082
rect 23919 13030 23929 13082
rect 23929 13030 23975 13082
rect 23679 13028 23735 13030
rect 23759 13028 23815 13030
rect 23839 13028 23895 13030
rect 23919 13028 23975 13030
rect 23679 11994 23735 11996
rect 23759 11994 23815 11996
rect 23839 11994 23895 11996
rect 23919 11994 23975 11996
rect 23679 11942 23725 11994
rect 23725 11942 23735 11994
rect 23759 11942 23789 11994
rect 23789 11942 23801 11994
rect 23801 11942 23815 11994
rect 23839 11942 23853 11994
rect 23853 11942 23865 11994
rect 23865 11942 23895 11994
rect 23919 11942 23929 11994
rect 23929 11942 23975 11994
rect 23679 11940 23735 11942
rect 23759 11940 23815 11942
rect 23839 11940 23895 11942
rect 23919 11940 23975 11942
rect 23679 10906 23735 10908
rect 23759 10906 23815 10908
rect 23839 10906 23895 10908
rect 23919 10906 23975 10908
rect 23679 10854 23725 10906
rect 23725 10854 23735 10906
rect 23759 10854 23789 10906
rect 23789 10854 23801 10906
rect 23801 10854 23815 10906
rect 23839 10854 23853 10906
rect 23853 10854 23865 10906
rect 23865 10854 23895 10906
rect 23919 10854 23929 10906
rect 23929 10854 23975 10906
rect 23679 10852 23735 10854
rect 23759 10852 23815 10854
rect 23839 10852 23895 10854
rect 23919 10852 23975 10854
rect 23679 9818 23735 9820
rect 23759 9818 23815 9820
rect 23839 9818 23895 9820
rect 23919 9818 23975 9820
rect 23679 9766 23725 9818
rect 23725 9766 23735 9818
rect 23759 9766 23789 9818
rect 23789 9766 23801 9818
rect 23801 9766 23815 9818
rect 23839 9766 23853 9818
rect 23853 9766 23865 9818
rect 23865 9766 23895 9818
rect 23919 9766 23929 9818
rect 23929 9766 23975 9818
rect 23679 9764 23735 9766
rect 23759 9764 23815 9766
rect 23839 9764 23895 9766
rect 23919 9764 23975 9766
rect 23679 8730 23735 8732
rect 23759 8730 23815 8732
rect 23839 8730 23895 8732
rect 23919 8730 23975 8732
rect 23679 8678 23725 8730
rect 23725 8678 23735 8730
rect 23759 8678 23789 8730
rect 23789 8678 23801 8730
rect 23801 8678 23815 8730
rect 23839 8678 23853 8730
rect 23853 8678 23865 8730
rect 23865 8678 23895 8730
rect 23919 8678 23929 8730
rect 23929 8678 23975 8730
rect 23679 8676 23735 8678
rect 23759 8676 23815 8678
rect 23839 8676 23895 8678
rect 23919 8676 23975 8678
rect 23679 7642 23735 7644
rect 23759 7642 23815 7644
rect 23839 7642 23895 7644
rect 23919 7642 23975 7644
rect 23679 7590 23725 7642
rect 23725 7590 23735 7642
rect 23759 7590 23789 7642
rect 23789 7590 23801 7642
rect 23801 7590 23815 7642
rect 23839 7590 23853 7642
rect 23853 7590 23865 7642
rect 23865 7590 23895 7642
rect 23919 7590 23929 7642
rect 23929 7590 23975 7642
rect 23679 7588 23735 7590
rect 23759 7588 23815 7590
rect 23839 7588 23895 7590
rect 23919 7588 23975 7590
rect 23679 6554 23735 6556
rect 23759 6554 23815 6556
rect 23839 6554 23895 6556
rect 23919 6554 23975 6556
rect 23679 6502 23725 6554
rect 23725 6502 23735 6554
rect 23759 6502 23789 6554
rect 23789 6502 23801 6554
rect 23801 6502 23815 6554
rect 23839 6502 23853 6554
rect 23853 6502 23865 6554
rect 23865 6502 23895 6554
rect 23919 6502 23929 6554
rect 23929 6502 23975 6554
rect 23679 6500 23735 6502
rect 23759 6500 23815 6502
rect 23839 6500 23895 6502
rect 23919 6500 23975 6502
rect 23679 5466 23735 5468
rect 23759 5466 23815 5468
rect 23839 5466 23895 5468
rect 23919 5466 23975 5468
rect 23679 5414 23725 5466
rect 23725 5414 23735 5466
rect 23759 5414 23789 5466
rect 23789 5414 23801 5466
rect 23801 5414 23815 5466
rect 23839 5414 23853 5466
rect 23853 5414 23865 5466
rect 23865 5414 23895 5466
rect 23919 5414 23929 5466
rect 23929 5414 23975 5466
rect 23679 5412 23735 5414
rect 23759 5412 23815 5414
rect 23839 5412 23895 5414
rect 23919 5412 23975 5414
rect 23679 4378 23735 4380
rect 23759 4378 23815 4380
rect 23839 4378 23895 4380
rect 23919 4378 23975 4380
rect 23679 4326 23725 4378
rect 23725 4326 23735 4378
rect 23759 4326 23789 4378
rect 23789 4326 23801 4378
rect 23801 4326 23815 4378
rect 23839 4326 23853 4378
rect 23853 4326 23865 4378
rect 23865 4326 23895 4378
rect 23919 4326 23929 4378
rect 23929 4326 23975 4378
rect 23679 4324 23735 4326
rect 23759 4324 23815 4326
rect 23839 4324 23895 4326
rect 23919 4324 23975 4326
rect 20350 3476 20352 3496
rect 20352 3476 20404 3496
rect 20404 3476 20406 3496
rect 20350 3440 20406 3476
rect 18694 2896 18750 2952
rect 20839 2746 20895 2748
rect 20919 2746 20975 2748
rect 20999 2746 21055 2748
rect 21079 2746 21135 2748
rect 20839 2694 20885 2746
rect 20885 2694 20895 2746
rect 20919 2694 20949 2746
rect 20949 2694 20961 2746
rect 20961 2694 20975 2746
rect 20999 2694 21013 2746
rect 21013 2694 21025 2746
rect 21025 2694 21055 2746
rect 21079 2694 21089 2746
rect 21089 2694 21135 2746
rect 20839 2692 20895 2694
rect 20919 2692 20975 2694
rect 20999 2692 21055 2694
rect 21079 2692 21135 2694
rect 23679 3290 23735 3292
rect 23759 3290 23815 3292
rect 23839 3290 23895 3292
rect 23919 3290 23975 3292
rect 23679 3238 23725 3290
rect 23725 3238 23735 3290
rect 23759 3238 23789 3290
rect 23789 3238 23801 3290
rect 23801 3238 23815 3290
rect 23839 3238 23853 3290
rect 23853 3238 23865 3290
rect 23865 3238 23895 3290
rect 23919 3238 23929 3290
rect 23929 3238 23975 3290
rect 23679 3236 23735 3238
rect 23759 3236 23815 3238
rect 23839 3236 23895 3238
rect 23919 3236 23975 3238
rect 23679 2202 23735 2204
rect 23759 2202 23815 2204
rect 23839 2202 23895 2204
rect 23919 2202 23975 2204
rect 23679 2150 23725 2202
rect 23725 2150 23735 2202
rect 23759 2150 23789 2202
rect 23789 2150 23801 2202
rect 23801 2150 23815 2202
rect 23839 2150 23853 2202
rect 23853 2150 23865 2202
rect 23865 2150 23895 2202
rect 23919 2150 23929 2202
rect 23929 2150 23975 2202
rect 23679 2148 23735 2150
rect 23759 2148 23815 2150
rect 23839 2148 23895 2150
rect 23919 2148 23975 2150
<< metal3 >>
rect 3786 22336 4102 22337
rect 3786 22272 3792 22336
rect 3856 22272 3872 22336
rect 3936 22272 3952 22336
rect 4016 22272 4032 22336
rect 4096 22272 4102 22336
rect 3786 22271 4102 22272
rect 9467 22336 9783 22337
rect 9467 22272 9473 22336
rect 9537 22272 9553 22336
rect 9617 22272 9633 22336
rect 9697 22272 9713 22336
rect 9777 22272 9783 22336
rect 9467 22271 9783 22272
rect 15148 22336 15464 22337
rect 15148 22272 15154 22336
rect 15218 22272 15234 22336
rect 15298 22272 15314 22336
rect 15378 22272 15394 22336
rect 15458 22272 15464 22336
rect 15148 22271 15464 22272
rect 20829 22336 21145 22337
rect 20829 22272 20835 22336
rect 20899 22272 20915 22336
rect 20979 22272 20995 22336
rect 21059 22272 21075 22336
rect 21139 22272 21145 22336
rect 20829 22271 21145 22272
rect 6626 21792 6942 21793
rect 6626 21728 6632 21792
rect 6696 21728 6712 21792
rect 6776 21728 6792 21792
rect 6856 21728 6872 21792
rect 6936 21728 6942 21792
rect 6626 21727 6942 21728
rect 12307 21792 12623 21793
rect 12307 21728 12313 21792
rect 12377 21728 12393 21792
rect 12457 21728 12473 21792
rect 12537 21728 12553 21792
rect 12617 21728 12623 21792
rect 12307 21727 12623 21728
rect 17988 21792 18304 21793
rect 17988 21728 17994 21792
rect 18058 21728 18074 21792
rect 18138 21728 18154 21792
rect 18218 21728 18234 21792
rect 18298 21728 18304 21792
rect 17988 21727 18304 21728
rect 23669 21792 23985 21793
rect 23669 21728 23675 21792
rect 23739 21728 23755 21792
rect 23819 21728 23835 21792
rect 23899 21728 23915 21792
rect 23979 21728 23985 21792
rect 23669 21727 23985 21728
rect 5441 21586 5507 21589
rect 16205 21586 16271 21589
rect 5441 21584 16271 21586
rect 5441 21528 5446 21584
rect 5502 21528 16210 21584
rect 16266 21528 16271 21584
rect 5441 21526 16271 21528
rect 5441 21523 5507 21526
rect 16205 21523 16271 21526
rect 3786 21248 4102 21249
rect 3786 21184 3792 21248
rect 3856 21184 3872 21248
rect 3936 21184 3952 21248
rect 4016 21184 4032 21248
rect 4096 21184 4102 21248
rect 3786 21183 4102 21184
rect 9467 21248 9783 21249
rect 9467 21184 9473 21248
rect 9537 21184 9553 21248
rect 9617 21184 9633 21248
rect 9697 21184 9713 21248
rect 9777 21184 9783 21248
rect 9467 21183 9783 21184
rect 15148 21248 15464 21249
rect 15148 21184 15154 21248
rect 15218 21184 15234 21248
rect 15298 21184 15314 21248
rect 15378 21184 15394 21248
rect 15458 21184 15464 21248
rect 15148 21183 15464 21184
rect 20829 21248 21145 21249
rect 20829 21184 20835 21248
rect 20899 21184 20915 21248
rect 20979 21184 20995 21248
rect 21059 21184 21075 21248
rect 21139 21184 21145 21248
rect 20829 21183 21145 21184
rect 13077 20772 13143 20773
rect 13077 20768 13124 20772
rect 13188 20770 13194 20772
rect 14457 20770 14523 20773
rect 14774 20770 14780 20772
rect 13077 20712 13082 20768
rect 13077 20708 13124 20712
rect 13188 20710 13234 20770
rect 14457 20768 14780 20770
rect 14457 20712 14462 20768
rect 14518 20712 14780 20768
rect 14457 20710 14780 20712
rect 13188 20708 13194 20710
rect 13077 20707 13143 20708
rect 14457 20707 14523 20710
rect 14774 20708 14780 20710
rect 14844 20708 14850 20772
rect 6626 20704 6942 20705
rect 6626 20640 6632 20704
rect 6696 20640 6712 20704
rect 6776 20640 6792 20704
rect 6856 20640 6872 20704
rect 6936 20640 6942 20704
rect 6626 20639 6942 20640
rect 12307 20704 12623 20705
rect 12307 20640 12313 20704
rect 12377 20640 12393 20704
rect 12457 20640 12473 20704
rect 12537 20640 12553 20704
rect 12617 20640 12623 20704
rect 12307 20639 12623 20640
rect 17988 20704 18304 20705
rect 17988 20640 17994 20704
rect 18058 20640 18074 20704
rect 18138 20640 18154 20704
rect 18218 20640 18234 20704
rect 18298 20640 18304 20704
rect 17988 20639 18304 20640
rect 23669 20704 23985 20705
rect 23669 20640 23675 20704
rect 23739 20640 23755 20704
rect 23819 20640 23835 20704
rect 23899 20640 23915 20704
rect 23979 20640 23985 20704
rect 23669 20639 23985 20640
rect 13353 20634 13419 20637
rect 17861 20634 17927 20637
rect 13353 20632 17927 20634
rect 13353 20576 13358 20632
rect 13414 20576 17866 20632
rect 17922 20576 17927 20632
rect 13353 20574 17927 20576
rect 13353 20571 13419 20574
rect 17861 20571 17927 20574
rect 13629 20362 13695 20365
rect 16665 20362 16731 20365
rect 13629 20360 16731 20362
rect 13629 20304 13634 20360
rect 13690 20304 16670 20360
rect 16726 20304 16731 20360
rect 13629 20302 16731 20304
rect 13629 20299 13695 20302
rect 16665 20299 16731 20302
rect 3786 20160 4102 20161
rect 3786 20096 3792 20160
rect 3856 20096 3872 20160
rect 3936 20096 3952 20160
rect 4016 20096 4032 20160
rect 4096 20096 4102 20160
rect 3786 20095 4102 20096
rect 9467 20160 9783 20161
rect 9467 20096 9473 20160
rect 9537 20096 9553 20160
rect 9617 20096 9633 20160
rect 9697 20096 9713 20160
rect 9777 20096 9783 20160
rect 9467 20095 9783 20096
rect 15148 20160 15464 20161
rect 15148 20096 15154 20160
rect 15218 20096 15234 20160
rect 15298 20096 15314 20160
rect 15378 20096 15394 20160
rect 15458 20096 15464 20160
rect 15148 20095 15464 20096
rect 20829 20160 21145 20161
rect 20829 20096 20835 20160
rect 20899 20096 20915 20160
rect 20979 20096 20995 20160
rect 21059 20096 21075 20160
rect 21139 20096 21145 20160
rect 20829 20095 21145 20096
rect 13261 19954 13327 19957
rect 15285 19954 15351 19957
rect 13261 19952 15351 19954
rect 13261 19896 13266 19952
rect 13322 19896 15290 19952
rect 15346 19896 15351 19952
rect 13261 19894 15351 19896
rect 13261 19891 13327 19894
rect 15285 19891 15351 19894
rect 15377 19818 15443 19821
rect 16849 19818 16915 19821
rect 15377 19816 16915 19818
rect 15377 19760 15382 19816
rect 15438 19760 16854 19816
rect 16910 19760 16915 19816
rect 15377 19758 16915 19760
rect 15377 19755 15443 19758
rect 16849 19755 16915 19758
rect 6626 19616 6942 19617
rect 6626 19552 6632 19616
rect 6696 19552 6712 19616
rect 6776 19552 6792 19616
rect 6856 19552 6872 19616
rect 6936 19552 6942 19616
rect 6626 19551 6942 19552
rect 12307 19616 12623 19617
rect 12307 19552 12313 19616
rect 12377 19552 12393 19616
rect 12457 19552 12473 19616
rect 12537 19552 12553 19616
rect 12617 19552 12623 19616
rect 12307 19551 12623 19552
rect 17988 19616 18304 19617
rect 17988 19552 17994 19616
rect 18058 19552 18074 19616
rect 18138 19552 18154 19616
rect 18218 19552 18234 19616
rect 18298 19552 18304 19616
rect 17988 19551 18304 19552
rect 23669 19616 23985 19617
rect 23669 19552 23675 19616
rect 23739 19552 23755 19616
rect 23819 19552 23835 19616
rect 23899 19552 23915 19616
rect 23979 19552 23985 19616
rect 23669 19551 23985 19552
rect 15745 19546 15811 19549
rect 17125 19546 17191 19549
rect 15745 19544 17191 19546
rect 15745 19488 15750 19544
rect 15806 19488 17130 19544
rect 17186 19488 17191 19544
rect 15745 19486 17191 19488
rect 15745 19483 15811 19486
rect 17125 19483 17191 19486
rect 15193 19410 15259 19413
rect 16757 19410 16823 19413
rect 15193 19408 16823 19410
rect 15193 19352 15198 19408
rect 15254 19352 16762 19408
rect 16818 19352 16823 19408
rect 15193 19350 16823 19352
rect 15193 19347 15259 19350
rect 16757 19347 16823 19350
rect 17309 19410 17375 19413
rect 17718 19410 17724 19412
rect 17309 19408 17724 19410
rect 17309 19352 17314 19408
rect 17370 19352 17724 19408
rect 17309 19350 17724 19352
rect 17309 19347 17375 19350
rect 17718 19348 17724 19350
rect 17788 19348 17794 19412
rect 3786 19072 4102 19073
rect 3786 19008 3792 19072
rect 3856 19008 3872 19072
rect 3936 19008 3952 19072
rect 4016 19008 4032 19072
rect 4096 19008 4102 19072
rect 3786 19007 4102 19008
rect 9467 19072 9783 19073
rect 9467 19008 9473 19072
rect 9537 19008 9553 19072
rect 9617 19008 9633 19072
rect 9697 19008 9713 19072
rect 9777 19008 9783 19072
rect 9467 19007 9783 19008
rect 15148 19072 15464 19073
rect 15148 19008 15154 19072
rect 15218 19008 15234 19072
rect 15298 19008 15314 19072
rect 15378 19008 15394 19072
rect 15458 19008 15464 19072
rect 15148 19007 15464 19008
rect 20829 19072 21145 19073
rect 20829 19008 20835 19072
rect 20899 19008 20915 19072
rect 20979 19008 20995 19072
rect 21059 19008 21075 19072
rect 21139 19008 21145 19072
rect 20829 19007 21145 19008
rect 6626 18528 6942 18529
rect 6626 18464 6632 18528
rect 6696 18464 6712 18528
rect 6776 18464 6792 18528
rect 6856 18464 6872 18528
rect 6936 18464 6942 18528
rect 6626 18463 6942 18464
rect 12307 18528 12623 18529
rect 12307 18464 12313 18528
rect 12377 18464 12393 18528
rect 12457 18464 12473 18528
rect 12537 18464 12553 18528
rect 12617 18464 12623 18528
rect 12307 18463 12623 18464
rect 17988 18528 18304 18529
rect 17988 18464 17994 18528
rect 18058 18464 18074 18528
rect 18138 18464 18154 18528
rect 18218 18464 18234 18528
rect 18298 18464 18304 18528
rect 17988 18463 18304 18464
rect 23669 18528 23985 18529
rect 23669 18464 23675 18528
rect 23739 18464 23755 18528
rect 23819 18464 23835 18528
rect 23899 18464 23915 18528
rect 23979 18464 23985 18528
rect 23669 18463 23985 18464
rect 20897 18186 20963 18189
rect 21398 18186 21404 18188
rect 20897 18184 21404 18186
rect 20897 18128 20902 18184
rect 20958 18128 21404 18184
rect 20897 18126 21404 18128
rect 20897 18123 20963 18126
rect 21398 18124 21404 18126
rect 21468 18124 21474 18188
rect 15745 18050 15811 18053
rect 16430 18050 16436 18052
rect 15745 18048 16436 18050
rect 15745 17992 15750 18048
rect 15806 17992 16436 18048
rect 15745 17990 16436 17992
rect 15745 17987 15811 17990
rect 16430 17988 16436 17990
rect 16500 17988 16506 18052
rect 3786 17984 4102 17985
rect 3786 17920 3792 17984
rect 3856 17920 3872 17984
rect 3936 17920 3952 17984
rect 4016 17920 4032 17984
rect 4096 17920 4102 17984
rect 3786 17919 4102 17920
rect 9467 17984 9783 17985
rect 9467 17920 9473 17984
rect 9537 17920 9553 17984
rect 9617 17920 9633 17984
rect 9697 17920 9713 17984
rect 9777 17920 9783 17984
rect 9467 17919 9783 17920
rect 15148 17984 15464 17985
rect 15148 17920 15154 17984
rect 15218 17920 15234 17984
rect 15298 17920 15314 17984
rect 15378 17920 15394 17984
rect 15458 17920 15464 17984
rect 15148 17919 15464 17920
rect 20829 17984 21145 17985
rect 20829 17920 20835 17984
rect 20899 17920 20915 17984
rect 20979 17920 20995 17984
rect 21059 17920 21075 17984
rect 21139 17920 21145 17984
rect 20829 17919 21145 17920
rect 6626 17440 6942 17441
rect 6626 17376 6632 17440
rect 6696 17376 6712 17440
rect 6776 17376 6792 17440
rect 6856 17376 6872 17440
rect 6936 17376 6942 17440
rect 6626 17375 6942 17376
rect 12307 17440 12623 17441
rect 12307 17376 12313 17440
rect 12377 17376 12393 17440
rect 12457 17376 12473 17440
rect 12537 17376 12553 17440
rect 12617 17376 12623 17440
rect 12307 17375 12623 17376
rect 17988 17440 18304 17441
rect 17988 17376 17994 17440
rect 18058 17376 18074 17440
rect 18138 17376 18154 17440
rect 18218 17376 18234 17440
rect 18298 17376 18304 17440
rect 17988 17375 18304 17376
rect 23669 17440 23985 17441
rect 23669 17376 23675 17440
rect 23739 17376 23755 17440
rect 23819 17376 23835 17440
rect 23899 17376 23915 17440
rect 23979 17376 23985 17440
rect 23669 17375 23985 17376
rect 3786 16896 4102 16897
rect 3786 16832 3792 16896
rect 3856 16832 3872 16896
rect 3936 16832 3952 16896
rect 4016 16832 4032 16896
rect 4096 16832 4102 16896
rect 3786 16831 4102 16832
rect 9467 16896 9783 16897
rect 9467 16832 9473 16896
rect 9537 16832 9553 16896
rect 9617 16832 9633 16896
rect 9697 16832 9713 16896
rect 9777 16832 9783 16896
rect 9467 16831 9783 16832
rect 15148 16896 15464 16897
rect 15148 16832 15154 16896
rect 15218 16832 15234 16896
rect 15298 16832 15314 16896
rect 15378 16832 15394 16896
rect 15458 16832 15464 16896
rect 15148 16831 15464 16832
rect 20829 16896 21145 16897
rect 20829 16832 20835 16896
rect 20899 16832 20915 16896
rect 20979 16832 20995 16896
rect 21059 16832 21075 16896
rect 21139 16832 21145 16896
rect 20829 16831 21145 16832
rect 16021 16826 16087 16829
rect 18965 16826 19031 16829
rect 16021 16824 19031 16826
rect 16021 16768 16026 16824
rect 16082 16768 18970 16824
rect 19026 16768 19031 16824
rect 16021 16766 19031 16768
rect 16021 16763 16087 16766
rect 18965 16763 19031 16766
rect 17769 16554 17835 16557
rect 18045 16554 18111 16557
rect 17769 16552 18111 16554
rect 17769 16496 17774 16552
rect 17830 16496 18050 16552
rect 18106 16496 18111 16552
rect 17769 16494 18111 16496
rect 17769 16491 17835 16494
rect 18045 16491 18111 16494
rect 6626 16352 6942 16353
rect 6626 16288 6632 16352
rect 6696 16288 6712 16352
rect 6776 16288 6792 16352
rect 6856 16288 6872 16352
rect 6936 16288 6942 16352
rect 6626 16287 6942 16288
rect 12307 16352 12623 16353
rect 12307 16288 12313 16352
rect 12377 16288 12393 16352
rect 12457 16288 12473 16352
rect 12537 16288 12553 16352
rect 12617 16288 12623 16352
rect 12307 16287 12623 16288
rect 17988 16352 18304 16353
rect 17988 16288 17994 16352
rect 18058 16288 18074 16352
rect 18138 16288 18154 16352
rect 18218 16288 18234 16352
rect 18298 16288 18304 16352
rect 17988 16287 18304 16288
rect 23669 16352 23985 16353
rect 23669 16288 23675 16352
rect 23739 16288 23755 16352
rect 23819 16288 23835 16352
rect 23899 16288 23915 16352
rect 23979 16288 23985 16352
rect 23669 16287 23985 16288
rect 18413 16146 18479 16149
rect 20805 16146 20871 16149
rect 22001 16146 22067 16149
rect 18413 16144 22067 16146
rect 18413 16088 18418 16144
rect 18474 16088 20810 16144
rect 20866 16088 22006 16144
rect 22062 16088 22067 16144
rect 18413 16086 22067 16088
rect 18413 16083 18479 16086
rect 20805 16083 20871 16086
rect 22001 16083 22067 16086
rect 18505 16010 18571 16013
rect 22093 16010 22159 16013
rect 18505 16008 22159 16010
rect 18505 15952 18510 16008
rect 18566 15952 22098 16008
rect 22154 15952 22159 16008
rect 18505 15950 22159 15952
rect 18505 15947 18571 15950
rect 22093 15947 22159 15950
rect 3786 15808 4102 15809
rect 3786 15744 3792 15808
rect 3856 15744 3872 15808
rect 3936 15744 3952 15808
rect 4016 15744 4032 15808
rect 4096 15744 4102 15808
rect 3786 15743 4102 15744
rect 9467 15808 9783 15809
rect 9467 15744 9473 15808
rect 9537 15744 9553 15808
rect 9617 15744 9633 15808
rect 9697 15744 9713 15808
rect 9777 15744 9783 15808
rect 9467 15743 9783 15744
rect 15148 15808 15464 15809
rect 15148 15744 15154 15808
rect 15218 15744 15234 15808
rect 15298 15744 15314 15808
rect 15378 15744 15394 15808
rect 15458 15744 15464 15808
rect 15148 15743 15464 15744
rect 20829 15808 21145 15809
rect 20829 15744 20835 15808
rect 20899 15744 20915 15808
rect 20979 15744 20995 15808
rect 21059 15744 21075 15808
rect 21139 15744 21145 15808
rect 20829 15743 21145 15744
rect 5257 15330 5323 15333
rect 5390 15330 5396 15332
rect 5257 15328 5396 15330
rect 5257 15272 5262 15328
rect 5318 15272 5396 15328
rect 5257 15270 5396 15272
rect 5257 15267 5323 15270
rect 5390 15268 5396 15270
rect 5460 15268 5466 15332
rect 6626 15264 6942 15265
rect 6626 15200 6632 15264
rect 6696 15200 6712 15264
rect 6776 15200 6792 15264
rect 6856 15200 6872 15264
rect 6936 15200 6942 15264
rect 6626 15199 6942 15200
rect 12307 15264 12623 15265
rect 12307 15200 12313 15264
rect 12377 15200 12393 15264
rect 12457 15200 12473 15264
rect 12537 15200 12553 15264
rect 12617 15200 12623 15264
rect 12307 15199 12623 15200
rect 17988 15264 18304 15265
rect 17988 15200 17994 15264
rect 18058 15200 18074 15264
rect 18138 15200 18154 15264
rect 18218 15200 18234 15264
rect 18298 15200 18304 15264
rect 17988 15199 18304 15200
rect 23669 15264 23985 15265
rect 23669 15200 23675 15264
rect 23739 15200 23755 15264
rect 23819 15200 23835 15264
rect 23899 15200 23915 15264
rect 23979 15200 23985 15264
rect 23669 15199 23985 15200
rect 2313 15058 2379 15061
rect 4981 15058 5047 15061
rect 7005 15058 7071 15061
rect 2313 15056 7071 15058
rect 2313 15000 2318 15056
rect 2374 15000 4986 15056
rect 5042 15000 7010 15056
rect 7066 15000 7071 15056
rect 2313 14998 7071 15000
rect 2313 14995 2379 14998
rect 4981 14995 5047 14998
rect 7005 14995 7071 14998
rect 3786 14720 4102 14721
rect 3786 14656 3792 14720
rect 3856 14656 3872 14720
rect 3936 14656 3952 14720
rect 4016 14656 4032 14720
rect 4096 14656 4102 14720
rect 3786 14655 4102 14656
rect 9467 14720 9783 14721
rect 9467 14656 9473 14720
rect 9537 14656 9553 14720
rect 9617 14656 9633 14720
rect 9697 14656 9713 14720
rect 9777 14656 9783 14720
rect 9467 14655 9783 14656
rect 15148 14720 15464 14721
rect 15148 14656 15154 14720
rect 15218 14656 15234 14720
rect 15298 14656 15314 14720
rect 15378 14656 15394 14720
rect 15458 14656 15464 14720
rect 15148 14655 15464 14656
rect 20829 14720 21145 14721
rect 20829 14656 20835 14720
rect 20899 14656 20915 14720
rect 20979 14656 20995 14720
rect 21059 14656 21075 14720
rect 21139 14656 21145 14720
rect 20829 14655 21145 14656
rect 16430 14588 16436 14652
rect 16500 14650 16506 14652
rect 19333 14650 19399 14653
rect 16500 14648 19399 14650
rect 16500 14592 19338 14648
rect 19394 14592 19399 14648
rect 16500 14590 19399 14592
rect 16500 14588 16506 14590
rect 19333 14587 19399 14590
rect 6626 14176 6942 14177
rect 6626 14112 6632 14176
rect 6696 14112 6712 14176
rect 6776 14112 6792 14176
rect 6856 14112 6872 14176
rect 6936 14112 6942 14176
rect 6626 14111 6942 14112
rect 12307 14176 12623 14177
rect 12307 14112 12313 14176
rect 12377 14112 12393 14176
rect 12457 14112 12473 14176
rect 12537 14112 12553 14176
rect 12617 14112 12623 14176
rect 12307 14111 12623 14112
rect 17988 14176 18304 14177
rect 17988 14112 17994 14176
rect 18058 14112 18074 14176
rect 18138 14112 18154 14176
rect 18218 14112 18234 14176
rect 18298 14112 18304 14176
rect 17988 14111 18304 14112
rect 23669 14176 23985 14177
rect 23669 14112 23675 14176
rect 23739 14112 23755 14176
rect 23819 14112 23835 14176
rect 23899 14112 23915 14176
rect 23979 14112 23985 14176
rect 23669 14111 23985 14112
rect 13077 14106 13143 14109
rect 15653 14106 15719 14109
rect 13077 14104 15719 14106
rect 13077 14048 13082 14104
rect 13138 14048 15658 14104
rect 15714 14048 15719 14104
rect 13077 14046 15719 14048
rect 13077 14043 13143 14046
rect 15653 14043 15719 14046
rect 17217 13970 17283 13973
rect 17174 13968 17283 13970
rect 17174 13912 17222 13968
rect 17278 13912 17283 13968
rect 17174 13907 17283 13912
rect 18229 13970 18295 13973
rect 19885 13970 19951 13973
rect 20989 13970 21055 13973
rect 18229 13968 21055 13970
rect 18229 13912 18234 13968
rect 18290 13912 19890 13968
rect 19946 13912 20994 13968
rect 21050 13912 21055 13968
rect 18229 13910 21055 13912
rect 18229 13907 18295 13910
rect 19885 13907 19951 13910
rect 20989 13907 21055 13910
rect 15929 13834 15995 13837
rect 16246 13834 16252 13836
rect 15929 13832 16252 13834
rect 15929 13776 15934 13832
rect 15990 13776 16252 13832
rect 15929 13774 16252 13776
rect 15929 13771 15995 13774
rect 16246 13772 16252 13774
rect 16316 13772 16322 13836
rect 3786 13632 4102 13633
rect 3786 13568 3792 13632
rect 3856 13568 3872 13632
rect 3936 13568 3952 13632
rect 4016 13568 4032 13632
rect 4096 13568 4102 13632
rect 3786 13567 4102 13568
rect 9467 13632 9783 13633
rect 9467 13568 9473 13632
rect 9537 13568 9553 13632
rect 9617 13568 9633 13632
rect 9697 13568 9713 13632
rect 9777 13568 9783 13632
rect 9467 13567 9783 13568
rect 15148 13632 15464 13633
rect 15148 13568 15154 13632
rect 15218 13568 15234 13632
rect 15298 13568 15314 13632
rect 15378 13568 15394 13632
rect 15458 13568 15464 13632
rect 15148 13567 15464 13568
rect 17174 13426 17234 13907
rect 22318 13772 22324 13836
rect 22388 13834 22394 13836
rect 22553 13834 22619 13837
rect 22388 13832 22619 13834
rect 22388 13776 22558 13832
rect 22614 13776 22619 13832
rect 22388 13774 22619 13776
rect 22388 13772 22394 13774
rect 22553 13771 22619 13774
rect 20829 13632 21145 13633
rect 20829 13568 20835 13632
rect 20899 13568 20915 13632
rect 20979 13568 20995 13632
rect 21059 13568 21075 13632
rect 21139 13568 21145 13632
rect 20829 13567 21145 13568
rect 17718 13500 17724 13564
rect 17788 13562 17794 13564
rect 19609 13562 19675 13565
rect 17788 13560 19675 13562
rect 17788 13504 19614 13560
rect 19670 13504 19675 13560
rect 17788 13502 19675 13504
rect 17788 13500 17794 13502
rect 19609 13499 19675 13502
rect 17309 13426 17375 13429
rect 17174 13424 17375 13426
rect 17174 13368 17314 13424
rect 17370 13368 17375 13424
rect 17174 13366 17375 13368
rect 17309 13363 17375 13366
rect 18597 13426 18663 13429
rect 22277 13426 22343 13429
rect 18597 13424 22343 13426
rect 18597 13368 18602 13424
rect 18658 13368 22282 13424
rect 22338 13368 22343 13424
rect 18597 13366 22343 13368
rect 18597 13363 18663 13366
rect 22277 13363 22343 13366
rect 17125 13290 17191 13293
rect 22737 13290 22803 13293
rect 17125 13288 22803 13290
rect 17125 13232 17130 13288
rect 17186 13232 22742 13288
rect 22798 13232 22803 13288
rect 17125 13230 22803 13232
rect 17125 13227 17191 13230
rect 22737 13227 22803 13230
rect 16941 13154 17007 13157
rect 17677 13154 17743 13157
rect 16941 13152 17743 13154
rect 16941 13096 16946 13152
rect 17002 13096 17682 13152
rect 17738 13096 17743 13152
rect 16941 13094 17743 13096
rect 16941 13091 17007 13094
rect 17677 13091 17743 13094
rect 19701 13154 19767 13157
rect 20345 13154 20411 13157
rect 19701 13152 20411 13154
rect 19701 13096 19706 13152
rect 19762 13096 20350 13152
rect 20406 13096 20411 13152
rect 19701 13094 20411 13096
rect 19701 13091 19767 13094
rect 20345 13091 20411 13094
rect 6626 13088 6942 13089
rect 6626 13024 6632 13088
rect 6696 13024 6712 13088
rect 6776 13024 6792 13088
rect 6856 13024 6872 13088
rect 6936 13024 6942 13088
rect 6626 13023 6942 13024
rect 12307 13088 12623 13089
rect 12307 13024 12313 13088
rect 12377 13024 12393 13088
rect 12457 13024 12473 13088
rect 12537 13024 12553 13088
rect 12617 13024 12623 13088
rect 12307 13023 12623 13024
rect 17988 13088 18304 13089
rect 17988 13024 17994 13088
rect 18058 13024 18074 13088
rect 18138 13024 18154 13088
rect 18218 13024 18234 13088
rect 18298 13024 18304 13088
rect 17988 13023 18304 13024
rect 23669 13088 23985 13089
rect 23669 13024 23675 13088
rect 23739 13024 23755 13088
rect 23819 13024 23835 13088
rect 23899 13024 23915 13088
rect 23979 13024 23985 13088
rect 23669 13023 23985 13024
rect 16113 13018 16179 13021
rect 17585 13018 17651 13021
rect 16113 13016 17651 13018
rect 16113 12960 16118 13016
rect 16174 12960 17590 13016
rect 17646 12960 17651 13016
rect 16113 12958 17651 12960
rect 16113 12955 16179 12958
rect 17585 12955 17651 12958
rect 15929 12882 15995 12885
rect 21265 12882 21331 12885
rect 15929 12880 21331 12882
rect 15929 12824 15934 12880
rect 15990 12824 21270 12880
rect 21326 12824 21331 12880
rect 15929 12822 21331 12824
rect 15929 12819 15995 12822
rect 21265 12819 21331 12822
rect 17401 12746 17467 12749
rect 17861 12746 17927 12749
rect 17401 12744 17927 12746
rect 17401 12688 17406 12744
rect 17462 12688 17866 12744
rect 17922 12688 17927 12744
rect 17401 12686 17927 12688
rect 17401 12683 17467 12686
rect 17861 12683 17927 12686
rect 20253 12610 20319 12613
rect 20253 12608 20730 12610
rect 20253 12552 20258 12608
rect 20314 12552 20730 12608
rect 20253 12550 20730 12552
rect 20253 12547 20319 12550
rect 3786 12544 4102 12545
rect 3786 12480 3792 12544
rect 3856 12480 3872 12544
rect 3936 12480 3952 12544
rect 4016 12480 4032 12544
rect 4096 12480 4102 12544
rect 3786 12479 4102 12480
rect 9467 12544 9783 12545
rect 9467 12480 9473 12544
rect 9537 12480 9553 12544
rect 9617 12480 9633 12544
rect 9697 12480 9713 12544
rect 9777 12480 9783 12544
rect 9467 12479 9783 12480
rect 15148 12544 15464 12545
rect 15148 12480 15154 12544
rect 15218 12480 15234 12544
rect 15298 12480 15314 12544
rect 15378 12480 15394 12544
rect 15458 12480 15464 12544
rect 15148 12479 15464 12480
rect 2773 12474 2839 12477
rect 3325 12474 3391 12477
rect 2773 12472 3391 12474
rect 2773 12416 2778 12472
rect 2834 12416 3330 12472
rect 3386 12416 3391 12472
rect 2773 12414 3391 12416
rect 2773 12411 2839 12414
rect 3325 12411 3391 12414
rect 13169 12340 13235 12341
rect 13118 12338 13124 12340
rect 13078 12278 13124 12338
rect 13188 12336 13235 12340
rect 13230 12280 13235 12336
rect 13118 12276 13124 12278
rect 13188 12276 13235 12280
rect 13169 12275 13235 12276
rect 14273 12202 14339 12205
rect 17217 12202 17283 12205
rect 14273 12200 17283 12202
rect 14273 12144 14278 12200
rect 14334 12144 17222 12200
rect 17278 12144 17283 12200
rect 14273 12142 17283 12144
rect 20670 12202 20730 12550
rect 20829 12544 21145 12545
rect 20829 12480 20835 12544
rect 20899 12480 20915 12544
rect 20979 12480 20995 12544
rect 21059 12480 21075 12544
rect 21139 12480 21145 12544
rect 20829 12479 21145 12480
rect 21541 12202 21607 12205
rect 20670 12200 21607 12202
rect 20670 12144 21546 12200
rect 21602 12144 21607 12200
rect 20670 12142 21607 12144
rect 14273 12139 14339 12142
rect 17217 12139 17283 12142
rect 21541 12139 21607 12142
rect 6626 12000 6942 12001
rect 6626 11936 6632 12000
rect 6696 11936 6712 12000
rect 6776 11936 6792 12000
rect 6856 11936 6872 12000
rect 6936 11936 6942 12000
rect 6626 11935 6942 11936
rect 12307 12000 12623 12001
rect 12307 11936 12313 12000
rect 12377 11936 12393 12000
rect 12457 11936 12473 12000
rect 12537 11936 12553 12000
rect 12617 11936 12623 12000
rect 12307 11935 12623 11936
rect 17988 12000 18304 12001
rect 17988 11936 17994 12000
rect 18058 11936 18074 12000
rect 18138 11936 18154 12000
rect 18218 11936 18234 12000
rect 18298 11936 18304 12000
rect 17988 11935 18304 11936
rect 23669 12000 23985 12001
rect 23669 11936 23675 12000
rect 23739 11936 23755 12000
rect 23819 11936 23835 12000
rect 23899 11936 23915 12000
rect 23979 11936 23985 12000
rect 23669 11935 23985 11936
rect 12617 11794 12683 11797
rect 14774 11794 14780 11796
rect 12617 11792 14780 11794
rect 12617 11736 12622 11792
rect 12678 11736 14780 11792
rect 12617 11734 14780 11736
rect 12617 11731 12683 11734
rect 14774 11732 14780 11734
rect 14844 11794 14850 11796
rect 15101 11794 15167 11797
rect 14844 11792 15167 11794
rect 14844 11736 15106 11792
rect 15162 11736 15167 11792
rect 14844 11734 15167 11736
rect 14844 11732 14850 11734
rect 15101 11731 15167 11734
rect 3786 11456 4102 11457
rect 3786 11392 3792 11456
rect 3856 11392 3872 11456
rect 3936 11392 3952 11456
rect 4016 11392 4032 11456
rect 4096 11392 4102 11456
rect 3786 11391 4102 11392
rect 9467 11456 9783 11457
rect 9467 11392 9473 11456
rect 9537 11392 9553 11456
rect 9617 11392 9633 11456
rect 9697 11392 9713 11456
rect 9777 11392 9783 11456
rect 9467 11391 9783 11392
rect 15148 11456 15464 11457
rect 15148 11392 15154 11456
rect 15218 11392 15234 11456
rect 15298 11392 15314 11456
rect 15378 11392 15394 11456
rect 15458 11392 15464 11456
rect 15148 11391 15464 11392
rect 20829 11456 21145 11457
rect 20829 11392 20835 11456
rect 20899 11392 20915 11456
rect 20979 11392 20995 11456
rect 21059 11392 21075 11456
rect 21139 11392 21145 11456
rect 20829 11391 21145 11392
rect 14733 11250 14799 11253
rect 14917 11250 14983 11253
rect 14733 11248 14983 11250
rect 14733 11192 14738 11248
rect 14794 11192 14922 11248
rect 14978 11192 14983 11248
rect 14733 11190 14983 11192
rect 14733 11187 14799 11190
rect 14917 11187 14983 11190
rect 18597 11250 18663 11253
rect 21173 11250 21239 11253
rect 18597 11248 21239 11250
rect 18597 11192 18602 11248
rect 18658 11192 21178 11248
rect 21234 11192 21239 11248
rect 18597 11190 21239 11192
rect 18597 11187 18663 11190
rect 21173 11187 21239 11190
rect 14273 11114 14339 11117
rect 14917 11114 14983 11117
rect 14273 11112 14983 11114
rect 14273 11056 14278 11112
rect 14334 11056 14922 11112
rect 14978 11056 14983 11112
rect 14273 11054 14983 11056
rect 14273 11051 14339 11054
rect 14917 11051 14983 11054
rect 18229 11114 18295 11117
rect 18505 11114 18571 11117
rect 18229 11112 18571 11114
rect 18229 11056 18234 11112
rect 18290 11056 18510 11112
rect 18566 11056 18571 11112
rect 18229 11054 18571 11056
rect 18229 11051 18295 11054
rect 18505 11051 18571 11054
rect 13077 10978 13143 10981
rect 14181 10978 14247 10981
rect 15561 10978 15627 10981
rect 13077 10976 15627 10978
rect 13077 10920 13082 10976
rect 13138 10920 14186 10976
rect 14242 10920 15566 10976
rect 15622 10920 15627 10976
rect 13077 10918 15627 10920
rect 13077 10915 13143 10918
rect 14181 10915 14247 10918
rect 15561 10915 15627 10918
rect 6626 10912 6942 10913
rect 6626 10848 6632 10912
rect 6696 10848 6712 10912
rect 6776 10848 6792 10912
rect 6856 10848 6872 10912
rect 6936 10848 6942 10912
rect 6626 10847 6942 10848
rect 12307 10912 12623 10913
rect 12307 10848 12313 10912
rect 12377 10848 12393 10912
rect 12457 10848 12473 10912
rect 12537 10848 12553 10912
rect 12617 10848 12623 10912
rect 12307 10847 12623 10848
rect 17988 10912 18304 10913
rect 17988 10848 17994 10912
rect 18058 10848 18074 10912
rect 18138 10848 18154 10912
rect 18218 10848 18234 10912
rect 18298 10848 18304 10912
rect 17988 10847 18304 10848
rect 23669 10912 23985 10913
rect 23669 10848 23675 10912
rect 23739 10848 23755 10912
rect 23819 10848 23835 10912
rect 23899 10848 23915 10912
rect 23979 10848 23985 10912
rect 23669 10847 23985 10848
rect 13445 10842 13511 10845
rect 13905 10842 13971 10845
rect 15101 10842 15167 10845
rect 13445 10840 15167 10842
rect 13445 10784 13450 10840
rect 13506 10784 13910 10840
rect 13966 10784 15106 10840
rect 15162 10784 15167 10840
rect 13445 10782 15167 10784
rect 13445 10779 13511 10782
rect 13905 10779 13971 10782
rect 15101 10779 15167 10782
rect 5390 10644 5396 10708
rect 5460 10706 5466 10708
rect 10501 10706 10567 10709
rect 5460 10704 10567 10706
rect 5460 10648 10506 10704
rect 10562 10648 10567 10704
rect 5460 10646 10567 10648
rect 5460 10644 5466 10646
rect 10501 10643 10567 10646
rect 18689 10706 18755 10709
rect 19057 10706 19123 10709
rect 18689 10704 19123 10706
rect 18689 10648 18694 10704
rect 18750 10648 19062 10704
rect 19118 10648 19123 10704
rect 18689 10646 19123 10648
rect 18689 10643 18755 10646
rect 19057 10643 19123 10646
rect 22318 10644 22324 10708
rect 22388 10706 22394 10708
rect 22645 10706 22711 10709
rect 22388 10704 22711 10706
rect 22388 10648 22650 10704
rect 22706 10648 22711 10704
rect 22388 10646 22711 10648
rect 22388 10644 22394 10646
rect 22645 10643 22711 10646
rect 7281 10572 7347 10573
rect 7230 10508 7236 10572
rect 7300 10570 7347 10572
rect 7300 10568 7392 10570
rect 7342 10512 7392 10568
rect 7300 10510 7392 10512
rect 7300 10508 7347 10510
rect 7281 10507 7347 10508
rect 3786 10368 4102 10369
rect 3786 10304 3792 10368
rect 3856 10304 3872 10368
rect 3936 10304 3952 10368
rect 4016 10304 4032 10368
rect 4096 10304 4102 10368
rect 3786 10303 4102 10304
rect 9467 10368 9783 10369
rect 9467 10304 9473 10368
rect 9537 10304 9553 10368
rect 9617 10304 9633 10368
rect 9697 10304 9713 10368
rect 9777 10304 9783 10368
rect 9467 10303 9783 10304
rect 15148 10368 15464 10369
rect 15148 10304 15154 10368
rect 15218 10304 15234 10368
rect 15298 10304 15314 10368
rect 15378 10304 15394 10368
rect 15458 10304 15464 10368
rect 15148 10303 15464 10304
rect 20829 10368 21145 10369
rect 20829 10304 20835 10368
rect 20899 10304 20915 10368
rect 20979 10304 20995 10368
rect 21059 10304 21075 10368
rect 21139 10304 21145 10368
rect 20829 10303 21145 10304
rect 5165 10026 5231 10029
rect 7005 10026 7071 10029
rect 5165 10024 7071 10026
rect 5165 9968 5170 10024
rect 5226 9968 7010 10024
rect 7066 9968 7071 10024
rect 5165 9966 7071 9968
rect 5165 9963 5231 9966
rect 7005 9963 7071 9966
rect 17493 10026 17559 10029
rect 17718 10026 17724 10028
rect 17493 10024 17724 10026
rect 17493 9968 17498 10024
rect 17554 9968 17724 10024
rect 17493 9966 17724 9968
rect 17493 9963 17559 9966
rect 17718 9964 17724 9966
rect 17788 9964 17794 10028
rect 10358 9828 10364 9892
rect 10428 9890 10434 9892
rect 10501 9890 10567 9893
rect 10428 9888 10567 9890
rect 10428 9832 10506 9888
rect 10562 9832 10567 9888
rect 10428 9830 10567 9832
rect 10428 9828 10434 9830
rect 10501 9827 10567 9830
rect 6626 9824 6942 9825
rect 6626 9760 6632 9824
rect 6696 9760 6712 9824
rect 6776 9760 6792 9824
rect 6856 9760 6872 9824
rect 6936 9760 6942 9824
rect 6626 9759 6942 9760
rect 12307 9824 12623 9825
rect 12307 9760 12313 9824
rect 12377 9760 12393 9824
rect 12457 9760 12473 9824
rect 12537 9760 12553 9824
rect 12617 9760 12623 9824
rect 12307 9759 12623 9760
rect 17988 9824 18304 9825
rect 17988 9760 17994 9824
rect 18058 9760 18074 9824
rect 18138 9760 18154 9824
rect 18218 9760 18234 9824
rect 18298 9760 18304 9824
rect 17988 9759 18304 9760
rect 23669 9824 23985 9825
rect 23669 9760 23675 9824
rect 23739 9760 23755 9824
rect 23819 9760 23835 9824
rect 23899 9760 23915 9824
rect 23979 9760 23985 9824
rect 23669 9759 23985 9760
rect 3509 9482 3575 9485
rect 5349 9482 5415 9485
rect 3509 9480 5415 9482
rect 3509 9424 3514 9480
rect 3570 9424 5354 9480
rect 5410 9424 5415 9480
rect 3509 9422 5415 9424
rect 3509 9419 3575 9422
rect 5349 9419 5415 9422
rect 5717 9482 5783 9485
rect 9121 9482 9187 9485
rect 9489 9482 9555 9485
rect 5717 9480 9555 9482
rect 5717 9424 5722 9480
rect 5778 9424 9126 9480
rect 9182 9424 9494 9480
rect 9550 9424 9555 9480
rect 5717 9422 9555 9424
rect 5717 9419 5783 9422
rect 9121 9419 9187 9422
rect 9489 9419 9555 9422
rect 5809 9346 5875 9349
rect 6637 9346 6703 9349
rect 5809 9344 6703 9346
rect 5809 9288 5814 9344
rect 5870 9288 6642 9344
rect 6698 9288 6703 9344
rect 5809 9286 6703 9288
rect 5809 9283 5875 9286
rect 6637 9283 6703 9286
rect 3786 9280 4102 9281
rect 3786 9216 3792 9280
rect 3856 9216 3872 9280
rect 3936 9216 3952 9280
rect 4016 9216 4032 9280
rect 4096 9216 4102 9280
rect 3786 9215 4102 9216
rect 9467 9280 9783 9281
rect 9467 9216 9473 9280
rect 9537 9216 9553 9280
rect 9617 9216 9633 9280
rect 9697 9216 9713 9280
rect 9777 9216 9783 9280
rect 9467 9215 9783 9216
rect 15148 9280 15464 9281
rect 15148 9216 15154 9280
rect 15218 9216 15234 9280
rect 15298 9216 15314 9280
rect 15378 9216 15394 9280
rect 15458 9216 15464 9280
rect 15148 9215 15464 9216
rect 20829 9280 21145 9281
rect 20829 9216 20835 9280
rect 20899 9216 20915 9280
rect 20979 9216 20995 9280
rect 21059 9216 21075 9280
rect 21139 9216 21145 9280
rect 20829 9215 21145 9216
rect 6626 8736 6942 8737
rect 6626 8672 6632 8736
rect 6696 8672 6712 8736
rect 6776 8672 6792 8736
rect 6856 8672 6872 8736
rect 6936 8672 6942 8736
rect 6626 8671 6942 8672
rect 12307 8736 12623 8737
rect 12307 8672 12313 8736
rect 12377 8672 12393 8736
rect 12457 8672 12473 8736
rect 12537 8672 12553 8736
rect 12617 8672 12623 8736
rect 12307 8671 12623 8672
rect 17988 8736 18304 8737
rect 17988 8672 17994 8736
rect 18058 8672 18074 8736
rect 18138 8672 18154 8736
rect 18218 8672 18234 8736
rect 18298 8672 18304 8736
rect 17988 8671 18304 8672
rect 23669 8736 23985 8737
rect 23669 8672 23675 8736
rect 23739 8672 23755 8736
rect 23819 8672 23835 8736
rect 23899 8672 23915 8736
rect 23979 8672 23985 8736
rect 23669 8671 23985 8672
rect 14733 8530 14799 8533
rect 18229 8530 18295 8533
rect 14733 8528 18295 8530
rect 14733 8472 14738 8528
rect 14794 8472 18234 8528
rect 18290 8472 18295 8528
rect 14733 8470 18295 8472
rect 14733 8467 14799 8470
rect 18229 8467 18295 8470
rect 16246 8332 16252 8396
rect 16316 8394 16322 8396
rect 22277 8394 22343 8397
rect 16316 8392 22343 8394
rect 16316 8336 22282 8392
rect 22338 8336 22343 8392
rect 16316 8334 22343 8336
rect 16316 8332 16322 8334
rect 22277 8331 22343 8334
rect 3786 8192 4102 8193
rect 3786 8128 3792 8192
rect 3856 8128 3872 8192
rect 3936 8128 3952 8192
rect 4016 8128 4032 8192
rect 4096 8128 4102 8192
rect 3786 8127 4102 8128
rect 9467 8192 9783 8193
rect 9467 8128 9473 8192
rect 9537 8128 9553 8192
rect 9617 8128 9633 8192
rect 9697 8128 9713 8192
rect 9777 8128 9783 8192
rect 9467 8127 9783 8128
rect 15148 8192 15464 8193
rect 15148 8128 15154 8192
rect 15218 8128 15234 8192
rect 15298 8128 15314 8192
rect 15378 8128 15394 8192
rect 15458 8128 15464 8192
rect 15148 8127 15464 8128
rect 20829 8192 21145 8193
rect 20829 8128 20835 8192
rect 20899 8128 20915 8192
rect 20979 8128 20995 8192
rect 21059 8128 21075 8192
rect 21139 8128 21145 8192
rect 20829 8127 21145 8128
rect 8477 7986 8543 7989
rect 14825 7986 14891 7989
rect 8477 7984 14891 7986
rect 8477 7928 8482 7984
rect 8538 7928 14830 7984
rect 14886 7928 14891 7984
rect 8477 7926 14891 7928
rect 8477 7923 8543 7926
rect 14825 7923 14891 7926
rect 6626 7648 6942 7649
rect 6626 7584 6632 7648
rect 6696 7584 6712 7648
rect 6776 7584 6792 7648
rect 6856 7584 6872 7648
rect 6936 7584 6942 7648
rect 6626 7583 6942 7584
rect 12307 7648 12623 7649
rect 12307 7584 12313 7648
rect 12377 7584 12393 7648
rect 12457 7584 12473 7648
rect 12537 7584 12553 7648
rect 12617 7584 12623 7648
rect 12307 7583 12623 7584
rect 17988 7648 18304 7649
rect 17988 7584 17994 7648
rect 18058 7584 18074 7648
rect 18138 7584 18154 7648
rect 18218 7584 18234 7648
rect 18298 7584 18304 7648
rect 17988 7583 18304 7584
rect 23669 7648 23985 7649
rect 23669 7584 23675 7648
rect 23739 7584 23755 7648
rect 23819 7584 23835 7648
rect 23899 7584 23915 7648
rect 23979 7584 23985 7648
rect 23669 7583 23985 7584
rect 11145 7306 11211 7309
rect 12893 7306 12959 7309
rect 11145 7304 12959 7306
rect 11145 7248 11150 7304
rect 11206 7248 12898 7304
rect 12954 7248 12959 7304
rect 11145 7246 12959 7248
rect 11145 7243 11211 7246
rect 12893 7243 12959 7246
rect 3786 7104 4102 7105
rect 3786 7040 3792 7104
rect 3856 7040 3872 7104
rect 3936 7040 3952 7104
rect 4016 7040 4032 7104
rect 4096 7040 4102 7104
rect 3786 7039 4102 7040
rect 9467 7104 9783 7105
rect 9467 7040 9473 7104
rect 9537 7040 9553 7104
rect 9617 7040 9633 7104
rect 9697 7040 9713 7104
rect 9777 7040 9783 7104
rect 9467 7039 9783 7040
rect 15148 7104 15464 7105
rect 15148 7040 15154 7104
rect 15218 7040 15234 7104
rect 15298 7040 15314 7104
rect 15378 7040 15394 7104
rect 15458 7040 15464 7104
rect 15148 7039 15464 7040
rect 20829 7104 21145 7105
rect 20829 7040 20835 7104
rect 20899 7040 20915 7104
rect 20979 7040 20995 7104
rect 21059 7040 21075 7104
rect 21139 7040 21145 7104
rect 20829 7039 21145 7040
rect 21398 6836 21404 6900
rect 21468 6898 21474 6900
rect 21541 6898 21607 6901
rect 21468 6896 21607 6898
rect 21468 6840 21546 6896
rect 21602 6840 21607 6896
rect 21468 6838 21607 6840
rect 21468 6836 21474 6838
rect 21541 6835 21607 6838
rect 5349 6762 5415 6765
rect 13629 6762 13695 6765
rect 5349 6760 13695 6762
rect 5349 6704 5354 6760
rect 5410 6704 13634 6760
rect 13690 6704 13695 6760
rect 5349 6702 13695 6704
rect 5349 6699 5415 6702
rect 13629 6699 13695 6702
rect 9949 6626 10015 6629
rect 10317 6626 10383 6629
rect 11973 6626 12039 6629
rect 12157 6626 12223 6629
rect 9949 6624 12223 6626
rect 9949 6568 9954 6624
rect 10010 6568 10322 6624
rect 10378 6568 11978 6624
rect 12034 6568 12162 6624
rect 12218 6568 12223 6624
rect 9949 6566 12223 6568
rect 9949 6563 10015 6566
rect 10317 6563 10383 6566
rect 11973 6563 12039 6566
rect 12157 6563 12223 6566
rect 6626 6560 6942 6561
rect 6626 6496 6632 6560
rect 6696 6496 6712 6560
rect 6776 6496 6792 6560
rect 6856 6496 6872 6560
rect 6936 6496 6942 6560
rect 6626 6495 6942 6496
rect 12307 6560 12623 6561
rect 12307 6496 12313 6560
rect 12377 6496 12393 6560
rect 12457 6496 12473 6560
rect 12537 6496 12553 6560
rect 12617 6496 12623 6560
rect 12307 6495 12623 6496
rect 17988 6560 18304 6561
rect 17988 6496 17994 6560
rect 18058 6496 18074 6560
rect 18138 6496 18154 6560
rect 18218 6496 18234 6560
rect 18298 6496 18304 6560
rect 17988 6495 18304 6496
rect 23669 6560 23985 6561
rect 23669 6496 23675 6560
rect 23739 6496 23755 6560
rect 23819 6496 23835 6560
rect 23899 6496 23915 6560
rect 23979 6496 23985 6560
rect 23669 6495 23985 6496
rect 8293 6490 8359 6493
rect 8937 6490 9003 6493
rect 8293 6488 9003 6490
rect 8293 6432 8298 6488
rect 8354 6432 8942 6488
rect 8998 6432 9003 6488
rect 8293 6430 9003 6432
rect 8293 6427 8359 6430
rect 8937 6427 9003 6430
rect 7649 6354 7715 6357
rect 8845 6354 8911 6357
rect 7649 6352 8911 6354
rect 7649 6296 7654 6352
rect 7710 6296 8850 6352
rect 8906 6296 8911 6352
rect 7649 6294 8911 6296
rect 7649 6291 7715 6294
rect 8845 6291 8911 6294
rect 17953 6354 18019 6357
rect 19149 6354 19215 6357
rect 17953 6352 19215 6354
rect 17953 6296 17958 6352
rect 18014 6296 19154 6352
rect 19210 6296 19215 6352
rect 17953 6294 19215 6296
rect 17953 6291 18019 6294
rect 19149 6291 19215 6294
rect 5165 6218 5231 6221
rect 12617 6218 12683 6221
rect 5165 6216 12683 6218
rect 5165 6160 5170 6216
rect 5226 6160 12622 6216
rect 12678 6160 12683 6216
rect 5165 6158 12683 6160
rect 5165 6155 5231 6158
rect 12617 6155 12683 6158
rect 3786 6016 4102 6017
rect 3786 5952 3792 6016
rect 3856 5952 3872 6016
rect 3936 5952 3952 6016
rect 4016 5952 4032 6016
rect 4096 5952 4102 6016
rect 3786 5951 4102 5952
rect 9467 6016 9783 6017
rect 9467 5952 9473 6016
rect 9537 5952 9553 6016
rect 9617 5952 9633 6016
rect 9697 5952 9713 6016
rect 9777 5952 9783 6016
rect 9467 5951 9783 5952
rect 15148 6016 15464 6017
rect 15148 5952 15154 6016
rect 15218 5952 15234 6016
rect 15298 5952 15314 6016
rect 15378 5952 15394 6016
rect 15458 5952 15464 6016
rect 15148 5951 15464 5952
rect 20829 6016 21145 6017
rect 20829 5952 20835 6016
rect 20899 5952 20915 6016
rect 20979 5952 20995 6016
rect 21059 5952 21075 6016
rect 21139 5952 21145 6016
rect 20829 5951 21145 5952
rect 11697 5946 11763 5949
rect 14825 5946 14891 5949
rect 11697 5944 14891 5946
rect 11697 5888 11702 5944
rect 11758 5888 14830 5944
rect 14886 5888 14891 5944
rect 11697 5886 14891 5888
rect 11697 5883 11763 5886
rect 14825 5883 14891 5886
rect 10133 5810 10199 5813
rect 10869 5810 10935 5813
rect 12249 5810 12315 5813
rect 10133 5808 12315 5810
rect 10133 5752 10138 5808
rect 10194 5752 10874 5808
rect 10930 5752 12254 5808
rect 12310 5752 12315 5808
rect 10133 5750 12315 5752
rect 14828 5810 14888 5883
rect 16021 5810 16087 5813
rect 14828 5808 16087 5810
rect 14828 5752 16026 5808
rect 16082 5752 16087 5808
rect 14828 5750 16087 5752
rect 10133 5747 10199 5750
rect 10869 5747 10935 5750
rect 12249 5747 12315 5750
rect 16021 5747 16087 5750
rect 9121 5538 9187 5541
rect 10358 5538 10364 5540
rect 9121 5536 10364 5538
rect 9121 5480 9126 5536
rect 9182 5480 10364 5536
rect 9121 5478 10364 5480
rect 9121 5475 9187 5478
rect 10358 5476 10364 5478
rect 10428 5476 10434 5540
rect 6626 5472 6942 5473
rect 6626 5408 6632 5472
rect 6696 5408 6712 5472
rect 6776 5408 6792 5472
rect 6856 5408 6872 5472
rect 6936 5408 6942 5472
rect 6626 5407 6942 5408
rect 12307 5472 12623 5473
rect 12307 5408 12313 5472
rect 12377 5408 12393 5472
rect 12457 5408 12473 5472
rect 12537 5408 12553 5472
rect 12617 5408 12623 5472
rect 12307 5407 12623 5408
rect 17988 5472 18304 5473
rect 17988 5408 17994 5472
rect 18058 5408 18074 5472
rect 18138 5408 18154 5472
rect 18218 5408 18234 5472
rect 18298 5408 18304 5472
rect 17988 5407 18304 5408
rect 23669 5472 23985 5473
rect 23669 5408 23675 5472
rect 23739 5408 23755 5472
rect 23819 5408 23835 5472
rect 23899 5408 23915 5472
rect 23979 5408 23985 5472
rect 23669 5407 23985 5408
rect 14273 5266 14339 5269
rect 16665 5266 16731 5269
rect 14273 5264 16731 5266
rect 14273 5208 14278 5264
rect 14334 5208 16670 5264
rect 16726 5208 16731 5264
rect 14273 5206 16731 5208
rect 14273 5203 14339 5206
rect 16665 5203 16731 5206
rect 6269 5130 6335 5133
rect 7230 5130 7236 5132
rect 6269 5128 7236 5130
rect 6269 5072 6274 5128
rect 6330 5072 7236 5128
rect 6269 5070 7236 5072
rect 6269 5067 6335 5070
rect 7230 5068 7236 5070
rect 7300 5130 7306 5132
rect 9673 5130 9739 5133
rect 7300 5128 9739 5130
rect 7300 5072 9678 5128
rect 9734 5072 9739 5128
rect 7300 5070 9739 5072
rect 7300 5068 7306 5070
rect 9673 5067 9739 5070
rect 14549 5130 14615 5133
rect 14825 5130 14891 5133
rect 14549 5128 14891 5130
rect 14549 5072 14554 5128
rect 14610 5072 14830 5128
rect 14886 5072 14891 5128
rect 14549 5070 14891 5072
rect 14549 5067 14615 5070
rect 14825 5067 14891 5070
rect 3786 4928 4102 4929
rect 3786 4864 3792 4928
rect 3856 4864 3872 4928
rect 3936 4864 3952 4928
rect 4016 4864 4032 4928
rect 4096 4864 4102 4928
rect 3786 4863 4102 4864
rect 9467 4928 9783 4929
rect 9467 4864 9473 4928
rect 9537 4864 9553 4928
rect 9617 4864 9633 4928
rect 9697 4864 9713 4928
rect 9777 4864 9783 4928
rect 9467 4863 9783 4864
rect 15148 4928 15464 4929
rect 15148 4864 15154 4928
rect 15218 4864 15234 4928
rect 15298 4864 15314 4928
rect 15378 4864 15394 4928
rect 15458 4864 15464 4928
rect 15148 4863 15464 4864
rect 20829 4928 21145 4929
rect 20829 4864 20835 4928
rect 20899 4864 20915 4928
rect 20979 4864 20995 4928
rect 21059 4864 21075 4928
rect 21139 4864 21145 4928
rect 20829 4863 21145 4864
rect 17718 4660 17724 4724
rect 17788 4722 17794 4724
rect 22093 4722 22159 4725
rect 17788 4720 22159 4722
rect 17788 4664 22098 4720
rect 22154 4664 22159 4720
rect 17788 4662 22159 4664
rect 17788 4660 17794 4662
rect 22093 4659 22159 4662
rect 6626 4384 6942 4385
rect 6626 4320 6632 4384
rect 6696 4320 6712 4384
rect 6776 4320 6792 4384
rect 6856 4320 6872 4384
rect 6936 4320 6942 4384
rect 6626 4319 6942 4320
rect 12307 4384 12623 4385
rect 12307 4320 12313 4384
rect 12377 4320 12393 4384
rect 12457 4320 12473 4384
rect 12537 4320 12553 4384
rect 12617 4320 12623 4384
rect 12307 4319 12623 4320
rect 17988 4384 18304 4385
rect 17988 4320 17994 4384
rect 18058 4320 18074 4384
rect 18138 4320 18154 4384
rect 18218 4320 18234 4384
rect 18298 4320 18304 4384
rect 17988 4319 18304 4320
rect 23669 4384 23985 4385
rect 23669 4320 23675 4384
rect 23739 4320 23755 4384
rect 23819 4320 23835 4384
rect 23899 4320 23915 4384
rect 23979 4320 23985 4384
rect 23669 4319 23985 4320
rect 8017 4178 8083 4181
rect 16113 4178 16179 4181
rect 8017 4176 16179 4178
rect 8017 4120 8022 4176
rect 8078 4120 16118 4176
rect 16174 4120 16179 4176
rect 8017 4118 16179 4120
rect 8017 4115 8083 4118
rect 16113 4115 16179 4118
rect 8661 4042 8727 4045
rect 11697 4042 11763 4045
rect 8661 4040 11763 4042
rect 8661 3984 8666 4040
rect 8722 3984 11702 4040
rect 11758 3984 11763 4040
rect 8661 3982 11763 3984
rect 8661 3979 8727 3982
rect 11697 3979 11763 3982
rect 3786 3840 4102 3841
rect 3786 3776 3792 3840
rect 3856 3776 3872 3840
rect 3936 3776 3952 3840
rect 4016 3776 4032 3840
rect 4096 3776 4102 3840
rect 3786 3775 4102 3776
rect 9467 3840 9783 3841
rect 9467 3776 9473 3840
rect 9537 3776 9553 3840
rect 9617 3776 9633 3840
rect 9697 3776 9713 3840
rect 9777 3776 9783 3840
rect 9467 3775 9783 3776
rect 15148 3840 15464 3841
rect 15148 3776 15154 3840
rect 15218 3776 15234 3840
rect 15298 3776 15314 3840
rect 15378 3776 15394 3840
rect 15458 3776 15464 3840
rect 15148 3775 15464 3776
rect 20829 3840 21145 3841
rect 20829 3776 20835 3840
rect 20899 3776 20915 3840
rect 20979 3776 20995 3840
rect 21059 3776 21075 3840
rect 21139 3776 21145 3840
rect 20829 3775 21145 3776
rect 4337 3770 4403 3773
rect 7649 3770 7715 3773
rect 4337 3768 7715 3770
rect 4337 3712 4342 3768
rect 4398 3712 7654 3768
rect 7710 3712 7715 3768
rect 4337 3710 7715 3712
rect 4337 3707 4403 3710
rect 7649 3707 7715 3710
rect 7189 3634 7255 3637
rect 16573 3634 16639 3637
rect 7189 3632 16639 3634
rect 7189 3576 7194 3632
rect 7250 3576 16578 3632
rect 16634 3576 16639 3632
rect 7189 3574 16639 3576
rect 7189 3571 7255 3574
rect 16573 3571 16639 3574
rect 3325 3498 3391 3501
rect 14825 3498 14891 3501
rect 16941 3498 17007 3501
rect 20345 3498 20411 3501
rect 3325 3496 17007 3498
rect 3325 3440 3330 3496
rect 3386 3440 14830 3496
rect 14886 3440 16946 3496
rect 17002 3440 17007 3496
rect 3325 3438 17007 3440
rect 3325 3435 3391 3438
rect 14825 3435 14891 3438
rect 16941 3435 17007 3438
rect 17864 3496 20411 3498
rect 17864 3440 20350 3496
rect 20406 3440 20411 3496
rect 17864 3438 20411 3440
rect 13629 3362 13695 3365
rect 17864 3362 17924 3438
rect 20345 3435 20411 3438
rect 13629 3360 17924 3362
rect 13629 3304 13634 3360
rect 13690 3304 17924 3360
rect 13629 3302 17924 3304
rect 13629 3299 13695 3302
rect 6626 3296 6942 3297
rect 6626 3232 6632 3296
rect 6696 3232 6712 3296
rect 6776 3232 6792 3296
rect 6856 3232 6872 3296
rect 6936 3232 6942 3296
rect 6626 3231 6942 3232
rect 12307 3296 12623 3297
rect 12307 3232 12313 3296
rect 12377 3232 12393 3296
rect 12457 3232 12473 3296
rect 12537 3232 12553 3296
rect 12617 3232 12623 3296
rect 12307 3231 12623 3232
rect 17988 3296 18304 3297
rect 17988 3232 17994 3296
rect 18058 3232 18074 3296
rect 18138 3232 18154 3296
rect 18218 3232 18234 3296
rect 18298 3232 18304 3296
rect 17988 3231 18304 3232
rect 23669 3296 23985 3297
rect 23669 3232 23675 3296
rect 23739 3232 23755 3296
rect 23819 3232 23835 3296
rect 23899 3232 23915 3296
rect 23979 3232 23985 3296
rect 23669 3231 23985 3232
rect 10961 3090 11027 3093
rect 17033 3090 17099 3093
rect 10961 3088 17099 3090
rect 10961 3032 10966 3088
rect 11022 3032 17038 3088
rect 17094 3032 17099 3088
rect 10961 3030 17099 3032
rect 10961 3027 11027 3030
rect 17033 3027 17099 3030
rect 5625 2954 5691 2957
rect 11053 2954 11119 2957
rect 5625 2952 11119 2954
rect 5625 2896 5630 2952
rect 5686 2896 11058 2952
rect 11114 2896 11119 2952
rect 5625 2894 11119 2896
rect 5625 2891 5691 2894
rect 11053 2891 11119 2894
rect 11237 2954 11303 2957
rect 18689 2954 18755 2957
rect 11237 2952 18755 2954
rect 11237 2896 11242 2952
rect 11298 2896 18694 2952
rect 18750 2896 18755 2952
rect 11237 2894 18755 2896
rect 11237 2891 11303 2894
rect 18689 2891 18755 2894
rect 3786 2752 4102 2753
rect 3786 2688 3792 2752
rect 3856 2688 3872 2752
rect 3936 2688 3952 2752
rect 4016 2688 4032 2752
rect 4096 2688 4102 2752
rect 3786 2687 4102 2688
rect 9467 2752 9783 2753
rect 9467 2688 9473 2752
rect 9537 2688 9553 2752
rect 9617 2688 9633 2752
rect 9697 2688 9713 2752
rect 9777 2688 9783 2752
rect 9467 2687 9783 2688
rect 15148 2752 15464 2753
rect 15148 2688 15154 2752
rect 15218 2688 15234 2752
rect 15298 2688 15314 2752
rect 15378 2688 15394 2752
rect 15458 2688 15464 2752
rect 15148 2687 15464 2688
rect 20829 2752 21145 2753
rect 20829 2688 20835 2752
rect 20899 2688 20915 2752
rect 20979 2688 20995 2752
rect 21059 2688 21075 2752
rect 21139 2688 21145 2752
rect 20829 2687 21145 2688
rect 6626 2208 6942 2209
rect 6626 2144 6632 2208
rect 6696 2144 6712 2208
rect 6776 2144 6792 2208
rect 6856 2144 6872 2208
rect 6936 2144 6942 2208
rect 6626 2143 6942 2144
rect 12307 2208 12623 2209
rect 12307 2144 12313 2208
rect 12377 2144 12393 2208
rect 12457 2144 12473 2208
rect 12537 2144 12553 2208
rect 12617 2144 12623 2208
rect 12307 2143 12623 2144
rect 17988 2208 18304 2209
rect 17988 2144 17994 2208
rect 18058 2144 18074 2208
rect 18138 2144 18154 2208
rect 18218 2144 18234 2208
rect 18298 2144 18304 2208
rect 17988 2143 18304 2144
rect 23669 2208 23985 2209
rect 23669 2144 23675 2208
rect 23739 2144 23755 2208
rect 23819 2144 23835 2208
rect 23899 2144 23915 2208
rect 23979 2144 23985 2208
rect 23669 2143 23985 2144
<< via3 >>
rect 3792 22332 3856 22336
rect 3792 22276 3796 22332
rect 3796 22276 3852 22332
rect 3852 22276 3856 22332
rect 3792 22272 3856 22276
rect 3872 22332 3936 22336
rect 3872 22276 3876 22332
rect 3876 22276 3932 22332
rect 3932 22276 3936 22332
rect 3872 22272 3936 22276
rect 3952 22332 4016 22336
rect 3952 22276 3956 22332
rect 3956 22276 4012 22332
rect 4012 22276 4016 22332
rect 3952 22272 4016 22276
rect 4032 22332 4096 22336
rect 4032 22276 4036 22332
rect 4036 22276 4092 22332
rect 4092 22276 4096 22332
rect 4032 22272 4096 22276
rect 9473 22332 9537 22336
rect 9473 22276 9477 22332
rect 9477 22276 9533 22332
rect 9533 22276 9537 22332
rect 9473 22272 9537 22276
rect 9553 22332 9617 22336
rect 9553 22276 9557 22332
rect 9557 22276 9613 22332
rect 9613 22276 9617 22332
rect 9553 22272 9617 22276
rect 9633 22332 9697 22336
rect 9633 22276 9637 22332
rect 9637 22276 9693 22332
rect 9693 22276 9697 22332
rect 9633 22272 9697 22276
rect 9713 22332 9777 22336
rect 9713 22276 9717 22332
rect 9717 22276 9773 22332
rect 9773 22276 9777 22332
rect 9713 22272 9777 22276
rect 15154 22332 15218 22336
rect 15154 22276 15158 22332
rect 15158 22276 15214 22332
rect 15214 22276 15218 22332
rect 15154 22272 15218 22276
rect 15234 22332 15298 22336
rect 15234 22276 15238 22332
rect 15238 22276 15294 22332
rect 15294 22276 15298 22332
rect 15234 22272 15298 22276
rect 15314 22332 15378 22336
rect 15314 22276 15318 22332
rect 15318 22276 15374 22332
rect 15374 22276 15378 22332
rect 15314 22272 15378 22276
rect 15394 22332 15458 22336
rect 15394 22276 15398 22332
rect 15398 22276 15454 22332
rect 15454 22276 15458 22332
rect 15394 22272 15458 22276
rect 20835 22332 20899 22336
rect 20835 22276 20839 22332
rect 20839 22276 20895 22332
rect 20895 22276 20899 22332
rect 20835 22272 20899 22276
rect 20915 22332 20979 22336
rect 20915 22276 20919 22332
rect 20919 22276 20975 22332
rect 20975 22276 20979 22332
rect 20915 22272 20979 22276
rect 20995 22332 21059 22336
rect 20995 22276 20999 22332
rect 20999 22276 21055 22332
rect 21055 22276 21059 22332
rect 20995 22272 21059 22276
rect 21075 22332 21139 22336
rect 21075 22276 21079 22332
rect 21079 22276 21135 22332
rect 21135 22276 21139 22332
rect 21075 22272 21139 22276
rect 6632 21788 6696 21792
rect 6632 21732 6636 21788
rect 6636 21732 6692 21788
rect 6692 21732 6696 21788
rect 6632 21728 6696 21732
rect 6712 21788 6776 21792
rect 6712 21732 6716 21788
rect 6716 21732 6772 21788
rect 6772 21732 6776 21788
rect 6712 21728 6776 21732
rect 6792 21788 6856 21792
rect 6792 21732 6796 21788
rect 6796 21732 6852 21788
rect 6852 21732 6856 21788
rect 6792 21728 6856 21732
rect 6872 21788 6936 21792
rect 6872 21732 6876 21788
rect 6876 21732 6932 21788
rect 6932 21732 6936 21788
rect 6872 21728 6936 21732
rect 12313 21788 12377 21792
rect 12313 21732 12317 21788
rect 12317 21732 12373 21788
rect 12373 21732 12377 21788
rect 12313 21728 12377 21732
rect 12393 21788 12457 21792
rect 12393 21732 12397 21788
rect 12397 21732 12453 21788
rect 12453 21732 12457 21788
rect 12393 21728 12457 21732
rect 12473 21788 12537 21792
rect 12473 21732 12477 21788
rect 12477 21732 12533 21788
rect 12533 21732 12537 21788
rect 12473 21728 12537 21732
rect 12553 21788 12617 21792
rect 12553 21732 12557 21788
rect 12557 21732 12613 21788
rect 12613 21732 12617 21788
rect 12553 21728 12617 21732
rect 17994 21788 18058 21792
rect 17994 21732 17998 21788
rect 17998 21732 18054 21788
rect 18054 21732 18058 21788
rect 17994 21728 18058 21732
rect 18074 21788 18138 21792
rect 18074 21732 18078 21788
rect 18078 21732 18134 21788
rect 18134 21732 18138 21788
rect 18074 21728 18138 21732
rect 18154 21788 18218 21792
rect 18154 21732 18158 21788
rect 18158 21732 18214 21788
rect 18214 21732 18218 21788
rect 18154 21728 18218 21732
rect 18234 21788 18298 21792
rect 18234 21732 18238 21788
rect 18238 21732 18294 21788
rect 18294 21732 18298 21788
rect 18234 21728 18298 21732
rect 23675 21788 23739 21792
rect 23675 21732 23679 21788
rect 23679 21732 23735 21788
rect 23735 21732 23739 21788
rect 23675 21728 23739 21732
rect 23755 21788 23819 21792
rect 23755 21732 23759 21788
rect 23759 21732 23815 21788
rect 23815 21732 23819 21788
rect 23755 21728 23819 21732
rect 23835 21788 23899 21792
rect 23835 21732 23839 21788
rect 23839 21732 23895 21788
rect 23895 21732 23899 21788
rect 23835 21728 23899 21732
rect 23915 21788 23979 21792
rect 23915 21732 23919 21788
rect 23919 21732 23975 21788
rect 23975 21732 23979 21788
rect 23915 21728 23979 21732
rect 3792 21244 3856 21248
rect 3792 21188 3796 21244
rect 3796 21188 3852 21244
rect 3852 21188 3856 21244
rect 3792 21184 3856 21188
rect 3872 21244 3936 21248
rect 3872 21188 3876 21244
rect 3876 21188 3932 21244
rect 3932 21188 3936 21244
rect 3872 21184 3936 21188
rect 3952 21244 4016 21248
rect 3952 21188 3956 21244
rect 3956 21188 4012 21244
rect 4012 21188 4016 21244
rect 3952 21184 4016 21188
rect 4032 21244 4096 21248
rect 4032 21188 4036 21244
rect 4036 21188 4092 21244
rect 4092 21188 4096 21244
rect 4032 21184 4096 21188
rect 9473 21244 9537 21248
rect 9473 21188 9477 21244
rect 9477 21188 9533 21244
rect 9533 21188 9537 21244
rect 9473 21184 9537 21188
rect 9553 21244 9617 21248
rect 9553 21188 9557 21244
rect 9557 21188 9613 21244
rect 9613 21188 9617 21244
rect 9553 21184 9617 21188
rect 9633 21244 9697 21248
rect 9633 21188 9637 21244
rect 9637 21188 9693 21244
rect 9693 21188 9697 21244
rect 9633 21184 9697 21188
rect 9713 21244 9777 21248
rect 9713 21188 9717 21244
rect 9717 21188 9773 21244
rect 9773 21188 9777 21244
rect 9713 21184 9777 21188
rect 15154 21244 15218 21248
rect 15154 21188 15158 21244
rect 15158 21188 15214 21244
rect 15214 21188 15218 21244
rect 15154 21184 15218 21188
rect 15234 21244 15298 21248
rect 15234 21188 15238 21244
rect 15238 21188 15294 21244
rect 15294 21188 15298 21244
rect 15234 21184 15298 21188
rect 15314 21244 15378 21248
rect 15314 21188 15318 21244
rect 15318 21188 15374 21244
rect 15374 21188 15378 21244
rect 15314 21184 15378 21188
rect 15394 21244 15458 21248
rect 15394 21188 15398 21244
rect 15398 21188 15454 21244
rect 15454 21188 15458 21244
rect 15394 21184 15458 21188
rect 20835 21244 20899 21248
rect 20835 21188 20839 21244
rect 20839 21188 20895 21244
rect 20895 21188 20899 21244
rect 20835 21184 20899 21188
rect 20915 21244 20979 21248
rect 20915 21188 20919 21244
rect 20919 21188 20975 21244
rect 20975 21188 20979 21244
rect 20915 21184 20979 21188
rect 20995 21244 21059 21248
rect 20995 21188 20999 21244
rect 20999 21188 21055 21244
rect 21055 21188 21059 21244
rect 20995 21184 21059 21188
rect 21075 21244 21139 21248
rect 21075 21188 21079 21244
rect 21079 21188 21135 21244
rect 21135 21188 21139 21244
rect 21075 21184 21139 21188
rect 13124 20768 13188 20772
rect 13124 20712 13138 20768
rect 13138 20712 13188 20768
rect 13124 20708 13188 20712
rect 14780 20708 14844 20772
rect 6632 20700 6696 20704
rect 6632 20644 6636 20700
rect 6636 20644 6692 20700
rect 6692 20644 6696 20700
rect 6632 20640 6696 20644
rect 6712 20700 6776 20704
rect 6712 20644 6716 20700
rect 6716 20644 6772 20700
rect 6772 20644 6776 20700
rect 6712 20640 6776 20644
rect 6792 20700 6856 20704
rect 6792 20644 6796 20700
rect 6796 20644 6852 20700
rect 6852 20644 6856 20700
rect 6792 20640 6856 20644
rect 6872 20700 6936 20704
rect 6872 20644 6876 20700
rect 6876 20644 6932 20700
rect 6932 20644 6936 20700
rect 6872 20640 6936 20644
rect 12313 20700 12377 20704
rect 12313 20644 12317 20700
rect 12317 20644 12373 20700
rect 12373 20644 12377 20700
rect 12313 20640 12377 20644
rect 12393 20700 12457 20704
rect 12393 20644 12397 20700
rect 12397 20644 12453 20700
rect 12453 20644 12457 20700
rect 12393 20640 12457 20644
rect 12473 20700 12537 20704
rect 12473 20644 12477 20700
rect 12477 20644 12533 20700
rect 12533 20644 12537 20700
rect 12473 20640 12537 20644
rect 12553 20700 12617 20704
rect 12553 20644 12557 20700
rect 12557 20644 12613 20700
rect 12613 20644 12617 20700
rect 12553 20640 12617 20644
rect 17994 20700 18058 20704
rect 17994 20644 17998 20700
rect 17998 20644 18054 20700
rect 18054 20644 18058 20700
rect 17994 20640 18058 20644
rect 18074 20700 18138 20704
rect 18074 20644 18078 20700
rect 18078 20644 18134 20700
rect 18134 20644 18138 20700
rect 18074 20640 18138 20644
rect 18154 20700 18218 20704
rect 18154 20644 18158 20700
rect 18158 20644 18214 20700
rect 18214 20644 18218 20700
rect 18154 20640 18218 20644
rect 18234 20700 18298 20704
rect 18234 20644 18238 20700
rect 18238 20644 18294 20700
rect 18294 20644 18298 20700
rect 18234 20640 18298 20644
rect 23675 20700 23739 20704
rect 23675 20644 23679 20700
rect 23679 20644 23735 20700
rect 23735 20644 23739 20700
rect 23675 20640 23739 20644
rect 23755 20700 23819 20704
rect 23755 20644 23759 20700
rect 23759 20644 23815 20700
rect 23815 20644 23819 20700
rect 23755 20640 23819 20644
rect 23835 20700 23899 20704
rect 23835 20644 23839 20700
rect 23839 20644 23895 20700
rect 23895 20644 23899 20700
rect 23835 20640 23899 20644
rect 23915 20700 23979 20704
rect 23915 20644 23919 20700
rect 23919 20644 23975 20700
rect 23975 20644 23979 20700
rect 23915 20640 23979 20644
rect 3792 20156 3856 20160
rect 3792 20100 3796 20156
rect 3796 20100 3852 20156
rect 3852 20100 3856 20156
rect 3792 20096 3856 20100
rect 3872 20156 3936 20160
rect 3872 20100 3876 20156
rect 3876 20100 3932 20156
rect 3932 20100 3936 20156
rect 3872 20096 3936 20100
rect 3952 20156 4016 20160
rect 3952 20100 3956 20156
rect 3956 20100 4012 20156
rect 4012 20100 4016 20156
rect 3952 20096 4016 20100
rect 4032 20156 4096 20160
rect 4032 20100 4036 20156
rect 4036 20100 4092 20156
rect 4092 20100 4096 20156
rect 4032 20096 4096 20100
rect 9473 20156 9537 20160
rect 9473 20100 9477 20156
rect 9477 20100 9533 20156
rect 9533 20100 9537 20156
rect 9473 20096 9537 20100
rect 9553 20156 9617 20160
rect 9553 20100 9557 20156
rect 9557 20100 9613 20156
rect 9613 20100 9617 20156
rect 9553 20096 9617 20100
rect 9633 20156 9697 20160
rect 9633 20100 9637 20156
rect 9637 20100 9693 20156
rect 9693 20100 9697 20156
rect 9633 20096 9697 20100
rect 9713 20156 9777 20160
rect 9713 20100 9717 20156
rect 9717 20100 9773 20156
rect 9773 20100 9777 20156
rect 9713 20096 9777 20100
rect 15154 20156 15218 20160
rect 15154 20100 15158 20156
rect 15158 20100 15214 20156
rect 15214 20100 15218 20156
rect 15154 20096 15218 20100
rect 15234 20156 15298 20160
rect 15234 20100 15238 20156
rect 15238 20100 15294 20156
rect 15294 20100 15298 20156
rect 15234 20096 15298 20100
rect 15314 20156 15378 20160
rect 15314 20100 15318 20156
rect 15318 20100 15374 20156
rect 15374 20100 15378 20156
rect 15314 20096 15378 20100
rect 15394 20156 15458 20160
rect 15394 20100 15398 20156
rect 15398 20100 15454 20156
rect 15454 20100 15458 20156
rect 15394 20096 15458 20100
rect 20835 20156 20899 20160
rect 20835 20100 20839 20156
rect 20839 20100 20895 20156
rect 20895 20100 20899 20156
rect 20835 20096 20899 20100
rect 20915 20156 20979 20160
rect 20915 20100 20919 20156
rect 20919 20100 20975 20156
rect 20975 20100 20979 20156
rect 20915 20096 20979 20100
rect 20995 20156 21059 20160
rect 20995 20100 20999 20156
rect 20999 20100 21055 20156
rect 21055 20100 21059 20156
rect 20995 20096 21059 20100
rect 21075 20156 21139 20160
rect 21075 20100 21079 20156
rect 21079 20100 21135 20156
rect 21135 20100 21139 20156
rect 21075 20096 21139 20100
rect 6632 19612 6696 19616
rect 6632 19556 6636 19612
rect 6636 19556 6692 19612
rect 6692 19556 6696 19612
rect 6632 19552 6696 19556
rect 6712 19612 6776 19616
rect 6712 19556 6716 19612
rect 6716 19556 6772 19612
rect 6772 19556 6776 19612
rect 6712 19552 6776 19556
rect 6792 19612 6856 19616
rect 6792 19556 6796 19612
rect 6796 19556 6852 19612
rect 6852 19556 6856 19612
rect 6792 19552 6856 19556
rect 6872 19612 6936 19616
rect 6872 19556 6876 19612
rect 6876 19556 6932 19612
rect 6932 19556 6936 19612
rect 6872 19552 6936 19556
rect 12313 19612 12377 19616
rect 12313 19556 12317 19612
rect 12317 19556 12373 19612
rect 12373 19556 12377 19612
rect 12313 19552 12377 19556
rect 12393 19612 12457 19616
rect 12393 19556 12397 19612
rect 12397 19556 12453 19612
rect 12453 19556 12457 19612
rect 12393 19552 12457 19556
rect 12473 19612 12537 19616
rect 12473 19556 12477 19612
rect 12477 19556 12533 19612
rect 12533 19556 12537 19612
rect 12473 19552 12537 19556
rect 12553 19612 12617 19616
rect 12553 19556 12557 19612
rect 12557 19556 12613 19612
rect 12613 19556 12617 19612
rect 12553 19552 12617 19556
rect 17994 19612 18058 19616
rect 17994 19556 17998 19612
rect 17998 19556 18054 19612
rect 18054 19556 18058 19612
rect 17994 19552 18058 19556
rect 18074 19612 18138 19616
rect 18074 19556 18078 19612
rect 18078 19556 18134 19612
rect 18134 19556 18138 19612
rect 18074 19552 18138 19556
rect 18154 19612 18218 19616
rect 18154 19556 18158 19612
rect 18158 19556 18214 19612
rect 18214 19556 18218 19612
rect 18154 19552 18218 19556
rect 18234 19612 18298 19616
rect 18234 19556 18238 19612
rect 18238 19556 18294 19612
rect 18294 19556 18298 19612
rect 18234 19552 18298 19556
rect 23675 19612 23739 19616
rect 23675 19556 23679 19612
rect 23679 19556 23735 19612
rect 23735 19556 23739 19612
rect 23675 19552 23739 19556
rect 23755 19612 23819 19616
rect 23755 19556 23759 19612
rect 23759 19556 23815 19612
rect 23815 19556 23819 19612
rect 23755 19552 23819 19556
rect 23835 19612 23899 19616
rect 23835 19556 23839 19612
rect 23839 19556 23895 19612
rect 23895 19556 23899 19612
rect 23835 19552 23899 19556
rect 23915 19612 23979 19616
rect 23915 19556 23919 19612
rect 23919 19556 23975 19612
rect 23975 19556 23979 19612
rect 23915 19552 23979 19556
rect 17724 19348 17788 19412
rect 3792 19068 3856 19072
rect 3792 19012 3796 19068
rect 3796 19012 3852 19068
rect 3852 19012 3856 19068
rect 3792 19008 3856 19012
rect 3872 19068 3936 19072
rect 3872 19012 3876 19068
rect 3876 19012 3932 19068
rect 3932 19012 3936 19068
rect 3872 19008 3936 19012
rect 3952 19068 4016 19072
rect 3952 19012 3956 19068
rect 3956 19012 4012 19068
rect 4012 19012 4016 19068
rect 3952 19008 4016 19012
rect 4032 19068 4096 19072
rect 4032 19012 4036 19068
rect 4036 19012 4092 19068
rect 4092 19012 4096 19068
rect 4032 19008 4096 19012
rect 9473 19068 9537 19072
rect 9473 19012 9477 19068
rect 9477 19012 9533 19068
rect 9533 19012 9537 19068
rect 9473 19008 9537 19012
rect 9553 19068 9617 19072
rect 9553 19012 9557 19068
rect 9557 19012 9613 19068
rect 9613 19012 9617 19068
rect 9553 19008 9617 19012
rect 9633 19068 9697 19072
rect 9633 19012 9637 19068
rect 9637 19012 9693 19068
rect 9693 19012 9697 19068
rect 9633 19008 9697 19012
rect 9713 19068 9777 19072
rect 9713 19012 9717 19068
rect 9717 19012 9773 19068
rect 9773 19012 9777 19068
rect 9713 19008 9777 19012
rect 15154 19068 15218 19072
rect 15154 19012 15158 19068
rect 15158 19012 15214 19068
rect 15214 19012 15218 19068
rect 15154 19008 15218 19012
rect 15234 19068 15298 19072
rect 15234 19012 15238 19068
rect 15238 19012 15294 19068
rect 15294 19012 15298 19068
rect 15234 19008 15298 19012
rect 15314 19068 15378 19072
rect 15314 19012 15318 19068
rect 15318 19012 15374 19068
rect 15374 19012 15378 19068
rect 15314 19008 15378 19012
rect 15394 19068 15458 19072
rect 15394 19012 15398 19068
rect 15398 19012 15454 19068
rect 15454 19012 15458 19068
rect 15394 19008 15458 19012
rect 20835 19068 20899 19072
rect 20835 19012 20839 19068
rect 20839 19012 20895 19068
rect 20895 19012 20899 19068
rect 20835 19008 20899 19012
rect 20915 19068 20979 19072
rect 20915 19012 20919 19068
rect 20919 19012 20975 19068
rect 20975 19012 20979 19068
rect 20915 19008 20979 19012
rect 20995 19068 21059 19072
rect 20995 19012 20999 19068
rect 20999 19012 21055 19068
rect 21055 19012 21059 19068
rect 20995 19008 21059 19012
rect 21075 19068 21139 19072
rect 21075 19012 21079 19068
rect 21079 19012 21135 19068
rect 21135 19012 21139 19068
rect 21075 19008 21139 19012
rect 6632 18524 6696 18528
rect 6632 18468 6636 18524
rect 6636 18468 6692 18524
rect 6692 18468 6696 18524
rect 6632 18464 6696 18468
rect 6712 18524 6776 18528
rect 6712 18468 6716 18524
rect 6716 18468 6772 18524
rect 6772 18468 6776 18524
rect 6712 18464 6776 18468
rect 6792 18524 6856 18528
rect 6792 18468 6796 18524
rect 6796 18468 6852 18524
rect 6852 18468 6856 18524
rect 6792 18464 6856 18468
rect 6872 18524 6936 18528
rect 6872 18468 6876 18524
rect 6876 18468 6932 18524
rect 6932 18468 6936 18524
rect 6872 18464 6936 18468
rect 12313 18524 12377 18528
rect 12313 18468 12317 18524
rect 12317 18468 12373 18524
rect 12373 18468 12377 18524
rect 12313 18464 12377 18468
rect 12393 18524 12457 18528
rect 12393 18468 12397 18524
rect 12397 18468 12453 18524
rect 12453 18468 12457 18524
rect 12393 18464 12457 18468
rect 12473 18524 12537 18528
rect 12473 18468 12477 18524
rect 12477 18468 12533 18524
rect 12533 18468 12537 18524
rect 12473 18464 12537 18468
rect 12553 18524 12617 18528
rect 12553 18468 12557 18524
rect 12557 18468 12613 18524
rect 12613 18468 12617 18524
rect 12553 18464 12617 18468
rect 17994 18524 18058 18528
rect 17994 18468 17998 18524
rect 17998 18468 18054 18524
rect 18054 18468 18058 18524
rect 17994 18464 18058 18468
rect 18074 18524 18138 18528
rect 18074 18468 18078 18524
rect 18078 18468 18134 18524
rect 18134 18468 18138 18524
rect 18074 18464 18138 18468
rect 18154 18524 18218 18528
rect 18154 18468 18158 18524
rect 18158 18468 18214 18524
rect 18214 18468 18218 18524
rect 18154 18464 18218 18468
rect 18234 18524 18298 18528
rect 18234 18468 18238 18524
rect 18238 18468 18294 18524
rect 18294 18468 18298 18524
rect 18234 18464 18298 18468
rect 23675 18524 23739 18528
rect 23675 18468 23679 18524
rect 23679 18468 23735 18524
rect 23735 18468 23739 18524
rect 23675 18464 23739 18468
rect 23755 18524 23819 18528
rect 23755 18468 23759 18524
rect 23759 18468 23815 18524
rect 23815 18468 23819 18524
rect 23755 18464 23819 18468
rect 23835 18524 23899 18528
rect 23835 18468 23839 18524
rect 23839 18468 23895 18524
rect 23895 18468 23899 18524
rect 23835 18464 23899 18468
rect 23915 18524 23979 18528
rect 23915 18468 23919 18524
rect 23919 18468 23975 18524
rect 23975 18468 23979 18524
rect 23915 18464 23979 18468
rect 21404 18124 21468 18188
rect 16436 17988 16500 18052
rect 3792 17980 3856 17984
rect 3792 17924 3796 17980
rect 3796 17924 3852 17980
rect 3852 17924 3856 17980
rect 3792 17920 3856 17924
rect 3872 17980 3936 17984
rect 3872 17924 3876 17980
rect 3876 17924 3932 17980
rect 3932 17924 3936 17980
rect 3872 17920 3936 17924
rect 3952 17980 4016 17984
rect 3952 17924 3956 17980
rect 3956 17924 4012 17980
rect 4012 17924 4016 17980
rect 3952 17920 4016 17924
rect 4032 17980 4096 17984
rect 4032 17924 4036 17980
rect 4036 17924 4092 17980
rect 4092 17924 4096 17980
rect 4032 17920 4096 17924
rect 9473 17980 9537 17984
rect 9473 17924 9477 17980
rect 9477 17924 9533 17980
rect 9533 17924 9537 17980
rect 9473 17920 9537 17924
rect 9553 17980 9617 17984
rect 9553 17924 9557 17980
rect 9557 17924 9613 17980
rect 9613 17924 9617 17980
rect 9553 17920 9617 17924
rect 9633 17980 9697 17984
rect 9633 17924 9637 17980
rect 9637 17924 9693 17980
rect 9693 17924 9697 17980
rect 9633 17920 9697 17924
rect 9713 17980 9777 17984
rect 9713 17924 9717 17980
rect 9717 17924 9773 17980
rect 9773 17924 9777 17980
rect 9713 17920 9777 17924
rect 15154 17980 15218 17984
rect 15154 17924 15158 17980
rect 15158 17924 15214 17980
rect 15214 17924 15218 17980
rect 15154 17920 15218 17924
rect 15234 17980 15298 17984
rect 15234 17924 15238 17980
rect 15238 17924 15294 17980
rect 15294 17924 15298 17980
rect 15234 17920 15298 17924
rect 15314 17980 15378 17984
rect 15314 17924 15318 17980
rect 15318 17924 15374 17980
rect 15374 17924 15378 17980
rect 15314 17920 15378 17924
rect 15394 17980 15458 17984
rect 15394 17924 15398 17980
rect 15398 17924 15454 17980
rect 15454 17924 15458 17980
rect 15394 17920 15458 17924
rect 20835 17980 20899 17984
rect 20835 17924 20839 17980
rect 20839 17924 20895 17980
rect 20895 17924 20899 17980
rect 20835 17920 20899 17924
rect 20915 17980 20979 17984
rect 20915 17924 20919 17980
rect 20919 17924 20975 17980
rect 20975 17924 20979 17980
rect 20915 17920 20979 17924
rect 20995 17980 21059 17984
rect 20995 17924 20999 17980
rect 20999 17924 21055 17980
rect 21055 17924 21059 17980
rect 20995 17920 21059 17924
rect 21075 17980 21139 17984
rect 21075 17924 21079 17980
rect 21079 17924 21135 17980
rect 21135 17924 21139 17980
rect 21075 17920 21139 17924
rect 6632 17436 6696 17440
rect 6632 17380 6636 17436
rect 6636 17380 6692 17436
rect 6692 17380 6696 17436
rect 6632 17376 6696 17380
rect 6712 17436 6776 17440
rect 6712 17380 6716 17436
rect 6716 17380 6772 17436
rect 6772 17380 6776 17436
rect 6712 17376 6776 17380
rect 6792 17436 6856 17440
rect 6792 17380 6796 17436
rect 6796 17380 6852 17436
rect 6852 17380 6856 17436
rect 6792 17376 6856 17380
rect 6872 17436 6936 17440
rect 6872 17380 6876 17436
rect 6876 17380 6932 17436
rect 6932 17380 6936 17436
rect 6872 17376 6936 17380
rect 12313 17436 12377 17440
rect 12313 17380 12317 17436
rect 12317 17380 12373 17436
rect 12373 17380 12377 17436
rect 12313 17376 12377 17380
rect 12393 17436 12457 17440
rect 12393 17380 12397 17436
rect 12397 17380 12453 17436
rect 12453 17380 12457 17436
rect 12393 17376 12457 17380
rect 12473 17436 12537 17440
rect 12473 17380 12477 17436
rect 12477 17380 12533 17436
rect 12533 17380 12537 17436
rect 12473 17376 12537 17380
rect 12553 17436 12617 17440
rect 12553 17380 12557 17436
rect 12557 17380 12613 17436
rect 12613 17380 12617 17436
rect 12553 17376 12617 17380
rect 17994 17436 18058 17440
rect 17994 17380 17998 17436
rect 17998 17380 18054 17436
rect 18054 17380 18058 17436
rect 17994 17376 18058 17380
rect 18074 17436 18138 17440
rect 18074 17380 18078 17436
rect 18078 17380 18134 17436
rect 18134 17380 18138 17436
rect 18074 17376 18138 17380
rect 18154 17436 18218 17440
rect 18154 17380 18158 17436
rect 18158 17380 18214 17436
rect 18214 17380 18218 17436
rect 18154 17376 18218 17380
rect 18234 17436 18298 17440
rect 18234 17380 18238 17436
rect 18238 17380 18294 17436
rect 18294 17380 18298 17436
rect 18234 17376 18298 17380
rect 23675 17436 23739 17440
rect 23675 17380 23679 17436
rect 23679 17380 23735 17436
rect 23735 17380 23739 17436
rect 23675 17376 23739 17380
rect 23755 17436 23819 17440
rect 23755 17380 23759 17436
rect 23759 17380 23815 17436
rect 23815 17380 23819 17436
rect 23755 17376 23819 17380
rect 23835 17436 23899 17440
rect 23835 17380 23839 17436
rect 23839 17380 23895 17436
rect 23895 17380 23899 17436
rect 23835 17376 23899 17380
rect 23915 17436 23979 17440
rect 23915 17380 23919 17436
rect 23919 17380 23975 17436
rect 23975 17380 23979 17436
rect 23915 17376 23979 17380
rect 3792 16892 3856 16896
rect 3792 16836 3796 16892
rect 3796 16836 3852 16892
rect 3852 16836 3856 16892
rect 3792 16832 3856 16836
rect 3872 16892 3936 16896
rect 3872 16836 3876 16892
rect 3876 16836 3932 16892
rect 3932 16836 3936 16892
rect 3872 16832 3936 16836
rect 3952 16892 4016 16896
rect 3952 16836 3956 16892
rect 3956 16836 4012 16892
rect 4012 16836 4016 16892
rect 3952 16832 4016 16836
rect 4032 16892 4096 16896
rect 4032 16836 4036 16892
rect 4036 16836 4092 16892
rect 4092 16836 4096 16892
rect 4032 16832 4096 16836
rect 9473 16892 9537 16896
rect 9473 16836 9477 16892
rect 9477 16836 9533 16892
rect 9533 16836 9537 16892
rect 9473 16832 9537 16836
rect 9553 16892 9617 16896
rect 9553 16836 9557 16892
rect 9557 16836 9613 16892
rect 9613 16836 9617 16892
rect 9553 16832 9617 16836
rect 9633 16892 9697 16896
rect 9633 16836 9637 16892
rect 9637 16836 9693 16892
rect 9693 16836 9697 16892
rect 9633 16832 9697 16836
rect 9713 16892 9777 16896
rect 9713 16836 9717 16892
rect 9717 16836 9773 16892
rect 9773 16836 9777 16892
rect 9713 16832 9777 16836
rect 15154 16892 15218 16896
rect 15154 16836 15158 16892
rect 15158 16836 15214 16892
rect 15214 16836 15218 16892
rect 15154 16832 15218 16836
rect 15234 16892 15298 16896
rect 15234 16836 15238 16892
rect 15238 16836 15294 16892
rect 15294 16836 15298 16892
rect 15234 16832 15298 16836
rect 15314 16892 15378 16896
rect 15314 16836 15318 16892
rect 15318 16836 15374 16892
rect 15374 16836 15378 16892
rect 15314 16832 15378 16836
rect 15394 16892 15458 16896
rect 15394 16836 15398 16892
rect 15398 16836 15454 16892
rect 15454 16836 15458 16892
rect 15394 16832 15458 16836
rect 20835 16892 20899 16896
rect 20835 16836 20839 16892
rect 20839 16836 20895 16892
rect 20895 16836 20899 16892
rect 20835 16832 20899 16836
rect 20915 16892 20979 16896
rect 20915 16836 20919 16892
rect 20919 16836 20975 16892
rect 20975 16836 20979 16892
rect 20915 16832 20979 16836
rect 20995 16892 21059 16896
rect 20995 16836 20999 16892
rect 20999 16836 21055 16892
rect 21055 16836 21059 16892
rect 20995 16832 21059 16836
rect 21075 16892 21139 16896
rect 21075 16836 21079 16892
rect 21079 16836 21135 16892
rect 21135 16836 21139 16892
rect 21075 16832 21139 16836
rect 6632 16348 6696 16352
rect 6632 16292 6636 16348
rect 6636 16292 6692 16348
rect 6692 16292 6696 16348
rect 6632 16288 6696 16292
rect 6712 16348 6776 16352
rect 6712 16292 6716 16348
rect 6716 16292 6772 16348
rect 6772 16292 6776 16348
rect 6712 16288 6776 16292
rect 6792 16348 6856 16352
rect 6792 16292 6796 16348
rect 6796 16292 6852 16348
rect 6852 16292 6856 16348
rect 6792 16288 6856 16292
rect 6872 16348 6936 16352
rect 6872 16292 6876 16348
rect 6876 16292 6932 16348
rect 6932 16292 6936 16348
rect 6872 16288 6936 16292
rect 12313 16348 12377 16352
rect 12313 16292 12317 16348
rect 12317 16292 12373 16348
rect 12373 16292 12377 16348
rect 12313 16288 12377 16292
rect 12393 16348 12457 16352
rect 12393 16292 12397 16348
rect 12397 16292 12453 16348
rect 12453 16292 12457 16348
rect 12393 16288 12457 16292
rect 12473 16348 12537 16352
rect 12473 16292 12477 16348
rect 12477 16292 12533 16348
rect 12533 16292 12537 16348
rect 12473 16288 12537 16292
rect 12553 16348 12617 16352
rect 12553 16292 12557 16348
rect 12557 16292 12613 16348
rect 12613 16292 12617 16348
rect 12553 16288 12617 16292
rect 17994 16348 18058 16352
rect 17994 16292 17998 16348
rect 17998 16292 18054 16348
rect 18054 16292 18058 16348
rect 17994 16288 18058 16292
rect 18074 16348 18138 16352
rect 18074 16292 18078 16348
rect 18078 16292 18134 16348
rect 18134 16292 18138 16348
rect 18074 16288 18138 16292
rect 18154 16348 18218 16352
rect 18154 16292 18158 16348
rect 18158 16292 18214 16348
rect 18214 16292 18218 16348
rect 18154 16288 18218 16292
rect 18234 16348 18298 16352
rect 18234 16292 18238 16348
rect 18238 16292 18294 16348
rect 18294 16292 18298 16348
rect 18234 16288 18298 16292
rect 23675 16348 23739 16352
rect 23675 16292 23679 16348
rect 23679 16292 23735 16348
rect 23735 16292 23739 16348
rect 23675 16288 23739 16292
rect 23755 16348 23819 16352
rect 23755 16292 23759 16348
rect 23759 16292 23815 16348
rect 23815 16292 23819 16348
rect 23755 16288 23819 16292
rect 23835 16348 23899 16352
rect 23835 16292 23839 16348
rect 23839 16292 23895 16348
rect 23895 16292 23899 16348
rect 23835 16288 23899 16292
rect 23915 16348 23979 16352
rect 23915 16292 23919 16348
rect 23919 16292 23975 16348
rect 23975 16292 23979 16348
rect 23915 16288 23979 16292
rect 3792 15804 3856 15808
rect 3792 15748 3796 15804
rect 3796 15748 3852 15804
rect 3852 15748 3856 15804
rect 3792 15744 3856 15748
rect 3872 15804 3936 15808
rect 3872 15748 3876 15804
rect 3876 15748 3932 15804
rect 3932 15748 3936 15804
rect 3872 15744 3936 15748
rect 3952 15804 4016 15808
rect 3952 15748 3956 15804
rect 3956 15748 4012 15804
rect 4012 15748 4016 15804
rect 3952 15744 4016 15748
rect 4032 15804 4096 15808
rect 4032 15748 4036 15804
rect 4036 15748 4092 15804
rect 4092 15748 4096 15804
rect 4032 15744 4096 15748
rect 9473 15804 9537 15808
rect 9473 15748 9477 15804
rect 9477 15748 9533 15804
rect 9533 15748 9537 15804
rect 9473 15744 9537 15748
rect 9553 15804 9617 15808
rect 9553 15748 9557 15804
rect 9557 15748 9613 15804
rect 9613 15748 9617 15804
rect 9553 15744 9617 15748
rect 9633 15804 9697 15808
rect 9633 15748 9637 15804
rect 9637 15748 9693 15804
rect 9693 15748 9697 15804
rect 9633 15744 9697 15748
rect 9713 15804 9777 15808
rect 9713 15748 9717 15804
rect 9717 15748 9773 15804
rect 9773 15748 9777 15804
rect 9713 15744 9777 15748
rect 15154 15804 15218 15808
rect 15154 15748 15158 15804
rect 15158 15748 15214 15804
rect 15214 15748 15218 15804
rect 15154 15744 15218 15748
rect 15234 15804 15298 15808
rect 15234 15748 15238 15804
rect 15238 15748 15294 15804
rect 15294 15748 15298 15804
rect 15234 15744 15298 15748
rect 15314 15804 15378 15808
rect 15314 15748 15318 15804
rect 15318 15748 15374 15804
rect 15374 15748 15378 15804
rect 15314 15744 15378 15748
rect 15394 15804 15458 15808
rect 15394 15748 15398 15804
rect 15398 15748 15454 15804
rect 15454 15748 15458 15804
rect 15394 15744 15458 15748
rect 20835 15804 20899 15808
rect 20835 15748 20839 15804
rect 20839 15748 20895 15804
rect 20895 15748 20899 15804
rect 20835 15744 20899 15748
rect 20915 15804 20979 15808
rect 20915 15748 20919 15804
rect 20919 15748 20975 15804
rect 20975 15748 20979 15804
rect 20915 15744 20979 15748
rect 20995 15804 21059 15808
rect 20995 15748 20999 15804
rect 20999 15748 21055 15804
rect 21055 15748 21059 15804
rect 20995 15744 21059 15748
rect 21075 15804 21139 15808
rect 21075 15748 21079 15804
rect 21079 15748 21135 15804
rect 21135 15748 21139 15804
rect 21075 15744 21139 15748
rect 5396 15268 5460 15332
rect 6632 15260 6696 15264
rect 6632 15204 6636 15260
rect 6636 15204 6692 15260
rect 6692 15204 6696 15260
rect 6632 15200 6696 15204
rect 6712 15260 6776 15264
rect 6712 15204 6716 15260
rect 6716 15204 6772 15260
rect 6772 15204 6776 15260
rect 6712 15200 6776 15204
rect 6792 15260 6856 15264
rect 6792 15204 6796 15260
rect 6796 15204 6852 15260
rect 6852 15204 6856 15260
rect 6792 15200 6856 15204
rect 6872 15260 6936 15264
rect 6872 15204 6876 15260
rect 6876 15204 6932 15260
rect 6932 15204 6936 15260
rect 6872 15200 6936 15204
rect 12313 15260 12377 15264
rect 12313 15204 12317 15260
rect 12317 15204 12373 15260
rect 12373 15204 12377 15260
rect 12313 15200 12377 15204
rect 12393 15260 12457 15264
rect 12393 15204 12397 15260
rect 12397 15204 12453 15260
rect 12453 15204 12457 15260
rect 12393 15200 12457 15204
rect 12473 15260 12537 15264
rect 12473 15204 12477 15260
rect 12477 15204 12533 15260
rect 12533 15204 12537 15260
rect 12473 15200 12537 15204
rect 12553 15260 12617 15264
rect 12553 15204 12557 15260
rect 12557 15204 12613 15260
rect 12613 15204 12617 15260
rect 12553 15200 12617 15204
rect 17994 15260 18058 15264
rect 17994 15204 17998 15260
rect 17998 15204 18054 15260
rect 18054 15204 18058 15260
rect 17994 15200 18058 15204
rect 18074 15260 18138 15264
rect 18074 15204 18078 15260
rect 18078 15204 18134 15260
rect 18134 15204 18138 15260
rect 18074 15200 18138 15204
rect 18154 15260 18218 15264
rect 18154 15204 18158 15260
rect 18158 15204 18214 15260
rect 18214 15204 18218 15260
rect 18154 15200 18218 15204
rect 18234 15260 18298 15264
rect 18234 15204 18238 15260
rect 18238 15204 18294 15260
rect 18294 15204 18298 15260
rect 18234 15200 18298 15204
rect 23675 15260 23739 15264
rect 23675 15204 23679 15260
rect 23679 15204 23735 15260
rect 23735 15204 23739 15260
rect 23675 15200 23739 15204
rect 23755 15260 23819 15264
rect 23755 15204 23759 15260
rect 23759 15204 23815 15260
rect 23815 15204 23819 15260
rect 23755 15200 23819 15204
rect 23835 15260 23899 15264
rect 23835 15204 23839 15260
rect 23839 15204 23895 15260
rect 23895 15204 23899 15260
rect 23835 15200 23899 15204
rect 23915 15260 23979 15264
rect 23915 15204 23919 15260
rect 23919 15204 23975 15260
rect 23975 15204 23979 15260
rect 23915 15200 23979 15204
rect 3792 14716 3856 14720
rect 3792 14660 3796 14716
rect 3796 14660 3852 14716
rect 3852 14660 3856 14716
rect 3792 14656 3856 14660
rect 3872 14716 3936 14720
rect 3872 14660 3876 14716
rect 3876 14660 3932 14716
rect 3932 14660 3936 14716
rect 3872 14656 3936 14660
rect 3952 14716 4016 14720
rect 3952 14660 3956 14716
rect 3956 14660 4012 14716
rect 4012 14660 4016 14716
rect 3952 14656 4016 14660
rect 4032 14716 4096 14720
rect 4032 14660 4036 14716
rect 4036 14660 4092 14716
rect 4092 14660 4096 14716
rect 4032 14656 4096 14660
rect 9473 14716 9537 14720
rect 9473 14660 9477 14716
rect 9477 14660 9533 14716
rect 9533 14660 9537 14716
rect 9473 14656 9537 14660
rect 9553 14716 9617 14720
rect 9553 14660 9557 14716
rect 9557 14660 9613 14716
rect 9613 14660 9617 14716
rect 9553 14656 9617 14660
rect 9633 14716 9697 14720
rect 9633 14660 9637 14716
rect 9637 14660 9693 14716
rect 9693 14660 9697 14716
rect 9633 14656 9697 14660
rect 9713 14716 9777 14720
rect 9713 14660 9717 14716
rect 9717 14660 9773 14716
rect 9773 14660 9777 14716
rect 9713 14656 9777 14660
rect 15154 14716 15218 14720
rect 15154 14660 15158 14716
rect 15158 14660 15214 14716
rect 15214 14660 15218 14716
rect 15154 14656 15218 14660
rect 15234 14716 15298 14720
rect 15234 14660 15238 14716
rect 15238 14660 15294 14716
rect 15294 14660 15298 14716
rect 15234 14656 15298 14660
rect 15314 14716 15378 14720
rect 15314 14660 15318 14716
rect 15318 14660 15374 14716
rect 15374 14660 15378 14716
rect 15314 14656 15378 14660
rect 15394 14716 15458 14720
rect 15394 14660 15398 14716
rect 15398 14660 15454 14716
rect 15454 14660 15458 14716
rect 15394 14656 15458 14660
rect 20835 14716 20899 14720
rect 20835 14660 20839 14716
rect 20839 14660 20895 14716
rect 20895 14660 20899 14716
rect 20835 14656 20899 14660
rect 20915 14716 20979 14720
rect 20915 14660 20919 14716
rect 20919 14660 20975 14716
rect 20975 14660 20979 14716
rect 20915 14656 20979 14660
rect 20995 14716 21059 14720
rect 20995 14660 20999 14716
rect 20999 14660 21055 14716
rect 21055 14660 21059 14716
rect 20995 14656 21059 14660
rect 21075 14716 21139 14720
rect 21075 14660 21079 14716
rect 21079 14660 21135 14716
rect 21135 14660 21139 14716
rect 21075 14656 21139 14660
rect 16436 14588 16500 14652
rect 6632 14172 6696 14176
rect 6632 14116 6636 14172
rect 6636 14116 6692 14172
rect 6692 14116 6696 14172
rect 6632 14112 6696 14116
rect 6712 14172 6776 14176
rect 6712 14116 6716 14172
rect 6716 14116 6772 14172
rect 6772 14116 6776 14172
rect 6712 14112 6776 14116
rect 6792 14172 6856 14176
rect 6792 14116 6796 14172
rect 6796 14116 6852 14172
rect 6852 14116 6856 14172
rect 6792 14112 6856 14116
rect 6872 14172 6936 14176
rect 6872 14116 6876 14172
rect 6876 14116 6932 14172
rect 6932 14116 6936 14172
rect 6872 14112 6936 14116
rect 12313 14172 12377 14176
rect 12313 14116 12317 14172
rect 12317 14116 12373 14172
rect 12373 14116 12377 14172
rect 12313 14112 12377 14116
rect 12393 14172 12457 14176
rect 12393 14116 12397 14172
rect 12397 14116 12453 14172
rect 12453 14116 12457 14172
rect 12393 14112 12457 14116
rect 12473 14172 12537 14176
rect 12473 14116 12477 14172
rect 12477 14116 12533 14172
rect 12533 14116 12537 14172
rect 12473 14112 12537 14116
rect 12553 14172 12617 14176
rect 12553 14116 12557 14172
rect 12557 14116 12613 14172
rect 12613 14116 12617 14172
rect 12553 14112 12617 14116
rect 17994 14172 18058 14176
rect 17994 14116 17998 14172
rect 17998 14116 18054 14172
rect 18054 14116 18058 14172
rect 17994 14112 18058 14116
rect 18074 14172 18138 14176
rect 18074 14116 18078 14172
rect 18078 14116 18134 14172
rect 18134 14116 18138 14172
rect 18074 14112 18138 14116
rect 18154 14172 18218 14176
rect 18154 14116 18158 14172
rect 18158 14116 18214 14172
rect 18214 14116 18218 14172
rect 18154 14112 18218 14116
rect 18234 14172 18298 14176
rect 18234 14116 18238 14172
rect 18238 14116 18294 14172
rect 18294 14116 18298 14172
rect 18234 14112 18298 14116
rect 23675 14172 23739 14176
rect 23675 14116 23679 14172
rect 23679 14116 23735 14172
rect 23735 14116 23739 14172
rect 23675 14112 23739 14116
rect 23755 14172 23819 14176
rect 23755 14116 23759 14172
rect 23759 14116 23815 14172
rect 23815 14116 23819 14172
rect 23755 14112 23819 14116
rect 23835 14172 23899 14176
rect 23835 14116 23839 14172
rect 23839 14116 23895 14172
rect 23895 14116 23899 14172
rect 23835 14112 23899 14116
rect 23915 14172 23979 14176
rect 23915 14116 23919 14172
rect 23919 14116 23975 14172
rect 23975 14116 23979 14172
rect 23915 14112 23979 14116
rect 16252 13772 16316 13836
rect 3792 13628 3856 13632
rect 3792 13572 3796 13628
rect 3796 13572 3852 13628
rect 3852 13572 3856 13628
rect 3792 13568 3856 13572
rect 3872 13628 3936 13632
rect 3872 13572 3876 13628
rect 3876 13572 3932 13628
rect 3932 13572 3936 13628
rect 3872 13568 3936 13572
rect 3952 13628 4016 13632
rect 3952 13572 3956 13628
rect 3956 13572 4012 13628
rect 4012 13572 4016 13628
rect 3952 13568 4016 13572
rect 4032 13628 4096 13632
rect 4032 13572 4036 13628
rect 4036 13572 4092 13628
rect 4092 13572 4096 13628
rect 4032 13568 4096 13572
rect 9473 13628 9537 13632
rect 9473 13572 9477 13628
rect 9477 13572 9533 13628
rect 9533 13572 9537 13628
rect 9473 13568 9537 13572
rect 9553 13628 9617 13632
rect 9553 13572 9557 13628
rect 9557 13572 9613 13628
rect 9613 13572 9617 13628
rect 9553 13568 9617 13572
rect 9633 13628 9697 13632
rect 9633 13572 9637 13628
rect 9637 13572 9693 13628
rect 9693 13572 9697 13628
rect 9633 13568 9697 13572
rect 9713 13628 9777 13632
rect 9713 13572 9717 13628
rect 9717 13572 9773 13628
rect 9773 13572 9777 13628
rect 9713 13568 9777 13572
rect 15154 13628 15218 13632
rect 15154 13572 15158 13628
rect 15158 13572 15214 13628
rect 15214 13572 15218 13628
rect 15154 13568 15218 13572
rect 15234 13628 15298 13632
rect 15234 13572 15238 13628
rect 15238 13572 15294 13628
rect 15294 13572 15298 13628
rect 15234 13568 15298 13572
rect 15314 13628 15378 13632
rect 15314 13572 15318 13628
rect 15318 13572 15374 13628
rect 15374 13572 15378 13628
rect 15314 13568 15378 13572
rect 15394 13628 15458 13632
rect 15394 13572 15398 13628
rect 15398 13572 15454 13628
rect 15454 13572 15458 13628
rect 15394 13568 15458 13572
rect 22324 13772 22388 13836
rect 20835 13628 20899 13632
rect 20835 13572 20839 13628
rect 20839 13572 20895 13628
rect 20895 13572 20899 13628
rect 20835 13568 20899 13572
rect 20915 13628 20979 13632
rect 20915 13572 20919 13628
rect 20919 13572 20975 13628
rect 20975 13572 20979 13628
rect 20915 13568 20979 13572
rect 20995 13628 21059 13632
rect 20995 13572 20999 13628
rect 20999 13572 21055 13628
rect 21055 13572 21059 13628
rect 20995 13568 21059 13572
rect 21075 13628 21139 13632
rect 21075 13572 21079 13628
rect 21079 13572 21135 13628
rect 21135 13572 21139 13628
rect 21075 13568 21139 13572
rect 17724 13500 17788 13564
rect 6632 13084 6696 13088
rect 6632 13028 6636 13084
rect 6636 13028 6692 13084
rect 6692 13028 6696 13084
rect 6632 13024 6696 13028
rect 6712 13084 6776 13088
rect 6712 13028 6716 13084
rect 6716 13028 6772 13084
rect 6772 13028 6776 13084
rect 6712 13024 6776 13028
rect 6792 13084 6856 13088
rect 6792 13028 6796 13084
rect 6796 13028 6852 13084
rect 6852 13028 6856 13084
rect 6792 13024 6856 13028
rect 6872 13084 6936 13088
rect 6872 13028 6876 13084
rect 6876 13028 6932 13084
rect 6932 13028 6936 13084
rect 6872 13024 6936 13028
rect 12313 13084 12377 13088
rect 12313 13028 12317 13084
rect 12317 13028 12373 13084
rect 12373 13028 12377 13084
rect 12313 13024 12377 13028
rect 12393 13084 12457 13088
rect 12393 13028 12397 13084
rect 12397 13028 12453 13084
rect 12453 13028 12457 13084
rect 12393 13024 12457 13028
rect 12473 13084 12537 13088
rect 12473 13028 12477 13084
rect 12477 13028 12533 13084
rect 12533 13028 12537 13084
rect 12473 13024 12537 13028
rect 12553 13084 12617 13088
rect 12553 13028 12557 13084
rect 12557 13028 12613 13084
rect 12613 13028 12617 13084
rect 12553 13024 12617 13028
rect 17994 13084 18058 13088
rect 17994 13028 17998 13084
rect 17998 13028 18054 13084
rect 18054 13028 18058 13084
rect 17994 13024 18058 13028
rect 18074 13084 18138 13088
rect 18074 13028 18078 13084
rect 18078 13028 18134 13084
rect 18134 13028 18138 13084
rect 18074 13024 18138 13028
rect 18154 13084 18218 13088
rect 18154 13028 18158 13084
rect 18158 13028 18214 13084
rect 18214 13028 18218 13084
rect 18154 13024 18218 13028
rect 18234 13084 18298 13088
rect 18234 13028 18238 13084
rect 18238 13028 18294 13084
rect 18294 13028 18298 13084
rect 18234 13024 18298 13028
rect 23675 13084 23739 13088
rect 23675 13028 23679 13084
rect 23679 13028 23735 13084
rect 23735 13028 23739 13084
rect 23675 13024 23739 13028
rect 23755 13084 23819 13088
rect 23755 13028 23759 13084
rect 23759 13028 23815 13084
rect 23815 13028 23819 13084
rect 23755 13024 23819 13028
rect 23835 13084 23899 13088
rect 23835 13028 23839 13084
rect 23839 13028 23895 13084
rect 23895 13028 23899 13084
rect 23835 13024 23899 13028
rect 23915 13084 23979 13088
rect 23915 13028 23919 13084
rect 23919 13028 23975 13084
rect 23975 13028 23979 13084
rect 23915 13024 23979 13028
rect 3792 12540 3856 12544
rect 3792 12484 3796 12540
rect 3796 12484 3852 12540
rect 3852 12484 3856 12540
rect 3792 12480 3856 12484
rect 3872 12540 3936 12544
rect 3872 12484 3876 12540
rect 3876 12484 3932 12540
rect 3932 12484 3936 12540
rect 3872 12480 3936 12484
rect 3952 12540 4016 12544
rect 3952 12484 3956 12540
rect 3956 12484 4012 12540
rect 4012 12484 4016 12540
rect 3952 12480 4016 12484
rect 4032 12540 4096 12544
rect 4032 12484 4036 12540
rect 4036 12484 4092 12540
rect 4092 12484 4096 12540
rect 4032 12480 4096 12484
rect 9473 12540 9537 12544
rect 9473 12484 9477 12540
rect 9477 12484 9533 12540
rect 9533 12484 9537 12540
rect 9473 12480 9537 12484
rect 9553 12540 9617 12544
rect 9553 12484 9557 12540
rect 9557 12484 9613 12540
rect 9613 12484 9617 12540
rect 9553 12480 9617 12484
rect 9633 12540 9697 12544
rect 9633 12484 9637 12540
rect 9637 12484 9693 12540
rect 9693 12484 9697 12540
rect 9633 12480 9697 12484
rect 9713 12540 9777 12544
rect 9713 12484 9717 12540
rect 9717 12484 9773 12540
rect 9773 12484 9777 12540
rect 9713 12480 9777 12484
rect 15154 12540 15218 12544
rect 15154 12484 15158 12540
rect 15158 12484 15214 12540
rect 15214 12484 15218 12540
rect 15154 12480 15218 12484
rect 15234 12540 15298 12544
rect 15234 12484 15238 12540
rect 15238 12484 15294 12540
rect 15294 12484 15298 12540
rect 15234 12480 15298 12484
rect 15314 12540 15378 12544
rect 15314 12484 15318 12540
rect 15318 12484 15374 12540
rect 15374 12484 15378 12540
rect 15314 12480 15378 12484
rect 15394 12540 15458 12544
rect 15394 12484 15398 12540
rect 15398 12484 15454 12540
rect 15454 12484 15458 12540
rect 15394 12480 15458 12484
rect 13124 12336 13188 12340
rect 13124 12280 13174 12336
rect 13174 12280 13188 12336
rect 13124 12276 13188 12280
rect 20835 12540 20899 12544
rect 20835 12484 20839 12540
rect 20839 12484 20895 12540
rect 20895 12484 20899 12540
rect 20835 12480 20899 12484
rect 20915 12540 20979 12544
rect 20915 12484 20919 12540
rect 20919 12484 20975 12540
rect 20975 12484 20979 12540
rect 20915 12480 20979 12484
rect 20995 12540 21059 12544
rect 20995 12484 20999 12540
rect 20999 12484 21055 12540
rect 21055 12484 21059 12540
rect 20995 12480 21059 12484
rect 21075 12540 21139 12544
rect 21075 12484 21079 12540
rect 21079 12484 21135 12540
rect 21135 12484 21139 12540
rect 21075 12480 21139 12484
rect 6632 11996 6696 12000
rect 6632 11940 6636 11996
rect 6636 11940 6692 11996
rect 6692 11940 6696 11996
rect 6632 11936 6696 11940
rect 6712 11996 6776 12000
rect 6712 11940 6716 11996
rect 6716 11940 6772 11996
rect 6772 11940 6776 11996
rect 6712 11936 6776 11940
rect 6792 11996 6856 12000
rect 6792 11940 6796 11996
rect 6796 11940 6852 11996
rect 6852 11940 6856 11996
rect 6792 11936 6856 11940
rect 6872 11996 6936 12000
rect 6872 11940 6876 11996
rect 6876 11940 6932 11996
rect 6932 11940 6936 11996
rect 6872 11936 6936 11940
rect 12313 11996 12377 12000
rect 12313 11940 12317 11996
rect 12317 11940 12373 11996
rect 12373 11940 12377 11996
rect 12313 11936 12377 11940
rect 12393 11996 12457 12000
rect 12393 11940 12397 11996
rect 12397 11940 12453 11996
rect 12453 11940 12457 11996
rect 12393 11936 12457 11940
rect 12473 11996 12537 12000
rect 12473 11940 12477 11996
rect 12477 11940 12533 11996
rect 12533 11940 12537 11996
rect 12473 11936 12537 11940
rect 12553 11996 12617 12000
rect 12553 11940 12557 11996
rect 12557 11940 12613 11996
rect 12613 11940 12617 11996
rect 12553 11936 12617 11940
rect 17994 11996 18058 12000
rect 17994 11940 17998 11996
rect 17998 11940 18054 11996
rect 18054 11940 18058 11996
rect 17994 11936 18058 11940
rect 18074 11996 18138 12000
rect 18074 11940 18078 11996
rect 18078 11940 18134 11996
rect 18134 11940 18138 11996
rect 18074 11936 18138 11940
rect 18154 11996 18218 12000
rect 18154 11940 18158 11996
rect 18158 11940 18214 11996
rect 18214 11940 18218 11996
rect 18154 11936 18218 11940
rect 18234 11996 18298 12000
rect 18234 11940 18238 11996
rect 18238 11940 18294 11996
rect 18294 11940 18298 11996
rect 18234 11936 18298 11940
rect 23675 11996 23739 12000
rect 23675 11940 23679 11996
rect 23679 11940 23735 11996
rect 23735 11940 23739 11996
rect 23675 11936 23739 11940
rect 23755 11996 23819 12000
rect 23755 11940 23759 11996
rect 23759 11940 23815 11996
rect 23815 11940 23819 11996
rect 23755 11936 23819 11940
rect 23835 11996 23899 12000
rect 23835 11940 23839 11996
rect 23839 11940 23895 11996
rect 23895 11940 23899 11996
rect 23835 11936 23899 11940
rect 23915 11996 23979 12000
rect 23915 11940 23919 11996
rect 23919 11940 23975 11996
rect 23975 11940 23979 11996
rect 23915 11936 23979 11940
rect 14780 11732 14844 11796
rect 3792 11452 3856 11456
rect 3792 11396 3796 11452
rect 3796 11396 3852 11452
rect 3852 11396 3856 11452
rect 3792 11392 3856 11396
rect 3872 11452 3936 11456
rect 3872 11396 3876 11452
rect 3876 11396 3932 11452
rect 3932 11396 3936 11452
rect 3872 11392 3936 11396
rect 3952 11452 4016 11456
rect 3952 11396 3956 11452
rect 3956 11396 4012 11452
rect 4012 11396 4016 11452
rect 3952 11392 4016 11396
rect 4032 11452 4096 11456
rect 4032 11396 4036 11452
rect 4036 11396 4092 11452
rect 4092 11396 4096 11452
rect 4032 11392 4096 11396
rect 9473 11452 9537 11456
rect 9473 11396 9477 11452
rect 9477 11396 9533 11452
rect 9533 11396 9537 11452
rect 9473 11392 9537 11396
rect 9553 11452 9617 11456
rect 9553 11396 9557 11452
rect 9557 11396 9613 11452
rect 9613 11396 9617 11452
rect 9553 11392 9617 11396
rect 9633 11452 9697 11456
rect 9633 11396 9637 11452
rect 9637 11396 9693 11452
rect 9693 11396 9697 11452
rect 9633 11392 9697 11396
rect 9713 11452 9777 11456
rect 9713 11396 9717 11452
rect 9717 11396 9773 11452
rect 9773 11396 9777 11452
rect 9713 11392 9777 11396
rect 15154 11452 15218 11456
rect 15154 11396 15158 11452
rect 15158 11396 15214 11452
rect 15214 11396 15218 11452
rect 15154 11392 15218 11396
rect 15234 11452 15298 11456
rect 15234 11396 15238 11452
rect 15238 11396 15294 11452
rect 15294 11396 15298 11452
rect 15234 11392 15298 11396
rect 15314 11452 15378 11456
rect 15314 11396 15318 11452
rect 15318 11396 15374 11452
rect 15374 11396 15378 11452
rect 15314 11392 15378 11396
rect 15394 11452 15458 11456
rect 15394 11396 15398 11452
rect 15398 11396 15454 11452
rect 15454 11396 15458 11452
rect 15394 11392 15458 11396
rect 20835 11452 20899 11456
rect 20835 11396 20839 11452
rect 20839 11396 20895 11452
rect 20895 11396 20899 11452
rect 20835 11392 20899 11396
rect 20915 11452 20979 11456
rect 20915 11396 20919 11452
rect 20919 11396 20975 11452
rect 20975 11396 20979 11452
rect 20915 11392 20979 11396
rect 20995 11452 21059 11456
rect 20995 11396 20999 11452
rect 20999 11396 21055 11452
rect 21055 11396 21059 11452
rect 20995 11392 21059 11396
rect 21075 11452 21139 11456
rect 21075 11396 21079 11452
rect 21079 11396 21135 11452
rect 21135 11396 21139 11452
rect 21075 11392 21139 11396
rect 6632 10908 6696 10912
rect 6632 10852 6636 10908
rect 6636 10852 6692 10908
rect 6692 10852 6696 10908
rect 6632 10848 6696 10852
rect 6712 10908 6776 10912
rect 6712 10852 6716 10908
rect 6716 10852 6772 10908
rect 6772 10852 6776 10908
rect 6712 10848 6776 10852
rect 6792 10908 6856 10912
rect 6792 10852 6796 10908
rect 6796 10852 6852 10908
rect 6852 10852 6856 10908
rect 6792 10848 6856 10852
rect 6872 10908 6936 10912
rect 6872 10852 6876 10908
rect 6876 10852 6932 10908
rect 6932 10852 6936 10908
rect 6872 10848 6936 10852
rect 12313 10908 12377 10912
rect 12313 10852 12317 10908
rect 12317 10852 12373 10908
rect 12373 10852 12377 10908
rect 12313 10848 12377 10852
rect 12393 10908 12457 10912
rect 12393 10852 12397 10908
rect 12397 10852 12453 10908
rect 12453 10852 12457 10908
rect 12393 10848 12457 10852
rect 12473 10908 12537 10912
rect 12473 10852 12477 10908
rect 12477 10852 12533 10908
rect 12533 10852 12537 10908
rect 12473 10848 12537 10852
rect 12553 10908 12617 10912
rect 12553 10852 12557 10908
rect 12557 10852 12613 10908
rect 12613 10852 12617 10908
rect 12553 10848 12617 10852
rect 17994 10908 18058 10912
rect 17994 10852 17998 10908
rect 17998 10852 18054 10908
rect 18054 10852 18058 10908
rect 17994 10848 18058 10852
rect 18074 10908 18138 10912
rect 18074 10852 18078 10908
rect 18078 10852 18134 10908
rect 18134 10852 18138 10908
rect 18074 10848 18138 10852
rect 18154 10908 18218 10912
rect 18154 10852 18158 10908
rect 18158 10852 18214 10908
rect 18214 10852 18218 10908
rect 18154 10848 18218 10852
rect 18234 10908 18298 10912
rect 18234 10852 18238 10908
rect 18238 10852 18294 10908
rect 18294 10852 18298 10908
rect 18234 10848 18298 10852
rect 23675 10908 23739 10912
rect 23675 10852 23679 10908
rect 23679 10852 23735 10908
rect 23735 10852 23739 10908
rect 23675 10848 23739 10852
rect 23755 10908 23819 10912
rect 23755 10852 23759 10908
rect 23759 10852 23815 10908
rect 23815 10852 23819 10908
rect 23755 10848 23819 10852
rect 23835 10908 23899 10912
rect 23835 10852 23839 10908
rect 23839 10852 23895 10908
rect 23895 10852 23899 10908
rect 23835 10848 23899 10852
rect 23915 10908 23979 10912
rect 23915 10852 23919 10908
rect 23919 10852 23975 10908
rect 23975 10852 23979 10908
rect 23915 10848 23979 10852
rect 5396 10644 5460 10708
rect 22324 10644 22388 10708
rect 7236 10568 7300 10572
rect 7236 10512 7286 10568
rect 7286 10512 7300 10568
rect 7236 10508 7300 10512
rect 3792 10364 3856 10368
rect 3792 10308 3796 10364
rect 3796 10308 3852 10364
rect 3852 10308 3856 10364
rect 3792 10304 3856 10308
rect 3872 10364 3936 10368
rect 3872 10308 3876 10364
rect 3876 10308 3932 10364
rect 3932 10308 3936 10364
rect 3872 10304 3936 10308
rect 3952 10364 4016 10368
rect 3952 10308 3956 10364
rect 3956 10308 4012 10364
rect 4012 10308 4016 10364
rect 3952 10304 4016 10308
rect 4032 10364 4096 10368
rect 4032 10308 4036 10364
rect 4036 10308 4092 10364
rect 4092 10308 4096 10364
rect 4032 10304 4096 10308
rect 9473 10364 9537 10368
rect 9473 10308 9477 10364
rect 9477 10308 9533 10364
rect 9533 10308 9537 10364
rect 9473 10304 9537 10308
rect 9553 10364 9617 10368
rect 9553 10308 9557 10364
rect 9557 10308 9613 10364
rect 9613 10308 9617 10364
rect 9553 10304 9617 10308
rect 9633 10364 9697 10368
rect 9633 10308 9637 10364
rect 9637 10308 9693 10364
rect 9693 10308 9697 10364
rect 9633 10304 9697 10308
rect 9713 10364 9777 10368
rect 9713 10308 9717 10364
rect 9717 10308 9773 10364
rect 9773 10308 9777 10364
rect 9713 10304 9777 10308
rect 15154 10364 15218 10368
rect 15154 10308 15158 10364
rect 15158 10308 15214 10364
rect 15214 10308 15218 10364
rect 15154 10304 15218 10308
rect 15234 10364 15298 10368
rect 15234 10308 15238 10364
rect 15238 10308 15294 10364
rect 15294 10308 15298 10364
rect 15234 10304 15298 10308
rect 15314 10364 15378 10368
rect 15314 10308 15318 10364
rect 15318 10308 15374 10364
rect 15374 10308 15378 10364
rect 15314 10304 15378 10308
rect 15394 10364 15458 10368
rect 15394 10308 15398 10364
rect 15398 10308 15454 10364
rect 15454 10308 15458 10364
rect 15394 10304 15458 10308
rect 20835 10364 20899 10368
rect 20835 10308 20839 10364
rect 20839 10308 20895 10364
rect 20895 10308 20899 10364
rect 20835 10304 20899 10308
rect 20915 10364 20979 10368
rect 20915 10308 20919 10364
rect 20919 10308 20975 10364
rect 20975 10308 20979 10364
rect 20915 10304 20979 10308
rect 20995 10364 21059 10368
rect 20995 10308 20999 10364
rect 20999 10308 21055 10364
rect 21055 10308 21059 10364
rect 20995 10304 21059 10308
rect 21075 10364 21139 10368
rect 21075 10308 21079 10364
rect 21079 10308 21135 10364
rect 21135 10308 21139 10364
rect 21075 10304 21139 10308
rect 17724 9964 17788 10028
rect 10364 9828 10428 9892
rect 6632 9820 6696 9824
rect 6632 9764 6636 9820
rect 6636 9764 6692 9820
rect 6692 9764 6696 9820
rect 6632 9760 6696 9764
rect 6712 9820 6776 9824
rect 6712 9764 6716 9820
rect 6716 9764 6772 9820
rect 6772 9764 6776 9820
rect 6712 9760 6776 9764
rect 6792 9820 6856 9824
rect 6792 9764 6796 9820
rect 6796 9764 6852 9820
rect 6852 9764 6856 9820
rect 6792 9760 6856 9764
rect 6872 9820 6936 9824
rect 6872 9764 6876 9820
rect 6876 9764 6932 9820
rect 6932 9764 6936 9820
rect 6872 9760 6936 9764
rect 12313 9820 12377 9824
rect 12313 9764 12317 9820
rect 12317 9764 12373 9820
rect 12373 9764 12377 9820
rect 12313 9760 12377 9764
rect 12393 9820 12457 9824
rect 12393 9764 12397 9820
rect 12397 9764 12453 9820
rect 12453 9764 12457 9820
rect 12393 9760 12457 9764
rect 12473 9820 12537 9824
rect 12473 9764 12477 9820
rect 12477 9764 12533 9820
rect 12533 9764 12537 9820
rect 12473 9760 12537 9764
rect 12553 9820 12617 9824
rect 12553 9764 12557 9820
rect 12557 9764 12613 9820
rect 12613 9764 12617 9820
rect 12553 9760 12617 9764
rect 17994 9820 18058 9824
rect 17994 9764 17998 9820
rect 17998 9764 18054 9820
rect 18054 9764 18058 9820
rect 17994 9760 18058 9764
rect 18074 9820 18138 9824
rect 18074 9764 18078 9820
rect 18078 9764 18134 9820
rect 18134 9764 18138 9820
rect 18074 9760 18138 9764
rect 18154 9820 18218 9824
rect 18154 9764 18158 9820
rect 18158 9764 18214 9820
rect 18214 9764 18218 9820
rect 18154 9760 18218 9764
rect 18234 9820 18298 9824
rect 18234 9764 18238 9820
rect 18238 9764 18294 9820
rect 18294 9764 18298 9820
rect 18234 9760 18298 9764
rect 23675 9820 23739 9824
rect 23675 9764 23679 9820
rect 23679 9764 23735 9820
rect 23735 9764 23739 9820
rect 23675 9760 23739 9764
rect 23755 9820 23819 9824
rect 23755 9764 23759 9820
rect 23759 9764 23815 9820
rect 23815 9764 23819 9820
rect 23755 9760 23819 9764
rect 23835 9820 23899 9824
rect 23835 9764 23839 9820
rect 23839 9764 23895 9820
rect 23895 9764 23899 9820
rect 23835 9760 23899 9764
rect 23915 9820 23979 9824
rect 23915 9764 23919 9820
rect 23919 9764 23975 9820
rect 23975 9764 23979 9820
rect 23915 9760 23979 9764
rect 3792 9276 3856 9280
rect 3792 9220 3796 9276
rect 3796 9220 3852 9276
rect 3852 9220 3856 9276
rect 3792 9216 3856 9220
rect 3872 9276 3936 9280
rect 3872 9220 3876 9276
rect 3876 9220 3932 9276
rect 3932 9220 3936 9276
rect 3872 9216 3936 9220
rect 3952 9276 4016 9280
rect 3952 9220 3956 9276
rect 3956 9220 4012 9276
rect 4012 9220 4016 9276
rect 3952 9216 4016 9220
rect 4032 9276 4096 9280
rect 4032 9220 4036 9276
rect 4036 9220 4092 9276
rect 4092 9220 4096 9276
rect 4032 9216 4096 9220
rect 9473 9276 9537 9280
rect 9473 9220 9477 9276
rect 9477 9220 9533 9276
rect 9533 9220 9537 9276
rect 9473 9216 9537 9220
rect 9553 9276 9617 9280
rect 9553 9220 9557 9276
rect 9557 9220 9613 9276
rect 9613 9220 9617 9276
rect 9553 9216 9617 9220
rect 9633 9276 9697 9280
rect 9633 9220 9637 9276
rect 9637 9220 9693 9276
rect 9693 9220 9697 9276
rect 9633 9216 9697 9220
rect 9713 9276 9777 9280
rect 9713 9220 9717 9276
rect 9717 9220 9773 9276
rect 9773 9220 9777 9276
rect 9713 9216 9777 9220
rect 15154 9276 15218 9280
rect 15154 9220 15158 9276
rect 15158 9220 15214 9276
rect 15214 9220 15218 9276
rect 15154 9216 15218 9220
rect 15234 9276 15298 9280
rect 15234 9220 15238 9276
rect 15238 9220 15294 9276
rect 15294 9220 15298 9276
rect 15234 9216 15298 9220
rect 15314 9276 15378 9280
rect 15314 9220 15318 9276
rect 15318 9220 15374 9276
rect 15374 9220 15378 9276
rect 15314 9216 15378 9220
rect 15394 9276 15458 9280
rect 15394 9220 15398 9276
rect 15398 9220 15454 9276
rect 15454 9220 15458 9276
rect 15394 9216 15458 9220
rect 20835 9276 20899 9280
rect 20835 9220 20839 9276
rect 20839 9220 20895 9276
rect 20895 9220 20899 9276
rect 20835 9216 20899 9220
rect 20915 9276 20979 9280
rect 20915 9220 20919 9276
rect 20919 9220 20975 9276
rect 20975 9220 20979 9276
rect 20915 9216 20979 9220
rect 20995 9276 21059 9280
rect 20995 9220 20999 9276
rect 20999 9220 21055 9276
rect 21055 9220 21059 9276
rect 20995 9216 21059 9220
rect 21075 9276 21139 9280
rect 21075 9220 21079 9276
rect 21079 9220 21135 9276
rect 21135 9220 21139 9276
rect 21075 9216 21139 9220
rect 6632 8732 6696 8736
rect 6632 8676 6636 8732
rect 6636 8676 6692 8732
rect 6692 8676 6696 8732
rect 6632 8672 6696 8676
rect 6712 8732 6776 8736
rect 6712 8676 6716 8732
rect 6716 8676 6772 8732
rect 6772 8676 6776 8732
rect 6712 8672 6776 8676
rect 6792 8732 6856 8736
rect 6792 8676 6796 8732
rect 6796 8676 6852 8732
rect 6852 8676 6856 8732
rect 6792 8672 6856 8676
rect 6872 8732 6936 8736
rect 6872 8676 6876 8732
rect 6876 8676 6932 8732
rect 6932 8676 6936 8732
rect 6872 8672 6936 8676
rect 12313 8732 12377 8736
rect 12313 8676 12317 8732
rect 12317 8676 12373 8732
rect 12373 8676 12377 8732
rect 12313 8672 12377 8676
rect 12393 8732 12457 8736
rect 12393 8676 12397 8732
rect 12397 8676 12453 8732
rect 12453 8676 12457 8732
rect 12393 8672 12457 8676
rect 12473 8732 12537 8736
rect 12473 8676 12477 8732
rect 12477 8676 12533 8732
rect 12533 8676 12537 8732
rect 12473 8672 12537 8676
rect 12553 8732 12617 8736
rect 12553 8676 12557 8732
rect 12557 8676 12613 8732
rect 12613 8676 12617 8732
rect 12553 8672 12617 8676
rect 17994 8732 18058 8736
rect 17994 8676 17998 8732
rect 17998 8676 18054 8732
rect 18054 8676 18058 8732
rect 17994 8672 18058 8676
rect 18074 8732 18138 8736
rect 18074 8676 18078 8732
rect 18078 8676 18134 8732
rect 18134 8676 18138 8732
rect 18074 8672 18138 8676
rect 18154 8732 18218 8736
rect 18154 8676 18158 8732
rect 18158 8676 18214 8732
rect 18214 8676 18218 8732
rect 18154 8672 18218 8676
rect 18234 8732 18298 8736
rect 18234 8676 18238 8732
rect 18238 8676 18294 8732
rect 18294 8676 18298 8732
rect 18234 8672 18298 8676
rect 23675 8732 23739 8736
rect 23675 8676 23679 8732
rect 23679 8676 23735 8732
rect 23735 8676 23739 8732
rect 23675 8672 23739 8676
rect 23755 8732 23819 8736
rect 23755 8676 23759 8732
rect 23759 8676 23815 8732
rect 23815 8676 23819 8732
rect 23755 8672 23819 8676
rect 23835 8732 23899 8736
rect 23835 8676 23839 8732
rect 23839 8676 23895 8732
rect 23895 8676 23899 8732
rect 23835 8672 23899 8676
rect 23915 8732 23979 8736
rect 23915 8676 23919 8732
rect 23919 8676 23975 8732
rect 23975 8676 23979 8732
rect 23915 8672 23979 8676
rect 16252 8332 16316 8396
rect 3792 8188 3856 8192
rect 3792 8132 3796 8188
rect 3796 8132 3852 8188
rect 3852 8132 3856 8188
rect 3792 8128 3856 8132
rect 3872 8188 3936 8192
rect 3872 8132 3876 8188
rect 3876 8132 3932 8188
rect 3932 8132 3936 8188
rect 3872 8128 3936 8132
rect 3952 8188 4016 8192
rect 3952 8132 3956 8188
rect 3956 8132 4012 8188
rect 4012 8132 4016 8188
rect 3952 8128 4016 8132
rect 4032 8188 4096 8192
rect 4032 8132 4036 8188
rect 4036 8132 4092 8188
rect 4092 8132 4096 8188
rect 4032 8128 4096 8132
rect 9473 8188 9537 8192
rect 9473 8132 9477 8188
rect 9477 8132 9533 8188
rect 9533 8132 9537 8188
rect 9473 8128 9537 8132
rect 9553 8188 9617 8192
rect 9553 8132 9557 8188
rect 9557 8132 9613 8188
rect 9613 8132 9617 8188
rect 9553 8128 9617 8132
rect 9633 8188 9697 8192
rect 9633 8132 9637 8188
rect 9637 8132 9693 8188
rect 9693 8132 9697 8188
rect 9633 8128 9697 8132
rect 9713 8188 9777 8192
rect 9713 8132 9717 8188
rect 9717 8132 9773 8188
rect 9773 8132 9777 8188
rect 9713 8128 9777 8132
rect 15154 8188 15218 8192
rect 15154 8132 15158 8188
rect 15158 8132 15214 8188
rect 15214 8132 15218 8188
rect 15154 8128 15218 8132
rect 15234 8188 15298 8192
rect 15234 8132 15238 8188
rect 15238 8132 15294 8188
rect 15294 8132 15298 8188
rect 15234 8128 15298 8132
rect 15314 8188 15378 8192
rect 15314 8132 15318 8188
rect 15318 8132 15374 8188
rect 15374 8132 15378 8188
rect 15314 8128 15378 8132
rect 15394 8188 15458 8192
rect 15394 8132 15398 8188
rect 15398 8132 15454 8188
rect 15454 8132 15458 8188
rect 15394 8128 15458 8132
rect 20835 8188 20899 8192
rect 20835 8132 20839 8188
rect 20839 8132 20895 8188
rect 20895 8132 20899 8188
rect 20835 8128 20899 8132
rect 20915 8188 20979 8192
rect 20915 8132 20919 8188
rect 20919 8132 20975 8188
rect 20975 8132 20979 8188
rect 20915 8128 20979 8132
rect 20995 8188 21059 8192
rect 20995 8132 20999 8188
rect 20999 8132 21055 8188
rect 21055 8132 21059 8188
rect 20995 8128 21059 8132
rect 21075 8188 21139 8192
rect 21075 8132 21079 8188
rect 21079 8132 21135 8188
rect 21135 8132 21139 8188
rect 21075 8128 21139 8132
rect 6632 7644 6696 7648
rect 6632 7588 6636 7644
rect 6636 7588 6692 7644
rect 6692 7588 6696 7644
rect 6632 7584 6696 7588
rect 6712 7644 6776 7648
rect 6712 7588 6716 7644
rect 6716 7588 6772 7644
rect 6772 7588 6776 7644
rect 6712 7584 6776 7588
rect 6792 7644 6856 7648
rect 6792 7588 6796 7644
rect 6796 7588 6852 7644
rect 6852 7588 6856 7644
rect 6792 7584 6856 7588
rect 6872 7644 6936 7648
rect 6872 7588 6876 7644
rect 6876 7588 6932 7644
rect 6932 7588 6936 7644
rect 6872 7584 6936 7588
rect 12313 7644 12377 7648
rect 12313 7588 12317 7644
rect 12317 7588 12373 7644
rect 12373 7588 12377 7644
rect 12313 7584 12377 7588
rect 12393 7644 12457 7648
rect 12393 7588 12397 7644
rect 12397 7588 12453 7644
rect 12453 7588 12457 7644
rect 12393 7584 12457 7588
rect 12473 7644 12537 7648
rect 12473 7588 12477 7644
rect 12477 7588 12533 7644
rect 12533 7588 12537 7644
rect 12473 7584 12537 7588
rect 12553 7644 12617 7648
rect 12553 7588 12557 7644
rect 12557 7588 12613 7644
rect 12613 7588 12617 7644
rect 12553 7584 12617 7588
rect 17994 7644 18058 7648
rect 17994 7588 17998 7644
rect 17998 7588 18054 7644
rect 18054 7588 18058 7644
rect 17994 7584 18058 7588
rect 18074 7644 18138 7648
rect 18074 7588 18078 7644
rect 18078 7588 18134 7644
rect 18134 7588 18138 7644
rect 18074 7584 18138 7588
rect 18154 7644 18218 7648
rect 18154 7588 18158 7644
rect 18158 7588 18214 7644
rect 18214 7588 18218 7644
rect 18154 7584 18218 7588
rect 18234 7644 18298 7648
rect 18234 7588 18238 7644
rect 18238 7588 18294 7644
rect 18294 7588 18298 7644
rect 18234 7584 18298 7588
rect 23675 7644 23739 7648
rect 23675 7588 23679 7644
rect 23679 7588 23735 7644
rect 23735 7588 23739 7644
rect 23675 7584 23739 7588
rect 23755 7644 23819 7648
rect 23755 7588 23759 7644
rect 23759 7588 23815 7644
rect 23815 7588 23819 7644
rect 23755 7584 23819 7588
rect 23835 7644 23899 7648
rect 23835 7588 23839 7644
rect 23839 7588 23895 7644
rect 23895 7588 23899 7644
rect 23835 7584 23899 7588
rect 23915 7644 23979 7648
rect 23915 7588 23919 7644
rect 23919 7588 23975 7644
rect 23975 7588 23979 7644
rect 23915 7584 23979 7588
rect 3792 7100 3856 7104
rect 3792 7044 3796 7100
rect 3796 7044 3852 7100
rect 3852 7044 3856 7100
rect 3792 7040 3856 7044
rect 3872 7100 3936 7104
rect 3872 7044 3876 7100
rect 3876 7044 3932 7100
rect 3932 7044 3936 7100
rect 3872 7040 3936 7044
rect 3952 7100 4016 7104
rect 3952 7044 3956 7100
rect 3956 7044 4012 7100
rect 4012 7044 4016 7100
rect 3952 7040 4016 7044
rect 4032 7100 4096 7104
rect 4032 7044 4036 7100
rect 4036 7044 4092 7100
rect 4092 7044 4096 7100
rect 4032 7040 4096 7044
rect 9473 7100 9537 7104
rect 9473 7044 9477 7100
rect 9477 7044 9533 7100
rect 9533 7044 9537 7100
rect 9473 7040 9537 7044
rect 9553 7100 9617 7104
rect 9553 7044 9557 7100
rect 9557 7044 9613 7100
rect 9613 7044 9617 7100
rect 9553 7040 9617 7044
rect 9633 7100 9697 7104
rect 9633 7044 9637 7100
rect 9637 7044 9693 7100
rect 9693 7044 9697 7100
rect 9633 7040 9697 7044
rect 9713 7100 9777 7104
rect 9713 7044 9717 7100
rect 9717 7044 9773 7100
rect 9773 7044 9777 7100
rect 9713 7040 9777 7044
rect 15154 7100 15218 7104
rect 15154 7044 15158 7100
rect 15158 7044 15214 7100
rect 15214 7044 15218 7100
rect 15154 7040 15218 7044
rect 15234 7100 15298 7104
rect 15234 7044 15238 7100
rect 15238 7044 15294 7100
rect 15294 7044 15298 7100
rect 15234 7040 15298 7044
rect 15314 7100 15378 7104
rect 15314 7044 15318 7100
rect 15318 7044 15374 7100
rect 15374 7044 15378 7100
rect 15314 7040 15378 7044
rect 15394 7100 15458 7104
rect 15394 7044 15398 7100
rect 15398 7044 15454 7100
rect 15454 7044 15458 7100
rect 15394 7040 15458 7044
rect 20835 7100 20899 7104
rect 20835 7044 20839 7100
rect 20839 7044 20895 7100
rect 20895 7044 20899 7100
rect 20835 7040 20899 7044
rect 20915 7100 20979 7104
rect 20915 7044 20919 7100
rect 20919 7044 20975 7100
rect 20975 7044 20979 7100
rect 20915 7040 20979 7044
rect 20995 7100 21059 7104
rect 20995 7044 20999 7100
rect 20999 7044 21055 7100
rect 21055 7044 21059 7100
rect 20995 7040 21059 7044
rect 21075 7100 21139 7104
rect 21075 7044 21079 7100
rect 21079 7044 21135 7100
rect 21135 7044 21139 7100
rect 21075 7040 21139 7044
rect 21404 6836 21468 6900
rect 6632 6556 6696 6560
rect 6632 6500 6636 6556
rect 6636 6500 6692 6556
rect 6692 6500 6696 6556
rect 6632 6496 6696 6500
rect 6712 6556 6776 6560
rect 6712 6500 6716 6556
rect 6716 6500 6772 6556
rect 6772 6500 6776 6556
rect 6712 6496 6776 6500
rect 6792 6556 6856 6560
rect 6792 6500 6796 6556
rect 6796 6500 6852 6556
rect 6852 6500 6856 6556
rect 6792 6496 6856 6500
rect 6872 6556 6936 6560
rect 6872 6500 6876 6556
rect 6876 6500 6932 6556
rect 6932 6500 6936 6556
rect 6872 6496 6936 6500
rect 12313 6556 12377 6560
rect 12313 6500 12317 6556
rect 12317 6500 12373 6556
rect 12373 6500 12377 6556
rect 12313 6496 12377 6500
rect 12393 6556 12457 6560
rect 12393 6500 12397 6556
rect 12397 6500 12453 6556
rect 12453 6500 12457 6556
rect 12393 6496 12457 6500
rect 12473 6556 12537 6560
rect 12473 6500 12477 6556
rect 12477 6500 12533 6556
rect 12533 6500 12537 6556
rect 12473 6496 12537 6500
rect 12553 6556 12617 6560
rect 12553 6500 12557 6556
rect 12557 6500 12613 6556
rect 12613 6500 12617 6556
rect 12553 6496 12617 6500
rect 17994 6556 18058 6560
rect 17994 6500 17998 6556
rect 17998 6500 18054 6556
rect 18054 6500 18058 6556
rect 17994 6496 18058 6500
rect 18074 6556 18138 6560
rect 18074 6500 18078 6556
rect 18078 6500 18134 6556
rect 18134 6500 18138 6556
rect 18074 6496 18138 6500
rect 18154 6556 18218 6560
rect 18154 6500 18158 6556
rect 18158 6500 18214 6556
rect 18214 6500 18218 6556
rect 18154 6496 18218 6500
rect 18234 6556 18298 6560
rect 18234 6500 18238 6556
rect 18238 6500 18294 6556
rect 18294 6500 18298 6556
rect 18234 6496 18298 6500
rect 23675 6556 23739 6560
rect 23675 6500 23679 6556
rect 23679 6500 23735 6556
rect 23735 6500 23739 6556
rect 23675 6496 23739 6500
rect 23755 6556 23819 6560
rect 23755 6500 23759 6556
rect 23759 6500 23815 6556
rect 23815 6500 23819 6556
rect 23755 6496 23819 6500
rect 23835 6556 23899 6560
rect 23835 6500 23839 6556
rect 23839 6500 23895 6556
rect 23895 6500 23899 6556
rect 23835 6496 23899 6500
rect 23915 6556 23979 6560
rect 23915 6500 23919 6556
rect 23919 6500 23975 6556
rect 23975 6500 23979 6556
rect 23915 6496 23979 6500
rect 3792 6012 3856 6016
rect 3792 5956 3796 6012
rect 3796 5956 3852 6012
rect 3852 5956 3856 6012
rect 3792 5952 3856 5956
rect 3872 6012 3936 6016
rect 3872 5956 3876 6012
rect 3876 5956 3932 6012
rect 3932 5956 3936 6012
rect 3872 5952 3936 5956
rect 3952 6012 4016 6016
rect 3952 5956 3956 6012
rect 3956 5956 4012 6012
rect 4012 5956 4016 6012
rect 3952 5952 4016 5956
rect 4032 6012 4096 6016
rect 4032 5956 4036 6012
rect 4036 5956 4092 6012
rect 4092 5956 4096 6012
rect 4032 5952 4096 5956
rect 9473 6012 9537 6016
rect 9473 5956 9477 6012
rect 9477 5956 9533 6012
rect 9533 5956 9537 6012
rect 9473 5952 9537 5956
rect 9553 6012 9617 6016
rect 9553 5956 9557 6012
rect 9557 5956 9613 6012
rect 9613 5956 9617 6012
rect 9553 5952 9617 5956
rect 9633 6012 9697 6016
rect 9633 5956 9637 6012
rect 9637 5956 9693 6012
rect 9693 5956 9697 6012
rect 9633 5952 9697 5956
rect 9713 6012 9777 6016
rect 9713 5956 9717 6012
rect 9717 5956 9773 6012
rect 9773 5956 9777 6012
rect 9713 5952 9777 5956
rect 15154 6012 15218 6016
rect 15154 5956 15158 6012
rect 15158 5956 15214 6012
rect 15214 5956 15218 6012
rect 15154 5952 15218 5956
rect 15234 6012 15298 6016
rect 15234 5956 15238 6012
rect 15238 5956 15294 6012
rect 15294 5956 15298 6012
rect 15234 5952 15298 5956
rect 15314 6012 15378 6016
rect 15314 5956 15318 6012
rect 15318 5956 15374 6012
rect 15374 5956 15378 6012
rect 15314 5952 15378 5956
rect 15394 6012 15458 6016
rect 15394 5956 15398 6012
rect 15398 5956 15454 6012
rect 15454 5956 15458 6012
rect 15394 5952 15458 5956
rect 20835 6012 20899 6016
rect 20835 5956 20839 6012
rect 20839 5956 20895 6012
rect 20895 5956 20899 6012
rect 20835 5952 20899 5956
rect 20915 6012 20979 6016
rect 20915 5956 20919 6012
rect 20919 5956 20975 6012
rect 20975 5956 20979 6012
rect 20915 5952 20979 5956
rect 20995 6012 21059 6016
rect 20995 5956 20999 6012
rect 20999 5956 21055 6012
rect 21055 5956 21059 6012
rect 20995 5952 21059 5956
rect 21075 6012 21139 6016
rect 21075 5956 21079 6012
rect 21079 5956 21135 6012
rect 21135 5956 21139 6012
rect 21075 5952 21139 5956
rect 10364 5476 10428 5540
rect 6632 5468 6696 5472
rect 6632 5412 6636 5468
rect 6636 5412 6692 5468
rect 6692 5412 6696 5468
rect 6632 5408 6696 5412
rect 6712 5468 6776 5472
rect 6712 5412 6716 5468
rect 6716 5412 6772 5468
rect 6772 5412 6776 5468
rect 6712 5408 6776 5412
rect 6792 5468 6856 5472
rect 6792 5412 6796 5468
rect 6796 5412 6852 5468
rect 6852 5412 6856 5468
rect 6792 5408 6856 5412
rect 6872 5468 6936 5472
rect 6872 5412 6876 5468
rect 6876 5412 6932 5468
rect 6932 5412 6936 5468
rect 6872 5408 6936 5412
rect 12313 5468 12377 5472
rect 12313 5412 12317 5468
rect 12317 5412 12373 5468
rect 12373 5412 12377 5468
rect 12313 5408 12377 5412
rect 12393 5468 12457 5472
rect 12393 5412 12397 5468
rect 12397 5412 12453 5468
rect 12453 5412 12457 5468
rect 12393 5408 12457 5412
rect 12473 5468 12537 5472
rect 12473 5412 12477 5468
rect 12477 5412 12533 5468
rect 12533 5412 12537 5468
rect 12473 5408 12537 5412
rect 12553 5468 12617 5472
rect 12553 5412 12557 5468
rect 12557 5412 12613 5468
rect 12613 5412 12617 5468
rect 12553 5408 12617 5412
rect 17994 5468 18058 5472
rect 17994 5412 17998 5468
rect 17998 5412 18054 5468
rect 18054 5412 18058 5468
rect 17994 5408 18058 5412
rect 18074 5468 18138 5472
rect 18074 5412 18078 5468
rect 18078 5412 18134 5468
rect 18134 5412 18138 5468
rect 18074 5408 18138 5412
rect 18154 5468 18218 5472
rect 18154 5412 18158 5468
rect 18158 5412 18214 5468
rect 18214 5412 18218 5468
rect 18154 5408 18218 5412
rect 18234 5468 18298 5472
rect 18234 5412 18238 5468
rect 18238 5412 18294 5468
rect 18294 5412 18298 5468
rect 18234 5408 18298 5412
rect 23675 5468 23739 5472
rect 23675 5412 23679 5468
rect 23679 5412 23735 5468
rect 23735 5412 23739 5468
rect 23675 5408 23739 5412
rect 23755 5468 23819 5472
rect 23755 5412 23759 5468
rect 23759 5412 23815 5468
rect 23815 5412 23819 5468
rect 23755 5408 23819 5412
rect 23835 5468 23899 5472
rect 23835 5412 23839 5468
rect 23839 5412 23895 5468
rect 23895 5412 23899 5468
rect 23835 5408 23899 5412
rect 23915 5468 23979 5472
rect 23915 5412 23919 5468
rect 23919 5412 23975 5468
rect 23975 5412 23979 5468
rect 23915 5408 23979 5412
rect 7236 5068 7300 5132
rect 3792 4924 3856 4928
rect 3792 4868 3796 4924
rect 3796 4868 3852 4924
rect 3852 4868 3856 4924
rect 3792 4864 3856 4868
rect 3872 4924 3936 4928
rect 3872 4868 3876 4924
rect 3876 4868 3932 4924
rect 3932 4868 3936 4924
rect 3872 4864 3936 4868
rect 3952 4924 4016 4928
rect 3952 4868 3956 4924
rect 3956 4868 4012 4924
rect 4012 4868 4016 4924
rect 3952 4864 4016 4868
rect 4032 4924 4096 4928
rect 4032 4868 4036 4924
rect 4036 4868 4092 4924
rect 4092 4868 4096 4924
rect 4032 4864 4096 4868
rect 9473 4924 9537 4928
rect 9473 4868 9477 4924
rect 9477 4868 9533 4924
rect 9533 4868 9537 4924
rect 9473 4864 9537 4868
rect 9553 4924 9617 4928
rect 9553 4868 9557 4924
rect 9557 4868 9613 4924
rect 9613 4868 9617 4924
rect 9553 4864 9617 4868
rect 9633 4924 9697 4928
rect 9633 4868 9637 4924
rect 9637 4868 9693 4924
rect 9693 4868 9697 4924
rect 9633 4864 9697 4868
rect 9713 4924 9777 4928
rect 9713 4868 9717 4924
rect 9717 4868 9773 4924
rect 9773 4868 9777 4924
rect 9713 4864 9777 4868
rect 15154 4924 15218 4928
rect 15154 4868 15158 4924
rect 15158 4868 15214 4924
rect 15214 4868 15218 4924
rect 15154 4864 15218 4868
rect 15234 4924 15298 4928
rect 15234 4868 15238 4924
rect 15238 4868 15294 4924
rect 15294 4868 15298 4924
rect 15234 4864 15298 4868
rect 15314 4924 15378 4928
rect 15314 4868 15318 4924
rect 15318 4868 15374 4924
rect 15374 4868 15378 4924
rect 15314 4864 15378 4868
rect 15394 4924 15458 4928
rect 15394 4868 15398 4924
rect 15398 4868 15454 4924
rect 15454 4868 15458 4924
rect 15394 4864 15458 4868
rect 20835 4924 20899 4928
rect 20835 4868 20839 4924
rect 20839 4868 20895 4924
rect 20895 4868 20899 4924
rect 20835 4864 20899 4868
rect 20915 4924 20979 4928
rect 20915 4868 20919 4924
rect 20919 4868 20975 4924
rect 20975 4868 20979 4924
rect 20915 4864 20979 4868
rect 20995 4924 21059 4928
rect 20995 4868 20999 4924
rect 20999 4868 21055 4924
rect 21055 4868 21059 4924
rect 20995 4864 21059 4868
rect 21075 4924 21139 4928
rect 21075 4868 21079 4924
rect 21079 4868 21135 4924
rect 21135 4868 21139 4924
rect 21075 4864 21139 4868
rect 17724 4660 17788 4724
rect 6632 4380 6696 4384
rect 6632 4324 6636 4380
rect 6636 4324 6692 4380
rect 6692 4324 6696 4380
rect 6632 4320 6696 4324
rect 6712 4380 6776 4384
rect 6712 4324 6716 4380
rect 6716 4324 6772 4380
rect 6772 4324 6776 4380
rect 6712 4320 6776 4324
rect 6792 4380 6856 4384
rect 6792 4324 6796 4380
rect 6796 4324 6852 4380
rect 6852 4324 6856 4380
rect 6792 4320 6856 4324
rect 6872 4380 6936 4384
rect 6872 4324 6876 4380
rect 6876 4324 6932 4380
rect 6932 4324 6936 4380
rect 6872 4320 6936 4324
rect 12313 4380 12377 4384
rect 12313 4324 12317 4380
rect 12317 4324 12373 4380
rect 12373 4324 12377 4380
rect 12313 4320 12377 4324
rect 12393 4380 12457 4384
rect 12393 4324 12397 4380
rect 12397 4324 12453 4380
rect 12453 4324 12457 4380
rect 12393 4320 12457 4324
rect 12473 4380 12537 4384
rect 12473 4324 12477 4380
rect 12477 4324 12533 4380
rect 12533 4324 12537 4380
rect 12473 4320 12537 4324
rect 12553 4380 12617 4384
rect 12553 4324 12557 4380
rect 12557 4324 12613 4380
rect 12613 4324 12617 4380
rect 12553 4320 12617 4324
rect 17994 4380 18058 4384
rect 17994 4324 17998 4380
rect 17998 4324 18054 4380
rect 18054 4324 18058 4380
rect 17994 4320 18058 4324
rect 18074 4380 18138 4384
rect 18074 4324 18078 4380
rect 18078 4324 18134 4380
rect 18134 4324 18138 4380
rect 18074 4320 18138 4324
rect 18154 4380 18218 4384
rect 18154 4324 18158 4380
rect 18158 4324 18214 4380
rect 18214 4324 18218 4380
rect 18154 4320 18218 4324
rect 18234 4380 18298 4384
rect 18234 4324 18238 4380
rect 18238 4324 18294 4380
rect 18294 4324 18298 4380
rect 18234 4320 18298 4324
rect 23675 4380 23739 4384
rect 23675 4324 23679 4380
rect 23679 4324 23735 4380
rect 23735 4324 23739 4380
rect 23675 4320 23739 4324
rect 23755 4380 23819 4384
rect 23755 4324 23759 4380
rect 23759 4324 23815 4380
rect 23815 4324 23819 4380
rect 23755 4320 23819 4324
rect 23835 4380 23899 4384
rect 23835 4324 23839 4380
rect 23839 4324 23895 4380
rect 23895 4324 23899 4380
rect 23835 4320 23899 4324
rect 23915 4380 23979 4384
rect 23915 4324 23919 4380
rect 23919 4324 23975 4380
rect 23975 4324 23979 4380
rect 23915 4320 23979 4324
rect 3792 3836 3856 3840
rect 3792 3780 3796 3836
rect 3796 3780 3852 3836
rect 3852 3780 3856 3836
rect 3792 3776 3856 3780
rect 3872 3836 3936 3840
rect 3872 3780 3876 3836
rect 3876 3780 3932 3836
rect 3932 3780 3936 3836
rect 3872 3776 3936 3780
rect 3952 3836 4016 3840
rect 3952 3780 3956 3836
rect 3956 3780 4012 3836
rect 4012 3780 4016 3836
rect 3952 3776 4016 3780
rect 4032 3836 4096 3840
rect 4032 3780 4036 3836
rect 4036 3780 4092 3836
rect 4092 3780 4096 3836
rect 4032 3776 4096 3780
rect 9473 3836 9537 3840
rect 9473 3780 9477 3836
rect 9477 3780 9533 3836
rect 9533 3780 9537 3836
rect 9473 3776 9537 3780
rect 9553 3836 9617 3840
rect 9553 3780 9557 3836
rect 9557 3780 9613 3836
rect 9613 3780 9617 3836
rect 9553 3776 9617 3780
rect 9633 3836 9697 3840
rect 9633 3780 9637 3836
rect 9637 3780 9693 3836
rect 9693 3780 9697 3836
rect 9633 3776 9697 3780
rect 9713 3836 9777 3840
rect 9713 3780 9717 3836
rect 9717 3780 9773 3836
rect 9773 3780 9777 3836
rect 9713 3776 9777 3780
rect 15154 3836 15218 3840
rect 15154 3780 15158 3836
rect 15158 3780 15214 3836
rect 15214 3780 15218 3836
rect 15154 3776 15218 3780
rect 15234 3836 15298 3840
rect 15234 3780 15238 3836
rect 15238 3780 15294 3836
rect 15294 3780 15298 3836
rect 15234 3776 15298 3780
rect 15314 3836 15378 3840
rect 15314 3780 15318 3836
rect 15318 3780 15374 3836
rect 15374 3780 15378 3836
rect 15314 3776 15378 3780
rect 15394 3836 15458 3840
rect 15394 3780 15398 3836
rect 15398 3780 15454 3836
rect 15454 3780 15458 3836
rect 15394 3776 15458 3780
rect 20835 3836 20899 3840
rect 20835 3780 20839 3836
rect 20839 3780 20895 3836
rect 20895 3780 20899 3836
rect 20835 3776 20899 3780
rect 20915 3836 20979 3840
rect 20915 3780 20919 3836
rect 20919 3780 20975 3836
rect 20975 3780 20979 3836
rect 20915 3776 20979 3780
rect 20995 3836 21059 3840
rect 20995 3780 20999 3836
rect 20999 3780 21055 3836
rect 21055 3780 21059 3836
rect 20995 3776 21059 3780
rect 21075 3836 21139 3840
rect 21075 3780 21079 3836
rect 21079 3780 21135 3836
rect 21135 3780 21139 3836
rect 21075 3776 21139 3780
rect 6632 3292 6696 3296
rect 6632 3236 6636 3292
rect 6636 3236 6692 3292
rect 6692 3236 6696 3292
rect 6632 3232 6696 3236
rect 6712 3292 6776 3296
rect 6712 3236 6716 3292
rect 6716 3236 6772 3292
rect 6772 3236 6776 3292
rect 6712 3232 6776 3236
rect 6792 3292 6856 3296
rect 6792 3236 6796 3292
rect 6796 3236 6852 3292
rect 6852 3236 6856 3292
rect 6792 3232 6856 3236
rect 6872 3292 6936 3296
rect 6872 3236 6876 3292
rect 6876 3236 6932 3292
rect 6932 3236 6936 3292
rect 6872 3232 6936 3236
rect 12313 3292 12377 3296
rect 12313 3236 12317 3292
rect 12317 3236 12373 3292
rect 12373 3236 12377 3292
rect 12313 3232 12377 3236
rect 12393 3292 12457 3296
rect 12393 3236 12397 3292
rect 12397 3236 12453 3292
rect 12453 3236 12457 3292
rect 12393 3232 12457 3236
rect 12473 3292 12537 3296
rect 12473 3236 12477 3292
rect 12477 3236 12533 3292
rect 12533 3236 12537 3292
rect 12473 3232 12537 3236
rect 12553 3292 12617 3296
rect 12553 3236 12557 3292
rect 12557 3236 12613 3292
rect 12613 3236 12617 3292
rect 12553 3232 12617 3236
rect 17994 3292 18058 3296
rect 17994 3236 17998 3292
rect 17998 3236 18054 3292
rect 18054 3236 18058 3292
rect 17994 3232 18058 3236
rect 18074 3292 18138 3296
rect 18074 3236 18078 3292
rect 18078 3236 18134 3292
rect 18134 3236 18138 3292
rect 18074 3232 18138 3236
rect 18154 3292 18218 3296
rect 18154 3236 18158 3292
rect 18158 3236 18214 3292
rect 18214 3236 18218 3292
rect 18154 3232 18218 3236
rect 18234 3292 18298 3296
rect 18234 3236 18238 3292
rect 18238 3236 18294 3292
rect 18294 3236 18298 3292
rect 18234 3232 18298 3236
rect 23675 3292 23739 3296
rect 23675 3236 23679 3292
rect 23679 3236 23735 3292
rect 23735 3236 23739 3292
rect 23675 3232 23739 3236
rect 23755 3292 23819 3296
rect 23755 3236 23759 3292
rect 23759 3236 23815 3292
rect 23815 3236 23819 3292
rect 23755 3232 23819 3236
rect 23835 3292 23899 3296
rect 23835 3236 23839 3292
rect 23839 3236 23895 3292
rect 23895 3236 23899 3292
rect 23835 3232 23899 3236
rect 23915 3292 23979 3296
rect 23915 3236 23919 3292
rect 23919 3236 23975 3292
rect 23975 3236 23979 3292
rect 23915 3232 23979 3236
rect 3792 2748 3856 2752
rect 3792 2692 3796 2748
rect 3796 2692 3852 2748
rect 3852 2692 3856 2748
rect 3792 2688 3856 2692
rect 3872 2748 3936 2752
rect 3872 2692 3876 2748
rect 3876 2692 3932 2748
rect 3932 2692 3936 2748
rect 3872 2688 3936 2692
rect 3952 2748 4016 2752
rect 3952 2692 3956 2748
rect 3956 2692 4012 2748
rect 4012 2692 4016 2748
rect 3952 2688 4016 2692
rect 4032 2748 4096 2752
rect 4032 2692 4036 2748
rect 4036 2692 4092 2748
rect 4092 2692 4096 2748
rect 4032 2688 4096 2692
rect 9473 2748 9537 2752
rect 9473 2692 9477 2748
rect 9477 2692 9533 2748
rect 9533 2692 9537 2748
rect 9473 2688 9537 2692
rect 9553 2748 9617 2752
rect 9553 2692 9557 2748
rect 9557 2692 9613 2748
rect 9613 2692 9617 2748
rect 9553 2688 9617 2692
rect 9633 2748 9697 2752
rect 9633 2692 9637 2748
rect 9637 2692 9693 2748
rect 9693 2692 9697 2748
rect 9633 2688 9697 2692
rect 9713 2748 9777 2752
rect 9713 2692 9717 2748
rect 9717 2692 9773 2748
rect 9773 2692 9777 2748
rect 9713 2688 9777 2692
rect 15154 2748 15218 2752
rect 15154 2692 15158 2748
rect 15158 2692 15214 2748
rect 15214 2692 15218 2748
rect 15154 2688 15218 2692
rect 15234 2748 15298 2752
rect 15234 2692 15238 2748
rect 15238 2692 15294 2748
rect 15294 2692 15298 2748
rect 15234 2688 15298 2692
rect 15314 2748 15378 2752
rect 15314 2692 15318 2748
rect 15318 2692 15374 2748
rect 15374 2692 15378 2748
rect 15314 2688 15378 2692
rect 15394 2748 15458 2752
rect 15394 2692 15398 2748
rect 15398 2692 15454 2748
rect 15454 2692 15458 2748
rect 15394 2688 15458 2692
rect 20835 2748 20899 2752
rect 20835 2692 20839 2748
rect 20839 2692 20895 2748
rect 20895 2692 20899 2748
rect 20835 2688 20899 2692
rect 20915 2748 20979 2752
rect 20915 2692 20919 2748
rect 20919 2692 20975 2748
rect 20975 2692 20979 2748
rect 20915 2688 20979 2692
rect 20995 2748 21059 2752
rect 20995 2692 20999 2748
rect 20999 2692 21055 2748
rect 21055 2692 21059 2748
rect 20995 2688 21059 2692
rect 21075 2748 21139 2752
rect 21075 2692 21079 2748
rect 21079 2692 21135 2748
rect 21135 2692 21139 2748
rect 21075 2688 21139 2692
rect 6632 2204 6696 2208
rect 6632 2148 6636 2204
rect 6636 2148 6692 2204
rect 6692 2148 6696 2204
rect 6632 2144 6696 2148
rect 6712 2204 6776 2208
rect 6712 2148 6716 2204
rect 6716 2148 6772 2204
rect 6772 2148 6776 2204
rect 6712 2144 6776 2148
rect 6792 2204 6856 2208
rect 6792 2148 6796 2204
rect 6796 2148 6852 2204
rect 6852 2148 6856 2204
rect 6792 2144 6856 2148
rect 6872 2204 6936 2208
rect 6872 2148 6876 2204
rect 6876 2148 6932 2204
rect 6932 2148 6936 2204
rect 6872 2144 6936 2148
rect 12313 2204 12377 2208
rect 12313 2148 12317 2204
rect 12317 2148 12373 2204
rect 12373 2148 12377 2204
rect 12313 2144 12377 2148
rect 12393 2204 12457 2208
rect 12393 2148 12397 2204
rect 12397 2148 12453 2204
rect 12453 2148 12457 2204
rect 12393 2144 12457 2148
rect 12473 2204 12537 2208
rect 12473 2148 12477 2204
rect 12477 2148 12533 2204
rect 12533 2148 12537 2204
rect 12473 2144 12537 2148
rect 12553 2204 12617 2208
rect 12553 2148 12557 2204
rect 12557 2148 12613 2204
rect 12613 2148 12617 2204
rect 12553 2144 12617 2148
rect 17994 2204 18058 2208
rect 17994 2148 17998 2204
rect 17998 2148 18054 2204
rect 18054 2148 18058 2204
rect 17994 2144 18058 2148
rect 18074 2204 18138 2208
rect 18074 2148 18078 2204
rect 18078 2148 18134 2204
rect 18134 2148 18138 2204
rect 18074 2144 18138 2148
rect 18154 2204 18218 2208
rect 18154 2148 18158 2204
rect 18158 2148 18214 2204
rect 18214 2148 18218 2204
rect 18154 2144 18218 2148
rect 18234 2204 18298 2208
rect 18234 2148 18238 2204
rect 18238 2148 18294 2204
rect 18294 2148 18298 2204
rect 18234 2144 18298 2148
rect 23675 2204 23739 2208
rect 23675 2148 23679 2204
rect 23679 2148 23735 2204
rect 23735 2148 23739 2204
rect 23675 2144 23739 2148
rect 23755 2204 23819 2208
rect 23755 2148 23759 2204
rect 23759 2148 23815 2204
rect 23815 2148 23819 2204
rect 23755 2144 23819 2148
rect 23835 2204 23899 2208
rect 23835 2148 23839 2204
rect 23839 2148 23895 2204
rect 23895 2148 23899 2204
rect 23835 2144 23899 2148
rect 23915 2204 23979 2208
rect 23915 2148 23919 2204
rect 23919 2148 23975 2204
rect 23975 2148 23979 2204
rect 23915 2144 23979 2148
<< metal4 >>
rect 3784 22336 4104 22352
rect 3784 22272 3792 22336
rect 3856 22272 3872 22336
rect 3936 22272 3952 22336
rect 4016 22272 4032 22336
rect 4096 22272 4104 22336
rect 3784 21248 4104 22272
rect 3784 21184 3792 21248
rect 3856 21184 3872 21248
rect 3936 21184 3952 21248
rect 4016 21184 4032 21248
rect 4096 21184 4104 21248
rect 3784 20160 4104 21184
rect 3784 20096 3792 20160
rect 3856 20096 3872 20160
rect 3936 20096 3952 20160
rect 4016 20096 4032 20160
rect 4096 20096 4104 20160
rect 3784 19072 4104 20096
rect 3784 19008 3792 19072
rect 3856 19008 3872 19072
rect 3936 19008 3952 19072
rect 4016 19008 4032 19072
rect 4096 19008 4104 19072
rect 3784 17984 4104 19008
rect 3784 17920 3792 17984
rect 3856 17920 3872 17984
rect 3936 17920 3952 17984
rect 4016 17920 4032 17984
rect 4096 17920 4104 17984
rect 3784 16896 4104 17920
rect 3784 16832 3792 16896
rect 3856 16832 3872 16896
rect 3936 16832 3952 16896
rect 4016 16832 4032 16896
rect 4096 16832 4104 16896
rect 3784 15808 4104 16832
rect 3784 15744 3792 15808
rect 3856 15744 3872 15808
rect 3936 15744 3952 15808
rect 4016 15744 4032 15808
rect 4096 15744 4104 15808
rect 3784 14720 4104 15744
rect 6624 21792 6944 22352
rect 6624 21728 6632 21792
rect 6696 21728 6712 21792
rect 6776 21728 6792 21792
rect 6856 21728 6872 21792
rect 6936 21728 6944 21792
rect 6624 20704 6944 21728
rect 6624 20640 6632 20704
rect 6696 20640 6712 20704
rect 6776 20640 6792 20704
rect 6856 20640 6872 20704
rect 6936 20640 6944 20704
rect 6624 19616 6944 20640
rect 6624 19552 6632 19616
rect 6696 19552 6712 19616
rect 6776 19552 6792 19616
rect 6856 19552 6872 19616
rect 6936 19552 6944 19616
rect 6624 18528 6944 19552
rect 6624 18464 6632 18528
rect 6696 18464 6712 18528
rect 6776 18464 6792 18528
rect 6856 18464 6872 18528
rect 6936 18464 6944 18528
rect 6624 17440 6944 18464
rect 6624 17376 6632 17440
rect 6696 17376 6712 17440
rect 6776 17376 6792 17440
rect 6856 17376 6872 17440
rect 6936 17376 6944 17440
rect 6624 16352 6944 17376
rect 6624 16288 6632 16352
rect 6696 16288 6712 16352
rect 6776 16288 6792 16352
rect 6856 16288 6872 16352
rect 6936 16288 6944 16352
rect 5395 15332 5461 15333
rect 5395 15268 5396 15332
rect 5460 15268 5461 15332
rect 5395 15267 5461 15268
rect 3784 14656 3792 14720
rect 3856 14656 3872 14720
rect 3936 14656 3952 14720
rect 4016 14656 4032 14720
rect 4096 14656 4104 14720
rect 3784 13632 4104 14656
rect 3784 13568 3792 13632
rect 3856 13568 3872 13632
rect 3936 13568 3952 13632
rect 4016 13568 4032 13632
rect 4096 13568 4104 13632
rect 3784 12544 4104 13568
rect 3784 12480 3792 12544
rect 3856 12480 3872 12544
rect 3936 12480 3952 12544
rect 4016 12480 4032 12544
rect 4096 12480 4104 12544
rect 3784 11456 4104 12480
rect 3784 11392 3792 11456
rect 3856 11392 3872 11456
rect 3936 11392 3952 11456
rect 4016 11392 4032 11456
rect 4096 11392 4104 11456
rect 3784 10368 4104 11392
rect 5398 10709 5458 15267
rect 6624 15264 6944 16288
rect 6624 15200 6632 15264
rect 6696 15200 6712 15264
rect 6776 15200 6792 15264
rect 6856 15200 6872 15264
rect 6936 15200 6944 15264
rect 6624 14176 6944 15200
rect 6624 14112 6632 14176
rect 6696 14112 6712 14176
rect 6776 14112 6792 14176
rect 6856 14112 6872 14176
rect 6936 14112 6944 14176
rect 6624 13088 6944 14112
rect 6624 13024 6632 13088
rect 6696 13024 6712 13088
rect 6776 13024 6792 13088
rect 6856 13024 6872 13088
rect 6936 13024 6944 13088
rect 6624 12000 6944 13024
rect 6624 11936 6632 12000
rect 6696 11936 6712 12000
rect 6776 11936 6792 12000
rect 6856 11936 6872 12000
rect 6936 11936 6944 12000
rect 6624 10912 6944 11936
rect 6624 10848 6632 10912
rect 6696 10848 6712 10912
rect 6776 10848 6792 10912
rect 6856 10848 6872 10912
rect 6936 10848 6944 10912
rect 5395 10708 5461 10709
rect 5395 10644 5396 10708
rect 5460 10644 5461 10708
rect 5395 10643 5461 10644
rect 3784 10304 3792 10368
rect 3856 10304 3872 10368
rect 3936 10304 3952 10368
rect 4016 10304 4032 10368
rect 4096 10304 4104 10368
rect 3784 9280 4104 10304
rect 3784 9216 3792 9280
rect 3856 9216 3872 9280
rect 3936 9216 3952 9280
rect 4016 9216 4032 9280
rect 4096 9216 4104 9280
rect 3784 8192 4104 9216
rect 3784 8128 3792 8192
rect 3856 8128 3872 8192
rect 3936 8128 3952 8192
rect 4016 8128 4032 8192
rect 4096 8128 4104 8192
rect 3784 7104 4104 8128
rect 3784 7040 3792 7104
rect 3856 7040 3872 7104
rect 3936 7040 3952 7104
rect 4016 7040 4032 7104
rect 4096 7040 4104 7104
rect 3784 6016 4104 7040
rect 3784 5952 3792 6016
rect 3856 5952 3872 6016
rect 3936 5952 3952 6016
rect 4016 5952 4032 6016
rect 4096 5952 4104 6016
rect 3784 4928 4104 5952
rect 3784 4864 3792 4928
rect 3856 4864 3872 4928
rect 3936 4864 3952 4928
rect 4016 4864 4032 4928
rect 4096 4864 4104 4928
rect 3784 3840 4104 4864
rect 3784 3776 3792 3840
rect 3856 3776 3872 3840
rect 3936 3776 3952 3840
rect 4016 3776 4032 3840
rect 4096 3776 4104 3840
rect 3784 2752 4104 3776
rect 3784 2688 3792 2752
rect 3856 2688 3872 2752
rect 3936 2688 3952 2752
rect 4016 2688 4032 2752
rect 4096 2688 4104 2752
rect 3784 2128 4104 2688
rect 6624 9824 6944 10848
rect 9465 22336 9785 22352
rect 9465 22272 9473 22336
rect 9537 22272 9553 22336
rect 9617 22272 9633 22336
rect 9697 22272 9713 22336
rect 9777 22272 9785 22336
rect 9465 21248 9785 22272
rect 9465 21184 9473 21248
rect 9537 21184 9553 21248
rect 9617 21184 9633 21248
rect 9697 21184 9713 21248
rect 9777 21184 9785 21248
rect 9465 20160 9785 21184
rect 9465 20096 9473 20160
rect 9537 20096 9553 20160
rect 9617 20096 9633 20160
rect 9697 20096 9713 20160
rect 9777 20096 9785 20160
rect 9465 19072 9785 20096
rect 9465 19008 9473 19072
rect 9537 19008 9553 19072
rect 9617 19008 9633 19072
rect 9697 19008 9713 19072
rect 9777 19008 9785 19072
rect 9465 17984 9785 19008
rect 9465 17920 9473 17984
rect 9537 17920 9553 17984
rect 9617 17920 9633 17984
rect 9697 17920 9713 17984
rect 9777 17920 9785 17984
rect 9465 16896 9785 17920
rect 9465 16832 9473 16896
rect 9537 16832 9553 16896
rect 9617 16832 9633 16896
rect 9697 16832 9713 16896
rect 9777 16832 9785 16896
rect 9465 15808 9785 16832
rect 9465 15744 9473 15808
rect 9537 15744 9553 15808
rect 9617 15744 9633 15808
rect 9697 15744 9713 15808
rect 9777 15744 9785 15808
rect 9465 14720 9785 15744
rect 9465 14656 9473 14720
rect 9537 14656 9553 14720
rect 9617 14656 9633 14720
rect 9697 14656 9713 14720
rect 9777 14656 9785 14720
rect 9465 13632 9785 14656
rect 9465 13568 9473 13632
rect 9537 13568 9553 13632
rect 9617 13568 9633 13632
rect 9697 13568 9713 13632
rect 9777 13568 9785 13632
rect 9465 12544 9785 13568
rect 9465 12480 9473 12544
rect 9537 12480 9553 12544
rect 9617 12480 9633 12544
rect 9697 12480 9713 12544
rect 9777 12480 9785 12544
rect 9465 11456 9785 12480
rect 9465 11392 9473 11456
rect 9537 11392 9553 11456
rect 9617 11392 9633 11456
rect 9697 11392 9713 11456
rect 9777 11392 9785 11456
rect 7235 10572 7301 10573
rect 7235 10508 7236 10572
rect 7300 10508 7301 10572
rect 7235 10507 7301 10508
rect 6624 9760 6632 9824
rect 6696 9760 6712 9824
rect 6776 9760 6792 9824
rect 6856 9760 6872 9824
rect 6936 9760 6944 9824
rect 6624 8736 6944 9760
rect 6624 8672 6632 8736
rect 6696 8672 6712 8736
rect 6776 8672 6792 8736
rect 6856 8672 6872 8736
rect 6936 8672 6944 8736
rect 6624 7648 6944 8672
rect 6624 7584 6632 7648
rect 6696 7584 6712 7648
rect 6776 7584 6792 7648
rect 6856 7584 6872 7648
rect 6936 7584 6944 7648
rect 6624 6560 6944 7584
rect 6624 6496 6632 6560
rect 6696 6496 6712 6560
rect 6776 6496 6792 6560
rect 6856 6496 6872 6560
rect 6936 6496 6944 6560
rect 6624 5472 6944 6496
rect 6624 5408 6632 5472
rect 6696 5408 6712 5472
rect 6776 5408 6792 5472
rect 6856 5408 6872 5472
rect 6936 5408 6944 5472
rect 6624 4384 6944 5408
rect 7238 5133 7298 10507
rect 9465 10368 9785 11392
rect 9465 10304 9473 10368
rect 9537 10304 9553 10368
rect 9617 10304 9633 10368
rect 9697 10304 9713 10368
rect 9777 10304 9785 10368
rect 9465 9280 9785 10304
rect 12305 21792 12625 22352
rect 12305 21728 12313 21792
rect 12377 21728 12393 21792
rect 12457 21728 12473 21792
rect 12537 21728 12553 21792
rect 12617 21728 12625 21792
rect 12305 20704 12625 21728
rect 15146 22336 15466 22352
rect 15146 22272 15154 22336
rect 15218 22272 15234 22336
rect 15298 22272 15314 22336
rect 15378 22272 15394 22336
rect 15458 22272 15466 22336
rect 15146 21248 15466 22272
rect 15146 21184 15154 21248
rect 15218 21184 15234 21248
rect 15298 21184 15314 21248
rect 15378 21184 15394 21248
rect 15458 21184 15466 21248
rect 13123 20772 13189 20773
rect 13123 20708 13124 20772
rect 13188 20708 13189 20772
rect 13123 20707 13189 20708
rect 14779 20772 14845 20773
rect 14779 20708 14780 20772
rect 14844 20708 14845 20772
rect 14779 20707 14845 20708
rect 12305 20640 12313 20704
rect 12377 20640 12393 20704
rect 12457 20640 12473 20704
rect 12537 20640 12553 20704
rect 12617 20640 12625 20704
rect 12305 19616 12625 20640
rect 12305 19552 12313 19616
rect 12377 19552 12393 19616
rect 12457 19552 12473 19616
rect 12537 19552 12553 19616
rect 12617 19552 12625 19616
rect 12305 18528 12625 19552
rect 12305 18464 12313 18528
rect 12377 18464 12393 18528
rect 12457 18464 12473 18528
rect 12537 18464 12553 18528
rect 12617 18464 12625 18528
rect 12305 17440 12625 18464
rect 12305 17376 12313 17440
rect 12377 17376 12393 17440
rect 12457 17376 12473 17440
rect 12537 17376 12553 17440
rect 12617 17376 12625 17440
rect 12305 16352 12625 17376
rect 12305 16288 12313 16352
rect 12377 16288 12393 16352
rect 12457 16288 12473 16352
rect 12537 16288 12553 16352
rect 12617 16288 12625 16352
rect 12305 15264 12625 16288
rect 12305 15200 12313 15264
rect 12377 15200 12393 15264
rect 12457 15200 12473 15264
rect 12537 15200 12553 15264
rect 12617 15200 12625 15264
rect 12305 14176 12625 15200
rect 12305 14112 12313 14176
rect 12377 14112 12393 14176
rect 12457 14112 12473 14176
rect 12537 14112 12553 14176
rect 12617 14112 12625 14176
rect 12305 13088 12625 14112
rect 12305 13024 12313 13088
rect 12377 13024 12393 13088
rect 12457 13024 12473 13088
rect 12537 13024 12553 13088
rect 12617 13024 12625 13088
rect 12305 12000 12625 13024
rect 13126 12341 13186 20707
rect 13123 12340 13189 12341
rect 13123 12276 13124 12340
rect 13188 12276 13189 12340
rect 13123 12275 13189 12276
rect 12305 11936 12313 12000
rect 12377 11936 12393 12000
rect 12457 11936 12473 12000
rect 12537 11936 12553 12000
rect 12617 11936 12625 12000
rect 12305 10912 12625 11936
rect 14782 11797 14842 20707
rect 15146 20160 15466 21184
rect 15146 20096 15154 20160
rect 15218 20096 15234 20160
rect 15298 20096 15314 20160
rect 15378 20096 15394 20160
rect 15458 20096 15466 20160
rect 15146 19072 15466 20096
rect 17986 21792 18306 22352
rect 17986 21728 17994 21792
rect 18058 21728 18074 21792
rect 18138 21728 18154 21792
rect 18218 21728 18234 21792
rect 18298 21728 18306 21792
rect 17986 20704 18306 21728
rect 17986 20640 17994 20704
rect 18058 20640 18074 20704
rect 18138 20640 18154 20704
rect 18218 20640 18234 20704
rect 18298 20640 18306 20704
rect 17986 19616 18306 20640
rect 17986 19552 17994 19616
rect 18058 19552 18074 19616
rect 18138 19552 18154 19616
rect 18218 19552 18234 19616
rect 18298 19552 18306 19616
rect 17723 19412 17789 19413
rect 17723 19348 17724 19412
rect 17788 19348 17789 19412
rect 17723 19347 17789 19348
rect 15146 19008 15154 19072
rect 15218 19008 15234 19072
rect 15298 19008 15314 19072
rect 15378 19008 15394 19072
rect 15458 19008 15466 19072
rect 15146 17984 15466 19008
rect 16435 18052 16501 18053
rect 16435 17988 16436 18052
rect 16500 17988 16501 18052
rect 16435 17987 16501 17988
rect 15146 17920 15154 17984
rect 15218 17920 15234 17984
rect 15298 17920 15314 17984
rect 15378 17920 15394 17984
rect 15458 17920 15466 17984
rect 15146 16896 15466 17920
rect 15146 16832 15154 16896
rect 15218 16832 15234 16896
rect 15298 16832 15314 16896
rect 15378 16832 15394 16896
rect 15458 16832 15466 16896
rect 15146 15808 15466 16832
rect 15146 15744 15154 15808
rect 15218 15744 15234 15808
rect 15298 15744 15314 15808
rect 15378 15744 15394 15808
rect 15458 15744 15466 15808
rect 15146 14720 15466 15744
rect 15146 14656 15154 14720
rect 15218 14656 15234 14720
rect 15298 14656 15314 14720
rect 15378 14656 15394 14720
rect 15458 14656 15466 14720
rect 15146 13632 15466 14656
rect 16438 14653 16498 17987
rect 16435 14652 16501 14653
rect 16435 14588 16436 14652
rect 16500 14588 16501 14652
rect 16435 14587 16501 14588
rect 16251 13836 16317 13837
rect 16251 13772 16252 13836
rect 16316 13772 16317 13836
rect 16251 13771 16317 13772
rect 15146 13568 15154 13632
rect 15218 13568 15234 13632
rect 15298 13568 15314 13632
rect 15378 13568 15394 13632
rect 15458 13568 15466 13632
rect 15146 12544 15466 13568
rect 15146 12480 15154 12544
rect 15218 12480 15234 12544
rect 15298 12480 15314 12544
rect 15378 12480 15394 12544
rect 15458 12480 15466 12544
rect 14779 11796 14845 11797
rect 14779 11732 14780 11796
rect 14844 11732 14845 11796
rect 14779 11731 14845 11732
rect 12305 10848 12313 10912
rect 12377 10848 12393 10912
rect 12457 10848 12473 10912
rect 12537 10848 12553 10912
rect 12617 10848 12625 10912
rect 10363 9892 10429 9893
rect 10363 9828 10364 9892
rect 10428 9828 10429 9892
rect 10363 9827 10429 9828
rect 9465 9216 9473 9280
rect 9537 9216 9553 9280
rect 9617 9216 9633 9280
rect 9697 9216 9713 9280
rect 9777 9216 9785 9280
rect 9465 8192 9785 9216
rect 9465 8128 9473 8192
rect 9537 8128 9553 8192
rect 9617 8128 9633 8192
rect 9697 8128 9713 8192
rect 9777 8128 9785 8192
rect 9465 7104 9785 8128
rect 9465 7040 9473 7104
rect 9537 7040 9553 7104
rect 9617 7040 9633 7104
rect 9697 7040 9713 7104
rect 9777 7040 9785 7104
rect 9465 6016 9785 7040
rect 9465 5952 9473 6016
rect 9537 5952 9553 6016
rect 9617 5952 9633 6016
rect 9697 5952 9713 6016
rect 9777 5952 9785 6016
rect 7235 5132 7301 5133
rect 7235 5068 7236 5132
rect 7300 5068 7301 5132
rect 7235 5067 7301 5068
rect 6624 4320 6632 4384
rect 6696 4320 6712 4384
rect 6776 4320 6792 4384
rect 6856 4320 6872 4384
rect 6936 4320 6944 4384
rect 6624 3296 6944 4320
rect 6624 3232 6632 3296
rect 6696 3232 6712 3296
rect 6776 3232 6792 3296
rect 6856 3232 6872 3296
rect 6936 3232 6944 3296
rect 6624 2208 6944 3232
rect 6624 2144 6632 2208
rect 6696 2144 6712 2208
rect 6776 2144 6792 2208
rect 6856 2144 6872 2208
rect 6936 2144 6944 2208
rect 6624 2128 6944 2144
rect 9465 4928 9785 5952
rect 10366 5541 10426 9827
rect 12305 9824 12625 10848
rect 12305 9760 12313 9824
rect 12377 9760 12393 9824
rect 12457 9760 12473 9824
rect 12537 9760 12553 9824
rect 12617 9760 12625 9824
rect 12305 8736 12625 9760
rect 12305 8672 12313 8736
rect 12377 8672 12393 8736
rect 12457 8672 12473 8736
rect 12537 8672 12553 8736
rect 12617 8672 12625 8736
rect 12305 7648 12625 8672
rect 12305 7584 12313 7648
rect 12377 7584 12393 7648
rect 12457 7584 12473 7648
rect 12537 7584 12553 7648
rect 12617 7584 12625 7648
rect 12305 6560 12625 7584
rect 12305 6496 12313 6560
rect 12377 6496 12393 6560
rect 12457 6496 12473 6560
rect 12537 6496 12553 6560
rect 12617 6496 12625 6560
rect 10363 5540 10429 5541
rect 10363 5476 10364 5540
rect 10428 5476 10429 5540
rect 10363 5475 10429 5476
rect 9465 4864 9473 4928
rect 9537 4864 9553 4928
rect 9617 4864 9633 4928
rect 9697 4864 9713 4928
rect 9777 4864 9785 4928
rect 9465 3840 9785 4864
rect 9465 3776 9473 3840
rect 9537 3776 9553 3840
rect 9617 3776 9633 3840
rect 9697 3776 9713 3840
rect 9777 3776 9785 3840
rect 9465 2752 9785 3776
rect 9465 2688 9473 2752
rect 9537 2688 9553 2752
rect 9617 2688 9633 2752
rect 9697 2688 9713 2752
rect 9777 2688 9785 2752
rect 9465 2128 9785 2688
rect 12305 5472 12625 6496
rect 12305 5408 12313 5472
rect 12377 5408 12393 5472
rect 12457 5408 12473 5472
rect 12537 5408 12553 5472
rect 12617 5408 12625 5472
rect 12305 4384 12625 5408
rect 12305 4320 12313 4384
rect 12377 4320 12393 4384
rect 12457 4320 12473 4384
rect 12537 4320 12553 4384
rect 12617 4320 12625 4384
rect 12305 3296 12625 4320
rect 12305 3232 12313 3296
rect 12377 3232 12393 3296
rect 12457 3232 12473 3296
rect 12537 3232 12553 3296
rect 12617 3232 12625 3296
rect 12305 2208 12625 3232
rect 12305 2144 12313 2208
rect 12377 2144 12393 2208
rect 12457 2144 12473 2208
rect 12537 2144 12553 2208
rect 12617 2144 12625 2208
rect 12305 2128 12625 2144
rect 15146 11456 15466 12480
rect 15146 11392 15154 11456
rect 15218 11392 15234 11456
rect 15298 11392 15314 11456
rect 15378 11392 15394 11456
rect 15458 11392 15466 11456
rect 15146 10368 15466 11392
rect 15146 10304 15154 10368
rect 15218 10304 15234 10368
rect 15298 10304 15314 10368
rect 15378 10304 15394 10368
rect 15458 10304 15466 10368
rect 15146 9280 15466 10304
rect 15146 9216 15154 9280
rect 15218 9216 15234 9280
rect 15298 9216 15314 9280
rect 15378 9216 15394 9280
rect 15458 9216 15466 9280
rect 15146 8192 15466 9216
rect 16254 8397 16314 13771
rect 17726 13565 17786 19347
rect 17986 18528 18306 19552
rect 17986 18464 17994 18528
rect 18058 18464 18074 18528
rect 18138 18464 18154 18528
rect 18218 18464 18234 18528
rect 18298 18464 18306 18528
rect 17986 17440 18306 18464
rect 17986 17376 17994 17440
rect 18058 17376 18074 17440
rect 18138 17376 18154 17440
rect 18218 17376 18234 17440
rect 18298 17376 18306 17440
rect 17986 16352 18306 17376
rect 17986 16288 17994 16352
rect 18058 16288 18074 16352
rect 18138 16288 18154 16352
rect 18218 16288 18234 16352
rect 18298 16288 18306 16352
rect 17986 15264 18306 16288
rect 17986 15200 17994 15264
rect 18058 15200 18074 15264
rect 18138 15200 18154 15264
rect 18218 15200 18234 15264
rect 18298 15200 18306 15264
rect 17986 14176 18306 15200
rect 17986 14112 17994 14176
rect 18058 14112 18074 14176
rect 18138 14112 18154 14176
rect 18218 14112 18234 14176
rect 18298 14112 18306 14176
rect 17723 13564 17789 13565
rect 17723 13500 17724 13564
rect 17788 13500 17789 13564
rect 17723 13499 17789 13500
rect 17986 13088 18306 14112
rect 17986 13024 17994 13088
rect 18058 13024 18074 13088
rect 18138 13024 18154 13088
rect 18218 13024 18234 13088
rect 18298 13024 18306 13088
rect 17986 12000 18306 13024
rect 17986 11936 17994 12000
rect 18058 11936 18074 12000
rect 18138 11936 18154 12000
rect 18218 11936 18234 12000
rect 18298 11936 18306 12000
rect 17986 10912 18306 11936
rect 17986 10848 17994 10912
rect 18058 10848 18074 10912
rect 18138 10848 18154 10912
rect 18218 10848 18234 10912
rect 18298 10848 18306 10912
rect 17723 10028 17789 10029
rect 17723 9964 17724 10028
rect 17788 9964 17789 10028
rect 17723 9963 17789 9964
rect 16251 8396 16317 8397
rect 16251 8332 16252 8396
rect 16316 8332 16317 8396
rect 16251 8331 16317 8332
rect 15146 8128 15154 8192
rect 15218 8128 15234 8192
rect 15298 8128 15314 8192
rect 15378 8128 15394 8192
rect 15458 8128 15466 8192
rect 15146 7104 15466 8128
rect 15146 7040 15154 7104
rect 15218 7040 15234 7104
rect 15298 7040 15314 7104
rect 15378 7040 15394 7104
rect 15458 7040 15466 7104
rect 15146 6016 15466 7040
rect 15146 5952 15154 6016
rect 15218 5952 15234 6016
rect 15298 5952 15314 6016
rect 15378 5952 15394 6016
rect 15458 5952 15466 6016
rect 15146 4928 15466 5952
rect 15146 4864 15154 4928
rect 15218 4864 15234 4928
rect 15298 4864 15314 4928
rect 15378 4864 15394 4928
rect 15458 4864 15466 4928
rect 15146 3840 15466 4864
rect 17726 4725 17786 9963
rect 17986 9824 18306 10848
rect 17986 9760 17994 9824
rect 18058 9760 18074 9824
rect 18138 9760 18154 9824
rect 18218 9760 18234 9824
rect 18298 9760 18306 9824
rect 17986 8736 18306 9760
rect 17986 8672 17994 8736
rect 18058 8672 18074 8736
rect 18138 8672 18154 8736
rect 18218 8672 18234 8736
rect 18298 8672 18306 8736
rect 17986 7648 18306 8672
rect 17986 7584 17994 7648
rect 18058 7584 18074 7648
rect 18138 7584 18154 7648
rect 18218 7584 18234 7648
rect 18298 7584 18306 7648
rect 17986 6560 18306 7584
rect 17986 6496 17994 6560
rect 18058 6496 18074 6560
rect 18138 6496 18154 6560
rect 18218 6496 18234 6560
rect 18298 6496 18306 6560
rect 17986 5472 18306 6496
rect 17986 5408 17994 5472
rect 18058 5408 18074 5472
rect 18138 5408 18154 5472
rect 18218 5408 18234 5472
rect 18298 5408 18306 5472
rect 17723 4724 17789 4725
rect 17723 4660 17724 4724
rect 17788 4660 17789 4724
rect 17723 4659 17789 4660
rect 15146 3776 15154 3840
rect 15218 3776 15234 3840
rect 15298 3776 15314 3840
rect 15378 3776 15394 3840
rect 15458 3776 15466 3840
rect 15146 2752 15466 3776
rect 15146 2688 15154 2752
rect 15218 2688 15234 2752
rect 15298 2688 15314 2752
rect 15378 2688 15394 2752
rect 15458 2688 15466 2752
rect 15146 2128 15466 2688
rect 17986 4384 18306 5408
rect 17986 4320 17994 4384
rect 18058 4320 18074 4384
rect 18138 4320 18154 4384
rect 18218 4320 18234 4384
rect 18298 4320 18306 4384
rect 17986 3296 18306 4320
rect 17986 3232 17994 3296
rect 18058 3232 18074 3296
rect 18138 3232 18154 3296
rect 18218 3232 18234 3296
rect 18298 3232 18306 3296
rect 17986 2208 18306 3232
rect 17986 2144 17994 2208
rect 18058 2144 18074 2208
rect 18138 2144 18154 2208
rect 18218 2144 18234 2208
rect 18298 2144 18306 2208
rect 17986 2128 18306 2144
rect 20827 22336 21147 22352
rect 20827 22272 20835 22336
rect 20899 22272 20915 22336
rect 20979 22272 20995 22336
rect 21059 22272 21075 22336
rect 21139 22272 21147 22336
rect 20827 21248 21147 22272
rect 20827 21184 20835 21248
rect 20899 21184 20915 21248
rect 20979 21184 20995 21248
rect 21059 21184 21075 21248
rect 21139 21184 21147 21248
rect 20827 20160 21147 21184
rect 20827 20096 20835 20160
rect 20899 20096 20915 20160
rect 20979 20096 20995 20160
rect 21059 20096 21075 20160
rect 21139 20096 21147 20160
rect 20827 19072 21147 20096
rect 20827 19008 20835 19072
rect 20899 19008 20915 19072
rect 20979 19008 20995 19072
rect 21059 19008 21075 19072
rect 21139 19008 21147 19072
rect 20827 17984 21147 19008
rect 23667 21792 23987 22352
rect 23667 21728 23675 21792
rect 23739 21728 23755 21792
rect 23819 21728 23835 21792
rect 23899 21728 23915 21792
rect 23979 21728 23987 21792
rect 23667 20704 23987 21728
rect 23667 20640 23675 20704
rect 23739 20640 23755 20704
rect 23819 20640 23835 20704
rect 23899 20640 23915 20704
rect 23979 20640 23987 20704
rect 23667 19616 23987 20640
rect 23667 19552 23675 19616
rect 23739 19552 23755 19616
rect 23819 19552 23835 19616
rect 23899 19552 23915 19616
rect 23979 19552 23987 19616
rect 23667 18528 23987 19552
rect 23667 18464 23675 18528
rect 23739 18464 23755 18528
rect 23819 18464 23835 18528
rect 23899 18464 23915 18528
rect 23979 18464 23987 18528
rect 21403 18188 21469 18189
rect 21403 18124 21404 18188
rect 21468 18124 21469 18188
rect 21403 18123 21469 18124
rect 20827 17920 20835 17984
rect 20899 17920 20915 17984
rect 20979 17920 20995 17984
rect 21059 17920 21075 17984
rect 21139 17920 21147 17984
rect 20827 16896 21147 17920
rect 20827 16832 20835 16896
rect 20899 16832 20915 16896
rect 20979 16832 20995 16896
rect 21059 16832 21075 16896
rect 21139 16832 21147 16896
rect 20827 15808 21147 16832
rect 20827 15744 20835 15808
rect 20899 15744 20915 15808
rect 20979 15744 20995 15808
rect 21059 15744 21075 15808
rect 21139 15744 21147 15808
rect 20827 14720 21147 15744
rect 20827 14656 20835 14720
rect 20899 14656 20915 14720
rect 20979 14656 20995 14720
rect 21059 14656 21075 14720
rect 21139 14656 21147 14720
rect 20827 13632 21147 14656
rect 20827 13568 20835 13632
rect 20899 13568 20915 13632
rect 20979 13568 20995 13632
rect 21059 13568 21075 13632
rect 21139 13568 21147 13632
rect 20827 12544 21147 13568
rect 20827 12480 20835 12544
rect 20899 12480 20915 12544
rect 20979 12480 20995 12544
rect 21059 12480 21075 12544
rect 21139 12480 21147 12544
rect 20827 11456 21147 12480
rect 20827 11392 20835 11456
rect 20899 11392 20915 11456
rect 20979 11392 20995 11456
rect 21059 11392 21075 11456
rect 21139 11392 21147 11456
rect 20827 10368 21147 11392
rect 20827 10304 20835 10368
rect 20899 10304 20915 10368
rect 20979 10304 20995 10368
rect 21059 10304 21075 10368
rect 21139 10304 21147 10368
rect 20827 9280 21147 10304
rect 20827 9216 20835 9280
rect 20899 9216 20915 9280
rect 20979 9216 20995 9280
rect 21059 9216 21075 9280
rect 21139 9216 21147 9280
rect 20827 8192 21147 9216
rect 20827 8128 20835 8192
rect 20899 8128 20915 8192
rect 20979 8128 20995 8192
rect 21059 8128 21075 8192
rect 21139 8128 21147 8192
rect 20827 7104 21147 8128
rect 20827 7040 20835 7104
rect 20899 7040 20915 7104
rect 20979 7040 20995 7104
rect 21059 7040 21075 7104
rect 21139 7040 21147 7104
rect 20827 6016 21147 7040
rect 21406 6901 21466 18123
rect 23667 17440 23987 18464
rect 23667 17376 23675 17440
rect 23739 17376 23755 17440
rect 23819 17376 23835 17440
rect 23899 17376 23915 17440
rect 23979 17376 23987 17440
rect 23667 16352 23987 17376
rect 23667 16288 23675 16352
rect 23739 16288 23755 16352
rect 23819 16288 23835 16352
rect 23899 16288 23915 16352
rect 23979 16288 23987 16352
rect 23667 15264 23987 16288
rect 23667 15200 23675 15264
rect 23739 15200 23755 15264
rect 23819 15200 23835 15264
rect 23899 15200 23915 15264
rect 23979 15200 23987 15264
rect 23667 14176 23987 15200
rect 23667 14112 23675 14176
rect 23739 14112 23755 14176
rect 23819 14112 23835 14176
rect 23899 14112 23915 14176
rect 23979 14112 23987 14176
rect 22323 13836 22389 13837
rect 22323 13772 22324 13836
rect 22388 13772 22389 13836
rect 22323 13771 22389 13772
rect 22326 10709 22386 13771
rect 23667 13088 23987 14112
rect 23667 13024 23675 13088
rect 23739 13024 23755 13088
rect 23819 13024 23835 13088
rect 23899 13024 23915 13088
rect 23979 13024 23987 13088
rect 23667 12000 23987 13024
rect 23667 11936 23675 12000
rect 23739 11936 23755 12000
rect 23819 11936 23835 12000
rect 23899 11936 23915 12000
rect 23979 11936 23987 12000
rect 23667 10912 23987 11936
rect 23667 10848 23675 10912
rect 23739 10848 23755 10912
rect 23819 10848 23835 10912
rect 23899 10848 23915 10912
rect 23979 10848 23987 10912
rect 22323 10708 22389 10709
rect 22323 10644 22324 10708
rect 22388 10644 22389 10708
rect 22323 10643 22389 10644
rect 23667 9824 23987 10848
rect 23667 9760 23675 9824
rect 23739 9760 23755 9824
rect 23819 9760 23835 9824
rect 23899 9760 23915 9824
rect 23979 9760 23987 9824
rect 23667 8736 23987 9760
rect 23667 8672 23675 8736
rect 23739 8672 23755 8736
rect 23819 8672 23835 8736
rect 23899 8672 23915 8736
rect 23979 8672 23987 8736
rect 23667 7648 23987 8672
rect 23667 7584 23675 7648
rect 23739 7584 23755 7648
rect 23819 7584 23835 7648
rect 23899 7584 23915 7648
rect 23979 7584 23987 7648
rect 21403 6900 21469 6901
rect 21403 6836 21404 6900
rect 21468 6836 21469 6900
rect 21403 6835 21469 6836
rect 20827 5952 20835 6016
rect 20899 5952 20915 6016
rect 20979 5952 20995 6016
rect 21059 5952 21075 6016
rect 21139 5952 21147 6016
rect 20827 4928 21147 5952
rect 20827 4864 20835 4928
rect 20899 4864 20915 4928
rect 20979 4864 20995 4928
rect 21059 4864 21075 4928
rect 21139 4864 21147 4928
rect 20827 3840 21147 4864
rect 20827 3776 20835 3840
rect 20899 3776 20915 3840
rect 20979 3776 20995 3840
rect 21059 3776 21075 3840
rect 21139 3776 21147 3840
rect 20827 2752 21147 3776
rect 20827 2688 20835 2752
rect 20899 2688 20915 2752
rect 20979 2688 20995 2752
rect 21059 2688 21075 2752
rect 21139 2688 21147 2752
rect 20827 2128 21147 2688
rect 23667 6560 23987 7584
rect 23667 6496 23675 6560
rect 23739 6496 23755 6560
rect 23819 6496 23835 6560
rect 23899 6496 23915 6560
rect 23979 6496 23987 6560
rect 23667 5472 23987 6496
rect 23667 5408 23675 5472
rect 23739 5408 23755 5472
rect 23819 5408 23835 5472
rect 23899 5408 23915 5472
rect 23979 5408 23987 5472
rect 23667 4384 23987 5408
rect 23667 4320 23675 4384
rect 23739 4320 23755 4384
rect 23819 4320 23835 4384
rect 23899 4320 23915 4384
rect 23979 4320 23987 4384
rect 23667 3296 23987 4320
rect 23667 3232 23675 3296
rect 23739 3232 23755 3296
rect 23819 3232 23835 3296
rect 23899 3232 23915 3296
rect 23979 3232 23987 3296
rect 23667 2208 23987 3232
rect 23667 2144 23675 2208
rect 23739 2144 23755 2208
rect 23819 2144 23835 2208
rect 23899 2144 23915 2208
rect 23979 2144 23987 2208
rect 23667 2128 23987 2144
use sky130_fd_sc_hd__diode_2  ANTENNA__372__A $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 9292 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__374__A
timestamp 1676037725
transform -1 0 12972 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__375__A
timestamp 1676037725
transform 1 0 15548 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__389__B
timestamp 1676037725
transform 1 0 7084 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__390__C
timestamp 1676037725
transform -1 0 4784 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__391__A
timestamp 1676037725
transform 1 0 9200 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__399__A
timestamp 1676037725
transform 1 0 16836 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__399__B
timestamp 1676037725
transform 1 0 16100 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__404__D
timestamp 1676037725
transform 1 0 3588 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__405__A
timestamp 1676037725
transform 1 0 11132 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__406__A0
timestamp 1676037725
transform -1 0 18124 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__408__A2
timestamp 1676037725
transform 1 0 11040 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__409__A2
timestamp 1676037725
transform 1 0 3312 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__422__A2
timestamp 1676037725
transform 1 0 3956 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__435__A
timestamp 1676037725
transform -1 0 14076 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__437__A2
timestamp 1676037725
transform -1 0 13708 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__437__B1
timestamp 1676037725
transform -1 0 14260 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__438__A2
timestamp 1676037725
transform 1 0 13340 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__438__B1
timestamp 1676037725
transform 1 0 15180 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__441__A
timestamp 1676037725
transform 1 0 13156 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__444__A
timestamp 1676037725
transform 1 0 14904 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__446__A
timestamp 1676037725
transform 1 0 12328 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__450__A1
timestamp 1676037725
transform 1 0 9568 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__450__B1
timestamp 1676037725
transform 1 0 11040 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__451__A1
timestamp 1676037725
transform 1 0 14260 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__451__B1
timestamp 1676037725
transform 1 0 14444 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__455__B
timestamp 1676037725
transform 1 0 13432 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__458__A1
timestamp 1676037725
transform 1 0 14352 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__463__B1
timestamp 1676037725
transform 1 0 13800 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__466__A
timestamp 1676037725
transform -1 0 15824 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__467__B
timestamp 1676037725
transform -1 0 21988 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__471__A
timestamp 1676037725
transform 1 0 18768 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__476__B1
timestamp 1676037725
transform 1 0 13064 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__477__A
timestamp 1676037725
transform 1 0 22632 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__480__A
timestamp 1676037725
transform -1 0 17756 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__480__B
timestamp 1676037725
transform 1 0 21436 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__482__B1
timestamp 1676037725
transform 1 0 12972 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__484__A
timestamp 1676037725
transform 1 0 16100 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__484__B
timestamp 1676037725
transform 1 0 14996 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__486__A
timestamp 1676037725
transform 1 0 14720 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__487__B
timestamp 1676037725
transform 1 0 20700 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__493__A
timestamp 1676037725
transform 1 0 16376 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__494__A
timestamp 1676037725
transform -1 0 19596 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__494__B
timestamp 1676037725
transform 1 0 18768 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__496__A2
timestamp 1676037725
transform 1 0 18492 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__497__A1
timestamp 1676037725
transform 1 0 15272 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__497__A2
timestamp 1676037725
transform 1 0 15824 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__497__B1
timestamp 1676037725
transform -1 0 14168 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__497__B2
timestamp 1676037725
transform 1 0 17940 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__498__A
timestamp 1676037725
transform 1 0 22816 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__498__B
timestamp 1676037725
transform -1 0 23368 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__499__A2
timestamp 1676037725
transform -1 0 21252 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__499__B1
timestamp 1676037725
transform -1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__502__C1
timestamp 1676037725
transform 1 0 11224 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__503__A
timestamp 1676037725
transform 1 0 11040 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__506__A1
timestamp 1676037725
transform 1 0 21160 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__506__A2
timestamp 1676037725
transform 1 0 21252 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__508__B
timestamp 1676037725
transform -1 0 21436 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__510__A
timestamp 1676037725
transform 1 0 20424 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__510__C
timestamp 1676037725
transform 1 0 19412 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__513__A1
timestamp 1676037725
transform 1 0 15916 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__514__B
timestamp 1676037725
transform 1 0 18308 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__515__A1
timestamp 1676037725
transform 1 0 20240 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__515__A2
timestamp 1676037725
transform 1 0 18492 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__516__A1
timestamp 1676037725
transform 1 0 15180 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__517__A
timestamp 1676037725
transform 1 0 15272 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__521__B1
timestamp 1676037725
transform -1 0 22540 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__521__C1
timestamp 1676037725
transform -1 0 22908 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__523__A
timestamp 1676037725
transform 1 0 20976 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__523__B
timestamp 1676037725
transform 1 0 20424 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__524__A
timestamp 1676037725
transform 1 0 23000 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__524__B
timestamp 1676037725
transform -1 0 23184 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__525__A1
timestamp 1676037725
transform -1 0 13156 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__526__A2
timestamp 1676037725
transform 1 0 22080 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__529__S
timestamp 1676037725
transform 1 0 16836 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__533__C
timestamp 1676037725
transform -1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__534__A2
timestamp 1676037725
transform 1 0 20976 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__535__B2
timestamp 1676037725
transform 1 0 20148 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__537__C1
timestamp 1676037725
transform 1 0 19228 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__539__A1
timestamp 1676037725
transform 1 0 15456 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__540__A3
timestamp 1676037725
transform 1 0 15088 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__541__B
timestamp 1676037725
transform -1 0 15824 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__544__A
timestamp 1676037725
transform 1 0 19964 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__546__C1
timestamp 1676037725
transform 1 0 22540 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__553__A2
timestamp 1676037725
transform -1 0 22172 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__555__B1
timestamp 1676037725
transform 1 0 22172 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__557__A1
timestamp 1676037725
transform 1 0 21988 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__557__B1
timestamp 1676037725
transform -1 0 23276 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__557__C1
timestamp 1676037725
transform 1 0 22724 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__560__A1
timestamp 1676037725
transform 1 0 18768 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__560__C1
timestamp 1676037725
transform 1 0 19412 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__564__B
timestamp 1676037725
transform 1 0 17296 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__565__A
timestamp 1676037725
transform 1 0 18308 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__566__A
timestamp 1676037725
transform -1 0 12604 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__567__A2
timestamp 1676037725
transform 1 0 20148 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__567__B1
timestamp 1676037725
transform 1 0 18860 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__567__B2
timestamp 1676037725
transform 1 0 20700 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__568__A1
timestamp 1676037725
transform 1 0 14260 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__568__A2
timestamp 1676037725
transform -1 0 11500 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__573__A
timestamp 1676037725
transform 1 0 11040 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__573__B
timestamp 1676037725
transform 1 0 13432 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__574__A1
timestamp 1676037725
transform 1 0 20056 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__576__A1
timestamp 1676037725
transform 1 0 18768 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__579__A1
timestamp 1676037725
transform 1 0 15824 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__580__A1
timestamp 1676037725
transform -1 0 17204 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__583__A
timestamp 1676037725
transform -1 0 14536 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__584__A
timestamp 1676037725
transform 1 0 18124 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__587__B1
timestamp 1676037725
transform 1 0 15548 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__589__A
timestamp 1676037725
transform 1 0 13616 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__589__B
timestamp 1676037725
transform 1 0 12052 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__590__A2
timestamp 1676037725
transform 1 0 16192 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__590__C1
timestamp 1676037725
transform 1 0 16744 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__591__A1
timestamp 1676037725
transform -1 0 16192 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__591__A2
timestamp 1676037725
transform 1 0 15456 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__592__A1
timestamp 1676037725
transform 1 0 16836 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__593__A
timestamp 1676037725
transform 1 0 13616 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__599__A1
timestamp 1676037725
transform 1 0 12696 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__601__C1
timestamp 1676037725
transform 1 0 18216 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__603__B1
timestamp 1676037725
transform 1 0 11040 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__605__B1
timestamp 1676037725
transform 1 0 14904 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__610__A
timestamp 1676037725
transform 1 0 15272 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__611__A1
timestamp 1676037725
transform 1 0 18768 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__612__B2
timestamp 1676037725
transform 1 0 20884 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__617__A1
timestamp 1676037725
transform -1 0 14996 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__622__A2
timestamp 1676037725
transform 1 0 16100 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__622__B1
timestamp 1676037725
transform 1 0 16468 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__624__A1
timestamp 1676037725
transform 1 0 16192 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__624__B1
timestamp 1676037725
transform 1 0 17572 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__629__A1
timestamp 1676037725
transform -1 0 14444 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__630__S
timestamp 1676037725
transform 1 0 11592 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__636__S
timestamp 1676037725
transform 1 0 11040 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__640__A1
timestamp 1676037725
transform -1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__641__A1_N
timestamp 1676037725
transform 1 0 17296 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__642__A2
timestamp 1676037725
transform -1 0 18032 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__645__A2
timestamp 1676037725
transform 1 0 11684 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__649__A1
timestamp 1676037725
transform 1 0 11132 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__650__A2
timestamp 1676037725
transform 1 0 14076 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__653__A
timestamp 1676037725
transform 1 0 5520 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__654__B1
timestamp 1676037725
transform 1 0 1748 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__660__A
timestamp 1676037725
transform 1 0 5888 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__661__B2
timestamp 1676037725
transform 1 0 7268 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__662__S
timestamp 1676037725
transform 1 0 12420 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__665__A2
timestamp 1676037725
transform 1 0 10396 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__666__A2
timestamp 1676037725
transform 1 0 11224 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__667__A1
timestamp 1676037725
transform -1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__667__A2
timestamp 1676037725
transform -1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__668__B1
timestamp 1676037725
transform 1 0 17388 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__669__A2
timestamp 1676037725
transform 1 0 16836 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__670__A2
timestamp 1676037725
transform 1 0 13524 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__673__A1
timestamp 1676037725
transform 1 0 10304 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__674__A1
timestamp 1676037725
transform 1 0 11224 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__675__S
timestamp 1676037725
transform 1 0 11684 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__678__A
timestamp 1676037725
transform 1 0 14812 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__678__B
timestamp 1676037725
transform 1 0 15364 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__679__A1
timestamp 1676037725
transform 1 0 9200 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__680__A
timestamp 1676037725
transform 1 0 9016 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__684__B
timestamp 1676037725
transform 1 0 3312 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__693__A1
timestamp 1676037725
transform 1 0 9660 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__699__A1
timestamp 1676037725
transform 1 0 11776 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__700__A1
timestamp 1676037725
transform 1 0 11040 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__703__B2
timestamp 1676037725
transform 1 0 5888 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__707__B1
timestamp 1676037725
transform 1 0 8464 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__712__A
timestamp 1676037725
transform 1 0 5980 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__712__B
timestamp 1676037725
transform 1 0 6532 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__713__A1
timestamp 1676037725
transform 1 0 7452 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__716__A3
timestamp 1676037725
transform 1 0 4508 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__718__A3
timestamp 1676037725
transform -1 0 1840 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__722__A2
timestamp 1676037725
transform 1 0 6532 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__722__A3
timestamp 1676037725
transform -1 0 1748 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__729__A1
timestamp 1676037725
transform 1 0 5888 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__736__B2
timestamp 1676037725
transform 1 0 4232 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__746__D
timestamp 1676037725
transform 1 0 8280 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__748__D
timestamp 1676037725
transform -1 0 10304 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__749__D
timestamp 1676037725
transform 1 0 10948 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__751__D
timestamp 1676037725
transform 1 0 10948 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__752__D
timestamp 1676037725
transform -1 0 11132 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__798__A
timestamp 1676037725
transform -1 0 1748 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A
timestamp 1676037725
transform 1 0 5796 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout16_A
timestamp 1676037725
transform -1 0 23368 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout17_A
timestamp 1676037725
transform 1 0 22540 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout24_A
timestamp 1676037725
transform -1 0 23276 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout45_A
timestamp 1676037725
transform 1 0 11684 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1676037725
transform -1 0 12144 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1676037725
transform -1 0 17112 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1676037725
transform -1 0 21528 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1676037725
transform -1 0 7176 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output5_A
timestamp 1676037725
transform 1 0 5888 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output8_A
timestamp 1676037725
transform 1 0 9108 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output10_A
timestamp 1676037725
transform -1 0 9844 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output11_A
timestamp 1676037725
transform 1 0 7820 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output12_A
timestamp 1676037725
transform 1 0 9108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1932 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2576 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36
timestamp 1676037725
transform 1 0 4416 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48
timestamp 1676037725
transform 1 0 5520 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1676037725
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1676037725
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65
timestamp 1676037725
transform 1 0 7084 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_75
timestamp 1676037725
transform 1 0 8004 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1676037725
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_89
timestamp 1676037725
transform 1 0 9292 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_96
timestamp 1676037725
transform 1 0 9936 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_103
timestamp 1676037725
transform 1 0 10580 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1676037725
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_113
timestamp 1676037725
transform 1 0 11500 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_120
timestamp 1676037725
transform 1 0 12144 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_127
timestamp 1676037725
transform 1 0 12788 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_134
timestamp 1676037725
transform 1 0 13432 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_146
timestamp 1676037725
transform 1 0 14536 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_153
timestamp 1676037725
transform 1 0 15180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_160
timestamp 1676037725
transform 1 0 15824 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1676037725
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1676037725
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_174
timestamp 1676037725
transform 1 0 17112 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_181
timestamp 1676037725
transform 1 0 17756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_188
timestamp 1676037725
transform 1 0 18400 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1676037725
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1676037725
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_202
timestamp 1676037725
transform 1 0 19688 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_209
timestamp 1676037725
transform 1 0 20332 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_216
timestamp 1676037725
transform 1 0 20976 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1676037725
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1676037725
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_230
timestamp 1676037725
transform 1 0 22264 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_237
timestamp 1676037725
transform 1 0 22908 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_243
timestamp 1676037725
transform 1 0 23460 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_7
timestamp 1676037725
transform 1 0 1748 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_17
timestamp 1676037725
transform 1 0 2668 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_27
timestamp 1676037725
transform 1 0 3588 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_39
timestamp 1676037725
transform 1 0 4692 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 1676037725
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_65
timestamp 1676037725
transform 1 0 7084 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_74
timestamp 1676037725
transform 1 0 7912 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_81
timestamp 1676037725
transform 1 0 8556 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_87
timestamp 1676037725
transform 1 0 9108 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_96
timestamp 1676037725
transform 1 0 9936 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_104
timestamp 1676037725
transform 1 0 10672 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1676037725
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_117
timestamp 1676037725
transform 1 0 11868 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_128
timestamp 1676037725
transform 1 0 12880 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_134
timestamp 1676037725
transform 1 0 13432 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_137
timestamp 1676037725
transform 1 0 13708 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_143
timestamp 1676037725
transform 1 0 14260 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_150 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14904 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_158
timestamp 1676037725
transform 1 0 15640 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_162
timestamp 1676037725
transform 1 0 16008 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_177
timestamp 1676037725
transform 1 0 17388 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_185
timestamp 1676037725
transform 1 0 18124 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_192
timestamp 1676037725
transform 1 0 18768 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_199
timestamp 1676037725
transform 1 0 19412 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_210
timestamp 1676037725
transform 1 0 20424 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1676037725
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1676037725
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_225
timestamp 1676037725
transform 1 0 21804 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_230
timestamp 1676037725
transform 1 0 22264 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_239
timestamp 1676037725
transform 1 0 23092 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_243
timestamp 1676037725
transform 1 0 23460 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_9
timestamp 1676037725
transform 1 0 1932 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1676037725
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_33
timestamp 1676037725
transform 1 0 4140 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_51
timestamp 1676037725
transform 1 0 5796 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_55
timestamp 1676037725
transform 1 0 6164 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_69
timestamp 1676037725
transform 1 0 7452 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp 1676037725
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_96
timestamp 1676037725
transform 1 0 9936 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_103
timestamp 1676037725
transform 1 0 10580 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_111
timestamp 1676037725
transform 1 0 11316 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_124
timestamp 1676037725
transform 1 0 12512 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1676037725
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_149
timestamp 1676037725
transform 1 0 14812 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_155
timestamp 1676037725
transform 1 0 15364 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_180
timestamp 1676037725
transform 1 0 17664 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_192
timestamp 1676037725
transform 1 0 18768 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1676037725
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_221
timestamp 1676037725
transform 1 0 21436 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_227
timestamp 1676037725
transform 1 0 21988 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_233
timestamp 1676037725
transform 1 0 22540 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_242
timestamp 1676037725
transform 1 0 23368 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_12
timestamp 1676037725
transform 1 0 2208 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_23
timestamp 1676037725
transform 1 0 3220 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_29
timestamp 1676037725
transform 1 0 3772 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_39
timestamp 1676037725
transform 1 0 4692 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_43
timestamp 1676037725
transform 1 0 5060 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1676037725
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1676037725
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_69
timestamp 1676037725
transform 1 0 7452 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_75
timestamp 1676037725
transform 1 0 8004 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_82
timestamp 1676037725
transform 1 0 8648 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_89
timestamp 1676037725
transform 1 0 9292 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_95
timestamp 1676037725
transform 1 0 9844 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_103
timestamp 1676037725
transform 1 0 10580 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 1676037725
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_113
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_123
timestamp 1676037725
transform 1 0 12420 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_129
timestamp 1676037725
transform 1 0 12972 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_135
timestamp 1676037725
transform 1 0 13524 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_141
timestamp 1676037725
transform 1 0 14076 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_147
timestamp 1676037725
transform 1 0 14628 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_155
timestamp 1676037725
transform 1 0 15364 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_164
timestamp 1676037725
transform 1 0 16192 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_173
timestamp 1676037725
transform 1 0 17020 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_179
timestamp 1676037725
transform 1 0 17572 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_185
timestamp 1676037725
transform 1 0 18124 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_196
timestamp 1676037725
transform 1 0 19136 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1676037725
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1676037725
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_225
timestamp 1676037725
transform 1 0 21804 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_231
timestamp 1676037725
transform 1 0 22356 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_237
timestamp 1676037725
transform 1 0 22908 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_243
timestamp 1676037725
transform 1 0 23460 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_9
timestamp 1676037725
transform 1 0 1932 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_20
timestamp 1676037725
transform 1 0 2944 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_26
timestamp 1676037725
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_33
timestamp 1676037725
transform 1 0 4140 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_43
timestamp 1676037725
transform 1 0 5060 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_49
timestamp 1676037725
transform 1 0 5612 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_53
timestamp 1676037725
transform 1 0 5980 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_71
timestamp 1676037725
transform 1 0 7636 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_78
timestamp 1676037725
transform 1 0 8280 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_93
timestamp 1676037725
transform 1 0 9660 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_105
timestamp 1676037725
transform 1 0 10764 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_109
timestamp 1676037725
transform 1 0 11132 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_112
timestamp 1676037725
transform 1 0 11408 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_120
timestamp 1676037725
transform 1 0 12144 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_127
timestamp 1676037725
transform 1 0 12788 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp 1676037725
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_145
timestamp 1676037725
transform 1 0 14444 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_151
timestamp 1676037725
transform 1 0 14996 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_157
timestamp 1676037725
transform 1 0 15548 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_163
timestamp 1676037725
transform 1 0 16100 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_172
timestamp 1676037725
transform 1 0 16928 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_178
timestamp 1676037725
transform 1 0 17480 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_184
timestamp 1676037725
transform 1 0 18032 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_194
timestamp 1676037725
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_197
timestamp 1676037725
transform 1 0 19228 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_206
timestamp 1676037725
transform 1 0 20056 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_213
timestamp 1676037725
transform 1 0 20700 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_219
timestamp 1676037725
transform 1 0 21252 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_240
timestamp 1676037725
transform 1 0 23184 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_16
timestamp 1676037725
transform 1 0 2576 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_26
timestamp 1676037725
transform 1 0 3496 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_34
timestamp 1676037725
transform 1 0 4232 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_46
timestamp 1676037725
transform 1 0 5336 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_5_53
timestamp 1676037725
transform 1 0 5980 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_66
timestamp 1676037725
transform 1 0 7176 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_83
timestamp 1676037725
transform 1 0 8740 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_89
timestamp 1676037725
transform 1 0 9292 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_95 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9844 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_107
timestamp 1676037725
transform 1 0 10948 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1676037725
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_121
timestamp 1676037725
transform 1 0 12236 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_125
timestamp 1676037725
transform 1 0 12604 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_131
timestamp 1676037725
transform 1 0 13156 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_137
timestamp 1676037725
transform 1 0 13708 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_143
timestamp 1676037725
transform 1 0 14260 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_154
timestamp 1676037725
transform 1 0 15272 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp 1676037725
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_5_189
timestamp 1676037725
transform 1 0 18492 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_197
timestamp 1676037725
transform 1 0 19228 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_207
timestamp 1676037725
transform 1 0 20148 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_216
timestamp 1676037725
transform 1 0 20976 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_222
timestamp 1676037725
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_225
timestamp 1676037725
transform 1 0 21804 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_229
timestamp 1676037725
transform 1 0 22172 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_238
timestamp 1676037725
transform 1 0 23000 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_7
timestamp 1676037725
transform 1 0 1748 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_15
timestamp 1676037725
transform 1 0 2484 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_26
timestamp 1676037725
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_36
timestamp 1676037725
transform 1 0 4416 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_40
timestamp 1676037725
transform 1 0 4784 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_57
timestamp 1676037725
transform 1 0 6348 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_63
timestamp 1676037725
transform 1 0 6900 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_67
timestamp 1676037725
transform 1 0 7268 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_71
timestamp 1676037725
transform 1 0 7636 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_81
timestamp 1676037725
transform 1 0 8556 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_90
timestamp 1676037725
transform 1 0 9384 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_105
timestamp 1676037725
transform 1 0 10764 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_111
timestamp 1676037725
transform 1 0 11316 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_123
timestamp 1676037725
transform 1 0 12420 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_134
timestamp 1676037725
transform 1 0 13432 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_149
timestamp 1676037725
transform 1 0 14812 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_156
timestamp 1676037725
transform 1 0 15456 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_165
timestamp 1676037725
transform 1 0 16284 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_169
timestamp 1676037725
transform 1 0 16652 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_184
timestamp 1676037725
transform 1 0 18032 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_193
timestamp 1676037725
transform 1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_197
timestamp 1676037725
transform 1 0 19228 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_212
timestamp 1676037725
transform 1 0 20608 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_224
timestamp 1676037725
transform 1 0 21712 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_6_238
timestamp 1676037725
transform 1 0 23000 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_9
timestamp 1676037725
transform 1 0 1932 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_27
timestamp 1676037725
transform 1 0 3588 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_41
timestamp 1676037725
transform 1 0 4876 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1676037725
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_66
timestamp 1676037725
transform 1 0 7176 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_74
timestamp 1676037725
transform 1 0 7912 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_83
timestamp 1676037725
transform 1 0 8740 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_95
timestamp 1676037725
transform 1 0 9844 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_103
timestamp 1676037725
transform 1 0 10580 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp 1676037725
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_121
timestamp 1676037725
transform 1 0 12236 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_133
timestamp 1676037725
transform 1 0 13340 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_143
timestamp 1676037725
transform 1 0 14260 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_149
timestamp 1676037725
transform 1 0 14812 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_159
timestamp 1676037725
transform 1 0 15732 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_165
timestamp 1676037725
transform 1 0 16284 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_173
timestamp 1676037725
transform 1 0 17020 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_181
timestamp 1676037725
transform 1 0 17756 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_191
timestamp 1676037725
transform 1 0 18676 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_211
timestamp 1676037725
transform 1 0 20516 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_220
timestamp 1676037725
transform 1 0 21344 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_225
timestamp 1676037725
transform 1 0 21804 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_233
timestamp 1676037725
transform 1 0 22540 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_242
timestamp 1676037725
transform 1 0 23368 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_9
timestamp 1676037725
transform 1 0 1932 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_17
timestamp 1676037725
transform 1 0 2668 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_26
timestamp 1676037725
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_39
timestamp 1676037725
transform 1 0 4692 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_57
timestamp 1676037725
transform 1 0 6348 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_82
timestamp 1676037725
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_89
timestamp 1676037725
transform 1 0 9292 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_97
timestamp 1676037725
transform 1 0 10028 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_103
timestamp 1676037725
transform 1 0 10580 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_109
timestamp 1676037725
transform 1 0 11132 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_112
timestamp 1676037725
transform 1 0 11408 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_118
timestamp 1676037725
transform 1 0 11960 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_130
timestamp 1676037725
transform 1 0 13064 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1676037725
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1676037725
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_146
timestamp 1676037725
transform 1 0 14536 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_153
timestamp 1676037725
transform 1 0 15180 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_159
timestamp 1676037725
transform 1 0 15732 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_165
timestamp 1676037725
transform 1 0 16284 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_168
timestamp 1676037725
transform 1 0 16560 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_172
timestamp 1676037725
transform 1 0 16928 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_175
timestamp 1676037725
transform 1 0 17204 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_181
timestamp 1676037725
transform 1 0 17756 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_194
timestamp 1676037725
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_197
timestamp 1676037725
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_213
timestamp 1676037725
transform 1 0 20700 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_219
timestamp 1676037725
transform 1 0 21252 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_226
timestamp 1676037725
transform 1 0 21896 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_235
timestamp 1676037725
transform 1 0 22724 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_8_241
timestamp 1676037725
transform 1 0 23276 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_12
timestamp 1676037725
transform 1 0 2208 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_24
timestamp 1676037725
transform 1 0 3312 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_31
timestamp 1676037725
transform 1 0 3956 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_39
timestamp 1676037725
transform 1 0 4692 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_49
timestamp 1676037725
transform 1 0 5612 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1676037725
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_66
timestamp 1676037725
transform 1 0 7176 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_81
timestamp 1676037725
transform 1 0 8556 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_92
timestamp 1676037725
transform 1 0 9568 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_101
timestamp 1676037725
transform 1 0 10396 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_107
timestamp 1676037725
transform 1 0 10948 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_110
timestamp 1676037725
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_122
timestamp 1676037725
transform 1 0 12328 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_132
timestamp 1676037725
transform 1 0 13248 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_9_140
timestamp 1676037725
transform 1 0 13984 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_155
timestamp 1676037725
transform 1 0 15364 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_163
timestamp 1676037725
transform 1 0 16100 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1676037725
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_169
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_175
timestamp 1676037725
transform 1 0 17204 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_192
timestamp 1676037725
transform 1 0 18768 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_209
timestamp 1676037725
transform 1 0 20332 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_218
timestamp 1676037725
transform 1 0 21160 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_9_225
timestamp 1676037725
transform 1 0 21804 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_239
timestamp 1676037725
transform 1 0 23092 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_243
timestamp 1676037725
transform 1 0 23460 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_15
timestamp 1676037725
transform 1 0 2484 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_25
timestamp 1676037725
transform 1 0 3404 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_41
timestamp 1676037725
transform 1 0 4876 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_53
timestamp 1676037725
transform 1 0 5980 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_68
timestamp 1676037725
transform 1 0 7360 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1676037725
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1676037725
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_89
timestamp 1676037725
transform 1 0 9292 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_97
timestamp 1676037725
transform 1 0 10028 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_110
timestamp 1676037725
transform 1 0 11224 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_114
timestamp 1676037725
transform 1 0 11592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_118
timestamp 1676037725
transform 1 0 11960 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_124
timestamp 1676037725
transform 1 0 12512 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_132
timestamp 1676037725
transform 1 0 13248 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 1676037725
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_141
timestamp 1676037725
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_157
timestamp 1676037725
transform 1 0 15548 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_164
timestamp 1676037725
transform 1 0 16192 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_185
timestamp 1676037725
transform 1 0 18124 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_191
timestamp 1676037725
transform 1 0 18676 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1676037725
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1676037725
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_202
timestamp 1676037725
transform 1 0 19688 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_210
timestamp 1676037725
transform 1 0 20424 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_217
timestamp 1676037725
transform 1 0 21068 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_223
timestamp 1676037725
transform 1 0 21620 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_239
timestamp 1676037725
transform 1 0 23092 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_243
timestamp 1676037725
transform 1 0 23460 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_9
timestamp 1676037725
transform 1 0 1932 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_20
timestamp 1676037725
transform 1 0 2944 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_31
timestamp 1676037725
transform 1 0 3956 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_39
timestamp 1676037725
transform 1 0 4692 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_49
timestamp 1676037725
transform 1 0 5612 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1676037725
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_70
timestamp 1676037725
transform 1 0 7544 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_82
timestamp 1676037725
transform 1 0 8648 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_88
timestamp 1676037725
transform 1 0 9200 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_94
timestamp 1676037725
transform 1 0 9752 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_101
timestamp 1676037725
transform 1 0 10396 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_107
timestamp 1676037725
transform 1 0 10948 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1676037725
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_113
timestamp 1676037725
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_122
timestamp 1676037725
transform 1 0 12328 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_132
timestamp 1676037725
transform 1 0 13248 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_11_154
timestamp 1676037725
transform 1 0 15272 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_160
timestamp 1676037725
transform 1 0 15824 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1676037725
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_169
timestamp 1676037725
transform 1 0 16652 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_175
timestamp 1676037725
transform 1 0 17204 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_188
timestamp 1676037725
transform 1 0 18400 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_204
timestamp 1676037725
transform 1 0 19872 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_210
timestamp 1676037725
transform 1 0 20424 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_216
timestamp 1676037725
transform 1 0 20976 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_221
timestamp 1676037725
transform 1 0 21436 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_225
timestamp 1676037725
transform 1 0 21804 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_229
timestamp 1676037725
transform 1 0 22172 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_237
timestamp 1676037725
transform 1 0 22908 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_243
timestamp 1676037725
transform 1 0 23460 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_7
timestamp 1676037725
transform 1 0 1748 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_17
timestamp 1676037725
transform 1 0 2668 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp 1676037725
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_37
timestamp 1676037725
transform 1 0 4508 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_47
timestamp 1676037725
transform 1 0 5428 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_55
timestamp 1676037725
transform 1 0 6164 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_63
timestamp 1676037725
transform 1 0 6900 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_75
timestamp 1676037725
transform 1 0 8004 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1676037725
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_89
timestamp 1676037725
transform 1 0 9292 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_98
timestamp 1676037725
transform 1 0 10120 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_109
timestamp 1676037725
transform 1 0 11132 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_117
timestamp 1676037725
transform 1 0 11868 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_125
timestamp 1676037725
transform 1 0 12604 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1676037725
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1676037725
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1676037725
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_148
timestamp 1676037725
transform 1 0 14720 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_159
timestamp 1676037725
transform 1 0 15732 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_167
timestamp 1676037725
transform 1 0 16468 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_177
timestamp 1676037725
transform 1 0 17388 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_188
timestamp 1676037725
transform 1 0 18400 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1676037725
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_197
timestamp 1676037725
transform 1 0 19228 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_212
timestamp 1676037725
transform 1 0 20608 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_224
timestamp 1676037725
transform 1 0 21712 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_230
timestamp 1676037725
transform 1 0 22264 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_236
timestamp 1676037725
transform 1 0 22816 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_242
timestamp 1676037725
transform 1 0 23368 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_3
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_11
timestamp 1676037725
transform 1 0 2116 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_21
timestamp 1676037725
transform 1 0 3036 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_32
timestamp 1676037725
transform 1 0 4048 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_42
timestamp 1676037725
transform 1 0 4968 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1676037725
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_61
timestamp 1676037725
transform 1 0 6716 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_67
timestamp 1676037725
transform 1 0 7268 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_79
timestamp 1676037725
transform 1 0 8372 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_91
timestamp 1676037725
transform 1 0 9476 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_100
timestamp 1676037725
transform 1 0 10304 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_106
timestamp 1676037725
transform 1 0 10856 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_110
timestamp 1676037725
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_113
timestamp 1676037725
transform 1 0 11500 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_119
timestamp 1676037725
transform 1 0 12052 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_131
timestamp 1676037725
transform 1 0 13156 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_140
timestamp 1676037725
transform 1 0 13984 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_146
timestamp 1676037725
transform 1 0 14536 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_152
timestamp 1676037725
transform 1 0 15088 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_158
timestamp 1676037725
transform 1 0 15640 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_164
timestamp 1676037725
transform 1 0 16192 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1676037725
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_180
timestamp 1676037725
transform 1 0 17664 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_192
timestamp 1676037725
transform 1 0 18768 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_196
timestamp 1676037725
transform 1 0 19136 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_203
timestamp 1676037725
transform 1 0 19780 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_214
timestamp 1676037725
transform 1 0 20792 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_220
timestamp 1676037725
transform 1 0 21344 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_225
timestamp 1676037725
transform 1 0 21804 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_234
timestamp 1676037725
transform 1 0 22632 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_240
timestamp 1676037725
transform 1 0 23184 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1676037725
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_7
timestamp 1676037725
transform 1 0 1748 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_16
timestamp 1676037725
transform 1 0 2576 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_26
timestamp 1676037725
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_29
timestamp 1676037725
transform 1 0 3772 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_33
timestamp 1676037725
transform 1 0 4140 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_36
timestamp 1676037725
transform 1 0 4416 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_48
timestamp 1676037725
transform 1 0 5520 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_54
timestamp 1676037725
transform 1 0 6072 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_62
timestamp 1676037725
transform 1 0 6808 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_66
timestamp 1676037725
transform 1 0 7176 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_69
timestamp 1676037725
transform 1 0 7452 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1676037725
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_85
timestamp 1676037725
transform 1 0 8924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_98
timestamp 1676037725
transform 1 0 10120 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_109
timestamp 1676037725
transform 1 0 11132 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_117
timestamp 1676037725
transform 1 0 11868 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_130
timestamp 1676037725
transform 1 0 13064 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_136
timestamp 1676037725
transform 1 0 13616 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_141
timestamp 1676037725
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_145
timestamp 1676037725
transform 1 0 14444 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_149
timestamp 1676037725
transform 1 0 14812 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_157
timestamp 1676037725
transform 1 0 15548 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_170
timestamp 1676037725
transform 1 0 16744 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_181
timestamp 1676037725
transform 1 0 17756 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_190
timestamp 1676037725
transform 1 0 18584 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_197
timestamp 1676037725
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_201
timestamp 1676037725
transform 1 0 19596 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_213
timestamp 1676037725
transform 1 0 20700 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_221
timestamp 1676037725
transform 1 0 21436 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_225
timestamp 1676037725
transform 1 0 21804 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_236
timestamp 1676037725
transform 1 0 22816 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_242
timestamp 1676037725
transform 1 0 23368 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_3
timestamp 1676037725
transform 1 0 1380 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_13
timestamp 1676037725
transform 1 0 2300 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_20
timestamp 1676037725
transform 1 0 2944 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_24
timestamp 1676037725
transform 1 0 3312 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_32
timestamp 1676037725
transform 1 0 4048 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_36
timestamp 1676037725
transform 1 0 4416 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_39
timestamp 1676037725
transform 1 0 4692 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_48
timestamp 1676037725
transform 1 0 5520 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_54
timestamp 1676037725
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_68
timestamp 1676037725
transform 1 0 7360 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_78
timestamp 1676037725
transform 1 0 8280 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_91
timestamp 1676037725
transform 1 0 9476 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_99
timestamp 1676037725
transform 1 0 10212 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_102
timestamp 1676037725
transform 1 0 10488 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_110
timestamp 1676037725
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_113
timestamp 1676037725
transform 1 0 11500 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_117
timestamp 1676037725
transform 1 0 11868 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_127
timestamp 1676037725
transform 1 0 12788 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_135
timestamp 1676037725
transform 1 0 13524 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_141
timestamp 1676037725
transform 1 0 14076 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_153
timestamp 1676037725
transform 1 0 15180 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_165
timestamp 1676037725
transform 1 0 16284 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_169
timestamp 1676037725
transform 1 0 16652 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_187
timestamp 1676037725
transform 1 0 18308 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_200
timestamp 1676037725
transform 1 0 19504 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_209
timestamp 1676037725
transform 1 0 20332 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_215
timestamp 1676037725
transform 1 0 20884 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_221
timestamp 1676037725
transform 1 0 21436 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_225
timestamp 1676037725
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_234
timestamp 1676037725
transform 1 0 22632 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_240
timestamp 1676037725
transform 1 0 23184 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1676037725
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_24
timestamp 1676037725
transform 1 0 3312 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1676037725
transform 1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_39
timestamp 1676037725
transform 1 0 4692 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_47
timestamp 1676037725
transform 1 0 5428 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_50
timestamp 1676037725
transform 1 0 5704 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_76
timestamp 1676037725
transform 1 0 8096 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1676037725
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_85
timestamp 1676037725
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_95
timestamp 1676037725
transform 1 0 9844 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_106
timestamp 1676037725
transform 1 0 10856 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_110
timestamp 1676037725
transform 1 0 11224 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_113
timestamp 1676037725
transform 1 0 11500 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_126
timestamp 1676037725
transform 1 0 12696 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_137
timestamp 1676037725
transform 1 0 13708 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1676037725
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_151
timestamp 1676037725
transform 1 0 14996 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_160
timestamp 1676037725
transform 1 0 15824 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_166
timestamp 1676037725
transform 1 0 16376 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_172
timestamp 1676037725
transform 1 0 16928 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_178
timestamp 1676037725
transform 1 0 17480 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_186
timestamp 1676037725
transform 1 0 18216 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1676037725
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_197
timestamp 1676037725
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_203
timestamp 1676037725
transform 1 0 19780 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_209
timestamp 1676037725
transform 1 0 20332 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_215
timestamp 1676037725
transform 1 0 20884 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_221
timestamp 1676037725
transform 1 0 21436 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_232
timestamp 1676037725
transform 1 0 22448 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_238
timestamp 1676037725
transform 1 0 23000 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1676037725
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_9
timestamp 1676037725
transform 1 0 1932 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_13
timestamp 1676037725
transform 1 0 2300 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_20
timestamp 1676037725
transform 1 0 2944 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_26
timestamp 1676037725
transform 1 0 3496 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_30
timestamp 1676037725
transform 1 0 3864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_36
timestamp 1676037725
transform 1 0 4416 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_48
timestamp 1676037725
transform 1 0 5520 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1676037725
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_57
timestamp 1676037725
transform 1 0 6348 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_61
timestamp 1676037725
transform 1 0 6716 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_69
timestamp 1676037725
transform 1 0 7452 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_78
timestamp 1676037725
transform 1 0 8280 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_91
timestamp 1676037725
transform 1 0 9476 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_101
timestamp 1676037725
transform 1 0 10396 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1676037725
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_113
timestamp 1676037725
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_121
timestamp 1676037725
transform 1 0 12236 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_129
timestamp 1676037725
transform 1 0 12972 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_144
timestamp 1676037725
transform 1 0 14352 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_150
timestamp 1676037725
transform 1 0 14904 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_156
timestamp 1676037725
transform 1 0 15456 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_162
timestamp 1676037725
transform 1 0 16008 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_17_169
timestamp 1676037725
transform 1 0 16652 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_175
timestamp 1676037725
transform 1 0 17204 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_183
timestamp 1676037725
transform 1 0 17940 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_189
timestamp 1676037725
transform 1 0 18492 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_195
timestamp 1676037725
transform 1 0 19044 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_206
timestamp 1676037725
transform 1 0 20056 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_212
timestamp 1676037725
transform 1 0 20608 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_218
timestamp 1676037725
transform 1 0 21160 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1676037725
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_225
timestamp 1676037725
transform 1 0 21804 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_234
timestamp 1676037725
transform 1 0 22632 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_241
timestamp 1676037725
transform 1 0 23276 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_3
timestamp 1676037725
transform 1 0 1380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_9
timestamp 1676037725
transform 1 0 1932 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_15
timestamp 1676037725
transform 1 0 2484 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_24
timestamp 1676037725
transform 1 0 3312 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1676037725
transform 1 0 3772 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_34
timestamp 1676037725
transform 1 0 4232 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_40
timestamp 1676037725
transform 1 0 4784 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_52
timestamp 1676037725
transform 1 0 5888 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_55
timestamp 1676037725
transform 1 0 6164 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_62
timestamp 1676037725
transform 1 0 6808 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_69
timestamp 1676037725
transform 1 0 7452 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_75
timestamp 1676037725
transform 1 0 8004 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_80
timestamp 1676037725
transform 1 0 8464 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_85
timestamp 1676037725
transform 1 0 8924 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_90
timestamp 1676037725
transform 1 0 9384 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_107
timestamp 1676037725
transform 1 0 10948 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_111
timestamp 1676037725
transform 1 0 11316 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_119
timestamp 1676037725
transform 1 0 12052 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_125
timestamp 1676037725
transform 1 0 12604 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_131
timestamp 1676037725
transform 1 0 13156 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1676037725
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1676037725
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_150
timestamp 1676037725
transform 1 0 14904 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_156
timestamp 1676037725
transform 1 0 15456 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_162
timestamp 1676037725
transform 1 0 16008 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_168
timestamp 1676037725
transform 1 0 16560 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_174
timestamp 1676037725
transform 1 0 17112 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_183
timestamp 1676037725
transform 1 0 17940 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1676037725
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1676037725
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1676037725
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_201
timestamp 1676037725
transform 1 0 19596 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_205
timestamp 1676037725
transform 1 0 19964 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_208
timestamp 1676037725
transform 1 0 20240 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_212
timestamp 1676037725
transform 1 0 20608 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_218
timestamp 1676037725
transform 1 0 21160 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_229
timestamp 1676037725
transform 1 0 22172 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_233
timestamp 1676037725
transform 1 0 22540 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_240
timestamp 1676037725
transform 1 0 23184 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_3
timestamp 1676037725
transform 1 0 1380 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_8
timestamp 1676037725
transform 1 0 1840 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_18
timestamp 1676037725
transform 1 0 2760 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_26
timestamp 1676037725
transform 1 0 3496 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_30
timestamp 1676037725
transform 1 0 3864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_36
timestamp 1676037725
transform 1 0 4416 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_47
timestamp 1676037725
transform 1 0 5428 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1676037725
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1676037725
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_61
timestamp 1676037725
transform 1 0 6716 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_72
timestamp 1676037725
transform 1 0 7728 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_79
timestamp 1676037725
transform 1 0 8372 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_90
timestamp 1676037725
transform 1 0 9384 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1676037725
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_113
timestamp 1676037725
transform 1 0 11500 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_125
timestamp 1676037725
transform 1 0 12604 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_133
timestamp 1676037725
transform 1 0 13340 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_148
timestamp 1676037725
transform 1 0 14720 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_152
timestamp 1676037725
transform 1 0 15088 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_155
timestamp 1676037725
transform 1 0 15364 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1676037725
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1676037725
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_179
timestamp 1676037725
transform 1 0 17572 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_185
timestamp 1676037725
transform 1 0 18124 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_191
timestamp 1676037725
transform 1 0 18676 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_207
timestamp 1676037725
transform 1 0 20148 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_215
timestamp 1676037725
transform 1 0 20884 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1676037725
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_225
timestamp 1676037725
transform 1 0 21804 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_229
timestamp 1676037725
transform 1 0 22172 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_238
timestamp 1676037725
transform 1 0 23000 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_20_3
timestamp 1676037725
transform 1 0 1380 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_18
timestamp 1676037725
transform 1 0 2760 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp 1676037725
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_29
timestamp 1676037725
transform 1 0 3772 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_33
timestamp 1676037725
transform 1 0 4140 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_39
timestamp 1676037725
transform 1 0 4692 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_49
timestamp 1676037725
transform 1 0 5612 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_61
timestamp 1676037725
transform 1 0 6716 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_81
timestamp 1676037725
transform 1 0 8556 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_85
timestamp 1676037725
transform 1 0 8924 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_91
timestamp 1676037725
transform 1 0 9476 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_106
timestamp 1676037725
transform 1 0 10856 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_112
timestamp 1676037725
transform 1 0 11408 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1676037725
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1676037725
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_150
timestamp 1676037725
transform 1 0 14904 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_159
timestamp 1676037725
transform 1 0 15732 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_169
timestamp 1676037725
transform 1 0 16652 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_180
timestamp 1676037725
transform 1 0 17664 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1676037725
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_197
timestamp 1676037725
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_206
timestamp 1676037725
transform 1 0 20056 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_217
timestamp 1676037725
transform 1 0 21068 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_227
timestamp 1676037725
transform 1 0 21988 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_241
timestamp 1676037725
transform 1 0 23276 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_3
timestamp 1676037725
transform 1 0 1380 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_7
timestamp 1676037725
transform 1 0 1748 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_12
timestamp 1676037725
transform 1 0 2208 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_32
timestamp 1676037725
transform 1 0 4048 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_40
timestamp 1676037725
transform 1 0 4784 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_52
timestamp 1676037725
transform 1 0 5888 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1676037725
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_71
timestamp 1676037725
transform 1 0 7636 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_93
timestamp 1676037725
transform 1 0 9660 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_100
timestamp 1676037725
transform 1 0 10304 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_109
timestamp 1676037725
transform 1 0 11132 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_113
timestamp 1676037725
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_117
timestamp 1676037725
transform 1 0 11868 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_125
timestamp 1676037725
transform 1 0 12604 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_128
timestamp 1676037725
transform 1 0 12880 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_142
timestamp 1676037725
transform 1 0 14168 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_153
timestamp 1676037725
transform 1 0 15180 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_164
timestamp 1676037725
transform 1 0 16192 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1676037725
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_173
timestamp 1676037725
transform 1 0 17020 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_179
timestamp 1676037725
transform 1 0 17572 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_187
timestamp 1676037725
transform 1 0 18308 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_21_202
timestamp 1676037725
transform 1 0 19688 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_208
timestamp 1676037725
transform 1 0 20240 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1676037725
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1676037725
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_225
timestamp 1676037725
transform 1 0 21804 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_239
timestamp 1676037725
transform 1 0 23092 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_243
timestamp 1676037725
transform 1 0 23460 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_3
timestamp 1676037725
transform 1 0 1380 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_9
timestamp 1676037725
transform 1 0 1932 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_15
timestamp 1676037725
transform 1 0 2484 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1676037725
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1676037725
transform 1 0 3772 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_40
timestamp 1676037725
transform 1 0 4784 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_48
timestamp 1676037725
transform 1 0 5520 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_58
timestamp 1676037725
transform 1 0 6440 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_69
timestamp 1676037725
transform 1 0 7452 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1676037725
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_85
timestamp 1676037725
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_94
timestamp 1676037725
transform 1 0 9752 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_102
timestamp 1676037725
transform 1 0 10488 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_112
timestamp 1676037725
transform 1 0 11408 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_118
timestamp 1676037725
transform 1 0 11960 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_126
timestamp 1676037725
transform 1 0 12696 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_136
timestamp 1676037725
transform 1 0 13616 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1676037725
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_152
timestamp 1676037725
transform 1 0 15088 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_22_167
timestamp 1676037725
transform 1 0 16468 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_173
timestamp 1676037725
transform 1 0 17020 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_181
timestamp 1676037725
transform 1 0 17756 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_193
timestamp 1676037725
transform 1 0 18860 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1676037725
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_206
timestamp 1676037725
transform 1 0 20056 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_212
timestamp 1676037725
transform 1 0 20608 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_218
timestamp 1676037725
transform 1 0 21160 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_227
timestamp 1676037725
transform 1 0 21988 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_237
timestamp 1676037725
transform 1 0 22908 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_243
timestamp 1676037725
transform 1 0 23460 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1676037725
transform 1 0 1380 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_12
timestamp 1676037725
transform 1 0 2208 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_16
timestamp 1676037725
transform 1 0 2576 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_36
timestamp 1676037725
transform 1 0 4416 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_47
timestamp 1676037725
transform 1 0 5428 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_51
timestamp 1676037725
transform 1 0 5796 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1676037725
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1676037725
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_63
timestamp 1676037725
transform 1 0 6900 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_94
timestamp 1676037725
transform 1 0 9752 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_100
timestamp 1676037725
transform 1 0 10304 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1676037725
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_113
timestamp 1676037725
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_117
timestamp 1676037725
transform 1 0 11868 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_134
timestamp 1676037725
transform 1 0 13432 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_144
timestamp 1676037725
transform 1 0 14352 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_152
timestamp 1676037725
transform 1 0 15088 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_156
timestamp 1676037725
transform 1 0 15456 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_163
timestamp 1676037725
transform 1 0 16100 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1676037725
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1676037725
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_173
timestamp 1676037725
transform 1 0 17020 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_185
timestamp 1676037725
transform 1 0 18124 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_191
timestamp 1676037725
transform 1 0 18676 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_194
timestamp 1676037725
transform 1 0 18952 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_205
timestamp 1676037725
transform 1 0 19964 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_218
timestamp 1676037725
transform 1 0 21160 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_225
timestamp 1676037725
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_235
timestamp 1676037725
transform 1 0 22724 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_241
timestamp 1676037725
transform 1 0 23276 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_24_3
timestamp 1676037725
transform 1 0 1380 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_9
timestamp 1676037725
transform 1 0 1932 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_16
timestamp 1676037725
transform 1 0 2576 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_26
timestamp 1676037725
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1676037725
transform 1 0 3772 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_37
timestamp 1676037725
transform 1 0 4508 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_41
timestamp 1676037725
transform 1 0 4876 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_58
timestamp 1676037725
transform 1 0 6440 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_70
timestamp 1676037725
transform 1 0 7544 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1676037725
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_85
timestamp 1676037725
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_103
timestamp 1676037725
transform 1 0 10580 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_119
timestamp 1676037725
transform 1 0 12052 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_132
timestamp 1676037725
transform 1 0 13248 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1676037725
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1676037725
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_146
timestamp 1676037725
transform 1 0 14536 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_159
timestamp 1676037725
transform 1 0 15732 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_165
timestamp 1676037725
transform 1 0 16284 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_173
timestamp 1676037725
transform 1 0 17020 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_187
timestamp 1676037725
transform 1 0 18308 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 1676037725
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1676037725
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_201
timestamp 1676037725
transform 1 0 19596 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_207
timestamp 1676037725
transform 1 0 20148 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_211
timestamp 1676037725
transform 1 0 20516 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_218
timestamp 1676037725
transform 1 0 21160 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_226
timestamp 1676037725
transform 1 0 21896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_231
timestamp 1676037725
transform 1 0 22356 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_237
timestamp 1676037725
transform 1 0 22908 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_243
timestamp 1676037725
transform 1 0 23460 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1676037725
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_15
timestamp 1676037725
transform 1 0 2484 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_36
timestamp 1676037725
transform 1 0 4416 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_48
timestamp 1676037725
transform 1 0 5520 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1676037725
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_69
timestamp 1676037725
transform 1 0 7452 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1676037725
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1676037725
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1676037725
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_113
timestamp 1676037725
transform 1 0 11500 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_121
timestamp 1676037725
transform 1 0 12236 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_147
timestamp 1676037725
transform 1 0 14628 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_153
timestamp 1676037725
transform 1 0 15180 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_159
timestamp 1676037725
transform 1 0 15732 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_165
timestamp 1676037725
transform 1 0 16284 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_169
timestamp 1676037725
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_177
timestamp 1676037725
transform 1 0 17388 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_185
timestamp 1676037725
transform 1 0 18124 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_192
timestamp 1676037725
transform 1 0 18768 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_200
timestamp 1676037725
transform 1 0 19504 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_206
timestamp 1676037725
transform 1 0 20056 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_218
timestamp 1676037725
transform 1 0 21160 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1676037725
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_229
timestamp 1676037725
transform 1 0 22172 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_235
timestamp 1676037725
transform 1 0 22724 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_243
timestamp 1676037725
transform 1 0 23460 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_3
timestamp 1676037725
transform 1 0 1380 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_9
timestamp 1676037725
transform 1 0 1932 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_26
timestamp 1676037725
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1676037725
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_41
timestamp 1676037725
transform 1 0 4876 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_61
timestamp 1676037725
transform 1 0 6716 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1676037725
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_85
timestamp 1676037725
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_106
timestamp 1676037725
transform 1 0 10856 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_114
timestamp 1676037725
transform 1 0 11592 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_121
timestamp 1676037725
transform 1 0 12236 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_132
timestamp 1676037725
transform 1 0 13248 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1676037725
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_141
timestamp 1676037725
transform 1 0 14076 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_152
timestamp 1676037725
transform 1 0 15088 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_163
timestamp 1676037725
transform 1 0 16100 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_169
timestamp 1676037725
transform 1 0 16652 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_173
timestamp 1676037725
transform 1 0 17020 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_182
timestamp 1676037725
transform 1 0 17848 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_190
timestamp 1676037725
transform 1 0 18584 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1676037725
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_197
timestamp 1676037725
transform 1 0 19228 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_203
timestamp 1676037725
transform 1 0 19780 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_212
timestamp 1676037725
transform 1 0 20608 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_218
timestamp 1676037725
transform 1 0 21160 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_226
timestamp 1676037725
transform 1 0 21896 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_232
timestamp 1676037725
transform 1 0 22448 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1676037725
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_15
timestamp 1676037725
transform 1 0 2484 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_36
timestamp 1676037725
transform 1 0 4416 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_48
timestamp 1676037725
transform 1 0 5520 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1676037725
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_69
timestamp 1676037725
transform 1 0 7452 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_77
timestamp 1676037725
transform 1 0 8188 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_80
timestamp 1676037725
transform 1 0 8464 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_103
timestamp 1676037725
transform 1 0 10580 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_109
timestamp 1676037725
transform 1 0 11132 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_113
timestamp 1676037725
transform 1 0 11500 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_121
timestamp 1676037725
transform 1 0 12236 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_132
timestamp 1676037725
transform 1 0 13248 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_147
timestamp 1676037725
transform 1 0 14628 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_157
timestamp 1676037725
transform 1 0 15548 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_163
timestamp 1676037725
transform 1 0 16100 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1676037725
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1676037725
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_175
timestamp 1676037725
transform 1 0 17204 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_179
timestamp 1676037725
transform 1 0 17572 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_186
timestamp 1676037725
transform 1 0 18216 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_203
timestamp 1676037725
transform 1 0 19780 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_209
timestamp 1676037725
transform 1 0 20332 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1676037725
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1676037725
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1676037725
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_237
timestamp 1676037725
transform 1 0 22908 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_243
timestamp 1676037725
transform 1 0 23460 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_3
timestamp 1676037725
transform 1 0 1380 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_9
timestamp 1676037725
transform 1 0 1932 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_26
timestamp 1676037725
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1676037725
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_41
timestamp 1676037725
transform 1 0 4876 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_49
timestamp 1676037725
transform 1 0 5612 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_66
timestamp 1676037725
transform 1 0 7176 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_78
timestamp 1676037725
transform 1 0 8280 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_85
timestamp 1676037725
transform 1 0 8924 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_103
timestamp 1676037725
transform 1 0 10580 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_115
timestamp 1676037725
transform 1 0 11684 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1676037725
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1676037725
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_141
timestamp 1676037725
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_146
timestamp 1676037725
transform 1 0 14536 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_152
timestamp 1676037725
transform 1 0 15088 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_158
timestamp 1676037725
transform 1 0 15640 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_168
timestamp 1676037725
transform 1 0 16560 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_174
timestamp 1676037725
transform 1 0 17112 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_181
timestamp 1676037725
transform 1 0 17756 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_188
timestamp 1676037725
transform 1 0 18400 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1676037725
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1676037725
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_204
timestamp 1676037725
transform 1 0 19872 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_216
timestamp 1676037725
transform 1 0 20976 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_222
timestamp 1676037725
transform 1 0 21528 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_229
timestamp 1676037725
transform 1 0 22172 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_235
timestamp 1676037725
transform 1 0 22724 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_243
timestamp 1676037725
transform 1 0 23460 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1676037725
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_15
timestamp 1676037725
transform 1 0 2484 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_35
timestamp 1676037725
transform 1 0 4324 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_47
timestamp 1676037725
transform 1 0 5428 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1676037725
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1676037725
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_69
timestamp 1676037725
transform 1 0 7452 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1676037725
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1676037725
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1676037725
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1676037725
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_125
timestamp 1676037725
transform 1 0 12604 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_136
timestamp 1676037725
transform 1 0 13616 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_148
timestamp 1676037725
transform 1 0 14720 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_154
timestamp 1676037725
transform 1 0 15272 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_160
timestamp 1676037725
transform 1 0 15824 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1676037725
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_169
timestamp 1676037725
transform 1 0 16652 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_175
timestamp 1676037725
transform 1 0 17204 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1676037725
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_193
timestamp 1676037725
transform 1 0 18860 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_199
timestamp 1676037725
transform 1 0 19412 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_211
timestamp 1676037725
transform 1 0 20516 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1676037725
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1676037725
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_225
timestamp 1676037725
transform 1 0 21804 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_235
timestamp 1676037725
transform 1 0 22724 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_243
timestamp 1676037725
transform 1 0 23460 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_3
timestamp 1676037725
transform 1 0 1380 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_9
timestamp 1676037725
transform 1 0 1932 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_26
timestamp 1676037725
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1676037725
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_41
timestamp 1676037725
transform 1 0 4876 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_49
timestamp 1676037725
transform 1 0 5612 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_53
timestamp 1676037725
transform 1 0 5980 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1676037725
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1676037725
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_85
timestamp 1676037725
transform 1 0 8924 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_103
timestamp 1676037725
transform 1 0 10580 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_115
timestamp 1676037725
transform 1 0 11684 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_127
timestamp 1676037725
transform 1 0 12788 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_136
timestamp 1676037725
transform 1 0 13616 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 1676037725
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_151
timestamp 1676037725
transform 1 0 14996 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_163
timestamp 1676037725
transform 1 0 16100 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_173
timestamp 1676037725
transform 1 0 17020 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_185
timestamp 1676037725
transform 1 0 18124 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1676037725
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_197
timestamp 1676037725
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_207
timestamp 1676037725
transform 1 0 20148 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_217
timestamp 1676037725
transform 1 0 21068 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_225
timestamp 1676037725
transform 1 0 21804 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_233
timestamp 1676037725
transform 1 0 22540 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_241
timestamp 1676037725
transform 1 0 23276 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1676037725
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_15
timestamp 1676037725
transform 1 0 2484 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_35
timestamp 1676037725
transform 1 0 4324 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_47
timestamp 1676037725
transform 1 0 5428 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1676037725
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_57
timestamp 1676037725
transform 1 0 6348 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_76
timestamp 1676037725
transform 1 0 8096 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_84
timestamp 1676037725
transform 1 0 8832 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_101
timestamp 1676037725
transform 1 0 10396 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_109
timestamp 1676037725
transform 1 0 11132 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1676037725
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1676037725
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_137
timestamp 1676037725
transform 1 0 13708 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_145
timestamp 1676037725
transform 1 0 14444 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_150
timestamp 1676037725
transform 1 0 14904 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_160
timestamp 1676037725
transform 1 0 15824 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_31_169
timestamp 1676037725
transform 1 0 16652 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_175
timestamp 1676037725
transform 1 0 17204 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_182
timestamp 1676037725
transform 1 0 17848 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_194
timestamp 1676037725
transform 1 0 18952 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_202
timestamp 1676037725
transform 1 0 19688 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_212
timestamp 1676037725
transform 1 0 20608 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_220
timestamp 1676037725
transform 1 0 21344 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1676037725
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_237
timestamp 1676037725
transform 1 0 22908 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_243
timestamp 1676037725
transform 1 0 23460 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_3
timestamp 1676037725
transform 1 0 1380 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_9
timestamp 1676037725
transform 1 0 1932 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_26
timestamp 1676037725
transform 1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1676037725
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_41
timestamp 1676037725
transform 1 0 4876 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_61
timestamp 1676037725
transform 1 0 6716 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_73
timestamp 1676037725
transform 1 0 7820 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_81
timestamp 1676037725
transform 1 0 8556 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_85
timestamp 1676037725
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_103
timestamp 1676037725
transform 1 0 10580 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_109
timestamp 1676037725
transform 1 0 11132 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_113
timestamp 1676037725
transform 1 0 11500 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_116
timestamp 1676037725
transform 1 0 11776 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_129
timestamp 1676037725
transform 1 0 12972 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_137
timestamp 1676037725
transform 1 0 13708 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_32_141
timestamp 1676037725
transform 1 0 14076 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_150
timestamp 1676037725
transform 1 0 14904 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_156
timestamp 1676037725
transform 1 0 15456 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_162
timestamp 1676037725
transform 1 0 16008 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_170
timestamp 1676037725
transform 1 0 16744 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_180
timestamp 1676037725
transform 1 0 17664 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_32_188
timestamp 1676037725
transform 1 0 18400 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_32_197
timestamp 1676037725
transform 1 0 19228 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_205
timestamp 1676037725
transform 1 0 19964 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_212
timestamp 1676037725
transform 1 0 20608 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_224
timestamp 1676037725
transform 1 0 21712 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_236
timestamp 1676037725
transform 1 0 22816 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1676037725
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_15
timestamp 1676037725
transform 1 0 2484 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_36
timestamp 1676037725
transform 1 0 4416 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_48
timestamp 1676037725
transform 1 0 5520 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1676037725
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1676037725
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_81
timestamp 1676037725
transform 1 0 8556 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_101
timestamp 1676037725
transform 1 0 10396 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_107
timestamp 1676037725
transform 1 0 10948 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1676037725
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_113
timestamp 1676037725
transform 1 0 11500 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_119
timestamp 1676037725
transform 1 0 12052 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_123
timestamp 1676037725
transform 1 0 12420 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_144
timestamp 1676037725
transform 1 0 14352 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_148
timestamp 1676037725
transform 1 0 14720 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_154
timestamp 1676037725
transform 1 0 15272 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_166
timestamp 1676037725
transform 1 0 16376 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_169
timestamp 1676037725
transform 1 0 16652 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_181
timestamp 1676037725
transform 1 0 17756 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_187
timestamp 1676037725
transform 1 0 18308 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_195
timestamp 1676037725
transform 1 0 19044 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_202
timestamp 1676037725
transform 1 0 19688 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_214
timestamp 1676037725
transform 1 0 20792 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_222
timestamp 1676037725
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1676037725
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_232
timestamp 1676037725
transform 1 0 22448 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_3
timestamp 1676037725
transform 1 0 1380 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_9
timestamp 1676037725
transform 1 0 1932 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_26
timestamp 1676037725
transform 1 0 3496 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_29
timestamp 1676037725
transform 1 0 3772 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_47
timestamp 1676037725
transform 1 0 5428 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_67
timestamp 1676037725
transform 1 0 7268 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_79
timestamp 1676037725
transform 1 0 8372 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1676037725
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_85
timestamp 1676037725
transform 1 0 8924 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_103
timestamp 1676037725
transform 1 0 10580 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_117
timestamp 1676037725
transform 1 0 11868 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_128
timestamp 1676037725
transform 1 0 12880 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_34_138
timestamp 1676037725
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_141
timestamp 1676037725
transform 1 0 14076 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_151
timestamp 1676037725
transform 1 0 14996 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_158
timestamp 1676037725
transform 1 0 15640 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_162
timestamp 1676037725
transform 1 0 16008 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_180
timestamp 1676037725
transform 1 0 17664 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_192
timestamp 1676037725
transform 1 0 18768 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1676037725
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_209
timestamp 1676037725
transform 1 0 20332 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_217
timestamp 1676037725
transform 1 0 21068 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_221
timestamp 1676037725
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_233
timestamp 1676037725
transform 1 0 22540 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_241
timestamp 1676037725
transform 1 0 23276 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1676037725
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_32
timestamp 1676037725
transform 1 0 4048 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 1676037725
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1676037725
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1676037725
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_81
timestamp 1676037725
transform 1 0 8556 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_101
timestamp 1676037725
transform 1 0 10396 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_107
timestamp 1676037725
transform 1 0 10948 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_110
timestamp 1676037725
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_113
timestamp 1676037725
transform 1 0 11500 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_122
timestamp 1676037725
transform 1 0 12328 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_132
timestamp 1676037725
transform 1 0 13248 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_136
timestamp 1676037725
transform 1 0 13616 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_143
timestamp 1676037725
transform 1 0 14260 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_147
timestamp 1676037725
transform 1 0 14628 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_155
timestamp 1676037725
transform 1 0 15364 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 1676037725
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_169
timestamp 1676037725
transform 1 0 16652 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_177
timestamp 1676037725
transform 1 0 17388 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_188
timestamp 1676037725
transform 1 0 18400 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_200
timestamp 1676037725
transform 1 0 19504 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_204
timestamp 1676037725
transform 1 0 19872 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_212
timestamp 1676037725
transform 1 0 20608 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_216
timestamp 1676037725
transform 1 0 20976 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_220
timestamp 1676037725
transform 1 0 21344 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1676037725
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_232
timestamp 1676037725
transform 1 0 22448 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1676037725
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1676037725
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1676037725
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1676037725
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1676037725
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_53
timestamp 1676037725
transform 1 0 5980 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_36_57
timestamp 1676037725
transform 1 0 6348 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_63
timestamp 1676037725
transform 1 0 6900 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_66
timestamp 1676037725
transform 1 0 7176 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_76
timestamp 1676037725
transform 1 0 8096 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_85
timestamp 1676037725
transform 1 0 8924 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_103
timestamp 1676037725
transform 1 0 10580 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_109
timestamp 1676037725
transform 1 0 11132 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_113
timestamp 1676037725
transform 1 0 11500 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_117
timestamp 1676037725
transform 1 0 11868 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_120
timestamp 1676037725
transform 1 0 12144 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_128
timestamp 1676037725
transform 1 0 12880 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_141
timestamp 1676037725
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_145
timestamp 1676037725
transform 1 0 14444 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_151
timestamp 1676037725
transform 1 0 14996 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_157
timestamp 1676037725
transform 1 0 15548 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_160
timestamp 1676037725
transform 1 0 15824 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_169
timestamp 1676037725
transform 1 0 16652 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_174
timestamp 1676037725
transform 1 0 17112 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_182
timestamp 1676037725
transform 1 0 17848 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_194
timestamp 1676037725
transform 1 0 18952 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1676037725
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_209
timestamp 1676037725
transform 1 0 20332 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_217
timestamp 1676037725
transform 1 0 21068 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_222
timestamp 1676037725
transform 1 0 21528 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_225
timestamp 1676037725
transform 1 0 21804 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_231
timestamp 1676037725
transform 1 0 22356 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_236
timestamp 1676037725
transform 1 0 22816 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 23828 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 23828 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 23828 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 23828 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 23828 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 23828 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 23828 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 23828 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 23828 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 23828 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 23828 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 23828 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 23828 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 23828 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 23828 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 23828 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1676037725
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1676037725
transform -1 0 23828 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1676037725
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1676037725
transform -1 0 23828 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1676037725
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1676037725
transform -1 0 23828 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1676037725
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1676037725
transform -1 0 23828 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1676037725
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1676037725
transform -1 0 23828 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1676037725
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1676037725
transform -1 0 23828 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1676037725
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1676037725
transform -1 0 23828 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1676037725
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1676037725
transform -1 0 23828 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1676037725
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1676037725
transform -1 0 23828 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1676037725
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1676037725
transform -1 0 23828 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1676037725
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1676037725
transform -1 0 23828 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1676037725
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1676037725
transform -1 0 23828 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1676037725
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1676037725
transform -1 0 23828 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1676037725
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1676037725
transform -1 0 23828 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1676037725
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1676037725
transform -1 0 23828 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1676037725
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1676037725
transform -1 0 23828 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1676037725
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1676037725
transform -1 0 23828 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1676037725
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1676037725
transform -1 0 23828 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1676037725
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1676037725
transform -1 0 23828 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1676037725
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1676037725
transform -1 0 23828 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1676037725
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1676037725
transform -1 0 23828 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1676037725
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1676037725
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1676037725
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1676037725
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1676037725
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1676037725
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1676037725
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1676037725
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1676037725
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1676037725
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1676037725
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1676037725
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1676037725
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1676037725
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1676037725
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1676037725
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1676037725
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1676037725
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1676037725
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1676037725
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1676037725
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1676037725
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1676037725
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1676037725
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1676037725
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1676037725
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1676037725
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1676037725
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1676037725
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1676037725
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1676037725
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1676037725
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1676037725
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1676037725
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1676037725
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1676037725
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1676037725
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1676037725
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1676037725
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1676037725
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1676037725
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1676037725
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1676037725
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1676037725
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1676037725
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1676037725
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1676037725
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1676037725
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1676037725
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1676037725
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1676037725
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1676037725
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1676037725
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1676037725
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1676037725
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1676037725
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1676037725
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1676037725
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1676037725
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1676037725
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1676037725
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1676037725
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1676037725
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1676037725
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1676037725
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1676037725
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1676037725
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1676037725
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1676037725
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1676037725
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1676037725
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1676037725
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1676037725
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1676037725
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1676037725
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1676037725
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1676037725
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1676037725
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1676037725
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1676037725
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1676037725
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1676037725
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1676037725
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1676037725
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1676037725
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1676037725
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1676037725
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1676037725
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1676037725
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1676037725
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1676037725
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1676037725
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1676037725
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1676037725
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1676037725
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1676037725
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1676037725
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1676037725
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1676037725
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1676037725
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1676037725
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1676037725
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1676037725
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1676037725
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1676037725
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1676037725
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1676037725
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1676037725
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1676037725
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1676037725
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1676037725
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1676037725
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1676037725
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1676037725
transform 1 0 6256 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1676037725
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1676037725
transform 1 0 11408 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1676037725
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1676037725
transform 1 0 16560 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1676037725
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1676037725
transform 1 0 21712 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__inv_6  _369_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4784 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _370_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 3956 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _371_
timestamp 1676037725
transform 1 0 5704 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _372_
timestamp 1676037725
transform -1 0 11132 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _373_
timestamp 1676037725
transform 1 0 15916 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _374_
timestamp 1676037725
transform 1 0 20424 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _375_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15732 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_8  _376_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7084 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__or2_4  _377_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5152 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _378_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3036 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or2_4  _379_
timestamp 1676037725
transform 1 0 6532 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _380_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 2576 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_4  _381_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3956 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__or3_4  _382_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5244 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _383_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 4416 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _384_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 4968 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _385_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 2300 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and2_4  _386_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 2944 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_4  _387_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5336 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nand2b_4  _388_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9108 0 1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_2  _389_
timestamp 1676037725
transform -1 0 2116 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand4b_4  _390_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1564 0 1 10880
box -38 -48 1786 592
use sky130_fd_sc_hd__nor3_4  _391_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 10948 0 1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_4  _392_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8648 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__or2_2  _393_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9016 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _394_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 2944 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _395_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 3496 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _396_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1748 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _397_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2024 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_4  _398_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 3588 0 -1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__and2_1  _399_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 16284 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3_4  _400_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 2668 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__nand3b_1  _401_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2116 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _402_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1656 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_4  _403_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11684 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__and4_4  _404_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4232 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _405_
timestamp 1676037725
transform 1 0 19964 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_2  _406_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 20148 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2_4  _407_
timestamp 1676037725
transform 1 0 2576 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _408_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 10672 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__a211oi_4  _409_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4876 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _410_
timestamp 1676037725
transform -1 0 11960 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_4  _411_
timestamp 1676037725
transform 1 0 8740 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nand2b_4  _412_
timestamp 1676037725
transform -1 0 7544 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__xor2_4  _413_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 8096 0 1 10880
box -38 -48 2062 592
use sky130_fd_sc_hd__nor2_1  _414_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 1932 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _415_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4324 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _416_
timestamp 1676037725
transform 1 0 4324 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and3_4  _417_
timestamp 1676037725
transform 1 0 6532 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_1  _418_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5244 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_4  _419_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5060 0 1 6528
box -38 -48 1326 592
use sky130_fd_sc_hd__a211o_4  _420_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 7636 0 1 4352
box -38 -48 1326 592
use sky130_fd_sc_hd__a31o_4  _421_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4508 0 1 3264
box -38 -48 1326 592
use sky130_fd_sc_hd__o221a_4  _422_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2024 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__a21oi_4  _423_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 8740 0 -1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _424_
timestamp 1676037725
transform -1 0 8556 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_1  _425_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 4692 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_2  _426_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 7452 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__o311ai_4  _427_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 17664 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__nor3_4  _428_
timestamp 1676037725
transform 1 0 6256 0 1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__or4_2  _429_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1840 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _430_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6992 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _431_
timestamp 1676037725
transform 1 0 5704 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_2  _432_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 5520 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _433_
timestamp 1676037725
transform 1 0 8372 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_4  _434_
timestamp 1676037725
transform -1 0 5888 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _435_
timestamp 1676037725
transform 1 0 20516 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_2  _436_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 20056 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a41oi_4  _437_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19412 0 1 3264
box -38 -48 2062 592
use sky130_fd_sc_hd__a41o_4  _438_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19504 0 -1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__nor2_1  _439_
timestamp 1676037725
transform -1 0 14904 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _440_
timestamp 1676037725
transform -1 0 15180 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _441_
timestamp 1676037725
transform -1 0 13800 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _442_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15916 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _443_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14260 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _444_
timestamp 1676037725
transform -1 0 13984 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _445_
timestamp 1676037725
transform -1 0 18860 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_4  _446_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 13156 0 -1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__nor3_2  _447_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11868 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_2  _448_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 7176 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _449_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9384 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _450_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 11868 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_2  _451_
timestamp 1676037725
transform -1 0 15272 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and3_4  _452_
timestamp 1676037725
transform 1 0 14904 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__or3_4  _453_
timestamp 1676037725
transform -1 0 12788 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _454_
timestamp 1676037725
transform -1 0 12236 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_4  _455_
timestamp 1676037725
transform 1 0 12236 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__clkinv_2  _456_
timestamp 1676037725
transform -1 0 21344 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_4  _457_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 15548 0 1 7616
box -38 -48 1326 592
use sky130_fd_sc_hd__a31o_2  _458_
timestamp 1676037725
transform -1 0 15364 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _459_
timestamp 1676037725
transform -1 0 13340 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_4  _460_
timestamp 1676037725
transform -1 0 18032 0 1 5440
box -38 -48 1326 592
use sky130_fd_sc_hd__nor2_4  _461_
timestamp 1676037725
transform -1 0 18952 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkinv_4  _462_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17756 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_4  _463_
timestamp 1676037725
transform -1 0 15272 0 -1 8704
box -38 -48 1326 592
use sky130_fd_sc_hd__o211a_4  _464_
timestamp 1676037725
transform -1 0 18492 0 -1 5440
box -38 -48 1326 592
use sky130_fd_sc_hd__nor2_8  _465_
timestamp 1676037725
transform 1 0 19044 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _466_
timestamp 1676037725
transform -1 0 14536 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _467_
timestamp 1676037725
transform 1 0 20884 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or3_4  _468_
timestamp 1676037725
transform 1 0 19504 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a2111o_4  _469_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16560 0 1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__and3_2  _470_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 18768 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or3_4  _471_
timestamp 1676037725
transform 1 0 19780 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_4  _472_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 20700 0 1 6528
box -38 -48 1326 592
use sky130_fd_sc_hd__a2bb2o_4  _473_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17296 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__nor2_2  _474_
timestamp 1676037725
transform -1 0 18584 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_2  _475_
timestamp 1676037725
transform 1 0 15088 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_4  _476_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11960 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _477_
timestamp 1676037725
transform 1 0 21528 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_4  _478_
timestamp 1676037725
transform 1 0 11776 0 1 13056
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_4  _479_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12604 0 -1 16320
box -38 -48 2062 592
use sky130_fd_sc_hd__nor2_1  _480_
timestamp 1676037725
transform -1 0 19688 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _481_
timestamp 1676037725
transform 1 0 21712 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_4  _482_
timestamp 1676037725
transform 1 0 13064 0 -1 11968
box -38 -48 1326 592
use sky130_fd_sc_hd__a21oi_1  _483_
timestamp 1676037725
transform -1 0 17204 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _484_
timestamp 1676037725
transform 1 0 14260 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _485_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16836 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _486_
timestamp 1676037725
transform 1 0 14260 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _487_
timestamp 1676037725
transform 1 0 19872 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o211ai_1  _488_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 17388 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _489_
timestamp 1676037725
transform -1 0 12052 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _490_
timestamp 1676037725
transform -1 0 11132 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _491_
timestamp 1676037725
transform 1 0 11684 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _492_
timestamp 1676037725
transform 1 0 12052 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _493_
timestamp 1676037725
transform 1 0 16560 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _494_
timestamp 1676037725
transform 1 0 16100 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or3_4  _495_
timestamp 1676037725
transform 1 0 17848 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _496_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 16376 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_4  _497_
timestamp 1676037725
transform -1 0 14720 0 -1 13056
box -38 -48 1326 592
use sky130_fd_sc_hd__nand2_2  _498_
timestamp 1676037725
transform -1 0 22448 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _499_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 21068 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _500_
timestamp 1676037725
transform -1 0 16652 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _501_
timestamp 1676037725
transform -1 0 10304 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_4  _502_
timestamp 1676037725
transform 1 0 9568 0 1 13056
box -38 -48 1326 592
use sky130_fd_sc_hd__inv_2  _503_
timestamp 1676037725
transform 1 0 12144 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_2  _504_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 19504 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _505_
timestamp 1676037725
transform 1 0 22356 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _506_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 20700 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _507_
timestamp 1676037725
transform 1 0 21528 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _508_
timestamp 1676037725
transform 1 0 21252 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _509_
timestamp 1676037725
transform 1 0 16928 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _510_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19412 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _511_
timestamp 1676037725
transform 1 0 19412 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _512_
timestamp 1676037725
transform 1 0 17112 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _513_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14352 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__and4_2  _514_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15548 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_4  _515_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 18400 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__a211o_1  _516_
timestamp 1676037725
transform -1 0 15180 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _517_
timestamp 1676037725
transform 1 0 15272 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _518_
timestamp 1676037725
transform 1 0 22908 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _519_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 23000 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _520_
timestamp 1676037725
transform -1 0 23000 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _521_
timestamp 1676037725
transform -1 0 23092 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _522_
timestamp 1676037725
transform -1 0 22632 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _523_
timestamp 1676037725
transform -1 0 21068 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _524_
timestamp 1676037725
transform -1 0 23276 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _525_
timestamp 1676037725
transform -1 0 21712 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _526_
timestamp 1676037725
transform -1 0 22632 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _527_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 22264 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _528_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 16192 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _529_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15640 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _530_
timestamp 1676037725
transform -1 0 22448 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _531_
timestamp 1676037725
transform 1 0 21620 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _532_
timestamp 1676037725
transform -1 0 21068 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _533_
timestamp 1676037725
transform -1 0 19872 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a311o_1  _534_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20424 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o32a_1  _535_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19872 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _536_
timestamp 1676037725
transform -1 0 19688 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _537_
timestamp 1676037725
transform 1 0 19780 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _538_
timestamp 1676037725
transform 1 0 18308 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _539_
timestamp 1676037725
transform 1 0 13984 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _540_
timestamp 1676037725
transform -1 0 13616 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _541_
timestamp 1676037725
transform -1 0 15640 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_4  _542_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 14352 0 -1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__a221o_1  _543_
timestamp 1676037725
transform 1 0 21988 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _544_
timestamp 1676037725
transform 1 0 19596 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _545_
timestamp 1676037725
transform 1 0 22080 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _546_
timestamp 1676037725
transform 1 0 21988 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _547_
timestamp 1676037725
transform 1 0 21988 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a22oi_4  _548_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16100 0 1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__o21a_1  _549_
timestamp 1676037725
transform -1 0 19780 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _550_
timestamp 1676037725
transform 1 0 21988 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _551_
timestamp 1676037725
transform -1 0 21160 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_1  _552_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 22724 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _553_
timestamp 1676037725
transform 1 0 22172 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_1  _554_
timestamp 1676037725
transform 1 0 20976 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _555_
timestamp 1676037725
transform 1 0 22356 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _556_
timestamp 1676037725
transform 1 0 21436 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_2  _557_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 23092 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__or3_1  _558_
timestamp 1676037725
transform 1 0 20700 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _559_
timestamp 1676037725
transform 1 0 20332 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _560_
timestamp 1676037725
transform 1 0 19320 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_4  _561_
timestamp 1676037725
transform 1 0 17020 0 -1 10880
box -38 -48 1326 592
use sky130_fd_sc_hd__a221o_1  _562_
timestamp 1676037725
transform 1 0 16836 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _563_
timestamp 1676037725
transform -1 0 17664 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _564_
timestamp 1676037725
transform 1 0 15364 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _565_
timestamp 1676037725
transform 1 0 16100 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _566_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 23184 0 1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__o22a_1  _567_
timestamp 1676037725
transform -1 0 18952 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _568_
timestamp 1676037725
transform 1 0 13064 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _569_
timestamp 1676037725
transform -1 0 17756 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _570_
timestamp 1676037725
transform 1 0 17204 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _571_
timestamp 1676037725
transform -1 0 17940 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _572_
timestamp 1676037725
transform 1 0 17204 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and3_4  _573_
timestamp 1676037725
transform 1 0 11868 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _574_
timestamp 1676037725
transform 1 0 19412 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_1  _575_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 17848 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _576_
timestamp 1676037725
transform 1 0 19044 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _577_
timestamp 1676037725
transform 1 0 14260 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _578_
timestamp 1676037725
transform 1 0 17664 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _579_
timestamp 1676037725
transform 1 0 16376 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _580_
timestamp 1676037725
transform 1 0 21068 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _581_
timestamp 1676037725
transform 1 0 20148 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _582_
timestamp 1676037725
transform 1 0 14904 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _583_
timestamp 1676037725
transform -1 0 14076 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _584_
timestamp 1676037725
transform -1 0 18952 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _585_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 17020 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a2111o_1  _586_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20332 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _587_
timestamp 1676037725
transform 1 0 15088 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _588_
timestamp 1676037725
transform 1 0 12604 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _589_
timestamp 1676037725
transform 1 0 11776 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _590_
timestamp 1676037725
transform 1 0 14260 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _591_
timestamp 1676037725
transform 1 0 14444 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o2111a_1  _592_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 15088 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__nor3_1  _593_
timestamp 1676037725
transform 1 0 14720 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _594_
timestamp 1676037725
transform -1 0 19780 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _595_
timestamp 1676037725
transform -1 0 13800 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _596_
timestamp 1676037725
transform -1 0 17664 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _597_
timestamp 1676037725
transform 1 0 18124 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _598_
timestamp 1676037725
transform 1 0 12604 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _599_
timestamp 1676037725
transform -1 0 12696 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _600_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 22264 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _601_
timestamp 1676037725
transform 1 0 18400 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_1  _602_
timestamp 1676037725
transform 1 0 14260 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _603_
timestamp 1676037725
transform 1 0 11316 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _604_
timestamp 1676037725
transform -1 0 12880 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _605_
timestamp 1676037725
transform -1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _606_
timestamp 1676037725
transform -1 0 13616 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _607_
timestamp 1676037725
transform 1 0 19412 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _608_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 16100 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _609_
timestamp 1676037725
transform -1 0 14904 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _610_
timestamp 1676037725
transform -1 0 15272 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _611_
timestamp 1676037725
transform -1 0 19780 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _612_
timestamp 1676037725
transform -1 0 20148 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _613_
timestamp 1676037725
transform 1 0 19136 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _614_
timestamp 1676037725
transform 1 0 20516 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _615_
timestamp 1676037725
transform 1 0 15640 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_1  _616_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15732 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _617_
timestamp 1676037725
transform 1 0 14720 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _618_
timestamp 1676037725
transform -1 0 18768 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _619_
timestamp 1676037725
transform 1 0 17664 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _620_
timestamp 1676037725
transform 1 0 17112 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _621_
timestamp 1676037725
transform 1 0 16468 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _622_
timestamp 1676037725
transform 1 0 16008 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _623_
timestamp 1676037725
transform 1 0 15456 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _624_
timestamp 1676037725
transform -1 0 14720 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _625_
timestamp 1676037725
transform -1 0 14904 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _626_
timestamp 1676037725
transform 1 0 14260 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _627_
timestamp 1676037725
transform 1 0 20056 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _628_
timestamp 1676037725
transform 1 0 17020 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _629_
timestamp 1676037725
transform 1 0 13432 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _630_
timestamp 1676037725
transform 1 0 12144 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _631_
timestamp 1676037725
transform -1 0 22448 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _632_
timestamp 1676037725
transform -1 0 21436 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _633_
timestamp 1676037725
transform -1 0 21344 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _634_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 20608 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _635_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 18400 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_4  _636_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10948 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _637_
timestamp 1676037725
transform 1 0 15732 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _638_
timestamp 1676037725
transform 1 0 8188 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _639_
timestamp 1676037725
transform -1 0 19136 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _640_
timestamp 1676037725
transform 1 0 16836 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _641_
timestamp 1676037725
transform 1 0 15640 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _642_
timestamp 1676037725
transform 1 0 16192 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _643_
timestamp 1676037725
transform 1 0 8740 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _644_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7728 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_1  _645_
timestamp 1676037725
transform 1 0 9200 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _646_
timestamp 1676037725
transform -1 0 9660 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _647_
timestamp 1676037725
transform -1 0 8556 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _648_
timestamp 1676037725
transform -1 0 10396 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _649_
timestamp 1676037725
transform -1 0 10764 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _650_
timestamp 1676037725
transform 1 0 14260 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _651_
timestamp 1676037725
transform 1 0 12788 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _652_
timestamp 1676037725
transform -1 0 11224 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _653_
timestamp 1676037725
transform 1 0 5060 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _654_
timestamp 1676037725
transform -1 0 2484 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _655_
timestamp 1676037725
transform 1 0 3312 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _656_
timestamp 1676037725
transform -1 0 8648 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _657_
timestamp 1676037725
transform -1 0 8188 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand3b_1  _658_
timestamp 1676037725
transform -1 0 8280 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _659_
timestamp 1676037725
transform -1 0 8648 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _660_
timestamp 1676037725
transform 1 0 7820 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _661_
timestamp 1676037725
transform 1 0 9108 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_4  _662_
timestamp 1676037725
transform 1 0 10120 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__a21o_2  _663_
timestamp 1676037725
transform -1 0 3496 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _664_
timestamp 1676037725
transform -1 0 10396 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _665_
timestamp 1676037725
transform 1 0 8924 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o2111a_1  _666_
timestamp 1676037725
transform -1 0 11224 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _667_
timestamp 1676037725
transform 1 0 18216 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _668_
timestamp 1676037725
transform 1 0 18032 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _669_
timestamp 1676037725
transform 1 0 15456 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _670_
timestamp 1676037725
transform 1 0 13708 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _671_
timestamp 1676037725
transform -1 0 13248 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _672_
timestamp 1676037725
transform -1 0 8372 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _673_
timestamp 1676037725
transform -1 0 11132 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_1  _674_
timestamp 1676037725
transform -1 0 11224 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_2  _675_
timestamp 1676037725
transform 1 0 10580 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__a41o_1  _676_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11684 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _677_
timestamp 1676037725
transform 1 0 10028 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _678_
timestamp 1676037725
transform 1 0 15180 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _679_
timestamp 1676037725
transform -1 0 10028 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _680_
timestamp 1676037725
transform -1 0 10304 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _681_
timestamp 1676037725
transform 1 0 8004 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _682_
timestamp 1676037725
transform -1 0 9844 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _683_
timestamp 1676037725
transform -1 0 10120 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _684_
timestamp 1676037725
transform -1 0 3312 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _685_
timestamp 1676037725
transform 1 0 3404 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _686_
timestamp 1676037725
transform -1 0 6900 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _687_
timestamp 1676037725
transform 1 0 6164 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _688_
timestamp 1676037725
transform 1 0 4784 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o21bai_1  _689_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14260 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _690_
timestamp 1676037725
transform 1 0 10580 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _691_
timestamp 1676037725
transform 1 0 10948 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _692_
timestamp 1676037725
transform 1 0 12420 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__o41a_1  _693_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 9936 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_1  _694_
timestamp 1676037725
transform 1 0 13064 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _695_
timestamp 1676037725
transform -1 0 13800 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _696_
timestamp 1676037725
transform 1 0 11684 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _697_
timestamp 1676037725
transform 1 0 10672 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _698_
timestamp 1676037725
transform -1 0 12420 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _699_
timestamp 1676037725
transform 1 0 11684 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _700_
timestamp 1676037725
transform 1 0 11684 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _701_
timestamp 1676037725
transform 1 0 3956 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _702_
timestamp 1676037725
transform 1 0 6808 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _703_
timestamp 1676037725
transform 1 0 6624 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _704_
timestamp 1676037725
transform -1 0 2576 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _705_
timestamp 1676037725
transform -1 0 2944 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _706_
timestamp 1676037725
transform 1 0 3956 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _707_
timestamp 1676037725
transform 1 0 8096 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _708_
timestamp 1676037725
transform 1 0 7084 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _709_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6164 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _710_
timestamp 1676037725
transform 1 0 5060 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _711_
timestamp 1676037725
transform -1 0 6440 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _712_
timestamp 1676037725
transform -1 0 7452 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _713_
timestamp 1676037725
transform -1 0 7452 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _714_
timestamp 1676037725
transform 1 0 8096 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _715_
timestamp 1676037725
transform -1 0 9752 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _716_
timestamp 1676037725
transform -1 0 4692 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _717_
timestamp 1676037725
transform -1 0 3496 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a31oi_1  _718_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 2484 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _719_
timestamp 1676037725
transform 1 0 1564 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _720_
timestamp 1676037725
transform 1 0 1564 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _721_
timestamp 1676037725
transform -1 0 2944 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _722_
timestamp 1676037725
transform -1 0 4048 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _723_
timestamp 1676037725
transform 1 0 3956 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _724_
timestamp 1676037725
transform -1 0 5428 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _725_
timestamp 1676037725
transform -1 0 3496 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _726_
timestamp 1676037725
transform -1 0 2208 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _727_
timestamp 1676037725
transform 1 0 2116 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _728_
timestamp 1676037725
transform 1 0 4232 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _729_
timestamp 1676037725
transform 1 0 6532 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _730_
timestamp 1676037725
transform 1 0 2024 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _731_
timestamp 1676037725
transform -1 0 2484 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _732_
timestamp 1676037725
transform -1 0 4784 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _733_
timestamp 1676037725
transform -1 0 12788 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o221ai_4  _734_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 8648 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__a32o_1  _735_
timestamp 1676037725
transform 1 0 12604 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _736_
timestamp 1676037725
transform 1 0 4784 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _737_
timestamp 1676037725
transform -1 0 6808 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _738_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 8096 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _739_
timestamp 1676037725
transform -1 0 6716 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _740_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2024 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _741_
timestamp 1676037725
transform -1 0 7176 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _742_
timestamp 1676037725
transform -1 0 10580 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _743_
timestamp 1676037725
transform -1 0 10396 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _744_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2668 0 -1 17408
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _745_
timestamp 1676037725
transform 1 0 2668 0 -1 15232
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _746_
timestamp 1676037725
transform 1 0 7084 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _747_
timestamp 1676037725
transform 1 0 9108 0 1 16320
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _748_
timestamp 1676037725
transform -1 0 9752 0 -1 15232
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _749_
timestamp 1676037725
transform 1 0 8832 0 -1 17408
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _750_
timestamp 1676037725
transform 1 0 8924 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _751_
timestamp 1676037725
transform 1 0 9108 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _752_
timestamp 1676037725
transform 1 0 9108 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _753_
timestamp 1676037725
transform 1 0 2024 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _754_
timestamp 1676037725
transform 1 0 2576 0 -1 18496
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _755_
timestamp 1676037725
transform 1 0 8188 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _756_
timestamp 1676037725
transform 1 0 4600 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _757_
timestamp 1676037725
transform 1 0 9108 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _758_
timestamp 1676037725
transform 1 0 9108 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _759_
timestamp 1676037725
transform 1 0 5796 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _760_
timestamp 1676037725
transform 1 0 9108 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _761_
timestamp 1676037725
transform 1 0 8924 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _762_
timestamp 1676037725
transform 1 0 4968 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _763_
timestamp 1676037725
transform -1 0 3496 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _764_
timestamp 1676037725
transform 1 0 2576 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _765_
timestamp 1676037725
transform 1 0 2484 0 -1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _766_
timestamp 1676037725
transform 1 0 2852 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _767_
timestamp 1676037725
transform -1 0 6716 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _768_
timestamp 1676037725
transform 1 0 2024 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _769_
timestamp 1676037725
transform -1 0 5428 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _770_
timestamp 1676037725
transform 1 0 2024 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_2  _798_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 4416 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6348 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1676037725
transform -1 0 4416 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1676037725
transform -1 0 4416 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1676037725
transform 1 0 7820 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1676037725
transform 1 0 7820 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_4  fanout13 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 14260 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout14
timestamp 1676037725
transform 1 0 15548 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 13248 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout16
timestamp 1676037725
transform -1 0 23184 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout17 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 22356 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout18
timestamp 1676037725
transform 1 0 22724 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout19
timestamp 1676037725
transform 1 0 15272 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout20
timestamp 1676037725
transform -1 0 21160 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout21
timestamp 1676037725
transform -1 0 20608 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout22
timestamp 1676037725
transform 1 0 21344 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout23
timestamp 1676037725
transform 1 0 20976 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout24 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19780 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout25
timestamp 1676037725
transform 1 0 22080 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout26
timestamp 1676037725
transform -1 0 15548 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout27
timestamp 1676037725
transform 1 0 13800 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  fanout28 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18768 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  fanout29
timestamp 1676037725
transform -1 0 10396 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout30
timestamp 1676037725
transform -1 0 4692 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout31
timestamp 1676037725
transform 1 0 2760 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout32
timestamp 1676037725
transform -1 0 3036 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  fanout33 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4324 0 -1 5440
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  fanout34
timestamp 1676037725
transform -1 0 3404 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout35
timestamp 1676037725
transform -1 0 5612 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout36
timestamp 1676037725
transform 1 0 6624 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout37
timestamp 1676037725
transform -1 0 3496 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  fanout38
timestamp 1676037725
transform 1 0 4784 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout39
timestamp 1676037725
transform 1 0 5060 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout40
timestamp 1676037725
transform 1 0 3956 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout41
timestamp 1676037725
transform -1 0 5428 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout42
timestamp 1676037725
transform 1 0 3956 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout43
timestamp 1676037725
transform -1 0 3496 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout44
timestamp 1676037725
transform -1 0 2760 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout45
timestamp 1676037725
transform 1 0 12420 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout46
timestamp 1676037725
transform 1 0 7820 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout47
timestamp 1676037725
transform -1 0 3496 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1676037725
transform 1 0 12512 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1676037725
transform 1 0 17480 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1676037725
transform -1 0 22816 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input4
timestamp 1676037725
transform 1 0 7544 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output5
timestamp 1676037725
transform 1 0 7452 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output6
timestamp 1676037725
transform -1 0 3496 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output7
timestamp 1676037725
transform -1 0 2576 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output8
timestamp 1676037725
transform -1 0 3588 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output9
timestamp 1676037725
transform -1 0 4692 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output10
timestamp 1676037725
transform -1 0 3496 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output11
timestamp 1676037725
transform -1 0 7084 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output12
timestamp 1676037725
transform -1 0 7084 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_48 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 10580 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_49
timestamp 1676037725
transform -1 0 9292 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_50
timestamp 1676037725
transform -1 0 8280 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_51
timestamp 1676037725
transform 1 0 7636 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_52
timestamp 1676037725
transform 1 0 8372 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_53
timestamp 1676037725
transform 1 0 9660 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_54
timestamp 1676037725
transform 1 0 10304 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_55
timestamp 1676037725
transform 1 0 10948 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_56
timestamp 1676037725
transform -1 0 12144 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_57
timestamp 1676037725
transform -1 0 12788 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_58
timestamp 1676037725
transform -1 0 13432 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_59
timestamp 1676037725
transform -1 0 14536 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_60
timestamp 1676037725
transform -1 0 15180 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_61
timestamp 1676037725
transform -1 0 15824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_62
timestamp 1676037725
transform -1 0 17112 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_63
timestamp 1676037725
transform -1 0 17756 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_64
timestamp 1676037725
transform -1 0 18400 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_65
timestamp 1676037725
transform -1 0 19688 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_66
timestamp 1676037725
transform -1 0 19412 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_67
timestamp 1676037725
transform -1 0 20332 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_68
timestamp 1676037725
transform -1 0 20976 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_69
timestamp 1676037725
transform -1 0 21068 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_70
timestamp 1676037725
transform -1 0 22264 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_71
timestamp 1676037725
transform -1 0 22264 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_72
timestamp 1676037725
transform -1 0 22908 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_73
timestamp 1676037725
transform -1 0 23092 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_74
timestamp 1676037725
transform 1 0 23092 0 1 3264
box -38 -48 314 592
<< labels >>
flabel metal2 s 2502 24200 2558 25000 0 FreeSans 224 90 0 0 clk
port 0 nsew signal input
flabel metal2 s 12438 24200 12494 25000 0 FreeSans 224 90 0 0 io_in[0]
port 1 nsew signal input
flabel metal2 s 17406 24200 17462 25000 0 FreeSans 224 90 0 0 io_in[1]
port 2 nsew signal input
flabel metal2 s 22374 24200 22430 25000 0 FreeSans 224 90 0 0 io_in[2]
port 3 nsew signal input
flabel metal2 s 6642 0 6698 800 0 FreeSans 224 90 0 0 io_oeb[0]
port 4 nsew signal tristate
flabel metal2 s 13082 0 13138 800 0 FreeSans 224 90 0 0 io_oeb[10]
port 5 nsew signal tristate
flabel metal2 s 13726 0 13782 800 0 FreeSans 224 90 0 0 io_oeb[11]
port 6 nsew signal tristate
flabel metal2 s 14370 0 14426 800 0 FreeSans 224 90 0 0 io_oeb[12]
port 7 nsew signal tristate
flabel metal2 s 15014 0 15070 800 0 FreeSans 224 90 0 0 io_oeb[13]
port 8 nsew signal tristate
flabel metal2 s 15658 0 15714 800 0 FreeSans 224 90 0 0 io_oeb[14]
port 9 nsew signal tristate
flabel metal2 s 16302 0 16358 800 0 FreeSans 224 90 0 0 io_oeb[15]
port 10 nsew signal tristate
flabel metal2 s 16946 0 17002 800 0 FreeSans 224 90 0 0 io_oeb[16]
port 11 nsew signal tristate
flabel metal2 s 17590 0 17646 800 0 FreeSans 224 90 0 0 io_oeb[17]
port 12 nsew signal tristate
flabel metal2 s 18234 0 18290 800 0 FreeSans 224 90 0 0 io_oeb[18]
port 13 nsew signal tristate
flabel metal2 s 18878 0 18934 800 0 FreeSans 224 90 0 0 io_oeb[19]
port 14 nsew signal tristate
flabel metal2 s 7286 0 7342 800 0 FreeSans 224 90 0 0 io_oeb[1]
port 15 nsew signal tristate
flabel metal2 s 19522 0 19578 800 0 FreeSans 224 90 0 0 io_oeb[20]
port 16 nsew signal tristate
flabel metal2 s 20166 0 20222 800 0 FreeSans 224 90 0 0 io_oeb[21]
port 17 nsew signal tristate
flabel metal2 s 20810 0 20866 800 0 FreeSans 224 90 0 0 io_oeb[22]
port 18 nsew signal tristate
flabel metal2 s 21454 0 21510 800 0 FreeSans 224 90 0 0 io_oeb[23]
port 19 nsew signal tristate
flabel metal2 s 22098 0 22154 800 0 FreeSans 224 90 0 0 io_oeb[24]
port 20 nsew signal tristate
flabel metal2 s 22742 0 22798 800 0 FreeSans 224 90 0 0 io_oeb[25]
port 21 nsew signal tristate
flabel metal2 s 23386 0 23442 800 0 FreeSans 224 90 0 0 io_oeb[26]
port 22 nsew signal tristate
flabel metal2 s 7930 0 7986 800 0 FreeSans 224 90 0 0 io_oeb[2]
port 23 nsew signal tristate
flabel metal2 s 8574 0 8630 800 0 FreeSans 224 90 0 0 io_oeb[3]
port 24 nsew signal tristate
flabel metal2 s 9218 0 9274 800 0 FreeSans 224 90 0 0 io_oeb[4]
port 25 nsew signal tristate
flabel metal2 s 9862 0 9918 800 0 FreeSans 224 90 0 0 io_oeb[5]
port 26 nsew signal tristate
flabel metal2 s 10506 0 10562 800 0 FreeSans 224 90 0 0 io_oeb[6]
port 27 nsew signal tristate
flabel metal2 s 11150 0 11206 800 0 FreeSans 224 90 0 0 io_oeb[7]
port 28 nsew signal tristate
flabel metal2 s 11794 0 11850 800 0 FreeSans 224 90 0 0 io_oeb[8]
port 29 nsew signal tristate
flabel metal2 s 12438 0 12494 800 0 FreeSans 224 90 0 0 io_oeb[9]
port 30 nsew signal tristate
flabel metal2 s 1490 0 1546 800 0 FreeSans 224 90 0 0 io_out[0]
port 31 nsew signal tristate
flabel metal2 s 2134 0 2190 800 0 FreeSans 224 90 0 0 io_out[1]
port 32 nsew signal tristate
flabel metal2 s 2778 0 2834 800 0 FreeSans 224 90 0 0 io_out[2]
port 33 nsew signal tristate
flabel metal2 s 3422 0 3478 800 0 FreeSans 224 90 0 0 io_out[3]
port 34 nsew signal tristate
flabel metal2 s 4066 0 4122 800 0 FreeSans 224 90 0 0 io_out[4]
port 35 nsew signal tristate
flabel metal2 s 4710 0 4766 800 0 FreeSans 224 90 0 0 io_out[5]
port 36 nsew signal tristate
flabel metal2 s 5354 0 5410 800 0 FreeSans 224 90 0 0 io_out[6]
port 37 nsew signal tristate
flabel metal2 s 5998 0 6054 800 0 FreeSans 224 90 0 0 io_out[7]
port 38 nsew signal tristate
flabel metal2 s 7470 24200 7526 25000 0 FreeSans 224 90 0 0 rst
port 39 nsew signal input
flabel metal4 s 3784 2128 4104 22352 0 FreeSans 1920 90 0 0 vccd1
port 40 nsew power bidirectional
flabel metal4 s 9465 2128 9785 22352 0 FreeSans 1920 90 0 0 vccd1
port 40 nsew power bidirectional
flabel metal4 s 15146 2128 15466 22352 0 FreeSans 1920 90 0 0 vccd1
port 40 nsew power bidirectional
flabel metal4 s 20827 2128 21147 22352 0 FreeSans 1920 90 0 0 vccd1
port 40 nsew power bidirectional
flabel metal4 s 6624 2128 6944 22352 0 FreeSans 1920 90 0 0 vssd1
port 41 nsew ground bidirectional
flabel metal4 s 12305 2128 12625 22352 0 FreeSans 1920 90 0 0 vssd1
port 41 nsew ground bidirectional
flabel metal4 s 17986 2128 18306 22352 0 FreeSans 1920 90 0 0 vssd1
port 41 nsew ground bidirectional
flabel metal4 s 23667 2128 23987 22352 0 FreeSans 1920 90 0 0 vssd1
port 41 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 25000 25000
<< end >>
