VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_vgatest
  CLASS BLOCK ;
  FOREIGN wrapped_vgatest ;
  ORIGIN 0.000 0.000 ;
  SIZE 375.000 BY 375.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 371.000 17.850 375.000 ;
    END
  END clk
  PIN io_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 371.000 187.040 375.000 187.640 ;
    END
  END io_in
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 371.000 79.490 375.000 ;
    END
  END io_out[0]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.030 371.000 110.310 375.000 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.850 371.000 141.130 375.000 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.670 371.000 171.950 375.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.490 371.000 202.770 375.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.310 371.000 233.590 375.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 371.000 264.410 375.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.950 371.000 295.230 375.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.770 371.000 326.050 375.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.590 371.000 356.870 375.000 ;
    END
  END io_out[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 371.000 48.670 375.000 ;
    END
  END rst
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 362.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 362.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 362.000 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 362.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 362.000 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 369.380 361.845 ;
      LAYER met1 ;
        RECT 3.290 10.640 369.380 362.000 ;
      LAYER met2 ;
        RECT 3.320 370.720 17.290 371.690 ;
        RECT 18.130 370.720 48.110 371.690 ;
        RECT 48.950 370.720 78.930 371.690 ;
        RECT 79.770 370.720 109.750 371.690 ;
        RECT 110.590 370.720 140.570 371.690 ;
        RECT 141.410 370.720 171.390 371.690 ;
        RECT 172.230 370.720 202.210 371.690 ;
        RECT 203.050 370.720 233.030 371.690 ;
        RECT 233.870 370.720 263.850 371.690 ;
        RECT 264.690 370.720 294.670 371.690 ;
        RECT 295.510 370.720 325.490 371.690 ;
        RECT 326.330 370.720 356.310 371.690 ;
        RECT 357.150 370.720 364.680 371.690 ;
        RECT 3.320 10.695 364.680 370.720 ;
      LAYER met3 ;
        RECT 3.745 188.040 371.000 361.925 ;
        RECT 3.745 186.640 370.600 188.040 ;
        RECT 3.745 10.715 371.000 186.640 ;
      LAYER met4 ;
        RECT 4.895 23.295 20.640 300.385 ;
        RECT 23.040 23.295 97.440 300.385 ;
        RECT 99.840 23.295 174.240 300.385 ;
        RECT 176.640 23.295 251.040 300.385 ;
        RECT 253.440 23.295 327.840 300.385 ;
        RECT 330.240 23.295 352.985 300.385 ;
  END
END wrapped_vgatest
END LIBRARY

