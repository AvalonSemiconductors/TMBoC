magic
tech sky130B
magscale 1 2
timestamp 1674824271
<< nwell >>
rect 1066 16581 18898 17147
rect 1066 15493 18898 16059
rect 1066 14405 18898 14971
rect 1066 13317 18898 13883
rect 1066 12229 18898 12795
rect 1066 11141 18898 11707
rect 1066 10053 18898 10619
rect 1066 8965 18898 9531
rect 1066 7877 18898 8443
rect 1066 6789 18898 7355
rect 1066 5701 18898 6267
rect 1066 4613 18898 5179
rect 1066 3525 18898 4091
rect 1066 2437 18898 3003
<< obsli1 >>
rect 1104 2159 18860 17425
<< obsm1 >>
rect 1104 2128 19019 17456
<< metal2 >>
rect 3330 19200 3386 20000
rect 9954 19200 10010 20000
rect 16578 19200 16634 20000
rect 1214 0 1270 800
rect 3698 0 3754 800
rect 6182 0 6238 800
rect 8666 0 8722 800
rect 11150 0 11206 800
rect 13634 0 13690 800
rect 16118 0 16174 800
rect 18602 0 18658 800
<< obsm2 >>
rect 1216 19144 3274 19258
rect 3442 19144 9898 19258
rect 10066 19144 16522 19258
rect 16690 19144 19013 19258
rect 1216 856 19013 19144
rect 1326 800 3642 856
rect 3810 800 6126 856
rect 6294 800 8610 856
rect 8778 800 11094 856
rect 11262 800 13578 856
rect 13746 800 16062 856
rect 16230 800 18546 856
rect 18714 800 19013 856
<< obsm3 >>
rect 3165 2143 19017 17441
<< metal4 >>
rect 3163 2128 3483 17456
rect 5382 2128 5702 17456
rect 7602 2128 7922 17456
rect 9821 2128 10141 17456
rect 12041 2128 12361 17456
rect 14260 2128 14580 17456
rect 16480 2128 16800 17456
rect 18699 2128 19019 17456
<< labels >>
rlabel metal2 s 3330 19200 3386 20000 6 clk
port 1 nsew signal input
rlabel metal2 s 16578 19200 16634 20000 6 io_in
port 2 nsew signal input
rlabel metal2 s 1214 0 1270 800 6 io_out[0]
port 3 nsew signal output
rlabel metal2 s 3698 0 3754 800 6 io_out[1]
port 4 nsew signal output
rlabel metal2 s 6182 0 6238 800 6 io_out[2]
port 5 nsew signal output
rlabel metal2 s 8666 0 8722 800 6 io_out[3]
port 6 nsew signal output
rlabel metal2 s 11150 0 11206 800 6 io_out[4]
port 7 nsew signal output
rlabel metal2 s 13634 0 13690 800 6 io_out[5]
port 8 nsew signal output
rlabel metal2 s 16118 0 16174 800 6 io_out[6]
port 9 nsew signal output
rlabel metal2 s 18602 0 18658 800 6 io_out[7]
port 10 nsew signal output
rlabel metal2 s 9954 19200 10010 20000 6 rst
port 11 nsew signal input
rlabel metal4 s 3163 2128 3483 17456 6 vccd1
port 12 nsew power bidirectional
rlabel metal4 s 7602 2128 7922 17456 6 vccd1
port 12 nsew power bidirectional
rlabel metal4 s 12041 2128 12361 17456 6 vccd1
port 12 nsew power bidirectional
rlabel metal4 s 16480 2128 16800 17456 6 vccd1
port 12 nsew power bidirectional
rlabel metal4 s 5382 2128 5702 17456 6 vssd1
port 13 nsew ground bidirectional
rlabel metal4 s 9821 2128 10141 17456 6 vssd1
port 13 nsew ground bidirectional
rlabel metal4 s 14260 2128 14580 17456 6 vssd1
port 13 nsew ground bidirectional
rlabel metal4 s 18699 2128 19019 17456 6 vssd1
port 13 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 20000 20000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1280348
string GDS_FILE /media/lucah/e6042058-84c8-448b-be8a-b40bc065b34b/TMBoC/openlane/Diceroll/runs/23_01_27_13_55/results/signoff/tt2_tholin_diceroll.magic.gds
string GDS_START 392556
<< end >>

