magic
tech sky130B
magscale 1 2
timestamp 1674824269
<< viali >>
rect 5825 17289 5859 17323
rect 16313 17289 16347 17323
rect 5120 17221 5154 17255
rect 12357 17221 12391 17255
rect 3065 17153 3099 17187
rect 6009 17153 6043 17187
rect 6745 17153 6779 17187
rect 9321 17153 9355 17187
rect 10057 17153 10091 17187
rect 10241 17153 10275 17187
rect 11069 17153 11103 17187
rect 11897 17153 11931 17187
rect 16865 17153 16899 17187
rect 5365 17085 5399 17119
rect 6929 17085 6963 17119
rect 17141 17085 17175 17119
rect 3249 17017 3283 17051
rect 10885 17017 10919 17051
rect 3985 16949 4019 16983
rect 6561 16949 6595 16983
rect 7389 16949 7423 16983
rect 9137 16949 9171 16983
rect 10425 16949 10459 16983
rect 11713 16949 11747 16983
rect 12909 16949 12943 16983
rect 2789 16745 2823 16779
rect 7205 16745 7239 16779
rect 9781 16745 9815 16779
rect 12633 16745 12667 16779
rect 10425 16609 10459 16643
rect 3157 16541 3191 16575
rect 5365 16541 5399 16575
rect 8585 16541 8619 16575
rect 2973 16473 3007 16507
rect 5632 16473 5666 16507
rect 8340 16473 8374 16507
rect 9873 16473 9907 16507
rect 10692 16473 10726 16507
rect 12265 16473 12299 16507
rect 12449 16473 12483 16507
rect 13093 16473 13127 16507
rect 3985 16405 4019 16439
rect 6745 16405 6779 16439
rect 11805 16405 11839 16439
rect 5825 16201 5859 16235
rect 6561 16201 6595 16235
rect 8217 16201 8251 16235
rect 10057 16201 10091 16235
rect 10701 16201 10735 16235
rect 4270 16133 4304 16167
rect 6745 16133 6779 16167
rect 6929 16133 6963 16167
rect 13982 16133 14016 16167
rect 6009 16065 6043 16099
rect 8033 16065 8067 16099
rect 8677 16065 8711 16099
rect 8944 16065 8978 16099
rect 10517 16065 10551 16099
rect 11897 16065 11931 16099
rect 12081 16065 12115 16099
rect 12173 16065 12207 16099
rect 12265 16065 12299 16099
rect 13001 16065 13035 16099
rect 13185 16065 13219 16099
rect 4537 15997 4571 16031
rect 7849 15997 7883 16031
rect 13093 15997 13127 16031
rect 13737 15997 13771 16031
rect 12541 15929 12575 15963
rect 3157 15861 3191 15895
rect 15117 15861 15151 15895
rect 12081 15657 12115 15691
rect 3433 15521 3467 15555
rect 3249 15453 3283 15487
rect 4169 15453 4203 15487
rect 4261 15453 4295 15487
rect 5273 15453 5307 15487
rect 7113 15453 7147 15487
rect 9505 15453 9539 15487
rect 12081 15453 12115 15487
rect 12265 15453 12299 15487
rect 12817 15453 12851 15487
rect 12909 15453 12943 15487
rect 5540 15385 5574 15419
rect 7380 15385 7414 15419
rect 9772 15385 9806 15419
rect 14565 15385 14599 15419
rect 14749 15385 14783 15419
rect 3065 15317 3099 15351
rect 3985 15317 4019 15351
rect 6653 15317 6687 15351
rect 8493 15317 8527 15351
rect 10885 15317 10919 15351
rect 14933 15317 14967 15351
rect 15761 15317 15795 15351
rect 4353 15113 4387 15147
rect 7481 15113 7515 15147
rect 9413 15113 9447 15147
rect 10241 15113 10275 15147
rect 15853 15113 15887 15147
rect 17141 15045 17175 15079
rect 2973 14977 3007 15011
rect 3229 14977 3263 15011
rect 6653 14977 6687 15011
rect 6837 14977 6871 15011
rect 7021 14977 7055 15011
rect 7665 14977 7699 15011
rect 9229 14977 9263 15011
rect 9873 14977 9907 15011
rect 10057 14977 10091 15011
rect 10885 14977 10919 15011
rect 12256 14977 12290 15011
rect 14096 14977 14130 15011
rect 16313 14977 16347 15011
rect 16957 14977 16991 15011
rect 17049 14977 17083 15011
rect 17233 14977 17267 15011
rect 11989 14909 12023 14943
rect 13829 14909 13863 14943
rect 17417 14909 17451 14943
rect 15209 14841 15243 14875
rect 5733 14773 5767 14807
rect 8677 14773 8711 14807
rect 10793 14773 10827 14807
rect 13369 14773 13403 14807
rect 16221 14773 16255 14807
rect 6469 14569 6503 14603
rect 12357 14569 12391 14603
rect 13185 14569 13219 14603
rect 5549 14501 5583 14535
rect 6101 14501 6135 14535
rect 14473 14501 14507 14535
rect 12817 14433 12851 14467
rect 16221 14433 16255 14467
rect 16405 14433 16439 14467
rect 17601 14433 17635 14467
rect 3249 14365 3283 14399
rect 4169 14365 4203 14399
rect 6009 14365 6043 14399
rect 6285 14365 6319 14399
rect 6929 14365 6963 14399
rect 9137 14365 9171 14399
rect 11069 14365 11103 14399
rect 11253 14365 11287 14399
rect 11713 14365 11747 14399
rect 11897 14365 11931 14399
rect 11989 14365 12023 14399
rect 12081 14365 12115 14399
rect 13277 14365 13311 14399
rect 14381 14365 14415 14399
rect 14657 14365 14691 14399
rect 16129 14365 16163 14399
rect 17116 14365 17150 14399
rect 4414 14297 4448 14331
rect 7174 14297 7208 14331
rect 9382 14297 9416 14331
rect 11161 14297 11195 14331
rect 17325 14297 17359 14331
rect 3433 14229 3467 14263
rect 8309 14229 8343 14263
rect 10517 14229 10551 14263
rect 14841 14229 14875 14263
rect 15761 14229 15795 14263
rect 16957 14229 16991 14263
rect 17233 14229 17267 14263
rect 3065 14025 3099 14059
rect 5371 14025 5405 14059
rect 7021 14025 7055 14059
rect 9229 14025 9263 14059
rect 9873 14025 9907 14059
rect 12633 14025 12667 14059
rect 14933 14025 14967 14059
rect 15945 14025 15979 14059
rect 17049 14025 17083 14059
rect 18061 14025 18095 14059
rect 5457 13957 5491 13991
rect 12541 13957 12575 13991
rect 2329 13889 2363 13923
rect 2513 13889 2547 13923
rect 4178 13889 4212 13923
rect 5273 13889 5307 13923
rect 5549 13889 5583 13923
rect 7297 13889 7331 13923
rect 7389 13889 7423 13923
rect 7481 13889 7515 13923
rect 7665 13889 7699 13923
rect 8585 13889 8619 13923
rect 8769 13889 8803 13923
rect 9045 13889 9079 13923
rect 10241 13889 10275 13923
rect 13737 13889 13771 13923
rect 14197 13889 14231 13923
rect 14381 13889 14415 13923
rect 14841 13889 14875 13923
rect 15025 13889 15059 13923
rect 16313 13889 16347 13923
rect 17417 13889 17451 13923
rect 17877 13889 17911 13923
rect 2605 13821 2639 13855
rect 4445 13821 4479 13855
rect 10057 13821 10091 13855
rect 10149 13821 10183 13855
rect 10333 13821 10367 13855
rect 12357 13821 12391 13855
rect 16221 13821 16255 13855
rect 2145 13753 2179 13787
rect 10885 13685 10919 13719
rect 13001 13685 13035 13719
rect 14381 13685 14415 13719
rect 16313 13685 16347 13719
rect 16865 13685 16899 13719
rect 17049 13685 17083 13719
rect 2421 13481 2455 13515
rect 3249 13481 3283 13515
rect 7573 13481 7607 13515
rect 9137 13481 9171 13515
rect 10057 13481 10091 13515
rect 18061 13481 18095 13515
rect 10149 13413 10183 13447
rect 10057 13345 10091 13379
rect 12265 13345 12299 13379
rect 2421 13277 2455 13311
rect 2697 13277 2731 13311
rect 5641 13277 5675 13311
rect 7481 13277 7515 13311
rect 7665 13277 7699 13311
rect 8401 13277 8435 13311
rect 8585 13277 8619 13311
rect 9321 13277 9355 13311
rect 9413 13277 9447 13311
rect 10333 13277 10367 13311
rect 10885 13277 10919 13311
rect 12173 13277 12207 13311
rect 14289 13277 14323 13311
rect 14545 13277 14579 13311
rect 16773 13277 16807 13311
rect 17601 13277 17635 13311
rect 18061 13277 18095 13311
rect 18245 13277 18279 13311
rect 2605 13209 2639 13243
rect 5908 13209 5942 13243
rect 10425 13209 10459 13243
rect 16589 13209 16623 13243
rect 16957 13209 16991 13243
rect 7021 13141 7055 13175
rect 8493 13141 8527 13175
rect 11069 13141 11103 13175
rect 12541 13141 12575 13175
rect 15669 13141 15703 13175
rect 17509 13141 17543 13175
rect 2697 12937 2731 12971
rect 5825 12937 5859 12971
rect 8309 12937 8343 12971
rect 10609 12937 10643 12971
rect 14197 12937 14231 12971
rect 14749 12937 14783 12971
rect 14933 12937 14967 12971
rect 10149 12869 10183 12903
rect 2237 12801 2271 12835
rect 2513 12801 2547 12835
rect 4730 12801 4764 12835
rect 6009 12801 6043 12835
rect 7205 12801 7239 12835
rect 9597 12801 9631 12835
rect 10333 12801 10367 12835
rect 10425 12801 10459 12835
rect 11713 12801 11747 12835
rect 11897 12801 11931 12835
rect 14930 12801 14964 12835
rect 15945 12801 15979 12835
rect 16129 12801 16163 12835
rect 17417 12801 17451 12835
rect 4997 12733 5031 12767
rect 7021 12733 7055 12767
rect 15301 12733 15335 12767
rect 15393 12733 15427 12767
rect 17325 12733 17359 12767
rect 2329 12665 2363 12699
rect 3617 12665 3651 12699
rect 17049 12665 17083 12699
rect 7389 12597 7423 12631
rect 10425 12597 10459 12631
rect 11069 12597 11103 12631
rect 11713 12597 11747 12631
rect 16037 12597 16071 12631
rect 2237 12393 2271 12427
rect 4261 12393 4295 12427
rect 6193 12393 6227 12427
rect 8585 12393 8619 12427
rect 9413 12393 9447 12427
rect 9597 12393 9631 12427
rect 11529 12393 11563 12427
rect 16497 12393 16531 12427
rect 17785 12393 17819 12427
rect 7021 12325 7055 12359
rect 9321 12257 9355 12291
rect 1777 12189 1811 12223
rect 2237 12189 2271 12223
rect 2421 12189 2455 12223
rect 2513 12189 2547 12223
rect 2973 12189 3007 12223
rect 4077 12189 4111 12223
rect 6377 12189 6411 12223
rect 6561 12189 6595 12223
rect 7297 12189 7331 12223
rect 7941 12189 7975 12223
rect 8309 12189 8343 12223
rect 8401 12189 8435 12223
rect 9229 12189 9263 12223
rect 10057 12189 10091 12223
rect 10701 12189 10735 12223
rect 11621 12189 11655 12223
rect 11897 12189 11931 12223
rect 12725 12189 12759 12223
rect 13001 12189 13035 12223
rect 14289 12189 14323 12223
rect 16681 12189 16715 12223
rect 17049 12189 17083 12223
rect 17509 12189 17543 12223
rect 7021 12121 7055 12155
rect 10793 12121 10827 12155
rect 14556 12121 14590 12155
rect 16773 12121 16807 12155
rect 16865 12121 16899 12155
rect 3157 12053 3191 12087
rect 7205 12053 7239 12087
rect 8033 12053 8067 12087
rect 8217 12053 8251 12087
rect 10241 12053 10275 12087
rect 10609 12053 10643 12087
rect 11345 12053 11379 12087
rect 12541 12053 12575 12087
rect 12909 12053 12943 12087
rect 15669 12053 15703 12087
rect 17969 12053 18003 12087
rect 6745 11849 6779 11883
rect 8401 11849 8435 11883
rect 8585 11849 8619 11883
rect 9413 11849 9447 11883
rect 10425 11849 10459 11883
rect 14565 11849 14599 11883
rect 15393 11849 15427 11883
rect 17509 11849 17543 11883
rect 6837 11781 6871 11815
rect 8309 11781 8343 11815
rect 11069 11781 11103 11815
rect 2789 11713 2823 11747
rect 3056 11713 3090 11747
rect 4896 11713 4930 11747
rect 6929 11713 6963 11747
rect 8217 11713 8251 11747
rect 9045 11713 9079 11747
rect 9229 11713 9263 11747
rect 10333 11713 10367 11747
rect 10517 11713 10551 11747
rect 10977 11713 11011 11747
rect 11161 11713 11195 11747
rect 11897 11713 11931 11747
rect 12541 11713 12575 11747
rect 12633 11713 12667 11747
rect 12817 11713 12851 11747
rect 13277 11713 13311 11747
rect 13461 11713 13495 11747
rect 14473 11713 14507 11747
rect 14657 11713 14691 11747
rect 15390 11713 15424 11747
rect 15761 11713 15795 11747
rect 16865 11713 16899 11747
rect 16957 11713 16991 11747
rect 17693 11713 17727 11747
rect 17877 11713 17911 11747
rect 4629 11645 4663 11679
rect 7113 11645 7147 11679
rect 8033 11645 8067 11679
rect 12081 11645 12115 11679
rect 15853 11645 15887 11679
rect 6009 11577 6043 11611
rect 12725 11577 12759 11611
rect 15209 11577 15243 11611
rect 4169 11509 4203 11543
rect 6561 11509 6595 11543
rect 9045 11509 9079 11543
rect 11713 11509 11747 11543
rect 13369 11509 13403 11543
rect 14013 11509 14047 11543
rect 17693 11509 17727 11543
rect 2881 11305 2915 11339
rect 3985 11305 4019 11339
rect 6101 11305 6135 11339
rect 7021 11305 7055 11339
rect 7665 11305 7699 11339
rect 10793 11305 10827 11339
rect 13277 11305 13311 11339
rect 17417 11305 17451 11339
rect 17693 11305 17727 11339
rect 6837 11237 6871 11271
rect 2513 11169 2547 11203
rect 4353 11169 4387 11203
rect 7941 11169 7975 11203
rect 8033 11169 8067 11203
rect 10425 11169 10459 11203
rect 13369 11169 13403 11203
rect 16037 11169 16071 11203
rect 17785 11169 17819 11203
rect 2697 11101 2731 11135
rect 4169 11101 4203 11135
rect 6101 11101 6135 11135
rect 6377 11101 6411 11135
rect 7849 11101 7883 11135
rect 8125 11101 8159 11135
rect 9321 11101 9355 11135
rect 9413 11101 9447 11135
rect 10609 11101 10643 11135
rect 12452 11079 12486 11113
rect 12541 11101 12575 11135
rect 12725 11101 12759 11135
rect 12817 11101 12851 11135
rect 13553 11101 13587 11135
rect 14565 11101 14599 11135
rect 14749 11101 14783 11135
rect 15393 11101 15427 11135
rect 15577 11101 15611 11135
rect 16221 11101 16255 11135
rect 16313 11101 16347 11135
rect 16405 11101 16439 11135
rect 16681 11101 16715 11135
rect 17601 11101 17635 11135
rect 6285 11033 6319 11067
rect 7005 11033 7039 11067
rect 7205 11033 7239 11067
rect 9137 11033 9171 11067
rect 12265 11033 12299 11067
rect 13277 11033 13311 11067
rect 16543 11033 16577 11067
rect 17877 11033 17911 11067
rect 5641 10965 5675 10999
rect 13737 10965 13771 10999
rect 14657 10965 14691 10999
rect 15577 10965 15611 10999
rect 3433 10761 3467 10795
rect 7941 10761 7975 10795
rect 9505 10761 9539 10795
rect 11805 10761 11839 10795
rect 12541 10761 12575 10795
rect 15393 10761 15427 10795
rect 17233 10761 17267 10795
rect 17417 10761 17451 10795
rect 9689 10693 9723 10727
rect 14280 10693 14314 10727
rect 18337 10693 18371 10727
rect 2605 10625 2639 10659
rect 3249 10625 3283 10659
rect 4169 10625 4203 10659
rect 4353 10625 4387 10659
rect 4997 10625 5031 10659
rect 5825 10625 5859 10659
rect 6009 10625 6043 10659
rect 6828 10625 6862 10659
rect 8401 10625 8435 10659
rect 8585 10625 8619 10659
rect 8677 10625 8711 10659
rect 9321 10625 9355 10659
rect 9413 10625 9447 10659
rect 10425 10625 10459 10659
rect 11713 10625 11747 10659
rect 11897 10625 11931 10659
rect 12817 10625 12851 10659
rect 13001 10625 13035 10659
rect 14013 10625 14047 10659
rect 15853 10625 15887 10659
rect 16037 10625 16071 10659
rect 17141 10625 17175 10659
rect 17969 10625 18003 10659
rect 3985 10557 4019 10591
rect 6561 10557 6595 10591
rect 10517 10557 10551 10591
rect 12725 10557 12759 10591
rect 12909 10557 12943 10591
rect 17049 10557 17083 10591
rect 17509 10557 17543 10591
rect 18153 10557 18187 10591
rect 10793 10489 10827 10523
rect 2789 10421 2823 10455
rect 4813 10421 4847 10455
rect 6009 10421 6043 10455
rect 8401 10421 8435 10455
rect 9137 10421 9171 10455
rect 16037 10421 16071 10455
rect 16865 10421 16899 10455
rect 18061 10421 18095 10455
rect 18337 10421 18371 10455
rect 3985 10217 4019 10251
rect 5733 10217 5767 10251
rect 7481 10217 7515 10251
rect 8585 10217 8619 10251
rect 10425 10217 10459 10251
rect 15117 10217 15151 10251
rect 15669 10217 15703 10251
rect 17049 10217 17083 10251
rect 17785 10217 17819 10251
rect 7849 10149 7883 10183
rect 13185 10149 13219 10183
rect 12909 10081 12943 10115
rect 17877 10081 17911 10115
rect 2329 10013 2363 10047
rect 2697 10013 2731 10047
rect 3157 10013 3191 10047
rect 7021 10013 7055 10047
rect 7665 10013 7699 10047
rect 7941 10013 7975 10047
rect 9137 10013 9171 10047
rect 11345 10013 11379 10047
rect 11621 10013 11655 10047
rect 12817 10013 12851 10047
rect 15298 10013 15332 10047
rect 15761 10013 15795 10047
rect 16681 10013 16715 10047
rect 16773 10013 16807 10047
rect 16865 10013 16899 10047
rect 17785 10013 17819 10047
rect 18061 10013 18095 10047
rect 2513 9945 2547 9979
rect 3341 9877 3375 9911
rect 11437 9877 11471 9911
rect 11805 9877 11839 9911
rect 13737 9877 13771 9911
rect 14381 9877 14415 9911
rect 15301 9877 15335 9911
rect 17601 9877 17635 9911
rect 8769 9673 8803 9707
rect 9781 9673 9815 9707
rect 3810 9605 3844 9639
rect 9413 9605 9447 9639
rect 9597 9605 9631 9639
rect 11989 9605 12023 9639
rect 13001 9605 13035 9639
rect 13705 9605 13739 9639
rect 13921 9605 13955 9639
rect 17785 9605 17819 9639
rect 4077 9537 4111 9571
rect 4537 9537 4571 9571
rect 4804 9537 4838 9571
rect 6745 9537 6779 9571
rect 7389 9537 7423 9571
rect 7645 9537 7679 9571
rect 10701 9537 10735 9571
rect 11713 9537 11747 9571
rect 11805 9537 11839 9571
rect 12817 9537 12851 9571
rect 13093 9537 13127 9571
rect 14657 9537 14691 9571
rect 14841 9537 14875 9571
rect 15761 9537 15795 9571
rect 15945 9537 15979 9571
rect 16865 9537 16899 9571
rect 17049 9537 17083 9571
rect 17509 9537 17543 9571
rect 10609 9469 10643 9503
rect 2697 9333 2731 9367
rect 5917 9333 5951 9367
rect 6837 9333 6871 9367
rect 10977 9333 11011 9367
rect 11713 9333 11747 9367
rect 12817 9333 12851 9367
rect 13553 9333 13587 9367
rect 13737 9333 13771 9367
rect 14657 9333 14691 9367
rect 15853 9333 15887 9367
rect 16957 9333 16991 9367
rect 4905 9129 4939 9163
rect 7757 9129 7791 9163
rect 9229 9129 9263 9163
rect 10701 9129 10735 9163
rect 14749 9129 14783 9163
rect 15301 9129 15335 9163
rect 16221 9129 16255 9163
rect 17233 9129 17267 9163
rect 5089 9061 5123 9095
rect 8309 9061 8343 9095
rect 10149 9061 10183 9095
rect 15853 9061 15887 9095
rect 16129 9061 16163 9095
rect 17325 9061 17359 9095
rect 10057 8993 10091 9027
rect 11345 8993 11379 9027
rect 15393 8993 15427 9027
rect 16313 8993 16347 9027
rect 5549 8925 5583 8959
rect 5733 8925 5767 8959
rect 7665 8925 7699 8959
rect 8493 8925 8527 8959
rect 9781 8925 9815 8959
rect 11897 8925 11931 8959
rect 12173 8925 12207 8959
rect 12357 8925 12391 8959
rect 12633 8925 12667 8959
rect 13185 8925 13219 8959
rect 13369 8925 13403 8959
rect 13461 8925 13495 8959
rect 13645 8925 13679 8959
rect 13737 8925 13771 8959
rect 14930 8925 14964 8959
rect 16589 8925 16623 8959
rect 17693 8925 17727 8959
rect 18153 8925 18187 8959
rect 4721 8857 4755 8891
rect 5641 8857 5675 8891
rect 6377 8857 6411 8891
rect 6561 8857 6595 8891
rect 4921 8789 4955 8823
rect 6193 8789 6227 8823
rect 11069 8789 11103 8823
rect 11161 8789 11195 8823
rect 12449 8789 12483 8823
rect 14933 8789 14967 8823
rect 16497 8789 16531 8823
rect 18245 8789 18279 8823
rect 4445 8585 4479 8619
rect 6561 8585 6595 8619
rect 6929 8585 6963 8619
rect 10977 8585 11011 8619
rect 12909 8585 12943 8619
rect 13185 8585 13219 8619
rect 8677 8517 8711 8551
rect 13068 8517 13102 8551
rect 14280 8517 14314 8551
rect 16957 8517 16991 8551
rect 2145 8449 2179 8483
rect 3065 8449 3099 8483
rect 3332 8449 3366 8483
rect 5089 8449 5123 8483
rect 8217 8449 8251 8483
rect 8309 8449 8343 8483
rect 9505 8449 9539 8483
rect 10609 8449 10643 8483
rect 11036 8449 11070 8483
rect 11713 8449 11747 8483
rect 12081 8449 12115 8483
rect 13553 8449 13587 8483
rect 16037 8449 16071 8483
rect 17601 8449 17635 8483
rect 17693 8449 17727 8483
rect 2053 8381 2087 8415
rect 4997 8381 5031 8415
rect 7021 8381 7055 8415
rect 7113 8381 7147 8415
rect 10517 8381 10551 8415
rect 12265 8381 12299 8415
rect 13277 8381 13311 8415
rect 14013 8381 14047 8415
rect 17785 8381 17819 8415
rect 2513 8313 2547 8347
rect 5457 8313 5491 8347
rect 8033 8313 8067 8347
rect 11805 8313 11839 8347
rect 15393 8313 15427 8347
rect 8493 8245 8527 8279
rect 9781 8245 9815 8279
rect 11161 8245 11195 8279
rect 16221 8245 16255 8279
rect 17417 8245 17451 8279
rect 2145 8041 2179 8075
rect 2605 8041 2639 8075
rect 6009 8041 6043 8075
rect 9597 8041 9631 8075
rect 12081 8041 12115 8075
rect 13553 8041 13587 8075
rect 17509 8041 17543 8075
rect 10333 7973 10367 8007
rect 1869 7905 1903 7939
rect 2789 7905 2823 7939
rect 2881 7905 2915 7939
rect 4261 7905 4295 7939
rect 4813 7905 4847 7939
rect 7941 7905 7975 7939
rect 9229 7905 9263 7939
rect 1777 7837 1811 7871
rect 2973 7837 3007 7871
rect 3065 7837 3099 7871
rect 4175 7837 4209 7871
rect 4353 7837 4387 7871
rect 4997 7837 5031 7871
rect 5181 7837 5215 7871
rect 5825 7837 5859 7871
rect 6561 7837 6595 7871
rect 6745 7837 6779 7871
rect 8309 7837 8343 7871
rect 8493 7837 8527 7871
rect 9413 7837 9447 7871
rect 10057 7837 10091 7871
rect 10149 7837 10183 7871
rect 11989 7837 12023 7871
rect 12173 7837 12207 7871
rect 13369 7837 13403 7871
rect 13553 7837 13587 7871
rect 16589 7837 16623 7871
rect 16773 7837 16807 7871
rect 17785 7837 17819 7871
rect 17877 7837 17911 7871
rect 17969 7837 18003 7871
rect 18153 7837 18187 7871
rect 8125 7769 8159 7803
rect 10333 7769 10367 7803
rect 10793 7769 10827 7803
rect 15853 7769 15887 7803
rect 6929 7701 6963 7735
rect 7481 7701 7515 7735
rect 8217 7701 8251 7735
rect 15761 7701 15795 7735
rect 16405 7701 16439 7735
rect 3433 7497 3467 7531
rect 4905 7497 4939 7531
rect 6009 7497 6043 7531
rect 7021 7497 7055 7531
rect 13093 7497 13127 7531
rect 16037 7497 16071 7531
rect 17233 7497 17267 7531
rect 4721 7429 4755 7463
rect 6745 7429 6779 7463
rect 11069 7429 11103 7463
rect 11958 7429 11992 7463
rect 14749 7429 14783 7463
rect 17693 7429 17727 7463
rect 2605 7361 2639 7395
rect 3617 7361 3651 7395
rect 3801 7361 3835 7395
rect 4537 7361 4571 7395
rect 5825 7361 5859 7395
rect 6009 7361 6043 7395
rect 7021 7361 7055 7395
rect 7849 7361 7883 7395
rect 8309 7361 8343 7395
rect 9413 7361 9447 7395
rect 9689 7361 9723 7395
rect 10977 7361 11011 7395
rect 11161 7361 11195 7395
rect 13553 7361 13587 7395
rect 14657 7361 14691 7395
rect 14933 7361 14967 7395
rect 15761 7361 15795 7395
rect 17601 7361 17635 7395
rect 2697 7293 2731 7327
rect 2973 7293 3007 7327
rect 8493 7293 8527 7327
rect 10517 7293 10551 7327
rect 11713 7293 11747 7327
rect 15393 7293 15427 7327
rect 15669 7293 15703 7327
rect 15878 7293 15912 7327
rect 17785 7293 17819 7327
rect 6929 7225 6963 7259
rect 7481 7225 7515 7259
rect 9505 7157 9539 7191
rect 9873 7157 9907 7191
rect 13737 7157 13771 7191
rect 14933 7157 14967 7191
rect 8401 6953 8435 6987
rect 16129 6953 16163 6987
rect 17233 6953 17267 6987
rect 17877 6953 17911 6987
rect 3985 6885 4019 6919
rect 2881 6817 2915 6851
rect 3157 6817 3191 6851
rect 3341 6817 3375 6851
rect 13645 6817 13679 6851
rect 14289 6817 14323 6851
rect 18153 6817 18187 6851
rect 2237 6749 2271 6783
rect 2421 6749 2455 6783
rect 3065 6749 3099 6783
rect 3249 6749 3283 6783
rect 5365 6749 5399 6783
rect 6285 6749 6319 6783
rect 6552 6749 6586 6783
rect 9137 6749 9171 6783
rect 9781 6749 9815 6783
rect 10037 6749 10071 6783
rect 11897 6749 11931 6783
rect 12449 6749 12483 6783
rect 12909 6749 12943 6783
rect 13737 6749 13771 6783
rect 16313 6749 16347 6783
rect 16405 6749 16439 6783
rect 17233 6749 17267 6783
rect 17417 6749 17451 6783
rect 17877 6749 17911 6783
rect 17969 6749 18003 6783
rect 2329 6681 2363 6715
rect 5098 6681 5132 6715
rect 8217 6681 8251 6715
rect 8433 6681 8467 6715
rect 13461 6681 13495 6715
rect 14534 6681 14568 6715
rect 16129 6681 16163 6715
rect 1777 6613 1811 6647
rect 7665 6613 7699 6647
rect 8585 6613 8619 6647
rect 9229 6613 9263 6647
rect 11161 6613 11195 6647
rect 12909 6613 12943 6647
rect 13737 6613 13771 6647
rect 15669 6613 15703 6647
rect 16589 6613 16623 6647
rect 17049 6613 17083 6647
rect 10977 6409 11011 6443
rect 11805 6409 11839 6443
rect 12725 6409 12759 6443
rect 15485 6409 15519 6443
rect 17049 6409 17083 6443
rect 18061 6409 18095 6443
rect 2789 6341 2823 6375
rect 7849 6341 7883 6375
rect 10057 6341 10091 6375
rect 10425 6341 10459 6375
rect 17693 6341 17727 6375
rect 2973 6273 3007 6307
rect 3065 6273 3099 6307
rect 3985 6273 4019 6307
rect 4169 6273 4203 6307
rect 4629 6273 4663 6307
rect 4896 6273 4930 6307
rect 6745 6273 6779 6307
rect 7665 6273 7699 6307
rect 8125 6273 8159 6307
rect 8309 6273 8343 6307
rect 9229 6273 9263 6307
rect 9413 6273 9447 6307
rect 10885 6273 10919 6307
rect 11713 6273 11747 6307
rect 11989 6273 12023 6307
rect 12725 6273 12759 6307
rect 12909 6273 12943 6307
rect 16865 6273 16899 6307
rect 17049 6273 17083 6307
rect 17509 6273 17543 6307
rect 17785 6273 17819 6307
rect 17877 6273 17911 6307
rect 8493 6205 8527 6239
rect 9137 6205 9171 6239
rect 9321 6205 9355 6239
rect 15025 6205 15059 6239
rect 2789 6137 2823 6171
rect 6009 6137 6043 6171
rect 15393 6137 15427 6171
rect 4169 6069 4203 6103
rect 6561 6069 6595 6103
rect 8953 6069 8987 6103
rect 11989 6069 12023 6103
rect 13461 6069 13495 6103
rect 16221 6069 16255 6103
rect 3985 5865 4019 5899
rect 7665 5865 7699 5899
rect 11437 5865 11471 5899
rect 12081 5865 12115 5899
rect 13737 5865 13771 5899
rect 15945 5865 15979 5899
rect 17601 5865 17635 5899
rect 17785 5865 17819 5899
rect 18245 5865 18279 5899
rect 3065 5797 3099 5831
rect 8309 5797 8343 5831
rect 16681 5797 16715 5831
rect 2329 5729 2363 5763
rect 4537 5729 4571 5763
rect 5273 5729 5307 5763
rect 7757 5729 7791 5763
rect 2789 5661 2823 5695
rect 3065 5661 3099 5695
rect 4721 5661 4755 5695
rect 4813 5661 4847 5695
rect 7021 5661 7055 5695
rect 7849 5661 7883 5695
rect 8309 5661 8343 5695
rect 8493 5661 8527 5695
rect 8585 5661 8619 5695
rect 9505 5661 9539 5695
rect 9781 5661 9815 5695
rect 10425 5661 10459 5695
rect 10609 5661 10643 5695
rect 10793 5661 10827 5695
rect 12265 5661 12299 5695
rect 12541 5661 12575 5695
rect 13093 5661 13127 5695
rect 13277 5661 13311 5695
rect 13553 5661 13587 5695
rect 15301 5661 15335 5695
rect 15485 5661 15519 5695
rect 15761 5661 15795 5695
rect 16957 5661 16991 5695
rect 2881 5593 2915 5627
rect 9597 5593 9631 5627
rect 10701 5593 10735 5627
rect 17417 5593 17451 5627
rect 4813 5525 4847 5559
rect 7481 5525 7515 5559
rect 9965 5525 9999 5559
rect 10977 5525 11011 5559
rect 12449 5525 12483 5559
rect 14841 5525 14875 5559
rect 16497 5525 16531 5559
rect 17617 5525 17651 5559
rect 2237 5321 2271 5355
rect 5457 5321 5491 5355
rect 5917 5321 5951 5355
rect 6929 5321 6963 5355
rect 10609 5321 10643 5355
rect 15301 5321 15335 5355
rect 18245 5321 18279 5355
rect 7849 5253 7883 5287
rect 9597 5253 9631 5287
rect 16129 5253 16163 5287
rect 16313 5253 16347 5287
rect 17601 5253 17635 5287
rect 3361 5185 3395 5219
rect 3617 5185 3651 5219
rect 4077 5185 4111 5219
rect 4333 5185 4367 5219
rect 6837 5185 6871 5219
rect 11161 5185 11195 5219
rect 11897 5185 11931 5219
rect 12153 5185 12187 5219
rect 13921 5185 13955 5219
rect 14188 5185 14222 5219
rect 16037 5185 16071 5219
rect 17233 5185 17267 5219
rect 6745 5117 6779 5151
rect 10885 5117 10919 5151
rect 7297 4981 7331 5015
rect 10977 4981 11011 5015
rect 13277 4981 13311 5015
rect 16313 4981 16347 5015
rect 17601 4981 17635 5015
rect 17785 4981 17819 5015
rect 2973 4777 3007 4811
rect 3341 4777 3375 4811
rect 4353 4777 4387 4811
rect 5273 4777 5307 4811
rect 6745 4777 6779 4811
rect 8585 4777 8619 4811
rect 9965 4777 9999 4811
rect 10793 4777 10827 4811
rect 14289 4777 14323 4811
rect 15853 4777 15887 4811
rect 16681 4777 16715 4811
rect 18153 4777 18187 4811
rect 10977 4709 11011 4743
rect 13737 4709 13771 4743
rect 15945 4709 15979 4743
rect 2881 4641 2915 4675
rect 7205 4641 7239 4675
rect 14448 4641 14482 4675
rect 14565 4641 14599 4675
rect 14933 4641 14967 4675
rect 3157 4573 3191 4607
rect 5549 4573 5583 4607
rect 6377 4573 6411 4607
rect 6561 4573 6595 4607
rect 7472 4573 7506 4607
rect 9137 4573 9171 4607
rect 9321 4573 9355 4607
rect 11437 4573 11471 4607
rect 16037 4573 16071 4607
rect 17749 4573 17783 4607
rect 17857 4573 17891 4607
rect 17969 4573 18003 4607
rect 9229 4505 9263 4539
rect 9949 4505 9983 4539
rect 10149 4505 10183 4539
rect 10609 4505 10643 4539
rect 10825 4505 10859 4539
rect 14657 4505 14691 4539
rect 15761 4505 15795 4539
rect 16665 4505 16699 4539
rect 16865 4505 16899 4539
rect 9781 4437 9815 4471
rect 11621 4437 11655 4471
rect 16497 4437 16531 4471
rect 8677 4233 8711 4267
rect 10701 4233 10735 4267
rect 13093 4233 13127 4267
rect 17233 4233 17267 4267
rect 5365 4165 5399 4199
rect 5549 4165 5583 4199
rect 11958 4165 11992 4199
rect 16865 4165 16899 4199
rect 17325 4165 17359 4199
rect 4537 4097 4571 4131
rect 5181 4097 5215 4131
rect 7481 4097 7515 4131
rect 8401 4097 8435 4131
rect 8769 4097 8803 4131
rect 9588 4097 9622 4131
rect 13921 4097 13955 4131
rect 14188 4097 14222 4131
rect 16129 4097 16163 4131
rect 16313 4097 16347 4131
rect 6561 4029 6595 4063
rect 7941 4029 7975 4063
rect 8585 4029 8619 4063
rect 9321 4029 9355 4063
rect 11713 4029 11747 4063
rect 16957 4029 16991 4063
rect 6929 3961 6963 3995
rect 16129 3961 16163 3995
rect 17049 3961 17083 3995
rect 4721 3893 4755 3927
rect 7021 3893 7055 3927
rect 7573 3893 7607 3927
rect 8401 3893 8435 3927
rect 15301 3893 15335 3927
rect 17877 3893 17911 3927
rect 8493 3689 8527 3723
rect 9505 3689 9539 3723
rect 17141 3689 17175 3723
rect 16497 3621 16531 3655
rect 7205 3553 7239 3587
rect 7665 3553 7699 3587
rect 5365 3485 5399 3519
rect 6193 3485 6227 3519
rect 6285 3485 6319 3519
rect 6469 3485 6503 3519
rect 6561 3485 6595 3519
rect 7573 3485 7607 3519
rect 8401 3485 8435 3519
rect 8585 3485 8619 3519
rect 9321 3485 9355 3519
rect 9965 3485 9999 3519
rect 10149 3485 10183 3519
rect 11253 3485 11287 3519
rect 12909 3485 12943 3519
rect 13001 3485 13035 3519
rect 13185 3485 13219 3519
rect 13277 3485 13311 3519
rect 14289 3485 14323 3519
rect 15485 3485 15519 3519
rect 16221 3485 16255 3519
rect 18061 3485 18095 3519
rect 5120 3417 5154 3451
rect 7849 3417 7883 3451
rect 16497 3417 16531 3451
rect 16957 3417 16991 3451
rect 17157 3417 17191 3451
rect 3985 3349 4019 3383
rect 6745 3349 6779 3383
rect 10057 3349 10091 3383
rect 11437 3349 11471 3383
rect 12173 3349 12207 3383
rect 12725 3349 12759 3383
rect 14473 3349 14507 3383
rect 15669 3349 15703 3383
rect 16313 3349 16347 3383
rect 17325 3349 17359 3383
rect 18245 3349 18279 3383
rect 6561 3145 6595 3179
rect 11161 3145 11195 3179
rect 13093 3145 13127 3179
rect 15393 3145 15427 3179
rect 17233 3145 17267 3179
rect 8002 3077 8036 3111
rect 16313 3077 16347 3111
rect 17325 3077 17359 3111
rect 18337 3077 18371 3111
rect 2789 3009 2823 3043
rect 3056 3009 3090 3043
rect 4629 3009 4663 3043
rect 4885 3009 4919 3043
rect 6745 3009 6779 3043
rect 6837 3009 6871 3043
rect 7021 3009 7055 3043
rect 7113 3009 7147 3043
rect 7757 3009 7791 3043
rect 9781 3009 9815 3043
rect 10048 3009 10082 3043
rect 11713 3009 11747 3043
rect 11969 3009 12003 3043
rect 14013 3009 14047 3043
rect 14280 3009 14314 3043
rect 15945 3009 15979 3043
rect 16129 3009 16163 3043
rect 18061 3009 18095 3043
rect 18153 3009 18187 3043
rect 17417 2941 17451 2975
rect 4169 2805 4203 2839
rect 6009 2805 6043 2839
rect 9137 2805 9171 2839
rect 16865 2805 16899 2839
rect 18061 2805 18095 2839
rect 5181 2601 5215 2635
rect 7573 2601 7607 2635
rect 10517 2601 10551 2635
rect 11805 2601 11839 2635
rect 13645 2601 13679 2635
rect 15669 2601 15703 2635
rect 17325 2601 17359 2635
rect 18153 2601 18187 2635
rect 6745 2533 6779 2567
rect 17693 2533 17727 2567
rect 14289 2465 14323 2499
rect 16221 2465 16255 2499
rect 1869 2397 1903 2431
rect 4261 2397 4295 2431
rect 5089 2397 5123 2431
rect 5273 2397 5307 2431
rect 6009 2397 6043 2431
rect 6561 2397 6595 2431
rect 7021 2397 7055 2431
rect 7481 2397 7515 2431
rect 7665 2397 7699 2431
rect 8585 2397 8619 2431
rect 9137 2397 9171 2431
rect 12265 2397 12299 2431
rect 16129 2397 16163 2431
rect 16313 2397 16347 2431
rect 17233 2397 17267 2431
rect 6929 2329 6963 2363
rect 9382 2329 9416 2363
rect 12532 2329 12566 2363
rect 14556 2329 14590 2363
rect 1685 2261 1719 2295
rect 4077 2261 4111 2295
rect 5825 2261 5859 2295
rect 8401 2261 8435 2295
<< metal1 >>
rect 1104 17434 19019 17456
rect 1104 17382 5388 17434
rect 5440 17382 5452 17434
rect 5504 17382 5516 17434
rect 5568 17382 5580 17434
rect 5632 17382 5644 17434
rect 5696 17382 9827 17434
rect 9879 17382 9891 17434
rect 9943 17382 9955 17434
rect 10007 17382 10019 17434
rect 10071 17382 10083 17434
rect 10135 17382 14266 17434
rect 14318 17382 14330 17434
rect 14382 17382 14394 17434
rect 14446 17382 14458 17434
rect 14510 17382 14522 17434
rect 14574 17382 18705 17434
rect 18757 17382 18769 17434
rect 18821 17382 18833 17434
rect 18885 17382 18897 17434
rect 18949 17382 18961 17434
rect 19013 17382 19019 17434
rect 1104 17360 19019 17382
rect 5813 17323 5871 17329
rect 5813 17289 5825 17323
rect 5859 17289 5871 17323
rect 5813 17283 5871 17289
rect 16301 17323 16359 17329
rect 16301 17289 16313 17323
rect 16347 17320 16359 17323
rect 16574 17320 16580 17332
rect 16347 17292 16580 17320
rect 16347 17289 16359 17292
rect 16301 17283 16359 17289
rect 5108 17255 5166 17261
rect 5108 17221 5120 17255
rect 5154 17252 5166 17255
rect 5828 17252 5856 17283
rect 16574 17280 16580 17292
rect 16632 17280 16638 17332
rect 12345 17255 12403 17261
rect 12345 17252 12357 17255
rect 5154 17224 5856 17252
rect 11072 17224 12357 17252
rect 5154 17221 5166 17224
rect 5108 17215 5166 17221
rect 2774 17144 2780 17196
rect 2832 17184 2838 17196
rect 3053 17187 3111 17193
rect 3053 17184 3065 17187
rect 2832 17156 3065 17184
rect 2832 17144 2838 17156
rect 3053 17153 3065 17156
rect 3099 17153 3111 17187
rect 3053 17147 3111 17153
rect 5997 17187 6055 17193
rect 5997 17153 6009 17187
rect 6043 17184 6055 17187
rect 6546 17184 6552 17196
rect 6043 17156 6552 17184
rect 6043 17153 6055 17156
rect 5997 17147 6055 17153
rect 6546 17144 6552 17156
rect 6604 17144 6610 17196
rect 6733 17187 6791 17193
rect 6733 17153 6745 17187
rect 6779 17184 6791 17187
rect 7190 17184 7196 17196
rect 6779 17156 7196 17184
rect 6779 17153 6791 17156
rect 6733 17147 6791 17153
rect 7190 17144 7196 17156
rect 7248 17144 7254 17196
rect 9306 17184 9312 17196
rect 9267 17156 9312 17184
rect 9306 17144 9312 17156
rect 9364 17144 9370 17196
rect 10045 17187 10103 17193
rect 10045 17153 10057 17187
rect 10091 17184 10103 17187
rect 10134 17184 10140 17196
rect 10091 17156 10140 17184
rect 10091 17153 10103 17156
rect 10045 17147 10103 17153
rect 10134 17144 10140 17156
rect 10192 17144 10198 17196
rect 10229 17187 10287 17193
rect 10229 17153 10241 17187
rect 10275 17153 10287 17187
rect 10229 17147 10287 17153
rect 5350 17116 5356 17128
rect 5311 17088 5356 17116
rect 5350 17076 5356 17088
rect 5408 17076 5414 17128
rect 6917 17119 6975 17125
rect 6917 17085 6929 17119
rect 6963 17116 6975 17119
rect 7098 17116 7104 17128
rect 6963 17088 7104 17116
rect 6963 17085 6975 17088
rect 6917 17079 6975 17085
rect 7098 17076 7104 17088
rect 7156 17076 7162 17128
rect 10244 17116 10272 17147
rect 10318 17144 10324 17196
rect 10376 17184 10382 17196
rect 11072 17193 11100 17224
rect 12345 17221 12357 17224
rect 12391 17221 12403 17255
rect 12345 17215 12403 17221
rect 11057 17187 11115 17193
rect 11057 17184 11069 17187
rect 10376 17156 11069 17184
rect 10376 17144 10382 17156
rect 11057 17153 11069 17156
rect 11103 17153 11115 17187
rect 11057 17147 11115 17153
rect 11885 17187 11943 17193
rect 11885 17153 11897 17187
rect 11931 17184 11943 17187
rect 12618 17184 12624 17196
rect 11931 17156 12624 17184
rect 11931 17153 11943 17156
rect 11885 17147 11943 17153
rect 12618 17144 12624 17156
rect 12676 17144 12682 17196
rect 16592 17184 16620 17280
rect 16853 17187 16911 17193
rect 16853 17184 16865 17187
rect 16592 17156 16865 17184
rect 16853 17153 16865 17156
rect 16899 17153 16911 17187
rect 16853 17147 16911 17153
rect 7392 17088 12434 17116
rect 3237 17051 3295 17057
rect 3237 17017 3249 17051
rect 3283 17048 3295 17051
rect 4246 17048 4252 17060
rect 3283 17020 4252 17048
rect 3283 17017 3295 17020
rect 3237 17011 3295 17017
rect 4246 17008 4252 17020
rect 4304 17008 4310 17060
rect 7392 16992 7420 17088
rect 9858 17008 9864 17060
rect 9916 17048 9922 17060
rect 10873 17051 10931 17057
rect 10873 17048 10885 17051
rect 9916 17020 10885 17048
rect 9916 17008 9922 17020
rect 10873 17017 10885 17020
rect 10919 17017 10931 17051
rect 10873 17011 10931 17017
rect 3970 16980 3976 16992
rect 3931 16952 3976 16980
rect 3970 16940 3976 16952
rect 4028 16940 4034 16992
rect 5994 16940 6000 16992
rect 6052 16980 6058 16992
rect 6549 16983 6607 16989
rect 6549 16980 6561 16983
rect 6052 16952 6561 16980
rect 6052 16940 6058 16952
rect 6549 16949 6561 16952
rect 6595 16949 6607 16983
rect 7374 16980 7380 16992
rect 7335 16952 7380 16980
rect 6549 16943 6607 16949
rect 7374 16940 7380 16952
rect 7432 16940 7438 16992
rect 8938 16940 8944 16992
rect 8996 16980 9002 16992
rect 9125 16983 9183 16989
rect 9125 16980 9137 16983
rect 8996 16952 9137 16980
rect 8996 16940 9002 16952
rect 9125 16949 9137 16952
rect 9171 16949 9183 16983
rect 9125 16943 9183 16949
rect 10413 16983 10471 16989
rect 10413 16949 10425 16983
rect 10459 16980 10471 16983
rect 10502 16980 10508 16992
rect 10459 16952 10508 16980
rect 10459 16949 10471 16952
rect 10413 16943 10471 16949
rect 10502 16940 10508 16952
rect 10560 16940 10566 16992
rect 10594 16940 10600 16992
rect 10652 16980 10658 16992
rect 11701 16983 11759 16989
rect 11701 16980 11713 16983
rect 10652 16952 11713 16980
rect 10652 16940 10658 16952
rect 11701 16949 11713 16952
rect 11747 16949 11759 16983
rect 12406 16980 12434 17088
rect 16942 17076 16948 17128
rect 17000 17116 17006 17128
rect 17129 17119 17187 17125
rect 17129 17116 17141 17119
rect 17000 17088 17141 17116
rect 17000 17076 17006 17088
rect 17129 17085 17141 17088
rect 17175 17085 17187 17119
rect 17129 17079 17187 17085
rect 12802 16980 12808 16992
rect 12406 16952 12808 16980
rect 11701 16943 11759 16949
rect 12802 16940 12808 16952
rect 12860 16980 12866 16992
rect 12897 16983 12955 16989
rect 12897 16980 12909 16983
rect 12860 16952 12909 16980
rect 12860 16940 12866 16952
rect 12897 16949 12909 16952
rect 12943 16949 12955 16983
rect 12897 16943 12955 16949
rect 1104 16890 18860 16912
rect 1104 16838 3169 16890
rect 3221 16838 3233 16890
rect 3285 16838 3297 16890
rect 3349 16838 3361 16890
rect 3413 16838 3425 16890
rect 3477 16838 7608 16890
rect 7660 16838 7672 16890
rect 7724 16838 7736 16890
rect 7788 16838 7800 16890
rect 7852 16838 7864 16890
rect 7916 16838 12047 16890
rect 12099 16838 12111 16890
rect 12163 16838 12175 16890
rect 12227 16838 12239 16890
rect 12291 16838 12303 16890
rect 12355 16838 16486 16890
rect 16538 16838 16550 16890
rect 16602 16838 16614 16890
rect 16666 16838 16678 16890
rect 16730 16838 16742 16890
rect 16794 16838 18860 16890
rect 1104 16816 18860 16838
rect 2774 16736 2780 16788
rect 2832 16776 2838 16788
rect 7190 16776 7196 16788
rect 2832 16748 2877 16776
rect 7151 16748 7196 16776
rect 2832 16736 2838 16748
rect 7190 16736 7196 16748
rect 7248 16736 7254 16788
rect 9769 16779 9827 16785
rect 9769 16745 9781 16779
rect 9815 16776 9827 16779
rect 10318 16776 10324 16788
rect 9815 16748 10324 16776
rect 9815 16745 9827 16748
rect 9769 16739 9827 16745
rect 10318 16736 10324 16748
rect 10376 16736 10382 16788
rect 12618 16776 12624 16788
rect 12579 16748 12624 16776
rect 12618 16736 12624 16748
rect 12676 16736 12682 16788
rect 10413 16643 10471 16649
rect 10413 16609 10425 16643
rect 10459 16609 10471 16643
rect 10413 16603 10471 16609
rect 3145 16575 3203 16581
rect 3145 16541 3157 16575
rect 3191 16572 3203 16575
rect 3970 16572 3976 16584
rect 3191 16544 3976 16572
rect 3191 16541 3203 16544
rect 3145 16535 3203 16541
rect 3970 16532 3976 16544
rect 4028 16532 4034 16584
rect 4982 16532 4988 16584
rect 5040 16572 5046 16584
rect 5350 16572 5356 16584
rect 5040 16544 5356 16572
rect 5040 16532 5046 16544
rect 5350 16532 5356 16544
rect 5408 16532 5414 16584
rect 8570 16572 8576 16584
rect 8531 16544 8576 16572
rect 8570 16532 8576 16544
rect 8628 16572 8634 16584
rect 10428 16572 10456 16603
rect 8628 16544 10456 16572
rect 8628 16532 8634 16544
rect 2961 16507 3019 16513
rect 2961 16473 2973 16507
rect 3007 16473 3019 16507
rect 2961 16467 3019 16473
rect 5620 16507 5678 16513
rect 5620 16473 5632 16507
rect 5666 16504 5678 16507
rect 5810 16504 5816 16516
rect 5666 16476 5816 16504
rect 5666 16473 5678 16476
rect 5620 16467 5678 16473
rect 2976 16436 3004 16467
rect 5810 16464 5816 16476
rect 5868 16464 5874 16516
rect 8328 16507 8386 16513
rect 8328 16473 8340 16507
rect 8374 16504 8386 16507
rect 9858 16504 9864 16516
rect 8374 16476 9720 16504
rect 9819 16476 9864 16504
rect 8374 16473 8386 16476
rect 8328 16467 8386 16473
rect 3694 16436 3700 16448
rect 2976 16408 3700 16436
rect 3694 16396 3700 16408
rect 3752 16436 3758 16448
rect 3973 16439 4031 16445
rect 3973 16436 3985 16439
rect 3752 16408 3985 16436
rect 3752 16396 3758 16408
rect 3973 16405 3985 16408
rect 4019 16405 4031 16439
rect 3973 16399 4031 16405
rect 6733 16439 6791 16445
rect 6733 16405 6745 16439
rect 6779 16436 6791 16439
rect 6914 16436 6920 16448
rect 6779 16408 6920 16436
rect 6779 16405 6791 16408
rect 6733 16399 6791 16405
rect 6914 16396 6920 16408
rect 6972 16396 6978 16448
rect 9692 16436 9720 16476
rect 9858 16464 9864 16476
rect 9916 16464 9922 16516
rect 10686 16513 10692 16516
rect 10680 16467 10692 16513
rect 10744 16504 10750 16516
rect 12253 16507 12311 16513
rect 10744 16476 10780 16504
rect 10686 16464 10692 16467
rect 10744 16464 10750 16476
rect 12253 16473 12265 16507
rect 12299 16473 12311 16507
rect 12253 16467 12311 16473
rect 12437 16507 12495 16513
rect 12437 16473 12449 16507
rect 12483 16504 12495 16507
rect 12802 16504 12808 16516
rect 12483 16476 12808 16504
rect 12483 16473 12495 16476
rect 12437 16467 12495 16473
rect 10594 16436 10600 16448
rect 9692 16408 10600 16436
rect 10594 16396 10600 16408
rect 10652 16396 10658 16448
rect 11793 16439 11851 16445
rect 11793 16405 11805 16439
rect 11839 16436 11851 16439
rect 12268 16436 12296 16467
rect 12802 16464 12808 16476
rect 12860 16504 12866 16516
rect 13081 16507 13139 16513
rect 13081 16504 13093 16507
rect 12860 16476 13093 16504
rect 12860 16464 12866 16476
rect 13081 16473 13093 16476
rect 13127 16473 13139 16507
rect 13081 16467 13139 16473
rect 11839 16408 12296 16436
rect 11839 16405 11851 16408
rect 11793 16399 11851 16405
rect 1104 16346 19019 16368
rect 1104 16294 5388 16346
rect 5440 16294 5452 16346
rect 5504 16294 5516 16346
rect 5568 16294 5580 16346
rect 5632 16294 5644 16346
rect 5696 16294 9827 16346
rect 9879 16294 9891 16346
rect 9943 16294 9955 16346
rect 10007 16294 10019 16346
rect 10071 16294 10083 16346
rect 10135 16294 14266 16346
rect 14318 16294 14330 16346
rect 14382 16294 14394 16346
rect 14446 16294 14458 16346
rect 14510 16294 14522 16346
rect 14574 16294 18705 16346
rect 18757 16294 18769 16346
rect 18821 16294 18833 16346
rect 18885 16294 18897 16346
rect 18949 16294 18961 16346
rect 19013 16294 19019 16346
rect 1104 16272 19019 16294
rect 5810 16232 5816 16244
rect 5771 16204 5816 16232
rect 5810 16192 5816 16204
rect 5868 16192 5874 16244
rect 6546 16232 6552 16244
rect 6507 16204 6552 16232
rect 6546 16192 6552 16204
rect 6604 16192 6610 16244
rect 7374 16232 7380 16244
rect 6748 16204 7380 16232
rect 4246 16124 4252 16176
rect 4304 16173 4310 16176
rect 6748 16173 6776 16204
rect 7374 16192 7380 16204
rect 7432 16192 7438 16244
rect 8205 16235 8263 16241
rect 8205 16201 8217 16235
rect 8251 16232 8263 16235
rect 9306 16232 9312 16244
rect 8251 16204 9312 16232
rect 8251 16201 8263 16204
rect 8205 16195 8263 16201
rect 9306 16192 9312 16204
rect 9364 16192 9370 16244
rect 10045 16235 10103 16241
rect 10045 16201 10057 16235
rect 10091 16232 10103 16235
rect 10226 16232 10232 16244
rect 10091 16204 10232 16232
rect 10091 16201 10103 16204
rect 10045 16195 10103 16201
rect 10226 16192 10232 16204
rect 10284 16192 10290 16244
rect 10686 16232 10692 16244
rect 10647 16204 10692 16232
rect 10686 16192 10692 16204
rect 10744 16192 10750 16244
rect 12434 16232 12440 16244
rect 12176 16204 12440 16232
rect 4304 16164 4316 16173
rect 6733 16167 6791 16173
rect 6733 16164 6745 16167
rect 4304 16136 4349 16164
rect 5828 16136 6745 16164
rect 4304 16127 4316 16136
rect 4304 16124 4310 16127
rect 3694 16056 3700 16108
rect 3752 16096 3758 16108
rect 5828 16096 5856 16136
rect 6733 16133 6745 16136
rect 6779 16133 6791 16167
rect 6914 16164 6920 16176
rect 6875 16136 6920 16164
rect 6733 16127 6791 16133
rect 6914 16124 6920 16136
rect 6972 16124 6978 16176
rect 8570 16124 8576 16176
rect 8628 16164 8634 16176
rect 9122 16164 9128 16176
rect 8628 16136 9128 16164
rect 8628 16124 8634 16136
rect 5994 16096 6000 16108
rect 3752 16068 5856 16096
rect 5955 16068 6000 16096
rect 3752 16056 3758 16068
rect 5994 16056 6000 16068
rect 6052 16056 6058 16108
rect 8018 16096 8024 16108
rect 7979 16068 8024 16096
rect 8018 16056 8024 16068
rect 8076 16056 8082 16108
rect 8680 16105 8708 16136
rect 9122 16124 9128 16136
rect 9180 16124 9186 16176
rect 8938 16105 8944 16108
rect 8665 16099 8723 16105
rect 8665 16065 8677 16099
rect 8711 16065 8723 16099
rect 8932 16096 8944 16105
rect 8899 16068 8944 16096
rect 8665 16059 8723 16065
rect 8932 16059 8944 16068
rect 8938 16056 8944 16059
rect 8996 16056 9002 16108
rect 10502 16096 10508 16108
rect 10463 16068 10508 16096
rect 10502 16056 10508 16068
rect 10560 16056 10566 16108
rect 11698 16056 11704 16108
rect 11756 16096 11762 16108
rect 12176 16105 12204 16204
rect 12434 16192 12440 16204
rect 12492 16232 12498 16244
rect 12492 16204 13216 16232
rect 12492 16192 12498 16204
rect 11885 16099 11943 16105
rect 11885 16096 11897 16099
rect 11756 16068 11897 16096
rect 11756 16056 11762 16068
rect 11885 16065 11897 16068
rect 11931 16065 11943 16099
rect 11885 16059 11943 16065
rect 12069 16099 12127 16105
rect 12069 16065 12081 16099
rect 12115 16065 12127 16099
rect 12069 16059 12127 16065
rect 12161 16099 12219 16105
rect 12161 16065 12173 16099
rect 12207 16065 12219 16099
rect 12161 16059 12219 16065
rect 4525 16031 4583 16037
rect 4525 15997 4537 16031
rect 4571 16028 4583 16031
rect 4982 16028 4988 16040
rect 4571 16000 4988 16028
rect 4571 15997 4583 16000
rect 4525 15991 4583 15997
rect 4982 15988 4988 16000
rect 5040 15988 5046 16040
rect 7098 15988 7104 16040
rect 7156 16028 7162 16040
rect 7837 16031 7895 16037
rect 7837 16028 7849 16031
rect 7156 16000 7849 16028
rect 7156 15988 7162 16000
rect 7837 15997 7849 16000
rect 7883 15997 7895 16031
rect 12084 16028 12112 16059
rect 12250 16056 12256 16108
rect 12308 16096 12314 16108
rect 13188 16105 13216 16204
rect 13970 16167 14028 16173
rect 13970 16164 13982 16167
rect 13280 16136 13982 16164
rect 12989 16099 13047 16105
rect 12989 16096 13001 16099
rect 12308 16068 13001 16096
rect 12308 16056 12314 16068
rect 12989 16065 13001 16068
rect 13035 16065 13047 16099
rect 12989 16059 13047 16065
rect 13173 16099 13231 16105
rect 13173 16065 13185 16099
rect 13219 16065 13231 16099
rect 13173 16059 13231 16065
rect 13081 16031 13139 16037
rect 13081 16028 13093 16031
rect 12084 16000 13093 16028
rect 7837 15991 7895 15997
rect 13081 15997 13093 16000
rect 13127 15997 13139 16031
rect 13081 15991 13139 15997
rect 11790 15920 11796 15972
rect 11848 15960 11854 15972
rect 12250 15960 12256 15972
rect 11848 15932 12256 15960
rect 11848 15920 11854 15932
rect 12250 15920 12256 15932
rect 12308 15920 12314 15972
rect 12529 15963 12587 15969
rect 12529 15929 12541 15963
rect 12575 15960 12587 15963
rect 13280 15960 13308 16136
rect 13970 16133 13982 16136
rect 14016 16133 14028 16167
rect 13970 16127 14028 16133
rect 13722 16028 13728 16040
rect 13683 16000 13728 16028
rect 13722 15988 13728 16000
rect 13780 15988 13786 16040
rect 12575 15932 13308 15960
rect 12575 15929 12587 15932
rect 12529 15923 12587 15929
rect 3050 15852 3056 15904
rect 3108 15892 3114 15904
rect 3145 15895 3203 15901
rect 3145 15892 3157 15895
rect 3108 15864 3157 15892
rect 3108 15852 3114 15864
rect 3145 15861 3157 15864
rect 3191 15861 3203 15895
rect 3145 15855 3203 15861
rect 3510 15852 3516 15904
rect 3568 15892 3574 15904
rect 8662 15892 8668 15904
rect 3568 15864 8668 15892
rect 3568 15852 3574 15864
rect 8662 15852 8668 15864
rect 8720 15852 8726 15904
rect 15105 15895 15163 15901
rect 15105 15861 15117 15895
rect 15151 15892 15163 15895
rect 17126 15892 17132 15904
rect 15151 15864 17132 15892
rect 15151 15861 15163 15864
rect 15105 15855 15163 15861
rect 17126 15852 17132 15864
rect 17184 15852 17190 15904
rect 1104 15802 18860 15824
rect 1104 15750 3169 15802
rect 3221 15750 3233 15802
rect 3285 15750 3297 15802
rect 3349 15750 3361 15802
rect 3413 15750 3425 15802
rect 3477 15750 7608 15802
rect 7660 15750 7672 15802
rect 7724 15750 7736 15802
rect 7788 15750 7800 15802
rect 7852 15750 7864 15802
rect 7916 15750 12047 15802
rect 12099 15750 12111 15802
rect 12163 15750 12175 15802
rect 12227 15750 12239 15802
rect 12291 15750 12303 15802
rect 12355 15750 16486 15802
rect 16538 15750 16550 15802
rect 16602 15750 16614 15802
rect 16666 15750 16678 15802
rect 16730 15750 16742 15802
rect 16794 15750 18860 15802
rect 1104 15728 18860 15750
rect 12069 15691 12127 15697
rect 12069 15657 12081 15691
rect 12115 15688 12127 15691
rect 12434 15688 12440 15700
rect 12115 15660 12440 15688
rect 12115 15657 12127 15660
rect 12069 15651 12127 15657
rect 12434 15648 12440 15660
rect 12492 15648 12498 15700
rect 3421 15555 3479 15561
rect 3421 15521 3433 15555
rect 3467 15552 3479 15555
rect 3467 15524 4292 15552
rect 3467 15521 3479 15524
rect 3421 15515 3479 15521
rect 4264 15496 4292 15524
rect 3050 15444 3056 15496
rect 3108 15484 3114 15496
rect 3237 15487 3295 15493
rect 3237 15484 3249 15487
rect 3108 15456 3249 15484
rect 3108 15444 3114 15456
rect 3237 15453 3249 15456
rect 3283 15453 3295 15487
rect 4154 15484 4160 15496
rect 4115 15456 4160 15484
rect 3237 15447 3295 15453
rect 4154 15444 4160 15456
rect 4212 15444 4218 15496
rect 4246 15444 4252 15496
rect 4304 15484 4310 15496
rect 4304 15456 4349 15484
rect 4304 15444 4310 15456
rect 4982 15444 4988 15496
rect 5040 15484 5046 15496
rect 5261 15487 5319 15493
rect 5261 15484 5273 15487
rect 5040 15456 5273 15484
rect 5040 15444 5046 15456
rect 5261 15453 5273 15456
rect 5307 15484 5319 15487
rect 7101 15487 7159 15493
rect 7101 15484 7113 15487
rect 5307 15456 7113 15484
rect 5307 15453 5319 15456
rect 5261 15447 5319 15453
rect 7101 15453 7113 15456
rect 7147 15453 7159 15487
rect 7101 15447 7159 15453
rect 9122 15444 9128 15496
rect 9180 15484 9186 15496
rect 9493 15487 9551 15493
rect 9493 15484 9505 15487
rect 9180 15456 9505 15484
rect 9180 15444 9186 15456
rect 9493 15453 9505 15456
rect 9539 15453 9551 15487
rect 9493 15447 9551 15453
rect 11422 15444 11428 15496
rect 11480 15484 11486 15496
rect 12069 15487 12127 15493
rect 12069 15484 12081 15487
rect 11480 15456 12081 15484
rect 11480 15444 11486 15456
rect 12069 15453 12081 15456
rect 12115 15453 12127 15487
rect 12069 15447 12127 15453
rect 12253 15487 12311 15493
rect 12253 15453 12265 15487
rect 12299 15484 12311 15487
rect 12805 15487 12863 15493
rect 12805 15484 12817 15487
rect 12299 15456 12817 15484
rect 12299 15453 12311 15456
rect 12253 15447 12311 15453
rect 12805 15453 12817 15456
rect 12851 15453 12863 15487
rect 12805 15447 12863 15453
rect 12897 15487 12955 15493
rect 12897 15453 12909 15487
rect 12943 15484 12955 15487
rect 13262 15484 13268 15496
rect 12943 15456 13268 15484
rect 12943 15453 12955 15456
rect 12897 15447 12955 15453
rect 5528 15419 5586 15425
rect 5528 15385 5540 15419
rect 5574 15416 5586 15419
rect 6454 15416 6460 15428
rect 5574 15388 6460 15416
rect 5574 15385 5586 15388
rect 5528 15379 5586 15385
rect 6454 15376 6460 15388
rect 6512 15376 6518 15428
rect 7368 15419 7426 15425
rect 7368 15385 7380 15419
rect 7414 15416 7426 15419
rect 7466 15416 7472 15428
rect 7414 15388 7472 15416
rect 7414 15385 7426 15388
rect 7368 15379 7426 15385
rect 7466 15376 7472 15388
rect 7524 15376 7530 15428
rect 9760 15419 9818 15425
rect 9760 15385 9772 15419
rect 9806 15385 9818 15419
rect 12084 15416 12112 15447
rect 13262 15444 13268 15456
rect 13320 15444 13326 15496
rect 14553 15419 14611 15425
rect 14553 15416 14565 15419
rect 12084 15388 14565 15416
rect 9760 15379 9818 15385
rect 14553 15385 14565 15388
rect 14599 15385 14611 15419
rect 14553 15379 14611 15385
rect 14737 15419 14795 15425
rect 14737 15385 14749 15419
rect 14783 15416 14795 15419
rect 15838 15416 15844 15428
rect 14783 15388 15844 15416
rect 14783 15385 14795 15388
rect 14737 15379 14795 15385
rect 2774 15308 2780 15360
rect 2832 15348 2838 15360
rect 3053 15351 3111 15357
rect 3053 15348 3065 15351
rect 2832 15320 3065 15348
rect 2832 15308 2838 15320
rect 3053 15317 3065 15320
rect 3099 15317 3111 15351
rect 3970 15348 3976 15360
rect 3931 15320 3976 15348
rect 3053 15311 3111 15317
rect 3970 15308 3976 15320
rect 4028 15308 4034 15360
rect 6641 15351 6699 15357
rect 6641 15317 6653 15351
rect 6687 15348 6699 15351
rect 6822 15348 6828 15360
rect 6687 15320 6828 15348
rect 6687 15317 6699 15320
rect 6641 15311 6699 15317
rect 6822 15308 6828 15320
rect 6880 15308 6886 15360
rect 8018 15308 8024 15360
rect 8076 15348 8082 15360
rect 8481 15351 8539 15357
rect 8481 15348 8493 15351
rect 8076 15320 8493 15348
rect 8076 15308 8082 15320
rect 8481 15317 8493 15320
rect 8527 15317 8539 15351
rect 8481 15311 8539 15317
rect 9674 15308 9680 15360
rect 9732 15348 9738 15360
rect 9784 15348 9812 15379
rect 15838 15376 15844 15388
rect 15896 15376 15902 15428
rect 10870 15348 10876 15360
rect 9732 15320 9812 15348
rect 10831 15320 10876 15348
rect 9732 15308 9738 15320
rect 10870 15308 10876 15320
rect 10928 15308 10934 15360
rect 14642 15308 14648 15360
rect 14700 15348 14706 15360
rect 14921 15351 14979 15357
rect 14921 15348 14933 15351
rect 14700 15320 14933 15348
rect 14700 15308 14706 15320
rect 14921 15317 14933 15320
rect 14967 15317 14979 15351
rect 15746 15348 15752 15360
rect 15707 15320 15752 15348
rect 14921 15311 14979 15317
rect 15746 15308 15752 15320
rect 15804 15308 15810 15360
rect 1104 15258 19019 15280
rect 1104 15206 5388 15258
rect 5440 15206 5452 15258
rect 5504 15206 5516 15258
rect 5568 15206 5580 15258
rect 5632 15206 5644 15258
rect 5696 15206 9827 15258
rect 9879 15206 9891 15258
rect 9943 15206 9955 15258
rect 10007 15206 10019 15258
rect 10071 15206 10083 15258
rect 10135 15206 14266 15258
rect 14318 15206 14330 15258
rect 14382 15206 14394 15258
rect 14446 15206 14458 15258
rect 14510 15206 14522 15258
rect 14574 15206 18705 15258
rect 18757 15206 18769 15258
rect 18821 15206 18833 15258
rect 18885 15206 18897 15258
rect 18949 15206 18961 15258
rect 19013 15206 19019 15258
rect 1104 15184 19019 15206
rect 4154 15104 4160 15156
rect 4212 15144 4218 15156
rect 4341 15147 4399 15153
rect 4341 15144 4353 15147
rect 4212 15116 4353 15144
rect 4212 15104 4218 15116
rect 4341 15113 4353 15116
rect 4387 15113 4399 15147
rect 7466 15144 7472 15156
rect 7427 15116 7472 15144
rect 4341 15107 4399 15113
rect 7466 15104 7472 15116
rect 7524 15104 7530 15156
rect 9401 15147 9459 15153
rect 9401 15113 9413 15147
rect 9447 15144 9459 15147
rect 9674 15144 9680 15156
rect 9447 15116 9680 15144
rect 9447 15113 9459 15116
rect 9401 15107 9459 15113
rect 9674 15104 9680 15116
rect 9732 15104 9738 15156
rect 10229 15147 10287 15153
rect 10229 15113 10241 15147
rect 10275 15113 10287 15147
rect 15838 15144 15844 15156
rect 15799 15116 15844 15144
rect 10229 15107 10287 15113
rect 4982 15076 4988 15088
rect 2976 15048 4988 15076
rect 2976 15017 3004 15048
rect 4982 15036 4988 15048
rect 5040 15036 5046 15088
rect 10244 15076 10272 15107
rect 15838 15104 15844 15116
rect 15896 15104 15902 15156
rect 13814 15076 13820 15088
rect 9232 15048 10272 15076
rect 11992 15048 13820 15076
rect 2961 15011 3019 15017
rect 2961 14977 2973 15011
rect 3007 14977 3019 15011
rect 2961 14971 3019 14977
rect 3050 14968 3056 15020
rect 3108 15008 3114 15020
rect 3217 15011 3275 15017
rect 3217 15008 3229 15011
rect 3108 14980 3229 15008
rect 3108 14968 3114 14980
rect 3217 14977 3229 14980
rect 3263 14977 3275 15011
rect 3217 14971 3275 14977
rect 4246 14968 4252 15020
rect 4304 15008 4310 15020
rect 6641 15011 6699 15017
rect 6641 15008 6653 15011
rect 4304 14980 6653 15008
rect 4304 14968 4310 14980
rect 6641 14977 6653 14980
rect 6687 14977 6699 15011
rect 6822 15008 6828 15020
rect 6783 14980 6828 15008
rect 6641 14971 6699 14977
rect 6656 14940 6684 14971
rect 6822 14968 6828 14980
rect 6880 14968 6886 15020
rect 9232 15017 9260 15048
rect 7009 15011 7067 15017
rect 7009 14977 7021 15011
rect 7055 15008 7067 15011
rect 7653 15011 7711 15017
rect 7653 15008 7665 15011
rect 7055 14980 7665 15008
rect 7055 14977 7067 14980
rect 7009 14971 7067 14977
rect 7653 14977 7665 14980
rect 7699 14977 7711 15011
rect 7653 14971 7711 14977
rect 9217 15011 9275 15017
rect 9217 14977 9229 15011
rect 9263 14977 9275 15011
rect 9217 14971 9275 14977
rect 9674 14968 9680 15020
rect 9732 15008 9738 15020
rect 9861 15011 9919 15017
rect 9861 15008 9873 15011
rect 9732 14980 9873 15008
rect 9732 14968 9738 14980
rect 9861 14977 9873 14980
rect 9907 14977 9919 15011
rect 9861 14971 9919 14977
rect 10045 15011 10103 15017
rect 10045 14977 10057 15011
rect 10091 15008 10103 15011
rect 10226 15008 10232 15020
rect 10091 14980 10232 15008
rect 10091 14977 10103 14980
rect 10045 14971 10103 14977
rect 10226 14968 10232 14980
rect 10284 14968 10290 15020
rect 10870 15008 10876 15020
rect 10831 14980 10876 15008
rect 10870 14968 10876 14980
rect 10928 14968 10934 15020
rect 7098 14940 7104 14952
rect 6656 14912 7104 14940
rect 7098 14900 7104 14912
rect 7156 14900 7162 14952
rect 9122 14900 9128 14952
rect 9180 14940 9186 14952
rect 11992 14949 12020 15048
rect 13814 15036 13820 15048
rect 13872 15036 13878 15088
rect 16316 15048 17080 15076
rect 12244 15011 12302 15017
rect 12244 14977 12256 15011
rect 12290 15008 12302 15011
rect 12526 15008 12532 15020
rect 12290 14980 12532 15008
rect 12290 14977 12302 14980
rect 12244 14971 12302 14977
rect 12526 14968 12532 14980
rect 12584 14968 12590 15020
rect 14084 15011 14142 15017
rect 14084 14977 14096 15011
rect 14130 15008 14142 15011
rect 14918 15008 14924 15020
rect 14130 14980 14924 15008
rect 14130 14977 14142 14980
rect 14084 14971 14142 14977
rect 14918 14968 14924 14980
rect 14976 14968 14982 15020
rect 16206 15008 16212 15020
rect 15212 14980 16212 15008
rect 11977 14943 12035 14949
rect 11977 14940 11989 14943
rect 9180 14912 11989 14940
rect 9180 14900 9186 14912
rect 11977 14909 11989 14912
rect 12023 14909 12035 14943
rect 13814 14940 13820 14952
rect 13775 14912 13820 14940
rect 11977 14903 12035 14909
rect 13814 14900 13820 14912
rect 13872 14900 13878 14952
rect 15212 14881 15240 14980
rect 16206 14968 16212 14980
rect 16264 15008 16270 15020
rect 16316 15017 16344 15048
rect 16301 15011 16359 15017
rect 16301 15008 16313 15011
rect 16264 14980 16313 15008
rect 16264 14968 16270 14980
rect 16301 14977 16313 14980
rect 16347 14977 16359 15011
rect 16942 15008 16948 15020
rect 16903 14980 16948 15008
rect 16301 14971 16359 14977
rect 16942 14968 16948 14980
rect 17000 14968 17006 15020
rect 17052 15017 17080 15048
rect 17126 15036 17132 15088
rect 17184 15076 17190 15088
rect 17184 15048 17229 15076
rect 17184 15036 17190 15048
rect 17037 15011 17095 15017
rect 17037 14977 17049 15011
rect 17083 14977 17095 15011
rect 17037 14971 17095 14977
rect 17221 15011 17279 15017
rect 17221 14977 17233 15011
rect 17267 15008 17279 15011
rect 17310 15008 17316 15020
rect 17267 14980 17316 15008
rect 17267 14977 17279 14980
rect 17221 14971 17279 14977
rect 15197 14875 15255 14881
rect 15197 14841 15209 14875
rect 15243 14841 15255 14875
rect 17236 14872 17264 14971
rect 17310 14968 17316 14980
rect 17368 14968 17374 15020
rect 17405 14943 17463 14949
rect 17405 14909 17417 14943
rect 17451 14940 17463 14943
rect 17678 14940 17684 14952
rect 17451 14912 17684 14940
rect 17451 14909 17463 14912
rect 17405 14903 17463 14909
rect 17678 14900 17684 14912
rect 17736 14900 17742 14952
rect 15197 14835 15255 14841
rect 15304 14844 17264 14872
rect 5721 14807 5779 14813
rect 5721 14773 5733 14807
rect 5767 14804 5779 14807
rect 5810 14804 5816 14816
rect 5767 14776 5816 14804
rect 5767 14773 5779 14776
rect 5721 14767 5779 14773
rect 5810 14764 5816 14776
rect 5868 14764 5874 14816
rect 8386 14764 8392 14816
rect 8444 14804 8450 14816
rect 8665 14807 8723 14813
rect 8665 14804 8677 14807
rect 8444 14776 8677 14804
rect 8444 14764 8450 14776
rect 8665 14773 8677 14776
rect 8711 14773 8723 14807
rect 10778 14804 10784 14816
rect 10739 14776 10784 14804
rect 8665 14767 8723 14773
rect 10778 14764 10784 14776
rect 10836 14764 10842 14816
rect 13262 14764 13268 14816
rect 13320 14804 13326 14816
rect 13357 14807 13415 14813
rect 13357 14804 13369 14807
rect 13320 14776 13369 14804
rect 13320 14764 13326 14776
rect 13357 14773 13369 14776
rect 13403 14804 13415 14807
rect 15304 14804 15332 14844
rect 13403 14776 15332 14804
rect 16209 14807 16267 14813
rect 13403 14773 13415 14776
rect 13357 14767 13415 14773
rect 16209 14773 16221 14807
rect 16255 14804 16267 14807
rect 16942 14804 16948 14816
rect 16255 14776 16948 14804
rect 16255 14773 16267 14776
rect 16209 14767 16267 14773
rect 16942 14764 16948 14776
rect 17000 14764 17006 14816
rect 1104 14714 18860 14736
rect 1104 14662 3169 14714
rect 3221 14662 3233 14714
rect 3285 14662 3297 14714
rect 3349 14662 3361 14714
rect 3413 14662 3425 14714
rect 3477 14662 7608 14714
rect 7660 14662 7672 14714
rect 7724 14662 7736 14714
rect 7788 14662 7800 14714
rect 7852 14662 7864 14714
rect 7916 14662 12047 14714
rect 12099 14662 12111 14714
rect 12163 14662 12175 14714
rect 12227 14662 12239 14714
rect 12291 14662 12303 14714
rect 12355 14662 16486 14714
rect 16538 14662 16550 14714
rect 16602 14662 16614 14714
rect 16666 14662 16678 14714
rect 16730 14662 16742 14714
rect 16794 14662 18860 14714
rect 1104 14640 18860 14662
rect 6454 14600 6460 14612
rect 6415 14572 6460 14600
rect 6454 14560 6460 14572
rect 6512 14560 6518 14612
rect 7098 14560 7104 14612
rect 7156 14600 7162 14612
rect 11698 14600 11704 14612
rect 7156 14572 11704 14600
rect 7156 14560 7162 14572
rect 11698 14560 11704 14572
rect 11756 14560 11762 14612
rect 12345 14603 12403 14609
rect 12345 14569 12357 14603
rect 12391 14600 12403 14603
rect 12526 14600 12532 14612
rect 12391 14572 12532 14600
rect 12391 14569 12403 14572
rect 12345 14563 12403 14569
rect 12526 14560 12532 14572
rect 12584 14560 12590 14612
rect 13173 14603 13231 14609
rect 13173 14569 13185 14603
rect 13219 14600 13231 14603
rect 16850 14600 16856 14612
rect 13219 14572 16856 14600
rect 13219 14569 13231 14572
rect 13173 14563 13231 14569
rect 16850 14560 16856 14572
rect 16908 14560 16914 14612
rect 5537 14535 5595 14541
rect 5537 14501 5549 14535
rect 5583 14532 5595 14535
rect 5718 14532 5724 14544
rect 5583 14504 5724 14532
rect 5583 14501 5595 14504
rect 5537 14495 5595 14501
rect 5718 14492 5724 14504
rect 5776 14532 5782 14544
rect 6089 14535 6147 14541
rect 6089 14532 6101 14535
rect 5776 14504 6101 14532
rect 5776 14492 5782 14504
rect 6089 14501 6101 14504
rect 6135 14501 6147 14535
rect 14461 14535 14519 14541
rect 14461 14532 14473 14535
rect 6089 14495 6147 14501
rect 11072 14504 14473 14532
rect 3237 14399 3295 14405
rect 3237 14365 3249 14399
rect 3283 14396 3295 14399
rect 3970 14396 3976 14408
rect 3283 14368 3976 14396
rect 3283 14365 3295 14368
rect 3237 14359 3295 14365
rect 3970 14356 3976 14368
rect 4028 14356 4034 14408
rect 4157 14399 4215 14405
rect 4157 14365 4169 14399
rect 4203 14396 4215 14399
rect 4982 14396 4988 14408
rect 4203 14368 4988 14396
rect 4203 14365 4215 14368
rect 4157 14359 4215 14365
rect 4982 14356 4988 14368
rect 5040 14356 5046 14408
rect 5994 14396 6000 14408
rect 5955 14368 6000 14396
rect 5994 14356 6000 14368
rect 6052 14356 6058 14408
rect 6270 14396 6276 14408
rect 6231 14368 6276 14396
rect 6270 14356 6276 14368
rect 6328 14356 6334 14408
rect 6917 14399 6975 14405
rect 6917 14365 6929 14399
rect 6963 14396 6975 14399
rect 8294 14396 8300 14408
rect 6963 14368 8300 14396
rect 6963 14365 6975 14368
rect 6917 14359 6975 14365
rect 8294 14356 8300 14368
rect 8352 14396 8358 14408
rect 9122 14396 9128 14408
rect 8352 14368 9128 14396
rect 8352 14356 8358 14368
rect 9122 14356 9128 14368
rect 9180 14356 9186 14408
rect 11072 14405 11100 14504
rect 14461 14501 14473 14504
rect 14507 14532 14519 14535
rect 15378 14532 15384 14544
rect 14507 14504 15384 14532
rect 14507 14501 14519 14504
rect 14461 14495 14519 14501
rect 15378 14492 15384 14504
rect 15436 14492 15442 14544
rect 12618 14464 12624 14476
rect 11256 14436 12624 14464
rect 11256 14405 11284 14436
rect 11057 14399 11115 14405
rect 11057 14365 11069 14399
rect 11103 14365 11115 14399
rect 11057 14359 11115 14365
rect 11241 14399 11299 14405
rect 11241 14365 11253 14399
rect 11287 14365 11299 14399
rect 11698 14396 11704 14408
rect 11659 14368 11704 14396
rect 11241 14359 11299 14365
rect 11698 14356 11704 14368
rect 11756 14356 11762 14408
rect 12084 14405 12112 14436
rect 12618 14424 12624 14436
rect 12676 14464 12682 14476
rect 12805 14467 12863 14473
rect 12805 14464 12817 14467
rect 12676 14436 12817 14464
rect 12676 14424 12682 14436
rect 12805 14433 12817 14436
rect 12851 14433 12863 14467
rect 16206 14464 16212 14476
rect 16167 14436 16212 14464
rect 12805 14427 12863 14433
rect 16206 14424 16212 14436
rect 16264 14424 16270 14476
rect 16390 14464 16396 14476
rect 16351 14436 16396 14464
rect 16390 14424 16396 14436
rect 16448 14424 16454 14476
rect 16942 14424 16948 14476
rect 17000 14464 17006 14476
rect 17402 14464 17408 14476
rect 17000 14436 17408 14464
rect 17000 14424 17006 14436
rect 17402 14424 17408 14436
rect 17460 14464 17466 14476
rect 17589 14467 17647 14473
rect 17589 14464 17601 14467
rect 17460 14436 17601 14464
rect 17460 14424 17466 14436
rect 17589 14433 17601 14436
rect 17635 14433 17647 14467
rect 17589 14427 17647 14433
rect 11885 14399 11943 14405
rect 11885 14365 11897 14399
rect 11931 14365 11943 14399
rect 11885 14359 11943 14365
rect 11977 14399 12035 14405
rect 11977 14365 11989 14399
rect 12023 14365 12035 14399
rect 11977 14359 12035 14365
rect 12069 14399 12127 14405
rect 12069 14365 12081 14399
rect 12115 14365 12127 14399
rect 13262 14396 13268 14408
rect 13223 14368 13268 14396
rect 12069 14359 12127 14365
rect 4402 14331 4460 14337
rect 4402 14328 4414 14331
rect 3436 14300 4414 14328
rect 3436 14269 3464 14300
rect 4402 14297 4414 14300
rect 4448 14297 4460 14331
rect 4402 14291 4460 14297
rect 7006 14288 7012 14340
rect 7064 14328 7070 14340
rect 7162 14331 7220 14337
rect 7162 14328 7174 14331
rect 7064 14300 7174 14328
rect 7064 14288 7070 14300
rect 7162 14297 7174 14300
rect 7208 14297 7220 14331
rect 7162 14291 7220 14297
rect 9214 14288 9220 14340
rect 9272 14328 9278 14340
rect 9370 14331 9428 14337
rect 9370 14328 9382 14331
rect 9272 14300 9382 14328
rect 9272 14288 9278 14300
rect 9370 14297 9382 14300
rect 9416 14297 9428 14331
rect 9370 14291 9428 14297
rect 10410 14288 10416 14340
rect 10468 14328 10474 14340
rect 11149 14331 11207 14337
rect 10468 14300 11100 14328
rect 10468 14288 10474 14300
rect 3421 14263 3479 14269
rect 3421 14229 3433 14263
rect 3467 14229 3479 14263
rect 3421 14223 3479 14229
rect 7926 14220 7932 14272
rect 7984 14260 7990 14272
rect 8297 14263 8355 14269
rect 8297 14260 8309 14263
rect 7984 14232 8309 14260
rect 7984 14220 7990 14232
rect 8297 14229 8309 14232
rect 8343 14229 8355 14263
rect 10502 14260 10508 14272
rect 10463 14232 10508 14260
rect 8297 14223 8355 14229
rect 10502 14220 10508 14232
rect 10560 14220 10566 14272
rect 11072 14260 11100 14300
rect 11149 14297 11161 14331
rect 11195 14328 11207 14331
rect 11900 14328 11928 14359
rect 11195 14300 11928 14328
rect 11195 14297 11207 14300
rect 11149 14291 11207 14297
rect 11992 14260 12020 14359
rect 13262 14356 13268 14368
rect 13320 14356 13326 14408
rect 14369 14399 14427 14405
rect 14369 14365 14381 14399
rect 14415 14365 14427 14399
rect 14642 14396 14648 14408
rect 14603 14368 14648 14396
rect 14369 14359 14427 14365
rect 14384 14328 14412 14359
rect 14642 14356 14648 14368
rect 14700 14356 14706 14408
rect 15838 14356 15844 14408
rect 15896 14396 15902 14408
rect 16117 14399 16175 14405
rect 16117 14396 16129 14399
rect 15896 14368 16129 14396
rect 15896 14356 15902 14368
rect 16117 14365 16129 14368
rect 16163 14365 16175 14399
rect 16224 14396 16252 14424
rect 17104 14399 17162 14405
rect 17104 14396 17116 14399
rect 16224 14368 17116 14396
rect 16117 14359 16175 14365
rect 17104 14365 17116 14368
rect 17150 14365 17162 14399
rect 17104 14359 17162 14365
rect 17310 14328 17316 14340
rect 14384 14300 15792 14328
rect 14090 14260 14096 14272
rect 11072 14232 14096 14260
rect 14090 14220 14096 14232
rect 14148 14220 14154 14272
rect 14826 14260 14832 14272
rect 14787 14232 14832 14260
rect 14826 14220 14832 14232
rect 14884 14220 14890 14272
rect 15764 14269 15792 14300
rect 17052 14300 17316 14328
rect 17052 14272 17080 14300
rect 17310 14288 17316 14300
rect 17368 14288 17374 14340
rect 15749 14263 15807 14269
rect 15749 14229 15761 14263
rect 15795 14260 15807 14263
rect 15838 14260 15844 14272
rect 15795 14232 15844 14260
rect 15795 14229 15807 14232
rect 15749 14223 15807 14229
rect 15838 14220 15844 14232
rect 15896 14220 15902 14272
rect 16942 14260 16948 14272
rect 16903 14232 16948 14260
rect 16942 14220 16948 14232
rect 17000 14220 17006 14272
rect 17034 14220 17040 14272
rect 17092 14220 17098 14272
rect 17126 14220 17132 14272
rect 17184 14260 17190 14272
rect 17221 14263 17279 14269
rect 17221 14260 17233 14263
rect 17184 14232 17233 14260
rect 17184 14220 17190 14232
rect 17221 14229 17233 14232
rect 17267 14229 17279 14263
rect 17221 14223 17279 14229
rect 1104 14170 19019 14192
rect 1104 14118 5388 14170
rect 5440 14118 5452 14170
rect 5504 14118 5516 14170
rect 5568 14118 5580 14170
rect 5632 14118 5644 14170
rect 5696 14118 9827 14170
rect 9879 14118 9891 14170
rect 9943 14118 9955 14170
rect 10007 14118 10019 14170
rect 10071 14118 10083 14170
rect 10135 14118 14266 14170
rect 14318 14118 14330 14170
rect 14382 14118 14394 14170
rect 14446 14118 14458 14170
rect 14510 14118 14522 14170
rect 14574 14118 18705 14170
rect 18757 14118 18769 14170
rect 18821 14118 18833 14170
rect 18885 14118 18897 14170
rect 18949 14118 18961 14170
rect 19013 14118 19019 14170
rect 1104 14096 19019 14118
rect 3053 14059 3111 14065
rect 3053 14056 3065 14059
rect 2746 14028 3065 14056
rect 2746 13932 2774 14028
rect 3053 14025 3065 14028
rect 3099 14025 3111 14059
rect 3053 14019 3111 14025
rect 5359 14059 5417 14065
rect 5359 14025 5371 14059
rect 5405 14056 5417 14059
rect 6270 14056 6276 14068
rect 5405 14028 6276 14056
rect 5405 14025 5417 14028
rect 5359 14019 5417 14025
rect 6270 14016 6276 14028
rect 6328 14016 6334 14068
rect 7006 14056 7012 14068
rect 6967 14028 7012 14056
rect 7006 14016 7012 14028
rect 7064 14016 7070 14068
rect 9214 14056 9220 14068
rect 9175 14028 9220 14056
rect 9214 14016 9220 14028
rect 9272 14016 9278 14068
rect 9674 14016 9680 14068
rect 9732 14056 9738 14068
rect 9861 14059 9919 14065
rect 9861 14056 9873 14059
rect 9732 14028 9873 14056
rect 9732 14016 9738 14028
rect 9861 14025 9873 14028
rect 9907 14025 9919 14059
rect 12618 14056 12624 14068
rect 12579 14028 12624 14056
rect 9861 14019 9919 14025
rect 12618 14016 12624 14028
rect 12676 14016 12682 14068
rect 14918 14056 14924 14068
rect 14879 14028 14924 14056
rect 14918 14016 14924 14028
rect 14976 14016 14982 14068
rect 15470 14016 15476 14068
rect 15528 14056 15534 14068
rect 15933 14059 15991 14065
rect 15933 14056 15945 14059
rect 15528 14028 15945 14056
rect 15528 14016 15534 14028
rect 15933 14025 15945 14028
rect 15979 14025 15991 14059
rect 15933 14019 15991 14025
rect 17037 14059 17095 14065
rect 17037 14025 17049 14059
rect 17083 14056 17095 14059
rect 17126 14056 17132 14068
rect 17083 14028 17132 14056
rect 17083 14025 17095 14028
rect 17037 14019 17095 14025
rect 17126 14016 17132 14028
rect 17184 14056 17190 14068
rect 17954 14056 17960 14068
rect 17184 14028 17960 14056
rect 17184 14016 17190 14028
rect 17954 14016 17960 14028
rect 18012 14016 18018 14068
rect 18049 14059 18107 14065
rect 18049 14025 18061 14059
rect 18095 14025 18107 14059
rect 18049 14019 18107 14025
rect 5445 13991 5503 13997
rect 5445 13988 5457 13991
rect 2314 13920 2320 13932
rect 2275 13892 2320 13920
rect 2314 13880 2320 13892
rect 2372 13880 2378 13932
rect 2501 13923 2559 13929
rect 2501 13889 2513 13923
rect 2547 13920 2559 13923
rect 2682 13920 2688 13932
rect 2547 13892 2688 13920
rect 2547 13889 2559 13892
rect 2501 13883 2559 13889
rect 2682 13880 2688 13892
rect 2740 13892 2774 13932
rect 3436 13960 5457 13988
rect 2740 13880 2746 13892
rect 2590 13852 2596 13864
rect 2503 13824 2596 13852
rect 2590 13812 2596 13824
rect 2648 13852 2654 13864
rect 3436 13852 3464 13960
rect 5445 13957 5457 13960
rect 5491 13988 5503 13991
rect 5994 13988 6000 14000
rect 5491 13960 6000 13988
rect 5491 13957 5503 13960
rect 5445 13951 5503 13957
rect 5994 13948 6000 13960
rect 6052 13948 6058 14000
rect 7098 13948 7104 14000
rect 7156 13988 7162 14000
rect 7156 13960 7696 13988
rect 7156 13948 7162 13960
rect 4154 13920 4160 13932
rect 4212 13929 4218 13932
rect 4124 13892 4160 13920
rect 4154 13880 4160 13892
rect 4212 13883 4224 13929
rect 4212 13880 4218 13883
rect 4338 13880 4344 13932
rect 4396 13920 4402 13932
rect 5261 13923 5319 13929
rect 5261 13920 5273 13923
rect 4396 13892 5273 13920
rect 4396 13880 4402 13892
rect 5261 13889 5273 13892
rect 5307 13889 5319 13923
rect 5261 13883 5319 13889
rect 5537 13923 5595 13929
rect 5537 13889 5549 13923
rect 5583 13920 5595 13923
rect 5718 13920 5724 13932
rect 5583 13892 5724 13920
rect 5583 13889 5595 13892
rect 5537 13883 5595 13889
rect 2648 13824 3464 13852
rect 4433 13855 4491 13861
rect 2648 13812 2654 13824
rect 4433 13821 4445 13855
rect 4479 13852 4491 13855
rect 4982 13852 4988 13864
rect 4479 13824 4988 13852
rect 4479 13821 4491 13824
rect 4433 13815 4491 13821
rect 4982 13812 4988 13824
rect 5040 13812 5046 13864
rect 5276 13852 5304 13883
rect 5718 13880 5724 13892
rect 5776 13880 5782 13932
rect 7190 13880 7196 13932
rect 7248 13920 7254 13932
rect 7285 13923 7343 13929
rect 7285 13920 7297 13923
rect 7248 13892 7297 13920
rect 7248 13880 7254 13892
rect 7285 13889 7297 13892
rect 7331 13889 7343 13923
rect 7285 13883 7343 13889
rect 7377 13923 7435 13929
rect 7377 13889 7389 13923
rect 7423 13889 7435 13923
rect 7377 13883 7435 13889
rect 5810 13852 5816 13864
rect 5276 13824 5816 13852
rect 5810 13812 5816 13824
rect 5868 13812 5874 13864
rect 7392 13852 7420 13883
rect 7466 13880 7472 13932
rect 7524 13920 7530 13932
rect 7668 13929 7696 13960
rect 8588 13960 9168 13988
rect 8588 13929 8616 13960
rect 7653 13923 7711 13929
rect 7524 13892 7569 13920
rect 7524 13880 7530 13892
rect 7653 13889 7665 13923
rect 7699 13889 7711 13923
rect 7653 13883 7711 13889
rect 8573 13923 8631 13929
rect 8573 13889 8585 13923
rect 8619 13889 8631 13923
rect 8754 13920 8760 13932
rect 8715 13892 8760 13920
rect 8573 13883 8631 13889
rect 8754 13880 8760 13892
rect 8812 13880 8818 13932
rect 9030 13920 9036 13932
rect 8991 13892 9036 13920
rect 9030 13880 9036 13892
rect 9088 13880 9094 13932
rect 9140 13920 9168 13960
rect 9306 13948 9312 14000
rect 9364 13988 9370 14000
rect 10318 13988 10324 14000
rect 9364 13960 10324 13988
rect 9364 13948 9370 13960
rect 10318 13948 10324 13960
rect 10376 13948 10382 14000
rect 12529 13991 12587 13997
rect 12529 13957 12541 13991
rect 12575 13988 12587 13991
rect 13262 13988 13268 14000
rect 12575 13960 13268 13988
rect 12575 13957 12587 13960
rect 12529 13951 12587 13957
rect 13262 13948 13268 13960
rect 13320 13948 13326 14000
rect 14200 13960 15056 13988
rect 14200 13932 14228 13960
rect 10229 13923 10287 13929
rect 9140 13892 10180 13920
rect 7300 13824 7420 13852
rect 8772 13852 8800 13880
rect 9950 13852 9956 13864
rect 8772 13824 9956 13852
rect 7300 13796 7328 13824
rect 9950 13812 9956 13824
rect 10008 13852 10014 13864
rect 10152 13861 10180 13892
rect 10229 13889 10241 13923
rect 10275 13920 10287 13923
rect 10778 13920 10784 13932
rect 10275 13892 10784 13920
rect 10275 13889 10287 13892
rect 10229 13883 10287 13889
rect 10778 13880 10784 13892
rect 10836 13880 10842 13932
rect 13725 13923 13783 13929
rect 10980 13892 13492 13920
rect 10045 13855 10103 13861
rect 10045 13852 10057 13855
rect 10008 13824 10057 13852
rect 10008 13812 10014 13824
rect 10045 13821 10057 13824
rect 10091 13821 10103 13855
rect 10045 13815 10103 13821
rect 10137 13855 10195 13861
rect 10137 13821 10149 13855
rect 10183 13821 10195 13855
rect 10318 13852 10324 13864
rect 10279 13824 10324 13852
rect 10137 13815 10195 13821
rect 2133 13787 2191 13793
rect 2133 13753 2145 13787
rect 2179 13784 2191 13787
rect 3050 13784 3056 13796
rect 2179 13756 3056 13784
rect 2179 13753 2191 13756
rect 2133 13747 2191 13753
rect 3050 13744 3056 13756
rect 3108 13744 3114 13796
rect 7282 13744 7288 13796
rect 7340 13744 7346 13796
rect 10152 13784 10180 13815
rect 10318 13812 10324 13824
rect 10376 13812 10382 13864
rect 10870 13852 10876 13864
rect 10428 13824 10876 13852
rect 10428 13784 10456 13824
rect 10870 13812 10876 13824
rect 10928 13812 10934 13864
rect 10152 13756 10456 13784
rect 8386 13676 8392 13728
rect 8444 13716 8450 13728
rect 9582 13716 9588 13728
rect 8444 13688 9588 13716
rect 8444 13676 8450 13688
rect 9582 13676 9588 13688
rect 9640 13716 9646 13728
rect 10873 13719 10931 13725
rect 10873 13716 10885 13719
rect 9640 13688 10885 13716
rect 9640 13676 9646 13688
rect 10873 13685 10885 13688
rect 10919 13716 10931 13719
rect 10980 13716 11008 13892
rect 12345 13855 12403 13861
rect 12345 13821 12357 13855
rect 12391 13821 12403 13855
rect 13464 13852 13492 13892
rect 13725 13889 13737 13923
rect 13771 13920 13783 13923
rect 14182 13920 14188 13932
rect 13771 13892 14188 13920
rect 13771 13889 13783 13892
rect 13725 13883 13783 13889
rect 14182 13880 14188 13892
rect 14240 13880 14246 13932
rect 14369 13923 14427 13929
rect 14369 13889 14381 13923
rect 14415 13920 14427 13923
rect 14642 13920 14648 13932
rect 14415 13892 14648 13920
rect 14415 13889 14427 13892
rect 14369 13883 14427 13889
rect 14642 13880 14648 13892
rect 14700 13880 14706 13932
rect 14826 13920 14832 13932
rect 14787 13892 14832 13920
rect 14826 13880 14832 13892
rect 14884 13880 14890 13932
rect 15028 13929 15056 13960
rect 16850 13948 16856 14000
rect 16908 13988 16914 14000
rect 17770 13988 17776 14000
rect 16908 13960 17776 13988
rect 16908 13948 16914 13960
rect 17770 13948 17776 13960
rect 17828 13988 17834 14000
rect 18064 13988 18092 14019
rect 17828 13960 18092 13988
rect 17828 13948 17834 13960
rect 15013 13923 15071 13929
rect 15013 13889 15025 13923
rect 15059 13889 15071 13923
rect 15013 13883 15071 13889
rect 16301 13923 16359 13929
rect 16301 13889 16313 13923
rect 16347 13889 16359 13923
rect 17402 13920 17408 13932
rect 17363 13892 17408 13920
rect 16301 13883 16359 13889
rect 15746 13852 15752 13864
rect 13464 13824 15752 13852
rect 12345 13815 12403 13821
rect 12360 13784 12388 13815
rect 15746 13812 15752 13824
rect 15804 13852 15810 13864
rect 16209 13855 16267 13861
rect 16209 13852 16221 13855
rect 15804 13824 16221 13852
rect 15804 13812 15810 13824
rect 16209 13821 16221 13824
rect 16255 13821 16267 13855
rect 16316 13852 16344 13883
rect 17402 13880 17408 13892
rect 17460 13920 17466 13932
rect 17865 13923 17923 13929
rect 17865 13920 17877 13923
rect 17460 13892 17877 13920
rect 17460 13880 17466 13892
rect 17865 13889 17877 13892
rect 17911 13889 17923 13923
rect 17865 13883 17923 13889
rect 18046 13852 18052 13864
rect 16316 13824 18052 13852
rect 16209 13815 16267 13821
rect 18046 13812 18052 13824
rect 18104 13812 18110 13864
rect 12434 13784 12440 13796
rect 12360 13756 12440 13784
rect 12434 13744 12440 13756
rect 12492 13744 12498 13796
rect 12986 13716 12992 13728
rect 10919 13688 11008 13716
rect 12947 13688 12992 13716
rect 10919 13685 10931 13688
rect 10873 13679 10931 13685
rect 12986 13676 12992 13688
rect 13044 13676 13050 13728
rect 14366 13716 14372 13728
rect 14327 13688 14372 13716
rect 14366 13676 14372 13688
rect 14424 13676 14430 13728
rect 16301 13719 16359 13725
rect 16301 13685 16313 13719
rect 16347 13716 16359 13719
rect 16390 13716 16396 13728
rect 16347 13688 16396 13716
rect 16347 13685 16359 13688
rect 16301 13679 16359 13685
rect 16390 13676 16396 13688
rect 16448 13716 16454 13728
rect 16853 13719 16911 13725
rect 16853 13716 16865 13719
rect 16448 13688 16865 13716
rect 16448 13676 16454 13688
rect 16853 13685 16865 13688
rect 16899 13685 16911 13719
rect 17034 13716 17040 13728
rect 16995 13688 17040 13716
rect 16853 13679 16911 13685
rect 17034 13676 17040 13688
rect 17092 13676 17098 13728
rect 1104 13626 18860 13648
rect 1104 13574 3169 13626
rect 3221 13574 3233 13626
rect 3285 13574 3297 13626
rect 3349 13574 3361 13626
rect 3413 13574 3425 13626
rect 3477 13574 7608 13626
rect 7660 13574 7672 13626
rect 7724 13574 7736 13626
rect 7788 13574 7800 13626
rect 7852 13574 7864 13626
rect 7916 13574 12047 13626
rect 12099 13574 12111 13626
rect 12163 13574 12175 13626
rect 12227 13574 12239 13626
rect 12291 13574 12303 13626
rect 12355 13574 16486 13626
rect 16538 13574 16550 13626
rect 16602 13574 16614 13626
rect 16666 13574 16678 13626
rect 16730 13574 16742 13626
rect 16794 13574 18860 13626
rect 1104 13552 18860 13574
rect 2314 13472 2320 13524
rect 2372 13512 2378 13524
rect 2409 13515 2467 13521
rect 2409 13512 2421 13515
rect 2372 13484 2421 13512
rect 2372 13472 2378 13484
rect 2409 13481 2421 13484
rect 2455 13481 2467 13515
rect 3237 13515 3295 13521
rect 3237 13512 3249 13515
rect 2409 13475 2467 13481
rect 2746 13484 3249 13512
rect 2746 13376 2774 13484
rect 3237 13481 3249 13484
rect 3283 13512 3295 13515
rect 4338 13512 4344 13524
rect 3283 13484 4344 13512
rect 3283 13481 3295 13484
rect 3237 13475 3295 13481
rect 4338 13472 4344 13484
rect 4396 13472 4402 13524
rect 7466 13472 7472 13524
rect 7524 13512 7530 13524
rect 7561 13515 7619 13521
rect 7561 13512 7573 13515
rect 7524 13484 7573 13512
rect 7524 13472 7530 13484
rect 7561 13481 7573 13484
rect 7607 13481 7619 13515
rect 9125 13515 9183 13521
rect 9125 13512 9137 13515
rect 7561 13475 7619 13481
rect 8312 13484 9137 13512
rect 7190 13404 7196 13456
rect 7248 13444 7254 13456
rect 8202 13444 8208 13456
rect 7248 13416 8208 13444
rect 7248 13404 7254 13416
rect 8202 13404 8208 13416
rect 8260 13444 8266 13456
rect 8312 13444 8340 13484
rect 9125 13481 9137 13484
rect 9171 13481 9183 13515
rect 9125 13475 9183 13481
rect 10045 13515 10103 13521
rect 10045 13481 10057 13515
rect 10091 13512 10103 13515
rect 10226 13512 10232 13524
rect 10091 13484 10232 13512
rect 10091 13481 10103 13484
rect 10045 13475 10103 13481
rect 10226 13472 10232 13484
rect 10284 13472 10290 13524
rect 18046 13512 18052 13524
rect 18007 13484 18052 13512
rect 18046 13472 18052 13484
rect 18104 13472 18110 13524
rect 8260 13416 8340 13444
rect 8260 13404 8266 13416
rect 9582 13404 9588 13456
rect 9640 13444 9646 13456
rect 10137 13447 10195 13453
rect 9640 13416 9996 13444
rect 9640 13404 9646 13416
rect 9968 13376 9996 13416
rect 10137 13413 10149 13447
rect 10183 13444 10195 13447
rect 10318 13444 10324 13456
rect 10183 13416 10324 13444
rect 10183 13413 10195 13416
rect 10137 13407 10195 13413
rect 10045 13379 10103 13385
rect 10045 13376 10057 13379
rect 2424 13348 2774 13376
rect 8582 13348 9674 13376
rect 9968 13348 10057 13376
rect 2222 13268 2228 13320
rect 2280 13308 2286 13320
rect 2424 13317 2452 13348
rect 2409 13311 2467 13317
rect 2409 13308 2421 13311
rect 2280 13280 2421 13308
rect 2280 13268 2286 13280
rect 2409 13277 2421 13280
rect 2455 13277 2467 13311
rect 2682 13308 2688 13320
rect 2643 13280 2688 13308
rect 2409 13271 2467 13277
rect 2682 13268 2688 13280
rect 2740 13268 2746 13320
rect 4982 13268 4988 13320
rect 5040 13308 5046 13320
rect 5629 13311 5687 13317
rect 5629 13308 5641 13311
rect 5040 13280 5641 13308
rect 5040 13268 5046 13280
rect 5629 13277 5641 13280
rect 5675 13277 5687 13311
rect 5629 13271 5687 13277
rect 7282 13268 7288 13320
rect 7340 13308 7346 13320
rect 7469 13311 7527 13317
rect 7469 13308 7481 13311
rect 7340 13280 7481 13308
rect 7340 13268 7346 13280
rect 7469 13277 7481 13280
rect 7515 13277 7527 13311
rect 7469 13271 7527 13277
rect 7653 13311 7711 13317
rect 7653 13277 7665 13311
rect 7699 13308 7711 13311
rect 7926 13308 7932 13320
rect 7699 13280 7932 13308
rect 7699 13277 7711 13280
rect 7653 13271 7711 13277
rect 7926 13268 7932 13280
rect 7984 13268 7990 13320
rect 8386 13308 8392 13320
rect 8347 13280 8392 13308
rect 8386 13268 8392 13280
rect 8444 13268 8450 13320
rect 8582 13317 8610 13348
rect 8573 13311 8631 13317
rect 8573 13277 8585 13311
rect 8619 13277 8631 13311
rect 8573 13271 8631 13277
rect 9309 13311 9367 13317
rect 9309 13277 9321 13311
rect 9355 13277 9367 13311
rect 9309 13271 9367 13277
rect 2590 13240 2596 13252
rect 2551 13212 2596 13240
rect 2590 13200 2596 13212
rect 2648 13200 2654 13252
rect 5902 13249 5908 13252
rect 5896 13203 5908 13249
rect 5960 13240 5966 13252
rect 7944 13240 7972 13268
rect 8938 13240 8944 13252
rect 5960 13212 5996 13240
rect 7944 13212 8944 13240
rect 5902 13200 5908 13203
rect 5960 13200 5966 13212
rect 8938 13200 8944 13212
rect 8996 13240 9002 13252
rect 9324 13240 9352 13271
rect 9398 13268 9404 13320
rect 9456 13308 9462 13320
rect 9646 13308 9674 13348
rect 10045 13345 10057 13348
rect 10091 13345 10103 13379
rect 10045 13339 10103 13345
rect 10152 13308 10180 13407
rect 10318 13404 10324 13416
rect 10376 13444 10382 13456
rect 10778 13444 10784 13456
rect 10376 13416 10784 13444
rect 10376 13404 10382 13416
rect 10778 13404 10784 13416
rect 10836 13404 10842 13456
rect 12250 13376 12256 13388
rect 12211 13348 12256 13376
rect 12250 13336 12256 13348
rect 12308 13336 12314 13388
rect 17034 13336 17040 13388
rect 17092 13376 17098 13388
rect 17092 13348 18276 13376
rect 17092 13336 17098 13348
rect 9456 13280 9501 13308
rect 9646 13280 10180 13308
rect 10321 13311 10379 13317
rect 9456 13268 9462 13280
rect 10321 13277 10333 13311
rect 10367 13308 10379 13311
rect 10502 13308 10508 13320
rect 10367 13280 10508 13308
rect 10367 13277 10379 13280
rect 10321 13271 10379 13277
rect 10502 13268 10508 13280
rect 10560 13268 10566 13320
rect 10594 13268 10600 13320
rect 10652 13308 10658 13320
rect 10873 13311 10931 13317
rect 10873 13308 10885 13311
rect 10652 13280 10885 13308
rect 10652 13268 10658 13280
rect 10873 13277 10885 13280
rect 10919 13277 10931 13311
rect 12158 13308 12164 13320
rect 12119 13280 12164 13308
rect 10873 13271 10931 13277
rect 12158 13268 12164 13280
rect 12216 13268 12222 13320
rect 13814 13268 13820 13320
rect 13872 13308 13878 13320
rect 14277 13311 14335 13317
rect 14277 13308 14289 13311
rect 13872 13280 14289 13308
rect 13872 13268 13878 13280
rect 14277 13277 14289 13280
rect 14323 13277 14335 13311
rect 14277 13271 14335 13277
rect 14366 13268 14372 13320
rect 14424 13308 14430 13320
rect 14533 13311 14591 13317
rect 14533 13308 14545 13311
rect 14424 13280 14545 13308
rect 14424 13268 14430 13280
rect 14533 13277 14545 13280
rect 14579 13277 14591 13311
rect 14533 13271 14591 13277
rect 16761 13311 16819 13317
rect 16761 13277 16773 13311
rect 16807 13308 16819 13311
rect 16850 13308 16856 13320
rect 16807 13280 16856 13308
rect 16807 13277 16819 13280
rect 16761 13271 16819 13277
rect 16850 13268 16856 13280
rect 16908 13268 16914 13320
rect 17402 13268 17408 13320
rect 17460 13308 17466 13320
rect 17589 13311 17647 13317
rect 17589 13308 17601 13311
rect 17460 13280 17601 13308
rect 17460 13268 17466 13280
rect 17589 13277 17601 13280
rect 17635 13277 17647 13311
rect 17589 13271 17647 13277
rect 17954 13268 17960 13320
rect 18012 13308 18018 13320
rect 18248 13317 18276 13348
rect 18049 13311 18107 13317
rect 18049 13308 18061 13311
rect 18012 13280 18061 13308
rect 18012 13268 18018 13280
rect 18049 13277 18061 13280
rect 18095 13277 18107 13311
rect 18049 13271 18107 13277
rect 18233 13311 18291 13317
rect 18233 13277 18245 13311
rect 18279 13277 18291 13311
rect 18233 13271 18291 13277
rect 8996 13212 9352 13240
rect 8996 13200 9002 13212
rect 9950 13200 9956 13252
rect 10008 13240 10014 13252
rect 10413 13243 10471 13249
rect 10413 13240 10425 13243
rect 10008 13212 10425 13240
rect 10008 13200 10014 13212
rect 10413 13209 10425 13212
rect 10459 13209 10471 13243
rect 16574 13240 16580 13252
rect 16535 13212 16580 13240
rect 10413 13203 10471 13209
rect 16574 13200 16580 13212
rect 16632 13200 16638 13252
rect 16945 13243 17003 13249
rect 16945 13209 16957 13243
rect 16991 13240 17003 13243
rect 17126 13240 17132 13252
rect 16991 13212 17132 13240
rect 16991 13209 17003 13212
rect 16945 13203 17003 13209
rect 7006 13172 7012 13184
rect 6967 13144 7012 13172
rect 7006 13132 7012 13144
rect 7064 13132 7070 13184
rect 8481 13175 8539 13181
rect 8481 13141 8493 13175
rect 8527 13172 8539 13175
rect 10962 13172 10968 13184
rect 8527 13144 10968 13172
rect 8527 13141 8539 13144
rect 8481 13135 8539 13141
rect 10962 13132 10968 13144
rect 11020 13132 11026 13184
rect 11057 13175 11115 13181
rect 11057 13141 11069 13175
rect 11103 13172 11115 13175
rect 11422 13172 11428 13184
rect 11103 13144 11428 13172
rect 11103 13141 11115 13144
rect 11057 13135 11115 13141
rect 11422 13132 11428 13144
rect 11480 13132 11486 13184
rect 12529 13175 12587 13181
rect 12529 13141 12541 13175
rect 12575 13172 12587 13175
rect 12710 13172 12716 13184
rect 12575 13144 12716 13172
rect 12575 13141 12587 13144
rect 12529 13135 12587 13141
rect 12710 13132 12716 13144
rect 12768 13132 12774 13184
rect 15654 13172 15660 13184
rect 15567 13144 15660 13172
rect 15654 13132 15660 13144
rect 15712 13172 15718 13184
rect 16960 13172 16988 13203
rect 17126 13200 17132 13212
rect 17184 13200 17190 13252
rect 17494 13172 17500 13184
rect 15712 13144 16988 13172
rect 17455 13144 17500 13172
rect 15712 13132 15718 13144
rect 17494 13132 17500 13144
rect 17552 13132 17558 13184
rect 1104 13082 19019 13104
rect 1104 13030 5388 13082
rect 5440 13030 5452 13082
rect 5504 13030 5516 13082
rect 5568 13030 5580 13082
rect 5632 13030 5644 13082
rect 5696 13030 9827 13082
rect 9879 13030 9891 13082
rect 9943 13030 9955 13082
rect 10007 13030 10019 13082
rect 10071 13030 10083 13082
rect 10135 13030 14266 13082
rect 14318 13030 14330 13082
rect 14382 13030 14394 13082
rect 14446 13030 14458 13082
rect 14510 13030 14522 13082
rect 14574 13030 18705 13082
rect 18757 13030 18769 13082
rect 18821 13030 18833 13082
rect 18885 13030 18897 13082
rect 18949 13030 18961 13082
rect 19013 13030 19019 13082
rect 1104 13008 19019 13030
rect 2685 12971 2743 12977
rect 2685 12937 2697 12971
rect 2731 12968 2743 12971
rect 4154 12968 4160 12980
rect 2731 12940 4160 12968
rect 2731 12937 2743 12940
rect 2685 12931 2743 12937
rect 4154 12928 4160 12940
rect 4212 12928 4218 12980
rect 5813 12971 5871 12977
rect 5813 12937 5825 12971
rect 5859 12968 5871 12971
rect 5902 12968 5908 12980
rect 5859 12940 5908 12968
rect 5859 12937 5871 12940
rect 5813 12931 5871 12937
rect 5902 12928 5908 12940
rect 5960 12928 5966 12980
rect 8294 12968 8300 12980
rect 8255 12940 8300 12968
rect 8294 12928 8300 12940
rect 8352 12928 8358 12980
rect 10594 12968 10600 12980
rect 10555 12940 10600 12968
rect 10594 12928 10600 12940
rect 10652 12928 10658 12980
rect 14182 12968 14188 12980
rect 14143 12940 14188 12968
rect 14182 12928 14188 12940
rect 14240 12928 14246 12980
rect 14642 12928 14648 12980
rect 14700 12968 14706 12980
rect 14737 12971 14795 12977
rect 14737 12968 14749 12971
rect 14700 12940 14749 12968
rect 14700 12928 14706 12940
rect 14737 12937 14749 12940
rect 14783 12937 14795 12971
rect 14737 12931 14795 12937
rect 14921 12971 14979 12977
rect 14921 12937 14933 12971
rect 14967 12937 14979 12971
rect 14921 12931 14979 12937
rect 2406 12900 2412 12912
rect 2240 12872 2412 12900
rect 2240 12841 2268 12872
rect 2406 12860 2412 12872
rect 2464 12900 2470 12912
rect 2590 12900 2596 12912
rect 2464 12872 2596 12900
rect 2464 12860 2470 12872
rect 2590 12860 2596 12872
rect 2648 12860 2654 12912
rect 9490 12860 9496 12912
rect 9548 12900 9554 12912
rect 10137 12903 10195 12909
rect 10137 12900 10149 12903
rect 9548 12872 10149 12900
rect 9548 12860 9554 12872
rect 10137 12869 10149 12872
rect 10183 12869 10195 12903
rect 12434 12900 12440 12912
rect 10137 12863 10195 12869
rect 11716 12872 12440 12900
rect 2225 12835 2283 12841
rect 2225 12801 2237 12835
rect 2271 12801 2283 12835
rect 2498 12832 2504 12844
rect 2459 12804 2504 12832
rect 2225 12795 2283 12801
rect 2498 12792 2504 12804
rect 2556 12792 2562 12844
rect 4246 12792 4252 12844
rect 4304 12832 4310 12844
rect 4718 12835 4776 12841
rect 4718 12832 4730 12835
rect 4304 12804 4730 12832
rect 4304 12792 4310 12804
rect 4718 12801 4730 12804
rect 4764 12801 4776 12835
rect 5994 12832 6000 12844
rect 5955 12804 6000 12832
rect 4718 12795 4776 12801
rect 5994 12792 6000 12804
rect 6052 12792 6058 12844
rect 7190 12832 7196 12844
rect 7151 12804 7196 12832
rect 7190 12792 7196 12804
rect 7248 12792 7254 12844
rect 9585 12835 9643 12841
rect 9585 12801 9597 12835
rect 9631 12832 9643 12835
rect 9674 12832 9680 12844
rect 9631 12804 9680 12832
rect 9631 12801 9643 12804
rect 9585 12795 9643 12801
rect 9674 12792 9680 12804
rect 9732 12792 9738 12844
rect 10318 12832 10324 12844
rect 10279 12804 10324 12832
rect 10318 12792 10324 12804
rect 10376 12792 10382 12844
rect 10413 12835 10471 12841
rect 10413 12801 10425 12835
rect 10459 12832 10471 12835
rect 11606 12832 11612 12844
rect 10459 12804 11612 12832
rect 10459 12801 10471 12804
rect 10413 12795 10471 12801
rect 4982 12724 4988 12776
rect 5040 12764 5046 12776
rect 7006 12764 7012 12776
rect 5040 12736 5133 12764
rect 6919 12736 7012 12764
rect 5040 12724 5046 12736
rect 7006 12724 7012 12736
rect 7064 12764 7070 12776
rect 10428 12764 10456 12795
rect 11606 12792 11612 12804
rect 11664 12792 11670 12844
rect 11716 12841 11744 12872
rect 12434 12860 12440 12872
rect 12492 12900 12498 12912
rect 13078 12900 13084 12912
rect 12492 12872 13084 12900
rect 12492 12860 12498 12872
rect 13078 12860 13084 12872
rect 13136 12860 13142 12912
rect 14090 12860 14096 12912
rect 14148 12900 14154 12912
rect 14936 12900 14964 12931
rect 15286 12900 15292 12912
rect 14148 12872 15292 12900
rect 14148 12860 14154 12872
rect 15286 12860 15292 12872
rect 15344 12860 15350 12912
rect 11701 12835 11759 12841
rect 11701 12801 11713 12835
rect 11747 12801 11759 12835
rect 11701 12795 11759 12801
rect 11885 12835 11943 12841
rect 11885 12801 11897 12835
rect 11931 12832 11943 12835
rect 12158 12832 12164 12844
rect 11931 12804 12164 12832
rect 11931 12801 11943 12804
rect 11885 12795 11943 12801
rect 11900 12764 11928 12795
rect 12158 12792 12164 12804
rect 12216 12792 12222 12844
rect 14918 12835 14976 12841
rect 14918 12801 14930 12835
rect 14964 12832 14976 12835
rect 15654 12832 15660 12844
rect 14964 12804 15660 12832
rect 14964 12801 14976 12804
rect 14918 12795 14976 12801
rect 15654 12792 15660 12804
rect 15712 12792 15718 12844
rect 15930 12832 15936 12844
rect 15891 12804 15936 12832
rect 15930 12792 15936 12804
rect 15988 12792 15994 12844
rect 16114 12832 16120 12844
rect 16075 12804 16120 12832
rect 16114 12792 16120 12804
rect 16172 12792 16178 12844
rect 16942 12792 16948 12844
rect 17000 12832 17006 12844
rect 17405 12835 17463 12841
rect 17405 12832 17417 12835
rect 17000 12804 17417 12832
rect 17000 12792 17006 12804
rect 17405 12801 17417 12804
rect 17451 12801 17463 12835
rect 17405 12795 17463 12801
rect 7064 12736 10456 12764
rect 10980 12736 11928 12764
rect 7064 12724 7070 12736
rect 2317 12699 2375 12705
rect 2317 12665 2329 12699
rect 2363 12696 2375 12699
rect 2590 12696 2596 12708
rect 2363 12668 2596 12696
rect 2363 12665 2375 12668
rect 2317 12659 2375 12665
rect 2590 12656 2596 12668
rect 2648 12696 2654 12708
rect 3605 12699 3663 12705
rect 3605 12696 3617 12699
rect 2648 12668 3617 12696
rect 2648 12656 2654 12668
rect 3605 12665 3617 12668
rect 3651 12665 3663 12699
rect 3605 12659 3663 12665
rect 4614 12588 4620 12640
rect 4672 12628 4678 12640
rect 5000 12628 5028 12724
rect 8202 12656 8208 12708
rect 8260 12696 8266 12708
rect 10980 12696 11008 12736
rect 12250 12724 12256 12776
rect 12308 12764 12314 12776
rect 15289 12767 15347 12773
rect 15289 12764 15301 12767
rect 12308 12736 15301 12764
rect 12308 12724 12314 12736
rect 15289 12733 15301 12736
rect 15335 12733 15347 12767
rect 15289 12727 15347 12733
rect 12802 12696 12808 12708
rect 8260 12668 11008 12696
rect 11072 12668 12808 12696
rect 8260 12656 8266 12668
rect 11072 12640 11100 12668
rect 12802 12656 12808 12668
rect 12860 12656 12866 12708
rect 15304 12696 15332 12727
rect 15378 12724 15384 12776
rect 15436 12764 15442 12776
rect 16022 12764 16028 12776
rect 15436 12736 16028 12764
rect 15436 12724 15442 12736
rect 16022 12724 16028 12736
rect 16080 12724 16086 12776
rect 16574 12724 16580 12776
rect 16632 12764 16638 12776
rect 17218 12764 17224 12776
rect 16632 12736 17224 12764
rect 16632 12724 16638 12736
rect 17218 12724 17224 12736
rect 17276 12764 17282 12776
rect 17313 12767 17371 12773
rect 17313 12764 17325 12767
rect 17276 12736 17325 12764
rect 17276 12724 17282 12736
rect 17313 12733 17325 12736
rect 17359 12733 17371 12767
rect 17313 12727 17371 12733
rect 17037 12699 17095 12705
rect 17037 12696 17049 12699
rect 15304 12668 17049 12696
rect 17037 12665 17049 12668
rect 17083 12665 17095 12699
rect 17037 12659 17095 12665
rect 7374 12628 7380 12640
rect 4672 12600 5028 12628
rect 7335 12600 7380 12628
rect 4672 12588 4678 12600
rect 7374 12588 7380 12600
rect 7432 12588 7438 12640
rect 10413 12631 10471 12637
rect 10413 12597 10425 12631
rect 10459 12628 10471 12631
rect 10502 12628 10508 12640
rect 10459 12600 10508 12628
rect 10459 12597 10471 12600
rect 10413 12591 10471 12597
rect 10502 12588 10508 12600
rect 10560 12628 10566 12640
rect 10778 12628 10784 12640
rect 10560 12600 10784 12628
rect 10560 12588 10566 12600
rect 10778 12588 10784 12600
rect 10836 12588 10842 12640
rect 11054 12628 11060 12640
rect 11015 12600 11060 12628
rect 11054 12588 11060 12600
rect 11112 12588 11118 12640
rect 11146 12588 11152 12640
rect 11204 12628 11210 12640
rect 11701 12631 11759 12637
rect 11701 12628 11713 12631
rect 11204 12600 11713 12628
rect 11204 12588 11210 12600
rect 11701 12597 11713 12600
rect 11747 12597 11759 12631
rect 11701 12591 11759 12597
rect 15746 12588 15752 12640
rect 15804 12628 15810 12640
rect 16025 12631 16083 12637
rect 16025 12628 16037 12631
rect 15804 12600 16037 12628
rect 15804 12588 15810 12600
rect 16025 12597 16037 12600
rect 16071 12597 16083 12631
rect 16025 12591 16083 12597
rect 1104 12538 18860 12560
rect 1104 12486 3169 12538
rect 3221 12486 3233 12538
rect 3285 12486 3297 12538
rect 3349 12486 3361 12538
rect 3413 12486 3425 12538
rect 3477 12486 7608 12538
rect 7660 12486 7672 12538
rect 7724 12486 7736 12538
rect 7788 12486 7800 12538
rect 7852 12486 7864 12538
rect 7916 12486 12047 12538
rect 12099 12486 12111 12538
rect 12163 12486 12175 12538
rect 12227 12486 12239 12538
rect 12291 12486 12303 12538
rect 12355 12486 16486 12538
rect 16538 12486 16550 12538
rect 16602 12486 16614 12538
rect 16666 12486 16678 12538
rect 16730 12486 16742 12538
rect 16794 12486 18860 12538
rect 1104 12464 18860 12486
rect 2225 12427 2283 12433
rect 2225 12393 2237 12427
rect 2271 12424 2283 12427
rect 2498 12424 2504 12436
rect 2271 12396 2504 12424
rect 2271 12393 2283 12396
rect 2225 12387 2283 12393
rect 2498 12384 2504 12396
rect 2556 12384 2562 12436
rect 4246 12424 4252 12436
rect 4207 12396 4252 12424
rect 4246 12384 4252 12396
rect 4304 12384 4310 12436
rect 5994 12384 6000 12436
rect 6052 12424 6058 12436
rect 6181 12427 6239 12433
rect 6181 12424 6193 12427
rect 6052 12396 6193 12424
rect 6052 12384 6058 12396
rect 6181 12393 6193 12396
rect 6227 12393 6239 12427
rect 6181 12387 6239 12393
rect 8573 12427 8631 12433
rect 8573 12393 8585 12427
rect 8619 12424 8631 12427
rect 9030 12424 9036 12436
rect 8619 12396 9036 12424
rect 8619 12393 8631 12396
rect 8573 12387 8631 12393
rect 9030 12384 9036 12396
rect 9088 12384 9094 12436
rect 9401 12427 9459 12433
rect 9401 12393 9413 12427
rect 9447 12393 9459 12427
rect 9401 12387 9459 12393
rect 7009 12359 7067 12365
rect 7009 12356 7021 12359
rect 6380 12328 7021 12356
rect 6380 12232 6408 12328
rect 7009 12325 7021 12328
rect 7055 12325 7067 12359
rect 7009 12319 7067 12325
rect 8202 12316 8208 12368
rect 8260 12356 8266 12368
rect 9416 12356 9444 12387
rect 9490 12384 9496 12436
rect 9548 12424 9554 12436
rect 9585 12427 9643 12433
rect 9585 12424 9597 12427
rect 9548 12396 9597 12424
rect 9548 12384 9554 12396
rect 9585 12393 9597 12396
rect 9631 12393 9643 12427
rect 9585 12387 9643 12393
rect 10042 12384 10048 12436
rect 10100 12424 10106 12436
rect 10686 12424 10692 12436
rect 10100 12396 10692 12424
rect 10100 12384 10106 12396
rect 10686 12384 10692 12396
rect 10744 12424 10750 12436
rect 11054 12424 11060 12436
rect 10744 12396 11060 12424
rect 10744 12384 10750 12396
rect 11054 12384 11060 12396
rect 11112 12384 11118 12436
rect 11514 12424 11520 12436
rect 11475 12396 11520 12424
rect 11514 12384 11520 12396
rect 11572 12384 11578 12436
rect 16114 12424 16120 12436
rect 13004 12396 16120 12424
rect 11532 12356 11560 12384
rect 8260 12328 11560 12356
rect 8260 12316 8266 12328
rect 6822 12248 6828 12300
rect 6880 12288 6886 12300
rect 9306 12288 9312 12300
rect 6880 12260 9312 12288
rect 6880 12248 6886 12260
rect 9306 12248 9312 12260
rect 9364 12248 9370 12300
rect 10870 12288 10876 12300
rect 10520 12260 10876 12288
rect 1765 12223 1823 12229
rect 1765 12189 1777 12223
rect 1811 12220 1823 12223
rect 2222 12220 2228 12232
rect 1811 12192 2228 12220
rect 1811 12189 1823 12192
rect 1765 12183 1823 12189
rect 2222 12180 2228 12192
rect 2280 12180 2286 12232
rect 2406 12220 2412 12232
rect 2367 12192 2412 12220
rect 2406 12180 2412 12192
rect 2464 12180 2470 12232
rect 2501 12223 2559 12229
rect 2501 12189 2513 12223
rect 2547 12220 2559 12223
rect 2590 12220 2596 12232
rect 2547 12192 2596 12220
rect 2547 12189 2559 12192
rect 2501 12183 2559 12189
rect 2590 12180 2596 12192
rect 2648 12180 2654 12232
rect 2866 12180 2872 12232
rect 2924 12220 2930 12232
rect 2961 12223 3019 12229
rect 2961 12220 2973 12223
rect 2924 12192 2973 12220
rect 2924 12180 2930 12192
rect 2961 12189 2973 12192
rect 3007 12189 3019 12223
rect 2961 12183 3019 12189
rect 3970 12180 3976 12232
rect 4028 12220 4034 12232
rect 4065 12223 4123 12229
rect 4065 12220 4077 12223
rect 4028 12192 4077 12220
rect 4028 12180 4034 12192
rect 4065 12189 4077 12192
rect 4111 12189 4123 12223
rect 6362 12220 6368 12232
rect 6323 12192 6368 12220
rect 4065 12183 4123 12189
rect 6362 12180 6368 12192
rect 6420 12180 6426 12232
rect 6549 12223 6607 12229
rect 6549 12189 6561 12223
rect 6595 12220 6607 12223
rect 7190 12220 7196 12232
rect 6595 12192 7196 12220
rect 6595 12189 6607 12192
rect 6549 12183 6607 12189
rect 7190 12180 7196 12192
rect 7248 12180 7254 12232
rect 7285 12223 7343 12229
rect 7285 12189 7297 12223
rect 7331 12220 7343 12223
rect 7374 12220 7380 12232
rect 7331 12192 7380 12220
rect 7331 12189 7343 12192
rect 7285 12183 7343 12189
rect 7374 12180 7380 12192
rect 7432 12220 7438 12232
rect 7926 12220 7932 12232
rect 7432 12192 7932 12220
rect 7432 12180 7438 12192
rect 7926 12180 7932 12192
rect 7984 12180 7990 12232
rect 8110 12180 8116 12232
rect 8168 12220 8174 12232
rect 8297 12223 8355 12229
rect 8297 12220 8309 12223
rect 8168 12192 8309 12220
rect 8168 12180 8174 12192
rect 8297 12189 8309 12192
rect 8343 12189 8355 12223
rect 8297 12183 8355 12189
rect 8386 12180 8392 12232
rect 8444 12220 8450 12232
rect 9214 12220 9220 12232
rect 8444 12192 8489 12220
rect 9175 12192 9220 12220
rect 8444 12180 8450 12192
rect 9214 12180 9220 12192
rect 9272 12180 9278 12232
rect 10045 12223 10103 12229
rect 10045 12189 10057 12223
rect 10091 12220 10103 12223
rect 10318 12220 10324 12232
rect 10091 12192 10324 12220
rect 10091 12189 10103 12192
rect 10045 12183 10103 12189
rect 10318 12180 10324 12192
rect 10376 12180 10382 12232
rect 10520 12164 10548 12260
rect 10870 12248 10876 12260
rect 10928 12248 10934 12300
rect 10962 12248 10968 12300
rect 11020 12288 11026 12300
rect 11238 12288 11244 12300
rect 11020 12260 11244 12288
rect 11020 12248 11026 12260
rect 11238 12248 11244 12260
rect 11296 12288 11302 12300
rect 11296 12260 11836 12288
rect 11296 12248 11302 12260
rect 10689 12223 10747 12229
rect 10689 12189 10701 12223
rect 10735 12220 10747 12223
rect 11146 12220 11152 12232
rect 10735 12192 11152 12220
rect 10735 12189 10747 12192
rect 10689 12183 10747 12189
rect 11146 12180 11152 12192
rect 11204 12180 11210 12232
rect 11609 12223 11667 12229
rect 11609 12189 11621 12223
rect 11655 12220 11667 12223
rect 11698 12220 11704 12232
rect 11655 12192 11704 12220
rect 11655 12189 11667 12192
rect 11609 12183 11667 12189
rect 11698 12180 11704 12192
rect 11756 12180 11762 12232
rect 11808 12220 11836 12260
rect 11885 12223 11943 12229
rect 11885 12220 11897 12223
rect 11808 12192 11897 12220
rect 11885 12189 11897 12192
rect 11931 12189 11943 12223
rect 12713 12223 12771 12229
rect 12713 12220 12725 12223
rect 11885 12183 11943 12189
rect 12406 12192 12725 12220
rect 7006 12152 7012 12164
rect 6967 12124 7012 12152
rect 7006 12112 7012 12124
rect 7064 12112 7070 12164
rect 10502 12152 10508 12164
rect 8220 12124 10508 12152
rect 3050 12044 3056 12096
rect 3108 12084 3114 12096
rect 3145 12087 3203 12093
rect 3145 12084 3157 12087
rect 3108 12056 3157 12084
rect 3108 12044 3114 12056
rect 3145 12053 3157 12056
rect 3191 12053 3203 12087
rect 3145 12047 3203 12053
rect 7098 12044 7104 12096
rect 7156 12084 7162 12096
rect 7193 12087 7251 12093
rect 7193 12084 7205 12087
rect 7156 12056 7205 12084
rect 7156 12044 7162 12056
rect 7193 12053 7205 12056
rect 7239 12084 7251 12087
rect 7282 12084 7288 12096
rect 7239 12056 7288 12084
rect 7239 12053 7251 12056
rect 7193 12047 7251 12053
rect 7282 12044 7288 12056
rect 7340 12084 7346 12096
rect 8018 12084 8024 12096
rect 7340 12056 8024 12084
rect 7340 12044 7346 12056
rect 8018 12044 8024 12056
rect 8076 12044 8082 12096
rect 8220 12093 8248 12124
rect 10502 12112 10508 12124
rect 10560 12112 10566 12164
rect 10781 12155 10839 12161
rect 10781 12121 10793 12155
rect 10827 12152 10839 12155
rect 11716 12152 11744 12180
rect 12406 12152 12434 12192
rect 12713 12189 12725 12192
rect 12759 12189 12771 12223
rect 12713 12183 12771 12189
rect 12802 12180 12808 12232
rect 12860 12220 12866 12232
rect 13004 12229 13032 12396
rect 16114 12384 16120 12396
rect 16172 12424 16178 12436
rect 16485 12427 16543 12433
rect 16485 12424 16497 12427
rect 16172 12396 16497 12424
rect 16172 12384 16178 12396
rect 16485 12393 16497 12396
rect 16531 12393 16543 12427
rect 17770 12424 17776 12436
rect 17731 12396 17776 12424
rect 16485 12387 16543 12393
rect 17770 12384 17776 12396
rect 17828 12384 17834 12436
rect 12989 12223 13047 12229
rect 12989 12220 13001 12223
rect 12860 12192 13001 12220
rect 12860 12180 12866 12192
rect 12989 12189 13001 12192
rect 13035 12189 13047 12223
rect 12989 12183 13047 12189
rect 13998 12180 14004 12232
rect 14056 12220 14062 12232
rect 14277 12223 14335 12229
rect 14277 12220 14289 12223
rect 14056 12192 14289 12220
rect 14056 12180 14062 12192
rect 14277 12189 14289 12192
rect 14323 12189 14335 12223
rect 16666 12220 16672 12232
rect 16627 12192 16672 12220
rect 14277 12183 14335 12189
rect 16666 12180 16672 12192
rect 16724 12180 16730 12232
rect 17037 12223 17095 12229
rect 17037 12189 17049 12223
rect 17083 12189 17095 12223
rect 17037 12183 17095 12189
rect 10827 12124 11376 12152
rect 11716 12124 12434 12152
rect 14544 12155 14602 12161
rect 10827 12121 10839 12124
rect 10781 12115 10839 12121
rect 8205 12087 8263 12093
rect 8205 12053 8217 12087
rect 8251 12053 8263 12087
rect 8205 12047 8263 12053
rect 8386 12044 8392 12096
rect 8444 12084 8450 12096
rect 10042 12084 10048 12096
rect 8444 12056 10048 12084
rect 8444 12044 8450 12056
rect 10042 12044 10048 12056
rect 10100 12044 10106 12096
rect 10226 12084 10232 12096
rect 10187 12056 10232 12084
rect 10226 12044 10232 12056
rect 10284 12044 10290 12096
rect 10410 12044 10416 12096
rect 10468 12084 10474 12096
rect 11348 12093 11376 12124
rect 14544 12121 14556 12155
rect 14590 12152 14602 12155
rect 14642 12152 14648 12164
rect 14590 12124 14648 12152
rect 14590 12121 14602 12124
rect 14544 12115 14602 12121
rect 14642 12112 14648 12124
rect 14700 12112 14706 12164
rect 15930 12152 15936 12164
rect 14752 12124 15936 12152
rect 10597 12087 10655 12093
rect 10597 12084 10609 12087
rect 10468 12056 10609 12084
rect 10468 12044 10474 12056
rect 10597 12053 10609 12056
rect 10643 12053 10655 12087
rect 10597 12047 10655 12053
rect 11333 12087 11391 12093
rect 11333 12053 11345 12087
rect 11379 12053 11391 12087
rect 12526 12084 12532 12096
rect 12487 12056 12532 12084
rect 11333 12047 11391 12053
rect 12526 12044 12532 12056
rect 12584 12044 12590 12096
rect 12618 12044 12624 12096
rect 12676 12084 12682 12096
rect 12897 12087 12955 12093
rect 12897 12084 12909 12087
rect 12676 12056 12909 12084
rect 12676 12044 12682 12056
rect 12897 12053 12909 12056
rect 12943 12084 12955 12087
rect 14752 12084 14780 12124
rect 15930 12112 15936 12124
rect 15988 12112 15994 12164
rect 16761 12155 16819 12161
rect 16761 12121 16773 12155
rect 16807 12121 16819 12155
rect 16761 12115 16819 12121
rect 12943 12056 14780 12084
rect 15657 12087 15715 12093
rect 12943 12053 12955 12056
rect 12897 12047 12955 12053
rect 15657 12053 15669 12087
rect 15703 12084 15715 12087
rect 16666 12084 16672 12096
rect 15703 12056 16672 12084
rect 15703 12053 15715 12056
rect 15657 12047 15715 12053
rect 16666 12044 16672 12056
rect 16724 12044 16730 12096
rect 16776 12084 16804 12115
rect 16850 12112 16856 12164
rect 16908 12152 16914 12164
rect 17052 12152 17080 12183
rect 17126 12180 17132 12232
rect 17184 12220 17190 12232
rect 17497 12223 17555 12229
rect 17497 12220 17509 12223
rect 17184 12192 17509 12220
rect 17184 12180 17190 12192
rect 17497 12189 17509 12192
rect 17543 12189 17555 12223
rect 17497 12183 17555 12189
rect 17218 12152 17224 12164
rect 16908 12124 16953 12152
rect 17052 12124 17224 12152
rect 16908 12112 16914 12124
rect 17218 12112 17224 12124
rect 17276 12112 17282 12164
rect 17034 12084 17040 12096
rect 16776 12056 17040 12084
rect 17034 12044 17040 12056
rect 17092 12044 17098 12096
rect 17954 12084 17960 12096
rect 17915 12056 17960 12084
rect 17954 12044 17960 12056
rect 18012 12044 18018 12096
rect 1104 11994 19019 12016
rect 1104 11942 5388 11994
rect 5440 11942 5452 11994
rect 5504 11942 5516 11994
rect 5568 11942 5580 11994
rect 5632 11942 5644 11994
rect 5696 11942 9827 11994
rect 9879 11942 9891 11994
rect 9943 11942 9955 11994
rect 10007 11942 10019 11994
rect 10071 11942 10083 11994
rect 10135 11942 14266 11994
rect 14318 11942 14330 11994
rect 14382 11942 14394 11994
rect 14446 11942 14458 11994
rect 14510 11942 14522 11994
rect 14574 11942 18705 11994
rect 18757 11942 18769 11994
rect 18821 11942 18833 11994
rect 18885 11942 18897 11994
rect 18949 11942 18961 11994
rect 19013 11942 19019 11994
rect 1104 11920 19019 11942
rect 6733 11883 6791 11889
rect 6733 11849 6745 11883
rect 6779 11880 6791 11883
rect 7926 11880 7932 11892
rect 6779 11852 7932 11880
rect 6779 11849 6791 11852
rect 6733 11843 6791 11849
rect 7926 11840 7932 11852
rect 7984 11880 7990 11892
rect 8389 11883 8447 11889
rect 8389 11880 8401 11883
rect 7984 11852 8401 11880
rect 7984 11840 7990 11852
rect 8389 11849 8401 11852
rect 8435 11849 8447 11883
rect 8389 11843 8447 11849
rect 8573 11883 8631 11889
rect 8573 11849 8585 11883
rect 8619 11880 8631 11883
rect 8754 11880 8760 11892
rect 8619 11852 8760 11880
rect 8619 11849 8631 11852
rect 8573 11843 8631 11849
rect 8754 11840 8760 11852
rect 8812 11840 8818 11892
rect 9214 11840 9220 11892
rect 9272 11880 9278 11892
rect 9401 11883 9459 11889
rect 9401 11880 9413 11883
rect 9272 11852 9413 11880
rect 9272 11840 9278 11852
rect 9401 11849 9413 11852
rect 9447 11849 9459 11883
rect 10410 11880 10416 11892
rect 10371 11852 10416 11880
rect 9401 11843 9459 11849
rect 10410 11840 10416 11852
rect 10468 11840 10474 11892
rect 12526 11840 12532 11892
rect 12584 11840 12590 11892
rect 14553 11883 14611 11889
rect 14553 11849 14565 11883
rect 14599 11880 14611 11883
rect 14642 11880 14648 11892
rect 14599 11852 14648 11880
rect 14599 11849 14611 11852
rect 14553 11843 14611 11849
rect 14642 11840 14648 11852
rect 14700 11840 14706 11892
rect 15286 11840 15292 11892
rect 15344 11880 15350 11892
rect 15381 11883 15439 11889
rect 15381 11880 15393 11883
rect 15344 11852 15393 11880
rect 15344 11840 15350 11852
rect 15381 11849 15393 11852
rect 15427 11849 15439 11883
rect 15381 11843 15439 11849
rect 15930 11840 15936 11892
rect 15988 11880 15994 11892
rect 17497 11883 17555 11889
rect 17497 11880 17509 11883
rect 15988 11852 17509 11880
rect 15988 11840 15994 11852
rect 17497 11849 17509 11852
rect 17543 11849 17555 11883
rect 17497 11843 17555 11849
rect 4614 11812 4620 11824
rect 2792 11784 4620 11812
rect 2792 11753 2820 11784
rect 4614 11772 4620 11784
rect 4672 11772 4678 11824
rect 6825 11815 6883 11821
rect 4816 11784 6776 11812
rect 3050 11753 3056 11756
rect 2777 11747 2835 11753
rect 2777 11713 2789 11747
rect 2823 11713 2835 11747
rect 3044 11744 3056 11753
rect 3011 11716 3056 11744
rect 2777 11707 2835 11713
rect 3044 11707 3056 11716
rect 3050 11704 3056 11707
rect 3108 11704 3114 11756
rect 3786 11704 3792 11756
rect 3844 11744 3850 11756
rect 4816 11744 4844 11784
rect 3844 11716 4844 11744
rect 4884 11747 4942 11753
rect 3844 11704 3850 11716
rect 4884 11713 4896 11747
rect 4930 11744 4942 11747
rect 6086 11744 6092 11756
rect 4930 11716 6092 11744
rect 4930 11713 4942 11716
rect 4884 11707 4942 11713
rect 6086 11704 6092 11716
rect 6144 11704 6150 11756
rect 6748 11744 6776 11784
rect 6825 11781 6837 11815
rect 6871 11812 6883 11815
rect 7098 11812 7104 11824
rect 6871 11784 7104 11812
rect 6871 11781 6883 11784
rect 6825 11775 6883 11781
rect 7098 11772 7104 11784
rect 7156 11772 7162 11824
rect 7282 11772 7288 11824
rect 7340 11812 7346 11824
rect 8297 11815 8355 11821
rect 8297 11812 8309 11815
rect 7340 11784 8309 11812
rect 7340 11772 7346 11784
rect 8297 11781 8309 11784
rect 8343 11781 8355 11815
rect 11054 11812 11060 11824
rect 8297 11775 8355 11781
rect 10336 11784 11060 11812
rect 6917 11747 6975 11753
rect 6917 11744 6929 11747
rect 6748 11716 6929 11744
rect 6917 11713 6929 11716
rect 6963 11744 6975 11747
rect 7006 11744 7012 11756
rect 6963 11716 7012 11744
rect 6963 11713 6975 11716
rect 6917 11707 6975 11713
rect 7006 11704 7012 11716
rect 7064 11704 7070 11756
rect 8202 11744 8208 11756
rect 8163 11716 8208 11744
rect 8202 11704 8208 11716
rect 8260 11704 8266 11756
rect 8570 11704 8576 11756
rect 8628 11744 8634 11756
rect 9033 11747 9091 11753
rect 9033 11744 9045 11747
rect 8628 11716 9045 11744
rect 8628 11704 8634 11716
rect 9033 11713 9045 11716
rect 9079 11713 9091 11747
rect 9214 11744 9220 11756
rect 9175 11716 9220 11744
rect 9033 11707 9091 11713
rect 9214 11704 9220 11716
rect 9272 11704 9278 11756
rect 9306 11704 9312 11756
rect 9364 11744 9370 11756
rect 10336 11753 10364 11784
rect 11054 11772 11060 11784
rect 11112 11772 11118 11824
rect 12544 11812 12572 11840
rect 12544 11784 13308 11812
rect 10321 11747 10379 11753
rect 10321 11744 10333 11747
rect 9364 11716 10333 11744
rect 9364 11704 9370 11716
rect 10321 11713 10333 11716
rect 10367 11713 10379 11747
rect 10502 11744 10508 11756
rect 10463 11716 10508 11744
rect 10321 11707 10379 11713
rect 10502 11704 10508 11716
rect 10560 11704 10566 11756
rect 10965 11747 11023 11753
rect 10965 11713 10977 11747
rect 11011 11713 11023 11747
rect 10965 11707 11023 11713
rect 11149 11747 11207 11753
rect 11149 11713 11161 11747
rect 11195 11713 11207 11747
rect 11149 11707 11207 11713
rect 4614 11676 4620 11688
rect 4575 11648 4620 11676
rect 4614 11636 4620 11648
rect 4672 11636 4678 11688
rect 7101 11679 7159 11685
rect 7101 11676 7113 11679
rect 6012 11648 7113 11676
rect 6012 11617 6040 11648
rect 7101 11645 7113 11648
rect 7147 11676 7159 11679
rect 8021 11679 8079 11685
rect 8021 11676 8033 11679
rect 7147 11648 8033 11676
rect 7147 11645 7159 11648
rect 7101 11639 7159 11645
rect 8021 11645 8033 11648
rect 8067 11676 8079 11679
rect 8110 11676 8116 11688
rect 8067 11648 8116 11676
rect 8067 11645 8079 11648
rect 8021 11639 8079 11645
rect 8110 11636 8116 11648
rect 8168 11676 8174 11688
rect 10980 11676 11008 11707
rect 8168 11648 11008 11676
rect 8168 11636 8174 11648
rect 5997 11611 6055 11617
rect 5997 11577 6009 11611
rect 6043 11577 6055 11611
rect 5997 11571 6055 11577
rect 9398 11568 9404 11620
rect 9456 11608 9462 11620
rect 11164 11608 11192 11707
rect 11606 11704 11612 11756
rect 11664 11744 11670 11756
rect 11885 11747 11943 11753
rect 11885 11744 11897 11747
rect 11664 11716 11897 11744
rect 11664 11704 11670 11716
rect 11885 11713 11897 11716
rect 11931 11744 11943 11747
rect 12529 11747 12587 11753
rect 12529 11744 12541 11747
rect 11931 11716 12541 11744
rect 11931 11713 11943 11716
rect 11885 11707 11943 11713
rect 12529 11713 12541 11716
rect 12575 11713 12587 11747
rect 12529 11707 12587 11713
rect 12618 11704 12624 11756
rect 12676 11744 12682 11756
rect 12802 11744 12808 11756
rect 12676 11716 12721 11744
rect 12763 11716 12808 11744
rect 12676 11704 12682 11716
rect 12802 11704 12808 11716
rect 12860 11704 12866 11756
rect 13280 11753 13308 11784
rect 13372 11784 15332 11812
rect 13265 11747 13323 11753
rect 13265 11713 13277 11747
rect 13311 11713 13323 11747
rect 13265 11707 13323 11713
rect 12069 11679 12127 11685
rect 12069 11676 12081 11679
rect 11900 11648 12081 11676
rect 11900 11620 11928 11648
rect 12069 11645 12081 11648
rect 12115 11645 12127 11679
rect 13372 11676 13400 11784
rect 13449 11747 13507 11753
rect 13449 11713 13461 11747
rect 13495 11713 13507 11747
rect 13449 11707 13507 11713
rect 14461 11747 14519 11753
rect 14461 11713 14473 11747
rect 14507 11713 14519 11747
rect 14461 11707 14519 11713
rect 14645 11747 14703 11753
rect 14645 11713 14657 11747
rect 14691 11744 14703 11747
rect 14691 11716 15240 11744
rect 14691 11713 14703 11716
rect 14645 11707 14703 11713
rect 12069 11639 12127 11645
rect 12176 11648 13400 11676
rect 9456 11580 11836 11608
rect 9456 11568 9462 11580
rect 4154 11540 4160 11552
rect 4115 11512 4160 11540
rect 4154 11500 4160 11512
rect 4212 11500 4218 11552
rect 6178 11500 6184 11552
rect 6236 11540 6242 11552
rect 6549 11543 6607 11549
rect 6549 11540 6561 11543
rect 6236 11512 6561 11540
rect 6236 11500 6242 11512
rect 6549 11509 6561 11512
rect 6595 11509 6607 11543
rect 6549 11503 6607 11509
rect 7006 11500 7012 11552
rect 7064 11540 7070 11552
rect 8570 11540 8576 11552
rect 7064 11512 8576 11540
rect 7064 11500 7070 11512
rect 8570 11500 8576 11512
rect 8628 11500 8634 11552
rect 8938 11500 8944 11552
rect 8996 11540 9002 11552
rect 9033 11543 9091 11549
rect 9033 11540 9045 11543
rect 8996 11512 9045 11540
rect 8996 11500 9002 11512
rect 9033 11509 9045 11512
rect 9079 11509 9091 11543
rect 11698 11540 11704 11552
rect 11659 11512 11704 11540
rect 9033 11503 9091 11509
rect 11698 11500 11704 11512
rect 11756 11500 11762 11552
rect 11808 11540 11836 11580
rect 11882 11568 11888 11620
rect 11940 11568 11946 11620
rect 12176 11540 12204 11648
rect 12434 11568 12440 11620
rect 12492 11608 12498 11620
rect 12713 11611 12771 11617
rect 12713 11608 12725 11611
rect 12492 11580 12725 11608
rect 12492 11568 12498 11580
rect 12713 11577 12725 11580
rect 12759 11608 12771 11611
rect 13464 11608 13492 11707
rect 12759 11580 13492 11608
rect 12759 11577 12771 11580
rect 12713 11571 12771 11577
rect 13354 11540 13360 11552
rect 11808 11512 12204 11540
rect 13315 11512 13360 11540
rect 13354 11500 13360 11512
rect 13412 11500 13418 11552
rect 14001 11543 14059 11549
rect 14001 11509 14013 11543
rect 14047 11540 14059 11543
rect 14182 11540 14188 11552
rect 14047 11512 14188 11540
rect 14047 11509 14059 11512
rect 14001 11503 14059 11509
rect 14182 11500 14188 11512
rect 14240 11540 14246 11552
rect 14476 11540 14504 11707
rect 15212 11617 15240 11716
rect 15197 11611 15255 11617
rect 15197 11577 15209 11611
rect 15243 11577 15255 11611
rect 15197 11571 15255 11577
rect 14826 11540 14832 11552
rect 14240 11512 14832 11540
rect 14240 11500 14246 11512
rect 14826 11500 14832 11512
rect 14884 11500 14890 11552
rect 15304 11540 15332 11784
rect 15580 11784 16436 11812
rect 15378 11747 15436 11753
rect 15378 11713 15390 11747
rect 15424 11744 15436 11747
rect 15580 11744 15608 11784
rect 16408 11756 16436 11784
rect 15746 11744 15752 11756
rect 15424 11716 15608 11744
rect 15707 11716 15752 11744
rect 15424 11713 15436 11716
rect 15378 11707 15436 11713
rect 15746 11704 15752 11716
rect 15804 11704 15810 11756
rect 16390 11704 16396 11756
rect 16448 11744 16454 11756
rect 16666 11744 16672 11756
rect 16448 11716 16672 11744
rect 16448 11704 16454 11716
rect 16666 11704 16672 11716
rect 16724 11744 16730 11756
rect 16853 11747 16911 11753
rect 16853 11744 16865 11747
rect 16724 11716 16865 11744
rect 16724 11704 16730 11716
rect 16853 11713 16865 11716
rect 16899 11713 16911 11747
rect 16853 11707 16911 11713
rect 16945 11747 17003 11753
rect 16945 11713 16957 11747
rect 16991 11744 17003 11747
rect 17586 11744 17592 11756
rect 16991 11716 17592 11744
rect 16991 11713 17003 11716
rect 16945 11707 17003 11713
rect 17586 11704 17592 11716
rect 17644 11744 17650 11756
rect 17681 11747 17739 11753
rect 17681 11744 17693 11747
rect 17644 11716 17693 11744
rect 17644 11704 17650 11716
rect 17681 11713 17693 11716
rect 17727 11713 17739 11747
rect 17681 11707 17739 11713
rect 17865 11747 17923 11753
rect 17865 11713 17877 11747
rect 17911 11744 17923 11747
rect 17954 11744 17960 11756
rect 17911 11716 17960 11744
rect 17911 11713 17923 11716
rect 17865 11707 17923 11713
rect 17954 11704 17960 11716
rect 18012 11704 18018 11756
rect 15841 11679 15899 11685
rect 15841 11676 15853 11679
rect 15764 11648 15853 11676
rect 15764 11620 15792 11648
rect 15841 11645 15853 11648
rect 15887 11676 15899 11679
rect 16022 11676 16028 11688
rect 15887 11648 16028 11676
rect 15887 11645 15899 11648
rect 15841 11639 15899 11645
rect 16022 11636 16028 11648
rect 16080 11636 16086 11688
rect 15746 11568 15752 11620
rect 15804 11568 15810 11620
rect 16206 11540 16212 11552
rect 15304 11512 16212 11540
rect 16206 11500 16212 11512
rect 16264 11540 16270 11552
rect 17494 11540 17500 11552
rect 16264 11512 17500 11540
rect 16264 11500 16270 11512
rect 17494 11500 17500 11512
rect 17552 11500 17558 11552
rect 17678 11540 17684 11552
rect 17639 11512 17684 11540
rect 17678 11500 17684 11512
rect 17736 11500 17742 11552
rect 1104 11450 18860 11472
rect 1104 11398 3169 11450
rect 3221 11398 3233 11450
rect 3285 11398 3297 11450
rect 3349 11398 3361 11450
rect 3413 11398 3425 11450
rect 3477 11398 7608 11450
rect 7660 11398 7672 11450
rect 7724 11398 7736 11450
rect 7788 11398 7800 11450
rect 7852 11398 7864 11450
rect 7916 11398 12047 11450
rect 12099 11398 12111 11450
rect 12163 11398 12175 11450
rect 12227 11398 12239 11450
rect 12291 11398 12303 11450
rect 12355 11398 16486 11450
rect 16538 11398 16550 11450
rect 16602 11398 16614 11450
rect 16666 11398 16678 11450
rect 16730 11398 16742 11450
rect 16794 11398 18860 11450
rect 1104 11376 18860 11398
rect 2866 11336 2872 11348
rect 2827 11308 2872 11336
rect 2866 11296 2872 11308
rect 2924 11296 2930 11348
rect 3970 11336 3976 11348
rect 3931 11308 3976 11336
rect 3970 11296 3976 11308
rect 4028 11296 4034 11348
rect 6086 11336 6092 11348
rect 6047 11308 6092 11336
rect 6086 11296 6092 11308
rect 6144 11296 6150 11348
rect 7006 11336 7012 11348
rect 6967 11308 7012 11336
rect 7006 11296 7012 11308
rect 7064 11296 7070 11348
rect 7190 11296 7196 11348
rect 7248 11336 7254 11348
rect 7653 11339 7711 11345
rect 7653 11336 7665 11339
rect 7248 11308 7665 11336
rect 7248 11296 7254 11308
rect 7653 11305 7665 11308
rect 7699 11305 7711 11339
rect 7653 11299 7711 11305
rect 10502 11296 10508 11348
rect 10560 11336 10566 11348
rect 10781 11339 10839 11345
rect 10781 11336 10793 11339
rect 10560 11308 10793 11336
rect 10560 11296 10566 11308
rect 10781 11305 10793 11308
rect 10827 11305 10839 11339
rect 10781 11299 10839 11305
rect 13170 11296 13176 11348
rect 13228 11336 13234 11348
rect 13265 11339 13323 11345
rect 13265 11336 13277 11339
rect 13228 11308 13277 11336
rect 13228 11296 13234 11308
rect 13265 11305 13277 11308
rect 13311 11305 13323 11339
rect 13265 11299 13323 11305
rect 16942 11296 16948 11348
rect 17000 11336 17006 11348
rect 17405 11339 17463 11345
rect 17405 11336 17417 11339
rect 17000 11308 17417 11336
rect 17000 11296 17006 11308
rect 17405 11305 17417 11308
rect 17451 11305 17463 11339
rect 17678 11336 17684 11348
rect 17639 11308 17684 11336
rect 17405 11299 17463 11305
rect 17678 11296 17684 11308
rect 17736 11296 17742 11348
rect 6825 11271 6883 11277
rect 6825 11237 6837 11271
rect 6871 11268 6883 11271
rect 8202 11268 8208 11280
rect 6871 11240 7328 11268
rect 6871 11237 6883 11240
rect 6825 11231 6883 11237
rect 2406 11160 2412 11212
rect 2464 11200 2470 11212
rect 2501 11203 2559 11209
rect 2501 11200 2513 11203
rect 2464 11172 2513 11200
rect 2464 11160 2470 11172
rect 2501 11169 2513 11172
rect 2547 11200 2559 11203
rect 4338 11200 4344 11212
rect 2547 11172 4016 11200
rect 4299 11172 4344 11200
rect 2547 11169 2559 11172
rect 2501 11163 2559 11169
rect 2685 11135 2743 11141
rect 2685 11101 2697 11135
rect 2731 11132 2743 11135
rect 3234 11132 3240 11144
rect 2731 11104 3240 11132
rect 2731 11101 2743 11104
rect 2685 11095 2743 11101
rect 3234 11092 3240 11104
rect 3292 11132 3298 11144
rect 3786 11132 3792 11144
rect 3292 11104 3792 11132
rect 3292 11092 3298 11104
rect 3786 11092 3792 11104
rect 3844 11092 3850 11144
rect 3988 11064 4016 11172
rect 4338 11160 4344 11172
rect 4396 11160 4402 11212
rect 7300 11144 7328 11240
rect 7944 11240 8208 11268
rect 7944 11209 7972 11240
rect 8202 11228 8208 11240
rect 8260 11228 8266 11280
rect 11698 11268 11704 11280
rect 9232 11240 11704 11268
rect 7929 11203 7987 11209
rect 7929 11169 7941 11203
rect 7975 11169 7987 11203
rect 7929 11163 7987 11169
rect 8021 11203 8079 11209
rect 8021 11169 8033 11203
rect 8067 11200 8079 11203
rect 8938 11200 8944 11212
rect 8067 11172 8944 11200
rect 8067 11169 8079 11172
rect 8021 11163 8079 11169
rect 8938 11160 8944 11172
rect 8996 11160 9002 11212
rect 4154 11132 4160 11144
rect 4115 11104 4160 11132
rect 4154 11092 4160 11104
rect 4212 11092 4218 11144
rect 6089 11135 6147 11141
rect 6089 11101 6101 11135
rect 6135 11132 6147 11135
rect 6178 11132 6184 11144
rect 6135 11104 6184 11132
rect 6135 11101 6147 11104
rect 6089 11095 6147 11101
rect 6178 11092 6184 11104
rect 6236 11092 6242 11144
rect 6362 11132 6368 11144
rect 6323 11104 6368 11132
rect 6362 11092 6368 11104
rect 6420 11092 6426 11144
rect 7282 11092 7288 11144
rect 7340 11132 7346 11144
rect 7837 11135 7895 11141
rect 7837 11132 7849 11135
rect 7340 11104 7849 11132
rect 7340 11092 7346 11104
rect 7837 11101 7849 11104
rect 7883 11101 7895 11135
rect 7837 11095 7895 11101
rect 8113 11135 8171 11141
rect 8113 11101 8125 11135
rect 8159 11132 8171 11135
rect 9232 11132 9260 11240
rect 11698 11228 11704 11240
rect 11756 11228 11762 11280
rect 12894 11268 12900 11280
rect 12406 11240 12900 11268
rect 10413 11203 10471 11209
rect 10413 11169 10425 11203
rect 10459 11200 10471 11203
rect 11882 11200 11888 11212
rect 10459 11172 11888 11200
rect 10459 11169 10471 11172
rect 10413 11163 10471 11169
rect 11882 11160 11888 11172
rect 11940 11200 11946 11212
rect 12406 11200 12434 11240
rect 12894 11228 12900 11240
rect 12952 11228 12958 11280
rect 17310 11268 17316 11280
rect 16132 11240 17316 11268
rect 11940 11172 12434 11200
rect 12728 11172 12940 11200
rect 11940 11160 11946 11172
rect 12728 11144 12756 11172
rect 8159 11104 9260 11132
rect 9309 11135 9367 11141
rect 8159 11101 8171 11104
rect 8113 11095 8171 11101
rect 9309 11101 9321 11135
rect 9355 11101 9367 11135
rect 9309 11095 9367 11101
rect 6273 11067 6331 11073
rect 3988 11036 4200 11064
rect 4172 11008 4200 11036
rect 6273 11033 6285 11067
rect 6319 11064 6331 11067
rect 6822 11064 6828 11076
rect 6319 11036 6828 11064
rect 6319 11033 6331 11036
rect 6273 11027 6331 11033
rect 6822 11024 6828 11036
rect 6880 11024 6886 11076
rect 6993 11067 7051 11073
rect 6993 11033 7005 11067
rect 7039 11064 7051 11067
rect 7193 11067 7251 11073
rect 7039 11036 7144 11064
rect 7039 11033 7051 11036
rect 6993 11027 7051 11033
rect 4154 10956 4160 11008
rect 4212 10956 4218 11008
rect 5629 10999 5687 11005
rect 5629 10965 5641 10999
rect 5675 10996 5687 10999
rect 5810 10996 5816 11008
rect 5675 10968 5816 10996
rect 5675 10965 5687 10968
rect 5629 10959 5687 10965
rect 5810 10956 5816 10968
rect 5868 10996 5874 11008
rect 6086 10996 6092 11008
rect 5868 10968 6092 10996
rect 5868 10956 5874 10968
rect 6086 10956 6092 10968
rect 6144 10956 6150 11008
rect 7116 10996 7144 11036
rect 7193 11033 7205 11067
rect 7239 11064 7251 11067
rect 8202 11064 8208 11076
rect 7239 11036 8208 11064
rect 7239 11033 7251 11036
rect 7193 11027 7251 11033
rect 8202 11024 8208 11036
rect 8260 11024 8266 11076
rect 8294 11024 8300 11076
rect 8352 11064 8358 11076
rect 9125 11067 9183 11073
rect 9125 11064 9137 11067
rect 8352 11036 9137 11064
rect 8352 11024 8358 11036
rect 9125 11033 9137 11036
rect 9171 11033 9183 11067
rect 9125 11027 9183 11033
rect 9324 11008 9352 11095
rect 9398 11092 9404 11144
rect 9456 11132 9462 11144
rect 10597 11135 10655 11141
rect 9456 11104 9501 11132
rect 9456 11092 9462 11104
rect 10597 11101 10609 11135
rect 10643 11132 10655 11135
rect 10778 11132 10784 11144
rect 10643 11104 10784 11132
rect 10643 11101 10655 11104
rect 10597 11095 10655 11101
rect 10778 11092 10784 11104
rect 10836 11092 10842 11144
rect 12440 11113 12498 11119
rect 12440 11079 12452 11113
rect 12486 11079 12498 11113
rect 12526 11092 12532 11144
rect 12584 11132 12590 11144
rect 12710 11132 12716 11144
rect 12584 11104 12629 11132
rect 12671 11104 12716 11132
rect 12584 11092 12590 11104
rect 12710 11092 12716 11104
rect 12768 11092 12774 11144
rect 12805 11135 12863 11141
rect 12805 11101 12817 11135
rect 12851 11101 12863 11135
rect 12912 11132 12940 11172
rect 12986 11160 12992 11212
rect 13044 11200 13050 11212
rect 13357 11203 13415 11209
rect 13357 11200 13369 11203
rect 13044 11172 13369 11200
rect 13044 11160 13050 11172
rect 13357 11169 13369 11172
rect 13403 11169 13415 11203
rect 14826 11200 14832 11212
rect 13357 11163 13415 11169
rect 14568 11172 14832 11200
rect 14568 11141 14596 11172
rect 14826 11160 14832 11172
rect 14884 11160 14890 11212
rect 16025 11203 16083 11209
rect 16025 11200 16037 11203
rect 15396 11172 16037 11200
rect 13541 11135 13599 11141
rect 13541 11132 13553 11135
rect 12912 11104 13553 11132
rect 12805 11095 12863 11101
rect 13541 11101 13553 11104
rect 13587 11101 13599 11135
rect 13541 11095 13599 11101
rect 14553 11135 14611 11141
rect 14553 11101 14565 11135
rect 14599 11101 14611 11135
rect 14734 11132 14740 11144
rect 14695 11104 14740 11132
rect 14553 11095 14611 11101
rect 12440 11076 12498 11079
rect 10704 11036 10916 11064
rect 8478 10996 8484 11008
rect 7116 10968 8484 10996
rect 8478 10956 8484 10968
rect 8536 10956 8542 11008
rect 9306 10996 9312 11008
rect 9219 10968 9312 10996
rect 9306 10956 9312 10968
rect 9364 10996 9370 11008
rect 10704 10996 10732 11036
rect 9364 10968 10732 10996
rect 10888 10996 10916 11036
rect 11882 11024 11888 11076
rect 11940 11064 11946 11076
rect 12253 11067 12311 11073
rect 12253 11064 12265 11067
rect 11940 11036 12265 11064
rect 11940 11024 11946 11036
rect 12253 11033 12265 11036
rect 12299 11033 12311 11067
rect 12253 11027 12311 11033
rect 12434 11024 12440 11076
rect 12492 11024 12498 11076
rect 12618 11024 12624 11076
rect 12676 11064 12682 11076
rect 12820 11064 12848 11095
rect 14734 11092 14740 11104
rect 14792 11092 14798 11144
rect 15194 11092 15200 11144
rect 15252 11132 15258 11144
rect 15396 11141 15424 11172
rect 16025 11169 16037 11172
rect 16071 11169 16083 11203
rect 16025 11163 16083 11169
rect 15381 11135 15439 11141
rect 15381 11132 15393 11135
rect 15252 11104 15393 11132
rect 15252 11092 15258 11104
rect 15381 11101 15393 11104
rect 15427 11101 15439 11135
rect 15381 11095 15439 11101
rect 15565 11135 15623 11141
rect 15565 11101 15577 11135
rect 15611 11132 15623 11135
rect 16132 11132 16160 11240
rect 17310 11228 17316 11240
rect 17368 11228 17374 11280
rect 16850 11200 16856 11212
rect 16316 11172 16856 11200
rect 16316 11141 16344 11172
rect 16850 11160 16856 11172
rect 16908 11200 16914 11212
rect 17402 11200 17408 11212
rect 16908 11172 17408 11200
rect 16908 11160 16914 11172
rect 17402 11160 17408 11172
rect 17460 11160 17466 11212
rect 17773 11203 17831 11209
rect 17773 11169 17785 11203
rect 17819 11200 17831 11203
rect 17954 11200 17960 11212
rect 17819 11172 17960 11200
rect 17819 11169 17831 11172
rect 17773 11163 17831 11169
rect 17954 11160 17960 11172
rect 18012 11160 18018 11212
rect 15611 11104 16160 11132
rect 16209 11135 16267 11141
rect 15611 11101 15623 11104
rect 15565 11095 15623 11101
rect 16209 11101 16221 11135
rect 16255 11101 16267 11135
rect 16209 11095 16267 11101
rect 16301 11135 16359 11141
rect 16301 11101 16313 11135
rect 16347 11101 16359 11135
rect 16301 11095 16359 11101
rect 13262 11064 13268 11076
rect 12676 11036 12848 11064
rect 13175 11036 13268 11064
rect 12676 11024 12682 11036
rect 13262 11024 13268 11036
rect 13320 11064 13326 11076
rect 16114 11064 16120 11076
rect 13320 11036 16120 11064
rect 13320 11024 13326 11036
rect 16114 11024 16120 11036
rect 16172 11024 16178 11076
rect 16224 11064 16252 11095
rect 16390 11092 16396 11144
rect 16448 11132 16454 11144
rect 16666 11132 16672 11144
rect 16448 11104 16493 11132
rect 16579 11104 16672 11132
rect 16448 11092 16454 11104
rect 16666 11092 16672 11104
rect 16724 11132 16730 11144
rect 17034 11132 17040 11144
rect 16724 11104 17040 11132
rect 16724 11092 16730 11104
rect 17034 11092 17040 11104
rect 17092 11092 17098 11144
rect 17586 11132 17592 11144
rect 17547 11104 17592 11132
rect 17586 11092 17592 11104
rect 17644 11092 17650 11144
rect 16531 11067 16589 11073
rect 16224 11036 16344 11064
rect 12802 10996 12808 11008
rect 10888 10968 12808 10996
rect 9364 10956 9370 10968
rect 12802 10956 12808 10968
rect 12860 10956 12866 11008
rect 13722 10996 13728 11008
rect 13683 10968 13728 10996
rect 13722 10956 13728 10968
rect 13780 10956 13786 11008
rect 14642 10996 14648 11008
rect 14603 10968 14648 10996
rect 14642 10956 14648 10968
rect 14700 10956 14706 11008
rect 15562 10996 15568 11008
rect 15523 10968 15568 10996
rect 15562 10956 15568 10968
rect 15620 10956 15626 11008
rect 16316 10996 16344 11036
rect 16531 11033 16543 11067
rect 16577 11064 16589 11067
rect 17126 11064 17132 11076
rect 16577 11036 17132 11064
rect 16577 11033 16589 11036
rect 16531 11027 16589 11033
rect 17126 11024 17132 11036
rect 17184 11024 17190 11076
rect 17494 11024 17500 11076
rect 17552 11064 17558 11076
rect 17865 11067 17923 11073
rect 17865 11064 17877 11067
rect 17552 11036 17877 11064
rect 17552 11024 17558 11036
rect 17865 11033 17877 11036
rect 17911 11033 17923 11067
rect 17865 11027 17923 11033
rect 17218 10996 17224 11008
rect 16316 10968 17224 10996
rect 17218 10956 17224 10968
rect 17276 10956 17282 11008
rect 1104 10906 19019 10928
rect 1104 10854 5388 10906
rect 5440 10854 5452 10906
rect 5504 10854 5516 10906
rect 5568 10854 5580 10906
rect 5632 10854 5644 10906
rect 5696 10854 9827 10906
rect 9879 10854 9891 10906
rect 9943 10854 9955 10906
rect 10007 10854 10019 10906
rect 10071 10854 10083 10906
rect 10135 10854 14266 10906
rect 14318 10854 14330 10906
rect 14382 10854 14394 10906
rect 14446 10854 14458 10906
rect 14510 10854 14522 10906
rect 14574 10854 18705 10906
rect 18757 10854 18769 10906
rect 18821 10854 18833 10906
rect 18885 10854 18897 10906
rect 18949 10854 18961 10906
rect 19013 10854 19019 10906
rect 1104 10832 19019 10854
rect 3421 10795 3479 10801
rect 3421 10761 3433 10795
rect 3467 10792 3479 10795
rect 7929 10795 7987 10801
rect 3467 10764 4200 10792
rect 3467 10761 3479 10764
rect 3421 10755 3479 10761
rect 2593 10659 2651 10665
rect 2593 10625 2605 10659
rect 2639 10656 2651 10659
rect 2774 10656 2780 10668
rect 2639 10628 2780 10656
rect 2639 10625 2651 10628
rect 2593 10619 2651 10625
rect 2774 10616 2780 10628
rect 2832 10616 2838 10668
rect 3234 10656 3240 10668
rect 3195 10628 3240 10656
rect 3234 10616 3240 10628
rect 3292 10616 3298 10668
rect 4172 10665 4200 10764
rect 7929 10761 7941 10795
rect 7975 10792 7987 10795
rect 9306 10792 9312 10804
rect 7975 10764 9312 10792
rect 7975 10761 7987 10764
rect 7929 10755 7987 10761
rect 9306 10752 9312 10764
rect 9364 10752 9370 10804
rect 9493 10795 9551 10801
rect 9493 10761 9505 10795
rect 9539 10792 9551 10795
rect 11514 10792 11520 10804
rect 9539 10764 11520 10792
rect 9539 10761 9551 10764
rect 9493 10755 9551 10761
rect 11514 10752 11520 10764
rect 11572 10752 11578 10804
rect 11790 10792 11796 10804
rect 11751 10764 11796 10792
rect 11790 10752 11796 10764
rect 11848 10752 11854 10804
rect 12529 10795 12587 10801
rect 12529 10761 12541 10795
rect 12575 10792 12587 10795
rect 12618 10792 12624 10804
rect 12575 10764 12624 10792
rect 12575 10761 12587 10764
rect 12529 10755 12587 10761
rect 12618 10752 12624 10764
rect 12676 10752 12682 10804
rect 12894 10752 12900 10804
rect 12952 10792 12958 10804
rect 15378 10792 15384 10804
rect 12952 10764 14780 10792
rect 15291 10764 15384 10792
rect 12952 10752 12958 10764
rect 8018 10724 8024 10736
rect 6012 10696 8024 10724
rect 4157 10659 4215 10665
rect 4157 10625 4169 10659
rect 4203 10656 4215 10659
rect 4246 10656 4252 10668
rect 4203 10628 4252 10656
rect 4203 10625 4215 10628
rect 4157 10619 4215 10625
rect 4246 10616 4252 10628
rect 4304 10616 4310 10668
rect 6012 10665 6040 10696
rect 8018 10684 8024 10696
rect 8076 10684 8082 10736
rect 8478 10684 8484 10736
rect 8536 10724 8542 10736
rect 8536 10696 8708 10724
rect 8536 10684 8542 10696
rect 4341 10659 4399 10665
rect 4341 10625 4353 10659
rect 4387 10656 4399 10659
rect 4985 10659 5043 10665
rect 4985 10656 4997 10659
rect 4387 10628 4997 10656
rect 4387 10625 4399 10628
rect 4341 10619 4399 10625
rect 4985 10625 4997 10628
rect 5031 10625 5043 10659
rect 4985 10619 5043 10625
rect 5813 10659 5871 10665
rect 5813 10625 5825 10659
rect 5859 10625 5871 10659
rect 5813 10619 5871 10625
rect 5997 10659 6055 10665
rect 5997 10625 6009 10659
rect 6043 10625 6055 10659
rect 5997 10619 6055 10625
rect 6816 10659 6874 10665
rect 6816 10625 6828 10659
rect 6862 10656 6874 10659
rect 7374 10656 7380 10668
rect 6862 10628 7380 10656
rect 6862 10625 6874 10628
rect 6816 10619 6874 10625
rect 3973 10591 4031 10597
rect 3973 10557 3985 10591
rect 4019 10588 4031 10591
rect 4430 10588 4436 10600
rect 4019 10560 4436 10588
rect 4019 10557 4031 10560
rect 3973 10551 4031 10557
rect 4430 10548 4436 10560
rect 4488 10548 4494 10600
rect 5828 10588 5856 10619
rect 7374 10616 7380 10628
rect 7432 10616 7438 10668
rect 8202 10616 8208 10668
rect 8260 10656 8266 10668
rect 8389 10659 8447 10665
rect 8389 10656 8401 10659
rect 8260 10628 8401 10656
rect 8260 10616 8266 10628
rect 8389 10625 8401 10628
rect 8435 10625 8447 10659
rect 8570 10656 8576 10668
rect 8531 10628 8576 10656
rect 8389 10619 8447 10625
rect 6086 10588 6092 10600
rect 5828 10560 6092 10588
rect 6086 10548 6092 10560
rect 6144 10548 6150 10600
rect 6546 10588 6552 10600
rect 6507 10560 6552 10588
rect 6546 10548 6552 10560
rect 6604 10548 6610 10600
rect 8404 10588 8432 10619
rect 8570 10616 8576 10628
rect 8628 10616 8634 10668
rect 8680 10665 8708 10696
rect 9214 10684 9220 10736
rect 9272 10724 9278 10736
rect 9677 10727 9735 10733
rect 9677 10724 9689 10727
rect 9272 10696 9689 10724
rect 9272 10684 9278 10696
rect 9677 10693 9689 10696
rect 9723 10693 9735 10727
rect 9677 10687 9735 10693
rect 14268 10727 14326 10733
rect 14268 10693 14280 10727
rect 14314 10724 14326 10727
rect 14642 10724 14648 10736
rect 14314 10696 14648 10724
rect 14314 10693 14326 10696
rect 14268 10687 14326 10693
rect 14642 10684 14648 10696
rect 14700 10684 14706 10736
rect 14752 10724 14780 10764
rect 15378 10752 15384 10764
rect 15436 10792 15442 10804
rect 17126 10792 17132 10804
rect 15436 10764 17132 10792
rect 15436 10752 15442 10764
rect 17126 10752 17132 10764
rect 17184 10792 17190 10804
rect 17221 10795 17279 10801
rect 17221 10792 17233 10795
rect 17184 10764 17233 10792
rect 17184 10752 17190 10764
rect 17221 10761 17233 10764
rect 17267 10761 17279 10795
rect 17402 10792 17408 10804
rect 17363 10764 17408 10792
rect 17221 10755 17279 10761
rect 17402 10752 17408 10764
rect 17460 10752 17466 10804
rect 16390 10724 16396 10736
rect 14752 10696 16396 10724
rect 16390 10684 16396 10696
rect 16448 10684 16454 10736
rect 17494 10684 17500 10736
rect 17552 10724 17558 10736
rect 18325 10727 18383 10733
rect 18325 10724 18337 10727
rect 17552 10696 18337 10724
rect 17552 10684 17558 10696
rect 18325 10693 18337 10696
rect 18371 10693 18383 10727
rect 18325 10687 18383 10693
rect 8665 10659 8723 10665
rect 8665 10625 8677 10659
rect 8711 10625 8723 10659
rect 9306 10656 9312 10668
rect 9267 10628 9312 10656
rect 8665 10619 8723 10625
rect 9306 10616 9312 10628
rect 9364 10616 9370 10668
rect 9401 10659 9459 10665
rect 9401 10625 9413 10659
rect 9447 10656 9459 10659
rect 9490 10656 9496 10668
rect 9447 10628 9496 10656
rect 9447 10625 9459 10628
rect 9401 10619 9459 10625
rect 9490 10616 9496 10628
rect 9548 10616 9554 10668
rect 10318 10616 10324 10668
rect 10376 10656 10382 10668
rect 10413 10659 10471 10665
rect 10413 10656 10425 10659
rect 10376 10628 10425 10656
rect 10376 10616 10382 10628
rect 10413 10625 10425 10628
rect 10459 10625 10471 10659
rect 11698 10656 11704 10668
rect 10413 10619 10471 10625
rect 10520 10628 11704 10656
rect 10336 10588 10364 10616
rect 10520 10597 10548 10628
rect 11698 10616 11704 10628
rect 11756 10616 11762 10668
rect 11885 10659 11943 10665
rect 11885 10625 11897 10659
rect 11931 10656 11943 10659
rect 12526 10656 12532 10668
rect 11931 10628 12532 10656
rect 11931 10625 11943 10628
rect 11885 10619 11943 10625
rect 8404 10560 10364 10588
rect 10505 10591 10563 10597
rect 10505 10557 10517 10591
rect 10551 10557 10563 10591
rect 11900 10588 11928 10619
rect 12526 10616 12532 10628
rect 12584 10616 12590 10668
rect 12802 10656 12808 10668
rect 12763 10628 12808 10656
rect 12802 10616 12808 10628
rect 12860 10616 12866 10668
rect 12986 10656 12992 10668
rect 12947 10628 12992 10656
rect 12986 10616 12992 10628
rect 13044 10616 13050 10668
rect 13998 10656 14004 10668
rect 13959 10628 14004 10656
rect 13998 10616 14004 10628
rect 14056 10616 14062 10668
rect 15838 10656 15844 10668
rect 14108 10628 15844 10656
rect 10505 10551 10563 10557
rect 10704 10560 11928 10588
rect 12713 10591 12771 10597
rect 8478 10480 8484 10532
rect 8536 10520 8542 10532
rect 10704 10520 10732 10560
rect 12713 10557 12725 10591
rect 12759 10557 12771 10591
rect 12894 10588 12900 10600
rect 12855 10560 12900 10588
rect 12713 10551 12771 10557
rect 8536 10492 10732 10520
rect 10781 10523 10839 10529
rect 8536 10480 8542 10492
rect 10781 10489 10793 10523
rect 10827 10520 10839 10523
rect 12728 10520 12756 10551
rect 12894 10548 12900 10560
rect 12952 10548 12958 10600
rect 14108 10588 14136 10628
rect 15838 10616 15844 10628
rect 15896 10616 15902 10668
rect 15930 10616 15936 10668
rect 15988 10656 15994 10668
rect 16025 10659 16083 10665
rect 16025 10656 16037 10659
rect 15988 10628 16037 10656
rect 15988 10616 15994 10628
rect 16025 10625 16037 10628
rect 16071 10625 16083 10659
rect 16025 10619 16083 10625
rect 16574 10616 16580 10668
rect 16632 10656 16638 10668
rect 17129 10659 17187 10665
rect 17129 10656 17141 10659
rect 16632 10628 17141 10656
rect 16632 10616 16638 10628
rect 17129 10625 17141 10628
rect 17175 10625 17187 10659
rect 17129 10619 17187 10625
rect 17586 10616 17592 10668
rect 17644 10656 17650 10668
rect 17957 10659 18015 10665
rect 17957 10656 17969 10659
rect 17644 10628 17969 10656
rect 17644 10616 17650 10628
rect 17957 10625 17969 10628
rect 18003 10625 18015 10659
rect 17957 10619 18015 10625
rect 17034 10588 17040 10600
rect 13004 10560 14136 10588
rect 16995 10560 17040 10588
rect 12802 10520 12808 10532
rect 10827 10492 12434 10520
rect 12715 10492 12808 10520
rect 10827 10489 10839 10492
rect 10781 10483 10839 10489
rect 2774 10412 2780 10464
rect 2832 10452 2838 10464
rect 4798 10452 4804 10464
rect 2832 10424 2877 10452
rect 4759 10424 4804 10452
rect 2832 10412 2838 10424
rect 4798 10412 4804 10424
rect 4856 10412 4862 10464
rect 5997 10455 6055 10461
rect 5997 10421 6009 10455
rect 6043 10452 6055 10455
rect 7466 10452 7472 10464
rect 6043 10424 7472 10452
rect 6043 10421 6055 10424
rect 5997 10415 6055 10421
rect 7466 10412 7472 10424
rect 7524 10412 7530 10464
rect 7926 10412 7932 10464
rect 7984 10452 7990 10464
rect 8389 10455 8447 10461
rect 8389 10452 8401 10455
rect 7984 10424 8401 10452
rect 7984 10412 7990 10424
rect 8389 10421 8401 10424
rect 8435 10421 8447 10455
rect 9122 10452 9128 10464
rect 9083 10424 9128 10452
rect 8389 10415 8447 10421
rect 9122 10412 9128 10424
rect 9180 10412 9186 10464
rect 12406 10452 12434 10492
rect 12802 10480 12808 10492
rect 12860 10520 12866 10532
rect 13004 10520 13032 10560
rect 17034 10548 17040 10560
rect 17092 10548 17098 10600
rect 17218 10548 17224 10600
rect 17276 10588 17282 10600
rect 17497 10591 17555 10597
rect 17497 10588 17509 10591
rect 17276 10560 17509 10588
rect 17276 10548 17282 10560
rect 17497 10557 17509 10560
rect 17543 10557 17555 10591
rect 17497 10551 17555 10557
rect 18046 10548 18052 10600
rect 18104 10588 18110 10600
rect 18141 10591 18199 10597
rect 18141 10588 18153 10591
rect 18104 10560 18153 10588
rect 18104 10548 18110 10560
rect 18141 10557 18153 10560
rect 18187 10557 18199 10591
rect 18141 10551 18199 10557
rect 12860 10492 13032 10520
rect 12860 10480 12866 10492
rect 13262 10452 13268 10464
rect 12406 10424 13268 10452
rect 13262 10412 13268 10424
rect 13320 10412 13326 10464
rect 16022 10452 16028 10464
rect 15983 10424 16028 10452
rect 16022 10412 16028 10424
rect 16080 10412 16086 10464
rect 16850 10452 16856 10464
rect 16811 10424 16856 10452
rect 16850 10412 16856 10424
rect 16908 10412 16914 10464
rect 17678 10412 17684 10464
rect 17736 10452 17742 10464
rect 18049 10455 18107 10461
rect 18049 10452 18061 10455
rect 17736 10424 18061 10452
rect 17736 10412 17742 10424
rect 18049 10421 18061 10424
rect 18095 10421 18107 10455
rect 18049 10415 18107 10421
rect 18138 10412 18144 10464
rect 18196 10452 18202 10464
rect 18325 10455 18383 10461
rect 18325 10452 18337 10455
rect 18196 10424 18337 10452
rect 18196 10412 18202 10424
rect 18325 10421 18337 10424
rect 18371 10421 18383 10455
rect 18325 10415 18383 10421
rect 1104 10362 18860 10384
rect 1104 10310 3169 10362
rect 3221 10310 3233 10362
rect 3285 10310 3297 10362
rect 3349 10310 3361 10362
rect 3413 10310 3425 10362
rect 3477 10310 7608 10362
rect 7660 10310 7672 10362
rect 7724 10310 7736 10362
rect 7788 10310 7800 10362
rect 7852 10310 7864 10362
rect 7916 10310 12047 10362
rect 12099 10310 12111 10362
rect 12163 10310 12175 10362
rect 12227 10310 12239 10362
rect 12291 10310 12303 10362
rect 12355 10310 16486 10362
rect 16538 10310 16550 10362
rect 16602 10310 16614 10362
rect 16666 10310 16678 10362
rect 16730 10310 16742 10362
rect 16794 10310 18860 10362
rect 1104 10288 18860 10310
rect 3694 10208 3700 10260
rect 3752 10248 3758 10260
rect 3973 10251 4031 10257
rect 3973 10248 3985 10251
rect 3752 10220 3985 10248
rect 3752 10208 3758 10220
rect 3973 10217 3985 10220
rect 4019 10217 4031 10251
rect 3973 10211 4031 10217
rect 5721 10251 5779 10257
rect 5721 10217 5733 10251
rect 5767 10248 5779 10251
rect 6546 10248 6552 10260
rect 5767 10220 6552 10248
rect 5767 10217 5779 10220
rect 5721 10211 5779 10217
rect 6546 10208 6552 10220
rect 6604 10208 6610 10260
rect 7374 10208 7380 10260
rect 7432 10248 7438 10260
rect 7469 10251 7527 10257
rect 7469 10248 7481 10251
rect 7432 10220 7481 10248
rect 7432 10208 7438 10220
rect 7469 10217 7481 10220
rect 7515 10217 7527 10251
rect 7469 10211 7527 10217
rect 8573 10251 8631 10257
rect 8573 10217 8585 10251
rect 8619 10248 8631 10251
rect 8662 10248 8668 10260
rect 8619 10220 8668 10248
rect 8619 10217 8631 10220
rect 8573 10211 8631 10217
rect 8662 10208 8668 10220
rect 8720 10208 8726 10260
rect 9674 10208 9680 10260
rect 9732 10248 9738 10260
rect 10413 10251 10471 10257
rect 10413 10248 10425 10251
rect 9732 10220 10425 10248
rect 9732 10208 9738 10220
rect 10413 10217 10425 10220
rect 10459 10217 10471 10251
rect 10413 10211 10471 10217
rect 11698 10208 11704 10260
rect 11756 10248 11762 10260
rect 11756 10220 13952 10248
rect 11756 10208 11762 10220
rect 7282 10140 7288 10192
rect 7340 10180 7346 10192
rect 7837 10183 7895 10189
rect 7837 10180 7849 10183
rect 7340 10152 7849 10180
rect 7340 10140 7346 10152
rect 7837 10149 7849 10152
rect 7883 10149 7895 10183
rect 7837 10143 7895 10149
rect 9692 10112 9720 10208
rect 11514 10140 11520 10192
rect 11572 10180 11578 10192
rect 13170 10180 13176 10192
rect 11572 10152 12434 10180
rect 13131 10152 13176 10180
rect 11572 10140 11578 10152
rect 7024 10084 9720 10112
rect 7024 10056 7052 10084
rect 10502 10072 10508 10124
rect 10560 10112 10566 10124
rect 12406 10112 12434 10152
rect 13170 10140 13176 10152
rect 13228 10140 13234 10192
rect 13924 10180 13952 10220
rect 14734 10208 14740 10260
rect 14792 10248 14798 10260
rect 15105 10251 15163 10257
rect 15105 10248 15117 10251
rect 14792 10220 15117 10248
rect 14792 10208 14798 10220
rect 15105 10217 15117 10220
rect 15151 10217 15163 10251
rect 15105 10211 15163 10217
rect 15562 10208 15568 10260
rect 15620 10248 15626 10260
rect 15657 10251 15715 10257
rect 15657 10248 15669 10251
rect 15620 10220 15669 10248
rect 15620 10208 15626 10220
rect 15657 10217 15669 10220
rect 15703 10217 15715 10251
rect 15657 10211 15715 10217
rect 17037 10251 17095 10257
rect 17037 10217 17049 10251
rect 17083 10248 17095 10251
rect 17494 10248 17500 10260
rect 17083 10220 17500 10248
rect 17083 10217 17095 10220
rect 17037 10211 17095 10217
rect 17494 10208 17500 10220
rect 17552 10208 17558 10260
rect 17770 10248 17776 10260
rect 17731 10220 17776 10248
rect 17770 10208 17776 10220
rect 17828 10208 17834 10260
rect 17862 10208 17868 10260
rect 17920 10208 17926 10260
rect 15470 10180 15476 10192
rect 13924 10152 15476 10180
rect 15470 10140 15476 10152
rect 15528 10140 15534 10192
rect 17880 10180 17908 10208
rect 16776 10152 17908 10180
rect 12897 10115 12955 10121
rect 12897 10112 12909 10115
rect 10560 10084 11652 10112
rect 12406 10084 12909 10112
rect 10560 10072 10566 10084
rect 2317 10047 2375 10053
rect 2317 10013 2329 10047
rect 2363 10044 2375 10047
rect 2685 10047 2743 10053
rect 2363 10016 2636 10044
rect 2363 10013 2375 10016
rect 2317 10007 2375 10013
rect 2498 9976 2504 9988
rect 2459 9948 2504 9976
rect 2498 9936 2504 9948
rect 2556 9936 2562 9988
rect 2608 9976 2636 10016
rect 2685 10013 2697 10047
rect 2731 10044 2743 10047
rect 3145 10047 3203 10053
rect 3145 10044 3157 10047
rect 2731 10016 3157 10044
rect 2731 10013 2743 10016
rect 2685 10007 2743 10013
rect 3145 10013 3157 10016
rect 3191 10013 3203 10047
rect 7006 10044 7012 10056
rect 6919 10016 7012 10044
rect 3145 10007 3203 10013
rect 7006 10004 7012 10016
rect 7064 10004 7070 10056
rect 7466 10004 7472 10056
rect 7524 10044 7530 10056
rect 7653 10047 7711 10053
rect 7653 10044 7665 10047
rect 7524 10016 7665 10044
rect 7524 10004 7530 10016
rect 7653 10013 7665 10016
rect 7699 10013 7711 10047
rect 7653 10007 7711 10013
rect 7929 10047 7987 10053
rect 7929 10013 7941 10047
rect 7975 10044 7987 10047
rect 8110 10044 8116 10056
rect 7975 10016 8116 10044
rect 7975 10013 7987 10016
rect 7929 10007 7987 10013
rect 8110 10004 8116 10016
rect 8168 10004 8174 10056
rect 8662 10004 8668 10056
rect 8720 10044 8726 10056
rect 9125 10047 9183 10053
rect 9125 10044 9137 10047
rect 8720 10016 9137 10044
rect 8720 10004 8726 10016
rect 9125 10013 9137 10016
rect 9171 10013 9183 10047
rect 11330 10044 11336 10056
rect 11291 10016 11336 10044
rect 9125 10007 9183 10013
rect 11330 10004 11336 10016
rect 11388 10004 11394 10056
rect 11624 10053 11652 10084
rect 12897 10081 12909 10084
rect 12943 10112 12955 10115
rect 15930 10112 15936 10124
rect 12943 10084 15936 10112
rect 12943 10081 12955 10084
rect 12897 10075 12955 10081
rect 15930 10072 15936 10084
rect 15988 10072 15994 10124
rect 16776 10112 16804 10152
rect 16684 10084 16804 10112
rect 11609 10047 11667 10053
rect 11609 10013 11621 10047
rect 11655 10013 11667 10047
rect 12802 10044 12808 10056
rect 12763 10016 12808 10044
rect 11609 10007 11667 10013
rect 12802 10004 12808 10016
rect 12860 10004 12866 10056
rect 15286 10047 15344 10053
rect 15286 10013 15298 10047
rect 15332 10044 15344 10047
rect 15378 10044 15384 10056
rect 15332 10016 15384 10044
rect 15332 10013 15344 10016
rect 15286 10007 15344 10013
rect 15378 10004 15384 10016
rect 15436 10004 15442 10056
rect 15746 10044 15752 10056
rect 15707 10016 15752 10044
rect 15746 10004 15752 10016
rect 15804 10004 15810 10056
rect 16684 10053 16712 10084
rect 17678 10072 17684 10124
rect 17736 10112 17742 10124
rect 17865 10115 17923 10121
rect 17865 10112 17877 10115
rect 17736 10084 17877 10112
rect 17736 10072 17742 10084
rect 17865 10081 17877 10084
rect 17911 10081 17923 10115
rect 17865 10075 17923 10081
rect 16669 10047 16727 10053
rect 16669 10013 16681 10047
rect 16715 10013 16727 10047
rect 16669 10007 16727 10013
rect 16761 10047 16819 10053
rect 16761 10013 16773 10047
rect 16807 10013 16819 10047
rect 16761 10007 16819 10013
rect 16853 10047 16911 10053
rect 16853 10013 16865 10047
rect 16899 10044 16911 10047
rect 17126 10044 17132 10056
rect 16899 10016 17132 10044
rect 16899 10013 16911 10016
rect 16853 10007 16911 10013
rect 3694 9976 3700 9988
rect 2608 9948 3700 9976
rect 3694 9936 3700 9948
rect 3752 9936 3758 9988
rect 8570 9936 8576 9988
rect 8628 9976 8634 9988
rect 9490 9976 9496 9988
rect 8628 9948 9496 9976
rect 8628 9936 8634 9948
rect 9490 9936 9496 9948
rect 9548 9936 9554 9988
rect 16776 9976 16804 10007
rect 17126 10004 17132 10016
rect 17184 10044 17190 10056
rect 17494 10044 17500 10056
rect 17184 10016 17500 10044
rect 17184 10004 17190 10016
rect 17494 10004 17500 10016
rect 17552 10004 17558 10056
rect 17586 10004 17592 10056
rect 17644 10044 17650 10056
rect 17773 10047 17831 10053
rect 17773 10044 17785 10047
rect 17644 10016 17785 10044
rect 17644 10004 17650 10016
rect 17773 10013 17785 10016
rect 17819 10013 17831 10047
rect 18046 10044 18052 10056
rect 18007 10016 18052 10044
rect 17773 10007 17831 10013
rect 18046 10004 18052 10016
rect 18104 10004 18110 10056
rect 17310 9976 17316 9988
rect 16776 9948 17316 9976
rect 17310 9936 17316 9948
rect 17368 9936 17374 9988
rect 3329 9911 3387 9917
rect 3329 9877 3341 9911
rect 3375 9908 3387 9911
rect 3602 9908 3608 9920
rect 3375 9880 3608 9908
rect 3375 9877 3387 9880
rect 3329 9871 3387 9877
rect 3602 9868 3608 9880
rect 3660 9868 3666 9920
rect 11422 9908 11428 9920
rect 11383 9880 11428 9908
rect 11422 9868 11428 9880
rect 11480 9868 11486 9920
rect 11606 9868 11612 9920
rect 11664 9908 11670 9920
rect 11793 9911 11851 9917
rect 11793 9908 11805 9911
rect 11664 9880 11805 9908
rect 11664 9868 11670 9880
rect 11793 9877 11805 9880
rect 11839 9877 11851 9911
rect 11793 9871 11851 9877
rect 13725 9911 13783 9917
rect 13725 9877 13737 9911
rect 13771 9908 13783 9911
rect 13814 9908 13820 9920
rect 13771 9880 13820 9908
rect 13771 9877 13783 9880
rect 13725 9871 13783 9877
rect 13814 9868 13820 9880
rect 13872 9908 13878 9920
rect 14369 9911 14427 9917
rect 14369 9908 14381 9911
rect 13872 9880 14381 9908
rect 13872 9868 13878 9880
rect 14369 9877 14381 9880
rect 14415 9908 14427 9911
rect 14826 9908 14832 9920
rect 14415 9880 14832 9908
rect 14415 9877 14427 9880
rect 14369 9871 14427 9877
rect 14826 9868 14832 9880
rect 14884 9868 14890 9920
rect 15289 9911 15347 9917
rect 15289 9877 15301 9911
rect 15335 9908 15347 9911
rect 15378 9908 15384 9920
rect 15335 9880 15384 9908
rect 15335 9877 15347 9880
rect 15289 9871 15347 9877
rect 15378 9868 15384 9880
rect 15436 9868 15442 9920
rect 17402 9868 17408 9920
rect 17460 9908 17466 9920
rect 17586 9908 17592 9920
rect 17460 9880 17592 9908
rect 17460 9868 17466 9880
rect 17586 9868 17592 9880
rect 17644 9868 17650 9920
rect 1104 9818 19019 9840
rect 1104 9766 5388 9818
rect 5440 9766 5452 9818
rect 5504 9766 5516 9818
rect 5568 9766 5580 9818
rect 5632 9766 5644 9818
rect 5696 9766 9827 9818
rect 9879 9766 9891 9818
rect 9943 9766 9955 9818
rect 10007 9766 10019 9818
rect 10071 9766 10083 9818
rect 10135 9766 14266 9818
rect 14318 9766 14330 9818
rect 14382 9766 14394 9818
rect 14446 9766 14458 9818
rect 14510 9766 14522 9818
rect 14574 9766 18705 9818
rect 18757 9766 18769 9818
rect 18821 9766 18833 9818
rect 18885 9766 18897 9818
rect 18949 9766 18961 9818
rect 19013 9766 19019 9818
rect 1104 9744 19019 9766
rect 8757 9707 8815 9713
rect 8757 9673 8769 9707
rect 8803 9673 8815 9707
rect 8757 9667 8815 9673
rect 9769 9707 9827 9713
rect 9769 9673 9781 9707
rect 9815 9704 9827 9707
rect 10318 9704 10324 9716
rect 9815 9676 10324 9704
rect 9815 9673 9827 9676
rect 9769 9667 9827 9673
rect 2774 9596 2780 9648
rect 2832 9636 2838 9648
rect 3798 9639 3856 9645
rect 3798 9636 3810 9639
rect 2832 9608 3810 9636
rect 2832 9596 2838 9608
rect 3798 9605 3810 9608
rect 3844 9605 3856 9639
rect 4614 9636 4620 9648
rect 4527 9608 4620 9636
rect 3798 9599 3856 9605
rect 4540 9577 4568 9608
rect 4614 9596 4620 9608
rect 4672 9636 4678 9648
rect 6546 9636 6552 9648
rect 4672 9608 6552 9636
rect 4672 9596 4678 9608
rect 6546 9596 6552 9608
rect 6604 9636 6610 9648
rect 8772 9636 8800 9667
rect 10318 9664 10324 9676
rect 10376 9664 10382 9716
rect 11422 9664 11428 9716
rect 11480 9704 11486 9716
rect 11480 9676 12434 9704
rect 11480 9664 11486 9676
rect 9214 9636 9220 9648
rect 6604 9608 7420 9636
rect 8772 9608 9220 9636
rect 6604 9596 6610 9608
rect 4798 9577 4804 9580
rect 4065 9571 4123 9577
rect 4065 9537 4077 9571
rect 4111 9568 4123 9571
rect 4525 9571 4583 9577
rect 4525 9568 4537 9571
rect 4111 9540 4537 9568
rect 4111 9537 4123 9540
rect 4065 9531 4123 9537
rect 4525 9537 4537 9540
rect 4571 9537 4583 9571
rect 4792 9568 4804 9577
rect 4759 9540 4804 9568
rect 4525 9531 4583 9537
rect 4792 9531 4804 9540
rect 4798 9528 4804 9531
rect 4856 9528 4862 9580
rect 6730 9568 6736 9580
rect 6691 9540 6736 9568
rect 6730 9528 6736 9540
rect 6788 9528 6794 9580
rect 7392 9577 7420 9608
rect 9214 9596 9220 9608
rect 9272 9636 9278 9648
rect 9401 9639 9459 9645
rect 9401 9636 9413 9639
rect 9272 9608 9413 9636
rect 9272 9596 9278 9608
rect 9401 9605 9413 9608
rect 9447 9605 9459 9639
rect 9582 9636 9588 9648
rect 9543 9608 9588 9636
rect 9401 9599 9459 9605
rect 9582 9596 9588 9608
rect 9640 9596 9646 9648
rect 11238 9636 11244 9648
rect 10704 9608 11244 9636
rect 7377 9571 7435 9577
rect 7377 9537 7389 9571
rect 7423 9537 7435 9571
rect 7377 9531 7435 9537
rect 7466 9528 7472 9580
rect 7524 9568 7530 9580
rect 10704 9577 10732 9608
rect 11238 9596 11244 9608
rect 11296 9596 11302 9648
rect 11330 9596 11336 9648
rect 11388 9636 11394 9648
rect 11974 9636 11980 9648
rect 11388 9608 11980 9636
rect 11388 9596 11394 9608
rect 11974 9596 11980 9608
rect 12032 9596 12038 9648
rect 12406 9636 12434 9676
rect 12820 9676 14044 9704
rect 12820 9636 12848 9676
rect 12986 9636 12992 9648
rect 12406 9608 12848 9636
rect 12947 9608 12992 9636
rect 12986 9596 12992 9608
rect 13044 9596 13050 9648
rect 13170 9596 13176 9648
rect 13228 9636 13234 9648
rect 13693 9639 13751 9645
rect 13693 9636 13705 9639
rect 13228 9608 13705 9636
rect 13228 9596 13234 9608
rect 13693 9605 13705 9608
rect 13739 9605 13751 9639
rect 13906 9636 13912 9648
rect 13867 9608 13912 9636
rect 13693 9599 13751 9605
rect 13906 9596 13912 9608
rect 13964 9596 13970 9648
rect 14016 9636 14044 9676
rect 16942 9636 16948 9648
rect 14016 9608 16948 9636
rect 7633 9571 7691 9577
rect 7633 9568 7645 9571
rect 7524 9540 7645 9568
rect 7524 9528 7530 9540
rect 7633 9537 7645 9540
rect 7679 9537 7691 9571
rect 7633 9531 7691 9537
rect 10689 9571 10747 9577
rect 10689 9537 10701 9571
rect 10735 9537 10747 9571
rect 10689 9531 10747 9537
rect 10778 9528 10784 9580
rect 10836 9568 10842 9580
rect 11701 9571 11759 9577
rect 11701 9568 11713 9571
rect 10836 9540 11713 9568
rect 10836 9528 10842 9540
rect 11701 9537 11713 9540
rect 11747 9537 11759 9571
rect 11701 9531 11759 9537
rect 11793 9571 11851 9577
rect 11793 9537 11805 9571
rect 11839 9537 11851 9571
rect 11793 9531 11851 9537
rect 10594 9500 10600 9512
rect 10555 9472 10600 9500
rect 10594 9460 10600 9472
rect 10652 9460 10658 9512
rect 11422 9460 11428 9512
rect 11480 9500 11486 9512
rect 11808 9500 11836 9531
rect 12342 9528 12348 9580
rect 12400 9568 12406 9580
rect 12805 9571 12863 9577
rect 12805 9568 12817 9571
rect 12400 9540 12817 9568
rect 12400 9528 12406 9540
rect 12805 9537 12817 9540
rect 12851 9537 12863 9571
rect 12805 9531 12863 9537
rect 13081 9571 13139 9577
rect 13081 9537 13093 9571
rect 13127 9568 13139 9571
rect 14645 9571 14703 9577
rect 13127 9540 13584 9568
rect 13127 9537 13139 9540
rect 13081 9531 13139 9537
rect 11480 9472 11836 9500
rect 11480 9460 11486 9472
rect 11054 9392 11060 9444
rect 11112 9432 11118 9444
rect 12342 9432 12348 9444
rect 11112 9404 12348 9432
rect 11112 9392 11118 9404
rect 12342 9392 12348 9404
rect 12400 9432 12406 9444
rect 13170 9432 13176 9444
rect 12400 9392 12434 9432
rect 1854 9324 1860 9376
rect 1912 9364 1918 9376
rect 2498 9364 2504 9376
rect 1912 9336 2504 9364
rect 1912 9324 1918 9336
rect 2498 9324 2504 9336
rect 2556 9364 2562 9376
rect 2685 9367 2743 9373
rect 2685 9364 2697 9367
rect 2556 9336 2697 9364
rect 2556 9324 2562 9336
rect 2685 9333 2697 9336
rect 2731 9333 2743 9367
rect 2685 9327 2743 9333
rect 4154 9324 4160 9376
rect 4212 9364 4218 9376
rect 5905 9367 5963 9373
rect 5905 9364 5917 9367
rect 4212 9336 5917 9364
rect 4212 9324 4218 9336
rect 5905 9333 5917 9336
rect 5951 9333 5963 9367
rect 5905 9327 5963 9333
rect 6825 9367 6883 9373
rect 6825 9333 6837 9367
rect 6871 9364 6883 9367
rect 8110 9364 8116 9376
rect 6871 9336 8116 9364
rect 6871 9333 6883 9336
rect 6825 9327 6883 9333
rect 8110 9324 8116 9336
rect 8168 9324 8174 9376
rect 10962 9364 10968 9376
rect 10923 9336 10968 9364
rect 10962 9324 10968 9336
rect 11020 9324 11026 9376
rect 11701 9367 11759 9373
rect 11701 9333 11713 9367
rect 11747 9364 11759 9367
rect 11790 9364 11796 9376
rect 11747 9336 11796 9364
rect 11747 9333 11759 9336
rect 11701 9327 11759 9333
rect 11790 9324 11796 9336
rect 11848 9324 11854 9376
rect 12406 9364 12434 9392
rect 12728 9404 13176 9432
rect 12728 9364 12756 9404
rect 13170 9392 13176 9404
rect 13228 9392 13234 9444
rect 13446 9432 13452 9444
rect 13372 9404 13452 9432
rect 12406 9336 12756 9364
rect 12805 9367 12863 9373
rect 12805 9333 12817 9367
rect 12851 9364 12863 9367
rect 13372 9364 13400 9404
rect 13446 9392 13452 9404
rect 13504 9392 13510 9444
rect 13556 9432 13584 9540
rect 14645 9537 14657 9571
rect 14691 9568 14703 9571
rect 14734 9568 14740 9580
rect 14691 9540 14740 9568
rect 14691 9537 14703 9540
rect 14645 9531 14703 9537
rect 14734 9528 14740 9540
rect 14792 9528 14798 9580
rect 14826 9528 14832 9580
rect 14884 9568 14890 9580
rect 15764 9577 15792 9608
rect 16942 9596 16948 9608
rect 17000 9596 17006 9648
rect 17770 9636 17776 9648
rect 17731 9608 17776 9636
rect 17770 9596 17776 9608
rect 17828 9596 17834 9648
rect 15749 9571 15807 9577
rect 14884 9540 14929 9568
rect 14884 9528 14890 9540
rect 15749 9537 15761 9571
rect 15795 9537 15807 9571
rect 15749 9531 15807 9537
rect 15930 9528 15936 9580
rect 15988 9568 15994 9580
rect 16758 9568 16764 9580
rect 15988 9540 16764 9568
rect 15988 9528 15994 9540
rect 16758 9528 16764 9540
rect 16816 9528 16822 9580
rect 16853 9571 16911 9577
rect 16853 9537 16865 9571
rect 16899 9537 16911 9571
rect 16853 9531 16911 9537
rect 17037 9571 17095 9577
rect 17037 9537 17049 9571
rect 17083 9537 17095 9571
rect 17494 9568 17500 9580
rect 17455 9540 17500 9568
rect 17037 9531 17095 9537
rect 15194 9432 15200 9444
rect 13556 9404 15200 9432
rect 13538 9364 13544 9376
rect 12851 9336 13400 9364
rect 13499 9336 13544 9364
rect 12851 9333 12863 9336
rect 12805 9327 12863 9333
rect 13538 9324 13544 9336
rect 13596 9324 13602 9376
rect 13740 9373 13768 9404
rect 15194 9392 15200 9404
rect 15252 9392 15258 9444
rect 16868 9432 16896 9531
rect 17052 9500 17080 9531
rect 17494 9528 17500 9540
rect 17552 9528 17558 9580
rect 18138 9500 18144 9512
rect 17052 9472 18144 9500
rect 18138 9460 18144 9472
rect 18196 9460 18202 9512
rect 18046 9432 18052 9444
rect 16868 9404 18052 9432
rect 18046 9392 18052 9404
rect 18104 9392 18110 9444
rect 13725 9367 13783 9373
rect 13725 9333 13737 9367
rect 13771 9333 13783 9367
rect 14642 9364 14648 9376
rect 14603 9336 14648 9364
rect 13725 9327 13783 9333
rect 14642 9324 14648 9336
rect 14700 9324 14706 9376
rect 15286 9324 15292 9376
rect 15344 9364 15350 9376
rect 15841 9367 15899 9373
rect 15841 9364 15853 9367
rect 15344 9336 15853 9364
rect 15344 9324 15350 9336
rect 15841 9333 15853 9336
rect 15887 9333 15899 9367
rect 16942 9364 16948 9376
rect 16903 9336 16948 9364
rect 15841 9327 15899 9333
rect 16942 9324 16948 9336
rect 17000 9324 17006 9376
rect 1104 9274 18860 9296
rect 1104 9222 3169 9274
rect 3221 9222 3233 9274
rect 3285 9222 3297 9274
rect 3349 9222 3361 9274
rect 3413 9222 3425 9274
rect 3477 9222 7608 9274
rect 7660 9222 7672 9274
rect 7724 9222 7736 9274
rect 7788 9222 7800 9274
rect 7852 9222 7864 9274
rect 7916 9222 12047 9274
rect 12099 9222 12111 9274
rect 12163 9222 12175 9274
rect 12227 9222 12239 9274
rect 12291 9222 12303 9274
rect 12355 9222 16486 9274
rect 16538 9222 16550 9274
rect 16602 9222 16614 9274
rect 16666 9222 16678 9274
rect 16730 9222 16742 9274
rect 16794 9222 18860 9274
rect 1104 9200 18860 9222
rect 4893 9163 4951 9169
rect 4893 9129 4905 9163
rect 4939 9160 4951 9163
rect 4982 9160 4988 9172
rect 4939 9132 4988 9160
rect 4939 9129 4951 9132
rect 4893 9123 4951 9129
rect 4982 9120 4988 9132
rect 5040 9120 5046 9172
rect 7745 9163 7803 9169
rect 7745 9129 7757 9163
rect 7791 9160 7803 9163
rect 8202 9160 8208 9172
rect 7791 9132 8208 9160
rect 7791 9129 7803 9132
rect 7745 9123 7803 9129
rect 8202 9120 8208 9132
rect 8260 9120 8266 9172
rect 9217 9163 9275 9169
rect 9217 9129 9229 9163
rect 9263 9160 9275 9163
rect 9582 9160 9588 9172
rect 9263 9132 9588 9160
rect 9263 9129 9275 9132
rect 9217 9123 9275 9129
rect 9582 9120 9588 9132
rect 9640 9120 9646 9172
rect 10594 9120 10600 9172
rect 10652 9160 10658 9172
rect 10689 9163 10747 9169
rect 10689 9160 10701 9163
rect 10652 9132 10701 9160
rect 10652 9120 10658 9132
rect 10689 9129 10701 9132
rect 10735 9129 10747 9163
rect 12894 9160 12900 9172
rect 10689 9123 10747 9129
rect 10980 9132 12900 9160
rect 5077 9095 5135 9101
rect 5077 9061 5089 9095
rect 5123 9092 5135 9095
rect 5902 9092 5908 9104
rect 5123 9064 5908 9092
rect 5123 9061 5135 9064
rect 5077 9055 5135 9061
rect 5902 9052 5908 9064
rect 5960 9092 5966 9104
rect 6822 9092 6828 9104
rect 5960 9064 6828 9092
rect 5960 9052 5966 9064
rect 6822 9052 6828 9064
rect 6880 9052 6886 9104
rect 8018 9052 8024 9104
rect 8076 9092 8082 9104
rect 8297 9095 8355 9101
rect 8297 9092 8309 9095
rect 8076 9064 8309 9092
rect 8076 9052 8082 9064
rect 8297 9061 8309 9064
rect 8343 9061 8355 9095
rect 8297 9055 8355 9061
rect 10137 9095 10195 9101
rect 10137 9061 10149 9095
rect 10183 9092 10195 9095
rect 10502 9092 10508 9104
rect 10183 9064 10508 9092
rect 10183 9061 10195 9064
rect 10137 9055 10195 9061
rect 10502 9052 10508 9064
rect 10560 9092 10566 9104
rect 10980 9092 11008 9132
rect 12894 9120 12900 9132
rect 12952 9120 12958 9172
rect 12986 9120 12992 9172
rect 13044 9160 13050 9172
rect 13906 9160 13912 9172
rect 13044 9132 13912 9160
rect 13044 9120 13050 9132
rect 13906 9120 13912 9132
rect 13964 9120 13970 9172
rect 14734 9160 14740 9172
rect 14695 9132 14740 9160
rect 14734 9120 14740 9132
rect 14792 9120 14798 9172
rect 15286 9160 15292 9172
rect 15247 9132 15292 9160
rect 15286 9120 15292 9132
rect 15344 9120 15350 9172
rect 16022 9120 16028 9172
rect 16080 9160 16086 9172
rect 16209 9163 16267 9169
rect 16209 9160 16221 9163
rect 16080 9132 16221 9160
rect 16080 9120 16086 9132
rect 16209 9129 16221 9132
rect 16255 9129 16267 9163
rect 16209 9123 16267 9129
rect 17034 9120 17040 9172
rect 17092 9160 17098 9172
rect 17221 9163 17279 9169
rect 17221 9160 17233 9163
rect 17092 9132 17233 9160
rect 17092 9120 17098 9132
rect 17221 9129 17233 9132
rect 17267 9160 17279 9163
rect 17770 9160 17776 9172
rect 17267 9132 17776 9160
rect 17267 9129 17279 9132
rect 17221 9123 17279 9129
rect 17770 9120 17776 9132
rect 17828 9120 17834 9172
rect 11514 9092 11520 9104
rect 10560 9064 11008 9092
rect 11072 9064 11520 9092
rect 10560 9052 10566 9064
rect 10045 9027 10103 9033
rect 10045 8993 10057 9027
rect 10091 9024 10103 9027
rect 10226 9024 10232 9036
rect 10091 8996 10232 9024
rect 10091 8993 10103 8996
rect 10045 8987 10103 8993
rect 10226 8984 10232 8996
rect 10284 9024 10290 9036
rect 11072 9024 11100 9064
rect 11514 9052 11520 9064
rect 11572 9052 11578 9104
rect 15841 9095 15899 9101
rect 15841 9092 15853 9095
rect 12176 9064 15853 9092
rect 10284 8996 11100 9024
rect 11333 9027 11391 9033
rect 10284 8984 10290 8996
rect 11333 8993 11345 9027
rect 11379 9024 11391 9027
rect 11422 9024 11428 9036
rect 11379 8996 11428 9024
rect 11379 8993 11391 8996
rect 11333 8987 11391 8993
rect 11422 8984 11428 8996
rect 11480 8984 11486 9036
rect 5074 8916 5080 8968
rect 5132 8916 5138 8968
rect 5537 8959 5595 8965
rect 5537 8925 5549 8959
rect 5583 8925 5595 8959
rect 5718 8956 5724 8968
rect 5679 8928 5724 8956
rect 5537 8919 5595 8925
rect 4709 8891 4767 8897
rect 4709 8857 4721 8891
rect 4755 8888 4767 8891
rect 5092 8888 5120 8916
rect 4755 8860 5120 8888
rect 4755 8857 4767 8860
rect 4709 8851 4767 8857
rect 4890 8780 4896 8832
rect 4948 8829 4954 8832
rect 4948 8823 4967 8829
rect 4955 8789 4967 8823
rect 5552 8820 5580 8919
rect 5718 8916 5724 8928
rect 5776 8916 5782 8968
rect 7653 8959 7711 8965
rect 7653 8925 7665 8959
rect 7699 8956 7711 8959
rect 8294 8956 8300 8968
rect 7699 8928 8300 8956
rect 7699 8925 7711 8928
rect 7653 8919 7711 8925
rect 8294 8916 8300 8928
rect 8352 8916 8358 8968
rect 8481 8959 8539 8965
rect 8481 8925 8493 8959
rect 8527 8956 8539 8959
rect 9122 8956 9128 8968
rect 8527 8928 9128 8956
rect 8527 8925 8539 8928
rect 8481 8919 8539 8925
rect 9122 8916 9128 8928
rect 9180 8916 9186 8968
rect 9306 8916 9312 8968
rect 9364 8956 9370 8968
rect 9769 8959 9827 8965
rect 9769 8956 9781 8959
rect 9364 8928 9781 8956
rect 9364 8916 9370 8928
rect 9769 8925 9781 8928
rect 9815 8925 9827 8959
rect 9769 8919 9827 8925
rect 10962 8916 10968 8968
rect 11020 8956 11026 8968
rect 11698 8956 11704 8968
rect 11020 8928 11704 8956
rect 11020 8916 11026 8928
rect 11698 8916 11704 8928
rect 11756 8956 11762 8968
rect 12176 8965 12204 9064
rect 15841 9061 15853 9064
rect 15887 9061 15899 9095
rect 16114 9092 16120 9104
rect 16075 9064 16120 9092
rect 15841 9055 15899 9061
rect 16114 9052 16120 9064
rect 16172 9052 16178 9104
rect 17310 9092 17316 9104
rect 17271 9064 17316 9092
rect 17310 9052 17316 9064
rect 17368 9052 17374 9104
rect 12250 8984 12256 9036
rect 12308 9024 12314 9036
rect 12308 8996 12388 9024
rect 12308 8984 12314 8996
rect 12360 8965 12388 8996
rect 12434 8984 12440 9036
rect 12492 9024 12498 9036
rect 12492 8996 13400 9024
rect 12492 8984 12498 8996
rect 13372 8965 13400 8996
rect 13538 8984 13544 9036
rect 13596 9024 13602 9036
rect 15381 9027 15439 9033
rect 15381 9024 15393 9027
rect 13596 8996 13768 9024
rect 13596 8984 13602 8996
rect 11885 8959 11943 8965
rect 11885 8956 11897 8959
rect 11756 8928 11897 8956
rect 11756 8916 11762 8928
rect 11885 8925 11897 8928
rect 11931 8925 11943 8959
rect 11885 8919 11943 8925
rect 12161 8959 12219 8965
rect 12161 8925 12173 8959
rect 12207 8925 12219 8959
rect 12161 8919 12219 8925
rect 12345 8959 12403 8965
rect 12345 8925 12357 8959
rect 12391 8925 12403 8959
rect 12345 8919 12403 8925
rect 12621 8959 12679 8965
rect 12621 8925 12633 8959
rect 12667 8956 12679 8959
rect 13173 8959 13231 8965
rect 13173 8956 13185 8959
rect 12667 8928 13185 8956
rect 12667 8925 12679 8928
rect 12621 8919 12679 8925
rect 13173 8925 13185 8928
rect 13219 8925 13231 8959
rect 13173 8919 13231 8925
rect 13357 8959 13415 8965
rect 13357 8925 13369 8959
rect 13403 8925 13415 8959
rect 13357 8919 13415 8925
rect 13449 8959 13507 8965
rect 13449 8925 13461 8959
rect 13495 8925 13507 8959
rect 13630 8956 13636 8968
rect 13591 8928 13636 8956
rect 13449 8919 13507 8925
rect 5629 8891 5687 8897
rect 5629 8857 5641 8891
rect 5675 8888 5687 8891
rect 6362 8888 6368 8900
rect 5675 8860 6368 8888
rect 5675 8857 5687 8860
rect 5629 8851 5687 8857
rect 6362 8848 6368 8860
rect 6420 8848 6426 8900
rect 6546 8888 6552 8900
rect 6507 8860 6552 8888
rect 6546 8848 6552 8860
rect 6604 8848 6610 8900
rect 9582 8848 9588 8900
rect 9640 8888 9646 8900
rect 11422 8888 11428 8900
rect 9640 8860 11428 8888
rect 9640 8848 9646 8860
rect 11422 8848 11428 8860
rect 11480 8848 11486 8900
rect 11790 8848 11796 8900
rect 11848 8888 11854 8900
rect 13464 8888 13492 8919
rect 13630 8916 13636 8928
rect 13688 8916 13694 8968
rect 13740 8965 13768 8996
rect 13832 8996 15393 9024
rect 13725 8959 13783 8965
rect 13725 8925 13737 8959
rect 13771 8925 13783 8959
rect 13725 8919 13783 8925
rect 11848 8860 13492 8888
rect 11848 8848 11854 8860
rect 5810 8820 5816 8832
rect 5552 8792 5816 8820
rect 4948 8783 4967 8789
rect 4948 8780 4954 8783
rect 5810 8780 5816 8792
rect 5868 8780 5874 8832
rect 6181 8823 6239 8829
rect 6181 8789 6193 8823
rect 6227 8820 6239 8823
rect 7098 8820 7104 8832
rect 6227 8792 7104 8820
rect 6227 8789 6239 8792
rect 6181 8783 6239 8789
rect 7098 8780 7104 8792
rect 7156 8780 7162 8832
rect 11054 8820 11060 8832
rect 11015 8792 11060 8820
rect 11054 8780 11060 8792
rect 11112 8780 11118 8832
rect 11149 8823 11207 8829
rect 11149 8789 11161 8823
rect 11195 8820 11207 8823
rect 11882 8820 11888 8832
rect 11195 8792 11888 8820
rect 11195 8789 11207 8792
rect 11149 8783 11207 8789
rect 11882 8780 11888 8792
rect 11940 8780 11946 8832
rect 12437 8823 12495 8829
rect 12437 8789 12449 8823
rect 12483 8820 12495 8823
rect 12526 8820 12532 8832
rect 12483 8792 12532 8820
rect 12483 8789 12495 8792
rect 12437 8783 12495 8789
rect 12526 8780 12532 8792
rect 12584 8780 12590 8832
rect 12894 8780 12900 8832
rect 12952 8820 12958 8832
rect 13832 8820 13860 8996
rect 15381 8993 15393 8996
rect 15427 9024 15439 9027
rect 15746 9024 15752 9036
rect 15427 8996 15752 9024
rect 15427 8993 15439 8996
rect 15381 8987 15439 8993
rect 15746 8984 15752 8996
rect 15804 8984 15810 9036
rect 16301 9027 16359 9033
rect 16301 8993 16313 9027
rect 16347 9024 16359 9027
rect 17494 9024 17500 9036
rect 16347 8996 17500 9024
rect 16347 8993 16359 8996
rect 16301 8987 16359 8993
rect 17494 8984 17500 8996
rect 17552 8984 17558 9036
rect 14918 8959 14976 8965
rect 14918 8925 14930 8959
rect 14964 8956 14976 8959
rect 15010 8956 15016 8968
rect 14964 8928 15016 8956
rect 14964 8925 14976 8928
rect 14918 8919 14976 8925
rect 15010 8916 15016 8928
rect 15068 8916 15074 8968
rect 16577 8959 16635 8965
rect 16577 8925 16589 8959
rect 16623 8956 16635 8959
rect 16942 8956 16948 8968
rect 16623 8928 16948 8956
rect 16623 8925 16635 8928
rect 16577 8919 16635 8925
rect 16942 8916 16948 8928
rect 17000 8916 17006 8968
rect 17126 8916 17132 8968
rect 17184 8956 17190 8968
rect 17678 8956 17684 8968
rect 17184 8928 17684 8956
rect 17184 8916 17190 8928
rect 17678 8916 17684 8928
rect 17736 8916 17742 8968
rect 18046 8916 18052 8968
rect 18104 8956 18110 8968
rect 18141 8959 18199 8965
rect 18141 8956 18153 8959
rect 18104 8928 18153 8956
rect 18104 8916 18110 8928
rect 18141 8925 18153 8928
rect 18187 8925 18199 8959
rect 18141 8919 18199 8925
rect 13906 8848 13912 8900
rect 13964 8888 13970 8900
rect 17586 8888 17592 8900
rect 13964 8860 17592 8888
rect 13964 8848 13970 8860
rect 17586 8848 17592 8860
rect 17644 8848 17650 8900
rect 12952 8792 13860 8820
rect 12952 8780 12958 8792
rect 13998 8780 14004 8832
rect 14056 8820 14062 8832
rect 14921 8823 14979 8829
rect 14921 8820 14933 8823
rect 14056 8792 14933 8820
rect 14056 8780 14062 8792
rect 14921 8789 14933 8792
rect 14967 8820 14979 8823
rect 15102 8820 15108 8832
rect 14967 8792 15108 8820
rect 14967 8789 14979 8792
rect 14921 8783 14979 8789
rect 15102 8780 15108 8792
rect 15160 8820 15166 8832
rect 15378 8820 15384 8832
rect 15160 8792 15384 8820
rect 15160 8780 15166 8792
rect 15378 8780 15384 8792
rect 15436 8780 15442 8832
rect 16485 8823 16543 8829
rect 16485 8789 16497 8823
rect 16531 8820 16543 8823
rect 17034 8820 17040 8832
rect 16531 8792 17040 8820
rect 16531 8789 16543 8792
rect 16485 8783 16543 8789
rect 17034 8780 17040 8792
rect 17092 8780 17098 8832
rect 18230 8820 18236 8832
rect 18191 8792 18236 8820
rect 18230 8780 18236 8792
rect 18288 8780 18294 8832
rect 1104 8730 19019 8752
rect 1104 8678 5388 8730
rect 5440 8678 5452 8730
rect 5504 8678 5516 8730
rect 5568 8678 5580 8730
rect 5632 8678 5644 8730
rect 5696 8678 9827 8730
rect 9879 8678 9891 8730
rect 9943 8678 9955 8730
rect 10007 8678 10019 8730
rect 10071 8678 10083 8730
rect 10135 8678 14266 8730
rect 14318 8678 14330 8730
rect 14382 8678 14394 8730
rect 14446 8678 14458 8730
rect 14510 8678 14522 8730
rect 14574 8678 18705 8730
rect 18757 8678 18769 8730
rect 18821 8678 18833 8730
rect 18885 8678 18897 8730
rect 18949 8678 18961 8730
rect 19013 8678 19019 8730
rect 1104 8656 19019 8678
rect 4430 8616 4436 8628
rect 4391 8588 4436 8616
rect 4430 8576 4436 8588
rect 4488 8576 4494 8628
rect 6546 8616 6552 8628
rect 6507 8588 6552 8616
rect 6546 8576 6552 8588
rect 6604 8576 6610 8628
rect 6822 8576 6828 8628
rect 6880 8616 6886 8628
rect 6917 8619 6975 8625
rect 6917 8616 6929 8619
rect 6880 8588 6929 8616
rect 6880 8576 6886 8588
rect 6917 8585 6929 8588
rect 6963 8585 6975 8619
rect 6917 8579 6975 8585
rect 9674 8576 9680 8628
rect 9732 8616 9738 8628
rect 10318 8616 10324 8628
rect 9732 8588 10324 8616
rect 9732 8576 9738 8588
rect 10318 8576 10324 8588
rect 10376 8616 10382 8628
rect 10965 8619 11023 8625
rect 10965 8616 10977 8619
rect 10376 8588 10977 8616
rect 10376 8576 10382 8588
rect 10965 8585 10977 8588
rect 11011 8616 11023 8619
rect 12250 8616 12256 8628
rect 11011 8588 12256 8616
rect 11011 8585 11023 8588
rect 10965 8579 11023 8585
rect 12250 8576 12256 8588
rect 12308 8576 12314 8628
rect 12897 8619 12955 8625
rect 12897 8616 12909 8619
rect 12406 8588 12909 8616
rect 4614 8548 4620 8560
rect 3068 8520 4620 8548
rect 2133 8483 2191 8489
rect 2133 8449 2145 8483
rect 2179 8480 2191 8483
rect 2590 8480 2596 8492
rect 2179 8452 2596 8480
rect 2179 8449 2191 8452
rect 2133 8443 2191 8449
rect 2590 8440 2596 8452
rect 2648 8440 2654 8492
rect 3068 8489 3096 8520
rect 4614 8508 4620 8520
rect 4672 8508 4678 8560
rect 6362 8508 6368 8560
rect 6420 8548 6426 8560
rect 6420 8520 8340 8548
rect 6420 8508 6426 8520
rect 3053 8483 3111 8489
rect 3053 8449 3065 8483
rect 3099 8449 3111 8483
rect 3053 8443 3111 8449
rect 3320 8483 3378 8489
rect 3320 8449 3332 8483
rect 3366 8480 3378 8483
rect 3602 8480 3608 8492
rect 3366 8452 3608 8480
rect 3366 8449 3378 8452
rect 3320 8443 3378 8449
rect 3602 8440 3608 8452
rect 3660 8440 3666 8492
rect 5074 8480 5080 8492
rect 5035 8452 5080 8480
rect 5074 8440 5080 8452
rect 5132 8440 5138 8492
rect 6012 8452 7144 8480
rect 6012 8424 6040 8452
rect 2038 8412 2044 8424
rect 1999 8384 2044 8412
rect 2038 8372 2044 8384
rect 2096 8372 2102 8424
rect 4982 8412 4988 8424
rect 4943 8384 4988 8412
rect 4982 8372 4988 8384
rect 5040 8372 5046 8424
rect 5994 8412 6000 8424
rect 5368 8384 6000 8412
rect 2501 8347 2559 8353
rect 2501 8313 2513 8347
rect 2547 8344 2559 8347
rect 5368 8344 5396 8384
rect 5994 8372 6000 8384
rect 6052 8372 6058 8424
rect 7116 8421 7144 8452
rect 8110 8440 8116 8492
rect 8168 8480 8174 8492
rect 8312 8489 8340 8520
rect 8478 8508 8484 8560
rect 8536 8548 8542 8560
rect 8665 8551 8723 8557
rect 8665 8548 8677 8551
rect 8536 8520 8677 8548
rect 8536 8508 8542 8520
rect 8665 8517 8677 8520
rect 8711 8517 8723 8551
rect 8665 8511 8723 8517
rect 9214 8508 9220 8560
rect 9272 8548 9278 8560
rect 12406 8548 12434 8588
rect 12897 8585 12909 8588
rect 12943 8585 12955 8619
rect 12897 8579 12955 8585
rect 13173 8619 13231 8625
rect 13173 8585 13185 8619
rect 13219 8616 13231 8619
rect 13354 8616 13360 8628
rect 13219 8588 13360 8616
rect 13219 8585 13231 8588
rect 13173 8579 13231 8585
rect 13354 8576 13360 8588
rect 13412 8576 13418 8628
rect 17218 8616 17224 8628
rect 14200 8588 17224 8616
rect 9272 8520 12434 8548
rect 13056 8551 13114 8557
rect 9272 8508 9278 8520
rect 13056 8517 13068 8551
rect 13102 8548 13114 8551
rect 14200 8548 14228 8588
rect 17218 8576 17224 8588
rect 17276 8576 17282 8628
rect 13102 8520 14228 8548
rect 14268 8551 14326 8557
rect 13102 8517 13114 8520
rect 13056 8511 13114 8517
rect 14268 8517 14280 8551
rect 14314 8548 14326 8551
rect 14642 8548 14648 8560
rect 14314 8520 14648 8548
rect 14314 8517 14326 8520
rect 14268 8511 14326 8517
rect 14642 8508 14648 8520
rect 14700 8508 14706 8560
rect 16945 8551 17003 8557
rect 16945 8517 16957 8551
rect 16991 8548 17003 8551
rect 17126 8548 17132 8560
rect 16991 8520 17132 8548
rect 16991 8517 17003 8520
rect 16945 8511 17003 8517
rect 17126 8508 17132 8520
rect 17184 8508 17190 8560
rect 8205 8483 8263 8489
rect 8205 8480 8217 8483
rect 8168 8452 8217 8480
rect 8168 8440 8174 8452
rect 8205 8449 8217 8452
rect 8251 8449 8263 8483
rect 8205 8443 8263 8449
rect 8297 8483 8355 8489
rect 8297 8449 8309 8483
rect 8343 8449 8355 8483
rect 8297 8443 8355 8449
rect 9030 8440 9036 8492
rect 9088 8480 9094 8492
rect 9493 8483 9551 8489
rect 9493 8480 9505 8483
rect 9088 8452 9505 8480
rect 9088 8440 9094 8452
rect 9493 8449 9505 8452
rect 9539 8449 9551 8483
rect 10594 8480 10600 8492
rect 10555 8452 10600 8480
rect 9493 8443 9551 8449
rect 10594 8440 10600 8452
rect 10652 8440 10658 8492
rect 11054 8489 11060 8492
rect 11024 8483 11060 8489
rect 11024 8449 11036 8483
rect 11024 8443 11060 8449
rect 11054 8440 11060 8443
rect 11112 8440 11118 8492
rect 11698 8480 11704 8492
rect 11659 8452 11704 8480
rect 11698 8440 11704 8452
rect 11756 8440 11762 8492
rect 11790 8440 11796 8492
rect 11848 8480 11854 8492
rect 12069 8483 12127 8489
rect 12069 8480 12081 8483
rect 11848 8452 12081 8480
rect 11848 8440 11854 8452
rect 12069 8449 12081 8452
rect 12115 8449 12127 8483
rect 12069 8443 12127 8449
rect 13541 8483 13599 8489
rect 13541 8449 13553 8483
rect 13587 8480 13599 8483
rect 13722 8480 13728 8492
rect 13587 8452 13728 8480
rect 13587 8449 13599 8452
rect 13541 8443 13599 8449
rect 13722 8440 13728 8452
rect 13780 8440 13786 8492
rect 16025 8483 16083 8489
rect 16025 8449 16037 8483
rect 16071 8480 16083 8483
rect 16206 8480 16212 8492
rect 16071 8452 16212 8480
rect 16071 8449 16083 8452
rect 16025 8443 16083 8449
rect 16206 8440 16212 8452
rect 16264 8480 16270 8492
rect 16850 8480 16856 8492
rect 16264 8452 16856 8480
rect 16264 8440 16270 8452
rect 16850 8440 16856 8452
rect 16908 8440 16914 8492
rect 17586 8480 17592 8492
rect 17547 8452 17592 8480
rect 17586 8440 17592 8452
rect 17644 8440 17650 8492
rect 17681 8483 17739 8489
rect 17681 8449 17693 8483
rect 17727 8480 17739 8483
rect 18230 8480 18236 8492
rect 17727 8452 18236 8480
rect 17727 8449 17739 8452
rect 17681 8443 17739 8449
rect 18230 8440 18236 8452
rect 18288 8440 18294 8492
rect 7009 8415 7067 8421
rect 7009 8381 7021 8415
rect 7055 8381 7067 8415
rect 7009 8375 7067 8381
rect 7101 8415 7159 8421
rect 7101 8381 7113 8415
rect 7147 8381 7159 8415
rect 10502 8412 10508 8424
rect 10463 8384 10508 8412
rect 7101 8375 7159 8381
rect 2547 8316 3096 8344
rect 2547 8313 2559 8316
rect 2501 8307 2559 8313
rect 3068 8276 3096 8316
rect 3988 8316 5396 8344
rect 5445 8347 5503 8353
rect 3988 8276 4016 8316
rect 5445 8313 5457 8347
rect 5491 8344 5503 8347
rect 5810 8344 5816 8356
rect 5491 8316 5816 8344
rect 5491 8313 5503 8316
rect 5445 8307 5503 8313
rect 5810 8304 5816 8316
rect 5868 8344 5874 8356
rect 6730 8344 6736 8356
rect 5868 8316 6736 8344
rect 5868 8304 5874 8316
rect 6730 8304 6736 8316
rect 6788 8304 6794 8356
rect 6914 8304 6920 8356
rect 6972 8344 6978 8356
rect 7024 8344 7052 8375
rect 10502 8372 10508 8384
rect 10560 8372 10566 8424
rect 11606 8372 11612 8424
rect 11664 8412 11670 8424
rect 12253 8415 12311 8421
rect 12253 8412 12265 8415
rect 11664 8384 12265 8412
rect 11664 8372 11670 8384
rect 12253 8381 12265 8384
rect 12299 8412 12311 8415
rect 12342 8412 12348 8424
rect 12299 8384 12348 8412
rect 12299 8381 12311 8384
rect 12253 8375 12311 8381
rect 12342 8372 12348 8384
rect 12400 8372 12406 8424
rect 13262 8372 13268 8424
rect 13320 8412 13326 8424
rect 13998 8412 14004 8424
rect 13320 8384 13365 8412
rect 13959 8384 14004 8412
rect 13320 8372 13326 8384
rect 13998 8372 14004 8384
rect 14056 8372 14062 8424
rect 17770 8412 17776 8424
rect 17731 8384 17776 8412
rect 17770 8372 17776 8384
rect 17828 8372 17834 8424
rect 6972 8316 7052 8344
rect 8021 8347 8079 8353
rect 6972 8304 6978 8316
rect 8021 8313 8033 8347
rect 8067 8344 8079 8347
rect 8570 8344 8576 8356
rect 8067 8316 8576 8344
rect 8067 8313 8079 8316
rect 8021 8307 8079 8313
rect 8570 8304 8576 8316
rect 8628 8304 8634 8356
rect 9398 8304 9404 8356
rect 9456 8344 9462 8356
rect 11793 8347 11851 8353
rect 11793 8344 11805 8347
rect 9456 8316 11805 8344
rect 9456 8304 9462 8316
rect 11793 8313 11805 8316
rect 11839 8313 11851 8347
rect 13814 8344 13820 8356
rect 11793 8307 11851 8313
rect 11900 8316 13820 8344
rect 3068 8248 4016 8276
rect 8481 8279 8539 8285
rect 8481 8245 8493 8279
rect 8527 8276 8539 8279
rect 9674 8276 9680 8288
rect 8527 8248 9680 8276
rect 8527 8245 8539 8248
rect 8481 8239 8539 8245
rect 9674 8236 9680 8248
rect 9732 8236 9738 8288
rect 9769 8279 9827 8285
rect 9769 8245 9781 8279
rect 9815 8276 9827 8279
rect 10318 8276 10324 8288
rect 9815 8248 10324 8276
rect 9815 8245 9827 8248
rect 9769 8239 9827 8245
rect 10318 8236 10324 8248
rect 10376 8236 10382 8288
rect 11146 8276 11152 8288
rect 11107 8248 11152 8276
rect 11146 8236 11152 8248
rect 11204 8236 11210 8288
rect 11514 8236 11520 8288
rect 11572 8276 11578 8288
rect 11900 8276 11928 8316
rect 13814 8304 13820 8316
rect 13872 8304 13878 8356
rect 15010 8304 15016 8356
rect 15068 8344 15074 8356
rect 15381 8347 15439 8353
rect 15381 8344 15393 8347
rect 15068 8316 15393 8344
rect 15068 8304 15074 8316
rect 15381 8313 15393 8316
rect 15427 8344 15439 8347
rect 17310 8344 17316 8356
rect 15427 8316 17316 8344
rect 15427 8313 15439 8316
rect 15381 8307 15439 8313
rect 17310 8304 17316 8316
rect 17368 8304 17374 8356
rect 11572 8248 11928 8276
rect 16209 8279 16267 8285
rect 11572 8236 11578 8248
rect 16209 8245 16221 8279
rect 16255 8276 16267 8279
rect 16390 8276 16396 8288
rect 16255 8248 16396 8276
rect 16255 8245 16267 8248
rect 16209 8239 16267 8245
rect 16390 8236 16396 8248
rect 16448 8236 16454 8288
rect 17402 8276 17408 8288
rect 17363 8248 17408 8276
rect 17402 8236 17408 8248
rect 17460 8236 17466 8288
rect 1104 8186 18860 8208
rect 1104 8134 3169 8186
rect 3221 8134 3233 8186
rect 3285 8134 3297 8186
rect 3349 8134 3361 8186
rect 3413 8134 3425 8186
rect 3477 8134 7608 8186
rect 7660 8134 7672 8186
rect 7724 8134 7736 8186
rect 7788 8134 7800 8186
rect 7852 8134 7864 8186
rect 7916 8134 12047 8186
rect 12099 8134 12111 8186
rect 12163 8134 12175 8186
rect 12227 8134 12239 8186
rect 12291 8134 12303 8186
rect 12355 8134 16486 8186
rect 16538 8134 16550 8186
rect 16602 8134 16614 8186
rect 16666 8134 16678 8186
rect 16730 8134 16742 8186
rect 16794 8134 18860 8186
rect 1104 8112 18860 8134
rect 2038 8032 2044 8084
rect 2096 8072 2102 8084
rect 2133 8075 2191 8081
rect 2133 8072 2145 8075
rect 2096 8044 2145 8072
rect 2096 8032 2102 8044
rect 2133 8041 2145 8044
rect 2179 8041 2191 8075
rect 2590 8072 2596 8084
rect 2551 8044 2596 8072
rect 2133 8035 2191 8041
rect 2590 8032 2596 8044
rect 2648 8032 2654 8084
rect 5997 8075 6055 8081
rect 5997 8041 6009 8075
rect 6043 8072 6055 8075
rect 6914 8072 6920 8084
rect 6043 8044 6920 8072
rect 6043 8041 6055 8044
rect 5997 8035 6055 8041
rect 6914 8032 6920 8044
rect 6972 8032 6978 8084
rect 9306 8032 9312 8084
rect 9364 8072 9370 8084
rect 9585 8075 9643 8081
rect 9585 8072 9597 8075
rect 9364 8044 9597 8072
rect 9364 8032 9370 8044
rect 9585 8041 9597 8044
rect 9631 8041 9643 8075
rect 9585 8035 9643 8041
rect 3050 8004 3056 8016
rect 2792 7976 3056 8004
rect 1854 7936 1860 7948
rect 1815 7908 1860 7936
rect 1854 7896 1860 7908
rect 1912 7896 1918 7948
rect 2792 7945 2820 7976
rect 3050 7964 3056 7976
rect 3108 8004 3114 8016
rect 4982 8004 4988 8016
rect 3108 7976 4988 8004
rect 3108 7964 3114 7976
rect 4982 7964 4988 7976
rect 5040 7964 5046 8016
rect 8294 7964 8300 8016
rect 8352 7964 8358 8016
rect 2777 7939 2835 7945
rect 2777 7905 2789 7939
rect 2823 7905 2835 7939
rect 2777 7899 2835 7905
rect 2869 7939 2927 7945
rect 2869 7905 2881 7939
rect 2915 7936 2927 7939
rect 4249 7939 4307 7945
rect 2915 7908 4108 7936
rect 2915 7905 2927 7908
rect 2869 7899 2927 7905
rect 1765 7871 1823 7877
rect 1765 7837 1777 7871
rect 1811 7837 1823 7871
rect 1765 7831 1823 7837
rect 2961 7871 3019 7877
rect 2961 7837 2973 7871
rect 3007 7837 3019 7871
rect 2961 7831 3019 7837
rect 3053 7871 3111 7877
rect 3053 7837 3065 7871
rect 3099 7868 3111 7871
rect 3418 7868 3424 7880
rect 3099 7840 3424 7868
rect 3099 7837 3111 7840
rect 3053 7831 3111 7837
rect 1780 7732 1808 7831
rect 2976 7800 3004 7831
rect 3418 7828 3424 7840
rect 3476 7828 3482 7880
rect 4080 7868 4108 7908
rect 4249 7905 4261 7939
rect 4295 7936 4307 7939
rect 4801 7939 4859 7945
rect 4801 7936 4813 7939
rect 4295 7908 4813 7936
rect 4295 7905 4307 7908
rect 4249 7899 4307 7905
rect 4801 7905 4813 7908
rect 4847 7936 4859 7939
rect 5074 7936 5080 7948
rect 4847 7908 5080 7936
rect 4847 7905 4859 7908
rect 4801 7899 4859 7905
rect 5074 7896 5080 7908
rect 5132 7896 5138 7948
rect 7929 7939 7987 7945
rect 7929 7905 7941 7939
rect 7975 7936 7987 7939
rect 8312 7936 8340 7964
rect 9214 7936 9220 7948
rect 7975 7908 9220 7936
rect 7975 7905 7987 7908
rect 7929 7899 7987 7905
rect 9214 7896 9220 7908
rect 9272 7896 9278 7948
rect 4154 7868 4160 7880
rect 4212 7877 4218 7880
rect 4080 7840 4160 7868
rect 4154 7828 4160 7840
rect 4212 7868 4221 7877
rect 4341 7871 4399 7877
rect 4212 7840 4257 7868
rect 4212 7831 4221 7840
rect 4341 7837 4353 7871
rect 4387 7837 4399 7871
rect 4341 7831 4399 7837
rect 4212 7828 4218 7831
rect 3970 7800 3976 7812
rect 2976 7772 3976 7800
rect 3970 7760 3976 7772
rect 4028 7800 4034 7812
rect 4356 7800 4384 7831
rect 4890 7828 4896 7880
rect 4948 7868 4954 7880
rect 4985 7871 5043 7877
rect 4985 7868 4997 7871
rect 4948 7840 4997 7868
rect 4948 7828 4954 7840
rect 4985 7837 4997 7840
rect 5031 7837 5043 7871
rect 4985 7831 5043 7837
rect 5169 7871 5227 7877
rect 5169 7837 5181 7871
rect 5215 7868 5227 7871
rect 5718 7868 5724 7880
rect 5215 7840 5724 7868
rect 5215 7837 5227 7840
rect 5169 7831 5227 7837
rect 5718 7828 5724 7840
rect 5776 7868 5782 7880
rect 5813 7871 5871 7877
rect 5813 7868 5825 7871
rect 5776 7840 5825 7868
rect 5776 7828 5782 7840
rect 5813 7837 5825 7840
rect 5859 7837 5871 7871
rect 5813 7831 5871 7837
rect 5994 7828 6000 7880
rect 6052 7868 6058 7880
rect 6549 7871 6607 7877
rect 6549 7868 6561 7871
rect 6052 7840 6561 7868
rect 6052 7828 6058 7840
rect 6549 7837 6561 7840
rect 6595 7837 6607 7871
rect 6730 7868 6736 7880
rect 6691 7840 6736 7868
rect 6549 7831 6607 7837
rect 6730 7828 6736 7840
rect 6788 7828 6794 7880
rect 6822 7828 6828 7880
rect 6880 7868 6886 7880
rect 8297 7871 8355 7877
rect 8297 7868 8309 7871
rect 6880 7840 8309 7868
rect 6880 7828 6886 7840
rect 8297 7837 8309 7840
rect 8343 7837 8355 7871
rect 8478 7868 8484 7880
rect 8439 7840 8484 7868
rect 8297 7831 8355 7837
rect 8478 7828 8484 7840
rect 8536 7828 8542 7880
rect 9398 7868 9404 7880
rect 9359 7840 9404 7868
rect 9398 7828 9404 7840
rect 9456 7828 9462 7880
rect 9600 7868 9628 8035
rect 11882 8032 11888 8084
rect 11940 8072 11946 8084
rect 12069 8075 12127 8081
rect 12069 8072 12081 8075
rect 11940 8044 12081 8072
rect 11940 8032 11946 8044
rect 12069 8041 12081 8044
rect 12115 8041 12127 8075
rect 12069 8035 12127 8041
rect 13262 8032 13268 8084
rect 13320 8072 13326 8084
rect 13541 8075 13599 8081
rect 13541 8072 13553 8075
rect 13320 8044 13553 8072
rect 13320 8032 13326 8044
rect 13541 8041 13553 8044
rect 13587 8041 13599 8075
rect 17494 8072 17500 8084
rect 17455 8044 17500 8072
rect 13541 8035 13599 8041
rect 17494 8032 17500 8044
rect 17552 8032 17558 8084
rect 9674 7964 9680 8016
rect 9732 8004 9738 8016
rect 10321 8007 10379 8013
rect 10321 8004 10333 8007
rect 9732 7976 10333 8004
rect 9732 7964 9738 7976
rect 10321 7973 10333 7976
rect 10367 7973 10379 8007
rect 10321 7967 10379 7973
rect 11606 7964 11612 8016
rect 11664 8004 11670 8016
rect 13906 8004 13912 8016
rect 11664 7976 13912 8004
rect 11664 7964 11670 7976
rect 13906 7964 13912 7976
rect 13964 7964 13970 8016
rect 11054 7896 11060 7948
rect 11112 7936 11118 7948
rect 13630 7936 13636 7948
rect 11112 7908 12204 7936
rect 11112 7896 11118 7908
rect 12176 7880 12204 7908
rect 13372 7908 13636 7936
rect 10045 7871 10103 7877
rect 10045 7868 10057 7871
rect 9600 7840 10057 7868
rect 10045 7837 10057 7840
rect 10091 7837 10103 7871
rect 10045 7831 10103 7837
rect 10137 7871 10195 7877
rect 10137 7837 10149 7871
rect 10183 7868 10195 7871
rect 11977 7871 12035 7877
rect 10183 7840 10916 7868
rect 10183 7837 10195 7840
rect 10137 7831 10195 7837
rect 8113 7803 8171 7809
rect 4028 7772 4384 7800
rect 6748 7772 7512 7800
rect 4028 7760 4034 7772
rect 6748 7744 6776 7772
rect 2958 7732 2964 7744
rect 1780 7704 2964 7732
rect 2958 7692 2964 7704
rect 3016 7692 3022 7744
rect 6730 7692 6736 7744
rect 6788 7692 6794 7744
rect 6914 7732 6920 7744
rect 6875 7704 6920 7732
rect 6914 7692 6920 7704
rect 6972 7692 6978 7744
rect 7484 7741 7512 7772
rect 8113 7769 8125 7803
rect 8159 7800 8171 7803
rect 8386 7800 8392 7812
rect 8159 7772 8392 7800
rect 8159 7769 8171 7772
rect 8113 7763 8171 7769
rect 8386 7760 8392 7772
rect 8444 7800 8450 7812
rect 9416 7800 9444 7828
rect 8444 7772 9444 7800
rect 8444 7760 8450 7772
rect 9490 7760 9496 7812
rect 9548 7800 9554 7812
rect 10152 7800 10180 7831
rect 10318 7800 10324 7812
rect 9548 7772 10180 7800
rect 10279 7772 10324 7800
rect 9548 7760 9554 7772
rect 10318 7760 10324 7772
rect 10376 7800 10382 7812
rect 10781 7803 10839 7809
rect 10781 7800 10793 7803
rect 10376 7772 10793 7800
rect 10376 7760 10382 7772
rect 10781 7769 10793 7772
rect 10827 7769 10839 7803
rect 10781 7763 10839 7769
rect 7469 7735 7527 7741
rect 7469 7701 7481 7735
rect 7515 7732 7527 7735
rect 7558 7732 7564 7744
rect 7515 7704 7564 7732
rect 7515 7701 7527 7704
rect 7469 7695 7527 7701
rect 7558 7692 7564 7704
rect 7616 7692 7622 7744
rect 8205 7735 8263 7741
rect 8205 7701 8217 7735
rect 8251 7732 8263 7735
rect 8754 7732 8760 7744
rect 8251 7704 8760 7732
rect 8251 7701 8263 7704
rect 8205 7695 8263 7701
rect 8754 7692 8760 7704
rect 8812 7732 8818 7744
rect 10226 7732 10232 7744
rect 8812 7704 10232 7732
rect 8812 7692 8818 7704
rect 10226 7692 10232 7704
rect 10284 7692 10290 7744
rect 10888 7732 10916 7840
rect 11977 7837 11989 7871
rect 12023 7837 12035 7871
rect 12158 7868 12164 7880
rect 12119 7840 12164 7868
rect 11977 7831 12035 7837
rect 11992 7800 12020 7831
rect 12158 7828 12164 7840
rect 12216 7828 12222 7880
rect 13372 7877 13400 7908
rect 13630 7896 13636 7908
rect 13688 7896 13694 7948
rect 15838 7896 15844 7948
rect 15896 7936 15902 7948
rect 18046 7936 18052 7948
rect 15896 7908 18052 7936
rect 15896 7896 15902 7908
rect 18046 7896 18052 7908
rect 18104 7936 18110 7948
rect 18104 7908 18197 7936
rect 18104 7896 18110 7908
rect 13357 7871 13415 7877
rect 13357 7837 13369 7871
rect 13403 7837 13415 7871
rect 13538 7868 13544 7880
rect 13499 7840 13544 7868
rect 13357 7831 13415 7837
rect 13538 7828 13544 7840
rect 13596 7828 13602 7880
rect 16577 7871 16635 7877
rect 16577 7837 16589 7871
rect 16623 7837 16635 7871
rect 16577 7831 16635 7837
rect 16761 7871 16819 7877
rect 16761 7837 16773 7871
rect 16807 7868 16819 7871
rect 16850 7868 16856 7880
rect 16807 7840 16856 7868
rect 16807 7837 16819 7840
rect 16761 7831 16819 7837
rect 12802 7800 12808 7812
rect 11992 7772 12808 7800
rect 12802 7760 12808 7772
rect 12860 7760 12866 7812
rect 15841 7803 15899 7809
rect 15841 7769 15853 7803
rect 15887 7800 15899 7803
rect 16022 7800 16028 7812
rect 15887 7772 16028 7800
rect 15887 7769 15899 7772
rect 15841 7763 15899 7769
rect 16022 7760 16028 7772
rect 16080 7760 16086 7812
rect 16592 7800 16620 7831
rect 16850 7828 16856 7840
rect 16908 7828 16914 7880
rect 17770 7868 17776 7880
rect 17731 7840 17776 7868
rect 17770 7828 17776 7840
rect 17828 7828 17834 7880
rect 17865 7871 17923 7877
rect 17865 7837 17877 7871
rect 17911 7837 17923 7871
rect 17865 7831 17923 7837
rect 17957 7871 18015 7877
rect 17957 7837 17969 7871
rect 18003 7868 18015 7871
rect 18064 7868 18092 7896
rect 18003 7840 18092 7868
rect 18141 7871 18199 7877
rect 18003 7837 18015 7840
rect 17957 7831 18015 7837
rect 18141 7837 18153 7871
rect 18187 7868 18199 7871
rect 18230 7868 18236 7880
rect 18187 7840 18236 7868
rect 18187 7837 18199 7840
rect 18141 7831 18199 7837
rect 16942 7800 16948 7812
rect 16592 7772 16948 7800
rect 16942 7760 16948 7772
rect 17000 7760 17006 7812
rect 13078 7732 13084 7744
rect 10888 7704 13084 7732
rect 13078 7692 13084 7704
rect 13136 7692 13142 7744
rect 15749 7735 15807 7741
rect 15749 7701 15761 7735
rect 15795 7732 15807 7735
rect 15930 7732 15936 7744
rect 15795 7704 15936 7732
rect 15795 7701 15807 7704
rect 15749 7695 15807 7701
rect 15930 7692 15936 7704
rect 15988 7692 15994 7744
rect 16393 7735 16451 7741
rect 16393 7701 16405 7735
rect 16439 7732 16451 7735
rect 17126 7732 17132 7744
rect 16439 7704 17132 7732
rect 16439 7701 16451 7704
rect 16393 7695 16451 7701
rect 17126 7692 17132 7704
rect 17184 7692 17190 7744
rect 17880 7732 17908 7831
rect 18230 7828 18236 7840
rect 18288 7828 18294 7880
rect 18138 7732 18144 7744
rect 17880 7704 18144 7732
rect 18138 7692 18144 7704
rect 18196 7692 18202 7744
rect 1104 7642 19019 7664
rect 1104 7590 5388 7642
rect 5440 7590 5452 7642
rect 5504 7590 5516 7642
rect 5568 7590 5580 7642
rect 5632 7590 5644 7642
rect 5696 7590 9827 7642
rect 9879 7590 9891 7642
rect 9943 7590 9955 7642
rect 10007 7590 10019 7642
rect 10071 7590 10083 7642
rect 10135 7590 14266 7642
rect 14318 7590 14330 7642
rect 14382 7590 14394 7642
rect 14446 7590 14458 7642
rect 14510 7590 14522 7642
rect 14574 7590 18705 7642
rect 18757 7590 18769 7642
rect 18821 7590 18833 7642
rect 18885 7590 18897 7642
rect 18949 7590 18961 7642
rect 19013 7590 19019 7642
rect 1104 7568 19019 7590
rect 3418 7528 3424 7540
rect 3379 7500 3424 7528
rect 3418 7488 3424 7500
rect 3476 7488 3482 7540
rect 4890 7528 4896 7540
rect 4851 7500 4896 7528
rect 4890 7488 4896 7500
rect 4948 7488 4954 7540
rect 5997 7531 6055 7537
rect 5997 7497 6009 7531
rect 6043 7528 6055 7531
rect 6822 7528 6828 7540
rect 6043 7500 6828 7528
rect 6043 7497 6055 7500
rect 5997 7491 6055 7497
rect 6822 7488 6828 7500
rect 6880 7488 6886 7540
rect 7009 7531 7067 7537
rect 7009 7497 7021 7531
rect 7055 7528 7067 7531
rect 7466 7528 7472 7540
rect 7055 7500 7472 7528
rect 7055 7497 7067 7500
rect 7009 7491 7067 7497
rect 7466 7488 7472 7500
rect 7524 7488 7530 7540
rect 7558 7488 7564 7540
rect 7616 7528 7622 7540
rect 7616 7500 10548 7528
rect 7616 7488 7622 7500
rect 2608 7432 3832 7460
rect 2608 7401 2636 7432
rect 3804 7401 3832 7432
rect 3970 7420 3976 7472
rect 4028 7460 4034 7472
rect 4709 7463 4767 7469
rect 4709 7460 4721 7463
rect 4028 7432 4721 7460
rect 4028 7420 4034 7432
rect 4709 7429 4721 7432
rect 4755 7429 4767 7463
rect 4709 7423 4767 7429
rect 5074 7420 5080 7472
rect 5132 7460 5138 7472
rect 6730 7460 6736 7472
rect 5132 7432 6736 7460
rect 5132 7420 5138 7432
rect 6730 7420 6736 7432
rect 6788 7420 6794 7472
rect 6914 7420 6920 7472
rect 6972 7460 6978 7472
rect 6972 7432 8340 7460
rect 6972 7420 6978 7432
rect 2593 7395 2651 7401
rect 2593 7361 2605 7395
rect 2639 7361 2651 7395
rect 3605 7395 3663 7401
rect 3605 7392 3617 7395
rect 2593 7355 2651 7361
rect 2792 7364 3617 7392
rect 2792 7336 2820 7364
rect 3605 7361 3617 7364
rect 3651 7361 3663 7395
rect 3605 7355 3663 7361
rect 3789 7395 3847 7401
rect 3789 7361 3801 7395
rect 3835 7392 3847 7395
rect 4430 7392 4436 7404
rect 3835 7364 4436 7392
rect 3835 7361 3847 7364
rect 3789 7355 3847 7361
rect 4430 7352 4436 7364
rect 4488 7352 4494 7404
rect 4525 7395 4583 7401
rect 4525 7361 4537 7395
rect 4571 7361 4583 7395
rect 4525 7355 4583 7361
rect 5813 7395 5871 7401
rect 5813 7361 5825 7395
rect 5859 7392 5871 7395
rect 5902 7392 5908 7404
rect 5859 7364 5908 7392
rect 5859 7361 5871 7364
rect 5813 7355 5871 7361
rect 2685 7327 2743 7333
rect 2685 7293 2697 7327
rect 2731 7324 2743 7327
rect 2774 7324 2780 7336
rect 2731 7296 2780 7324
rect 2731 7293 2743 7296
rect 2685 7287 2743 7293
rect 2774 7284 2780 7296
rect 2832 7324 2838 7336
rect 2961 7327 3019 7333
rect 2832 7296 2925 7324
rect 2832 7284 2838 7296
rect 2961 7293 2973 7327
rect 3007 7324 3019 7327
rect 3050 7324 3056 7336
rect 3007 7296 3056 7324
rect 3007 7293 3019 7296
rect 2961 7287 3019 7293
rect 3050 7284 3056 7296
rect 3108 7284 3114 7336
rect 4154 7284 4160 7336
rect 4212 7324 4218 7336
rect 4540 7324 4568 7355
rect 5902 7352 5908 7364
rect 5960 7352 5966 7404
rect 5994 7352 6000 7404
rect 6052 7392 6058 7404
rect 7009 7395 7067 7401
rect 6052 7364 6097 7392
rect 6052 7352 6058 7364
rect 7009 7361 7021 7395
rect 7055 7392 7067 7395
rect 7282 7392 7288 7404
rect 7055 7364 7288 7392
rect 7055 7361 7067 7364
rect 7009 7355 7067 7361
rect 7282 7352 7288 7364
rect 7340 7352 7346 7404
rect 8312 7401 8340 7432
rect 7837 7395 7895 7401
rect 7837 7361 7849 7395
rect 7883 7392 7895 7395
rect 8297 7395 8355 7401
rect 7883 7364 8248 7392
rect 7883 7361 7895 7364
rect 7837 7355 7895 7361
rect 4212 7296 4568 7324
rect 4212 7284 4218 7296
rect 6546 7284 6552 7336
rect 6604 7324 6610 7336
rect 6604 7296 7512 7324
rect 6604 7284 6610 7296
rect 7484 7265 7512 7296
rect 8018 7284 8024 7336
rect 8076 7284 8082 7336
rect 6917 7259 6975 7265
rect 6917 7225 6929 7259
rect 6963 7225 6975 7259
rect 6917 7219 6975 7225
rect 7469 7259 7527 7265
rect 7469 7225 7481 7259
rect 7515 7225 7527 7259
rect 7469 7219 7527 7225
rect 8220 7256 8248 7364
rect 8297 7361 8309 7395
rect 8343 7361 8355 7395
rect 8297 7355 8355 7361
rect 9401 7395 9459 7401
rect 9401 7361 9413 7395
rect 9447 7392 9459 7395
rect 9490 7392 9496 7404
rect 9447 7364 9496 7392
rect 9447 7361 9459 7364
rect 9401 7355 9459 7361
rect 9490 7352 9496 7364
rect 9548 7352 9554 7404
rect 9674 7392 9680 7404
rect 9635 7364 9680 7392
rect 9674 7352 9680 7364
rect 9732 7352 9738 7404
rect 8478 7324 8484 7336
rect 8439 7296 8484 7324
rect 8478 7284 8484 7296
rect 8536 7284 8542 7336
rect 10520 7333 10548 7500
rect 12158 7488 12164 7540
rect 12216 7528 12222 7540
rect 13081 7531 13139 7537
rect 13081 7528 13093 7531
rect 12216 7500 13093 7528
rect 12216 7488 12222 7500
rect 13081 7497 13093 7500
rect 13127 7528 13139 7531
rect 15838 7528 15844 7540
rect 13127 7500 15844 7528
rect 13127 7497 13139 7500
rect 13081 7491 13139 7497
rect 15838 7488 15844 7500
rect 15896 7488 15902 7540
rect 16022 7528 16028 7540
rect 15983 7500 16028 7528
rect 16022 7488 16028 7500
rect 16080 7488 16086 7540
rect 17218 7528 17224 7540
rect 17179 7500 17224 7528
rect 17218 7488 17224 7500
rect 17276 7488 17282 7540
rect 11057 7463 11115 7469
rect 11057 7429 11069 7463
rect 11103 7460 11115 7463
rect 11946 7463 12004 7469
rect 11946 7460 11958 7463
rect 11103 7432 11958 7460
rect 11103 7429 11115 7432
rect 11057 7423 11115 7429
rect 11946 7429 11958 7432
rect 11992 7429 12004 7463
rect 11946 7423 12004 7429
rect 14737 7463 14795 7469
rect 14737 7429 14749 7463
rect 14783 7460 14795 7463
rect 17681 7463 17739 7469
rect 14783 7432 16712 7460
rect 14783 7429 14795 7432
rect 14737 7423 14795 7429
rect 10965 7395 11023 7401
rect 10965 7361 10977 7395
rect 11011 7361 11023 7395
rect 11146 7392 11152 7404
rect 11107 7364 11152 7392
rect 10965 7355 11023 7361
rect 10505 7327 10563 7333
rect 10505 7293 10517 7327
rect 10551 7324 10563 7327
rect 10980 7324 11008 7355
rect 11146 7352 11152 7364
rect 11204 7352 11210 7404
rect 13538 7392 13544 7404
rect 13499 7364 13544 7392
rect 13538 7352 13544 7364
rect 13596 7352 13602 7404
rect 13814 7352 13820 7404
rect 13872 7392 13878 7404
rect 14645 7395 14703 7401
rect 14645 7392 14657 7395
rect 13872 7364 14657 7392
rect 13872 7352 13878 7364
rect 14645 7361 14657 7364
rect 14691 7361 14703 7395
rect 14645 7355 14703 7361
rect 14921 7395 14979 7401
rect 14921 7361 14933 7395
rect 14967 7392 14979 7395
rect 15749 7395 15807 7401
rect 15749 7392 15761 7395
rect 14967 7364 15761 7392
rect 14967 7361 14979 7364
rect 14921 7355 14979 7361
rect 15749 7361 15761 7364
rect 15795 7392 15807 7395
rect 16114 7392 16120 7404
rect 15795 7364 16120 7392
rect 15795 7361 15807 7364
rect 15749 7355 15807 7361
rect 16114 7352 16120 7364
rect 16172 7352 16178 7404
rect 11606 7324 11612 7336
rect 10551 7296 11612 7324
rect 10551 7293 10563 7296
rect 10505 7287 10563 7293
rect 11606 7284 11612 7296
rect 11664 7284 11670 7336
rect 11701 7327 11759 7333
rect 11701 7293 11713 7327
rect 11747 7293 11759 7327
rect 11701 7287 11759 7293
rect 9030 7256 9036 7268
rect 8220 7228 9036 7256
rect 6932 7188 6960 7219
rect 7926 7188 7932 7200
rect 6932 7160 7932 7188
rect 7926 7148 7932 7160
rect 7984 7148 7990 7200
rect 8110 7148 8116 7200
rect 8168 7188 8174 7200
rect 8220 7188 8248 7228
rect 9030 7216 9036 7228
rect 9088 7216 9094 7268
rect 9674 7216 9680 7268
rect 9732 7256 9738 7268
rect 11716 7256 11744 7287
rect 15194 7284 15200 7336
rect 15252 7324 15258 7336
rect 15381 7327 15439 7333
rect 15381 7324 15393 7327
rect 15252 7296 15393 7324
rect 15252 7284 15258 7296
rect 15381 7293 15393 7296
rect 15427 7293 15439 7327
rect 15381 7287 15439 7293
rect 15657 7327 15715 7333
rect 15657 7293 15669 7327
rect 15703 7293 15715 7327
rect 15657 7287 15715 7293
rect 9732 7228 11744 7256
rect 15672 7256 15700 7287
rect 15838 7284 15844 7336
rect 15896 7333 15902 7336
rect 15896 7327 15924 7333
rect 15912 7293 15924 7327
rect 16684 7324 16712 7432
rect 17681 7429 17693 7463
rect 17727 7460 17739 7463
rect 18046 7460 18052 7472
rect 17727 7432 18052 7460
rect 17727 7429 17739 7432
rect 17681 7423 17739 7429
rect 18046 7420 18052 7432
rect 18104 7420 18110 7472
rect 17589 7395 17647 7401
rect 17589 7361 17601 7395
rect 17635 7392 17647 7395
rect 17954 7392 17960 7404
rect 17635 7364 17960 7392
rect 17635 7361 17647 7364
rect 17589 7355 17647 7361
rect 17954 7352 17960 7364
rect 18012 7352 18018 7404
rect 17402 7324 17408 7336
rect 16684 7296 17408 7324
rect 15896 7287 15924 7293
rect 15896 7284 15902 7287
rect 17402 7284 17408 7296
rect 17460 7324 17466 7336
rect 17773 7327 17831 7333
rect 17773 7324 17785 7327
rect 17460 7296 17785 7324
rect 17460 7284 17466 7296
rect 17773 7293 17785 7296
rect 17819 7293 17831 7327
rect 17773 7287 17831 7293
rect 18230 7256 18236 7268
rect 15672 7228 18236 7256
rect 9732 7216 9738 7228
rect 18230 7216 18236 7228
rect 18288 7216 18294 7268
rect 8168 7160 8248 7188
rect 8168 7148 8174 7160
rect 8662 7148 8668 7200
rect 8720 7188 8726 7200
rect 9493 7191 9551 7197
rect 9493 7188 9505 7191
rect 8720 7160 9505 7188
rect 8720 7148 8726 7160
rect 9493 7157 9505 7160
rect 9539 7157 9551 7191
rect 9858 7188 9864 7200
rect 9819 7160 9864 7188
rect 9493 7151 9551 7157
rect 9858 7148 9864 7160
rect 9916 7148 9922 7200
rect 13722 7188 13728 7200
rect 13683 7160 13728 7188
rect 13722 7148 13728 7160
rect 13780 7148 13786 7200
rect 13814 7148 13820 7200
rect 13872 7188 13878 7200
rect 14921 7191 14979 7197
rect 14921 7188 14933 7191
rect 13872 7160 14933 7188
rect 13872 7148 13878 7160
rect 14921 7157 14933 7160
rect 14967 7157 14979 7191
rect 14921 7151 14979 7157
rect 17586 7148 17592 7200
rect 17644 7188 17650 7200
rect 17862 7188 17868 7200
rect 17644 7160 17868 7188
rect 17644 7148 17650 7160
rect 17862 7148 17868 7160
rect 17920 7148 17926 7200
rect 1104 7098 18860 7120
rect 1104 7046 3169 7098
rect 3221 7046 3233 7098
rect 3285 7046 3297 7098
rect 3349 7046 3361 7098
rect 3413 7046 3425 7098
rect 3477 7046 7608 7098
rect 7660 7046 7672 7098
rect 7724 7046 7736 7098
rect 7788 7046 7800 7098
rect 7852 7046 7864 7098
rect 7916 7046 12047 7098
rect 12099 7046 12111 7098
rect 12163 7046 12175 7098
rect 12227 7046 12239 7098
rect 12291 7046 12303 7098
rect 12355 7046 16486 7098
rect 16538 7046 16550 7098
rect 16602 7046 16614 7098
rect 16666 7046 16678 7098
rect 16730 7046 16742 7098
rect 16794 7046 18860 7098
rect 1104 7024 18860 7046
rect 8386 6984 8392 6996
rect 8347 6956 8392 6984
rect 8386 6944 8392 6956
rect 8444 6944 8450 6996
rect 16114 6984 16120 6996
rect 16075 6956 16120 6984
rect 16114 6944 16120 6956
rect 16172 6944 16178 6996
rect 17218 6984 17224 6996
rect 17179 6956 17224 6984
rect 17218 6944 17224 6956
rect 17276 6944 17282 6996
rect 17865 6987 17923 6993
rect 17865 6953 17877 6987
rect 17911 6984 17923 6987
rect 17954 6984 17960 6996
rect 17911 6956 17960 6984
rect 17911 6953 17923 6956
rect 17865 6947 17923 6953
rect 17954 6944 17960 6956
rect 18012 6944 18018 6996
rect 3973 6919 4031 6925
rect 3973 6916 3985 6919
rect 3160 6888 3985 6916
rect 2869 6851 2927 6857
rect 2869 6848 2881 6851
rect 2424 6820 2881 6848
rect 2222 6780 2228 6792
rect 2183 6752 2228 6780
rect 2222 6740 2228 6752
rect 2280 6740 2286 6792
rect 2424 6789 2452 6820
rect 2869 6817 2881 6820
rect 2915 6817 2927 6851
rect 2869 6811 2927 6817
rect 2958 6808 2964 6860
rect 3016 6848 3022 6860
rect 3160 6857 3188 6888
rect 3973 6885 3985 6888
rect 4019 6885 4031 6919
rect 3973 6879 4031 6885
rect 3145 6851 3203 6857
rect 3145 6848 3157 6851
rect 3016 6820 3157 6848
rect 3016 6808 3022 6820
rect 3145 6817 3157 6820
rect 3191 6817 3203 6851
rect 3145 6811 3203 6817
rect 3329 6851 3387 6857
rect 3329 6817 3341 6851
rect 3375 6848 3387 6851
rect 3694 6848 3700 6860
rect 3375 6820 3700 6848
rect 3375 6817 3387 6820
rect 3329 6811 3387 6817
rect 3694 6808 3700 6820
rect 3752 6808 3758 6860
rect 13633 6851 13691 6857
rect 13633 6817 13645 6851
rect 13679 6848 13691 6851
rect 13814 6848 13820 6860
rect 13679 6820 13820 6848
rect 13679 6817 13691 6820
rect 13633 6811 13691 6817
rect 13814 6808 13820 6820
rect 13872 6808 13878 6860
rect 13998 6808 14004 6860
rect 14056 6848 14062 6860
rect 14277 6851 14335 6857
rect 14277 6848 14289 6851
rect 14056 6820 14289 6848
rect 14056 6808 14062 6820
rect 14277 6817 14289 6820
rect 14323 6817 14335 6851
rect 16022 6848 16028 6860
rect 14277 6811 14335 6817
rect 15304 6820 16028 6848
rect 2409 6783 2467 6789
rect 2409 6749 2421 6783
rect 2455 6749 2467 6783
rect 2409 6743 2467 6749
rect 2774 6740 2780 6792
rect 2832 6780 2838 6792
rect 3050 6780 3056 6792
rect 2832 6752 3056 6780
rect 2832 6740 2838 6752
rect 3050 6740 3056 6752
rect 3108 6740 3114 6792
rect 3234 6780 3240 6792
rect 3195 6752 3240 6780
rect 3234 6740 3240 6752
rect 3292 6740 3298 6792
rect 4614 6740 4620 6792
rect 4672 6780 4678 6792
rect 6546 6789 6552 6792
rect 5353 6783 5411 6789
rect 5353 6780 5365 6783
rect 4672 6752 5365 6780
rect 4672 6740 4678 6752
rect 5353 6749 5365 6752
rect 5399 6780 5411 6783
rect 6273 6783 6331 6789
rect 6273 6780 6285 6783
rect 5399 6752 6285 6780
rect 5399 6749 5411 6752
rect 5353 6743 5411 6749
rect 6273 6749 6285 6752
rect 6319 6749 6331 6783
rect 6540 6780 6552 6789
rect 6507 6752 6552 6780
rect 6273 6743 6331 6749
rect 6540 6743 6552 6752
rect 6546 6740 6552 6743
rect 6604 6740 6610 6792
rect 9122 6780 9128 6792
rect 8128 6752 8984 6780
rect 9083 6752 9128 6780
rect 2317 6715 2375 6721
rect 2317 6681 2329 6715
rect 2363 6712 2375 6715
rect 5086 6715 5144 6721
rect 5086 6712 5098 6715
rect 2363 6684 5098 6712
rect 2363 6681 2375 6684
rect 2317 6675 2375 6681
rect 5086 6681 5098 6684
rect 5132 6681 5144 6715
rect 5086 6675 5144 6681
rect 6086 6672 6092 6724
rect 6144 6712 6150 6724
rect 8128 6712 8156 6752
rect 6144 6684 8156 6712
rect 8205 6715 8263 6721
rect 6144 6672 6150 6684
rect 8205 6681 8217 6715
rect 8251 6712 8263 6715
rect 8294 6712 8300 6724
rect 8251 6684 8300 6712
rect 8251 6681 8263 6684
rect 8205 6675 8263 6681
rect 8294 6672 8300 6684
rect 8352 6672 8358 6724
rect 8421 6715 8479 6721
rect 8421 6681 8433 6715
rect 8467 6712 8479 6715
rect 8754 6712 8760 6724
rect 8467 6684 8760 6712
rect 8467 6681 8479 6684
rect 8421 6675 8479 6681
rect 8754 6672 8760 6684
rect 8812 6672 8818 6724
rect 8956 6712 8984 6752
rect 9122 6740 9128 6752
rect 9180 6740 9186 6792
rect 9674 6740 9680 6792
rect 9732 6780 9738 6792
rect 9769 6783 9827 6789
rect 9769 6780 9781 6783
rect 9732 6752 9781 6780
rect 9732 6740 9738 6752
rect 9769 6749 9781 6752
rect 9815 6749 9827 6783
rect 9769 6743 9827 6749
rect 9858 6740 9864 6792
rect 9916 6780 9922 6792
rect 10025 6783 10083 6789
rect 10025 6780 10037 6783
rect 9916 6752 10037 6780
rect 9916 6740 9922 6752
rect 10025 6749 10037 6752
rect 10071 6749 10083 6783
rect 11885 6783 11943 6789
rect 11885 6780 11897 6783
rect 10025 6743 10083 6749
rect 10704 6752 11897 6780
rect 10704 6724 10732 6752
rect 11885 6749 11897 6752
rect 11931 6749 11943 6783
rect 11885 6743 11943 6749
rect 12437 6783 12495 6789
rect 12437 6749 12449 6783
rect 12483 6749 12495 6783
rect 12437 6743 12495 6749
rect 12897 6783 12955 6789
rect 12897 6749 12909 6783
rect 12943 6780 12955 6783
rect 13538 6780 13544 6792
rect 12943 6752 13544 6780
rect 12943 6749 12955 6752
rect 12897 6743 12955 6749
rect 10318 6712 10324 6724
rect 8956 6684 10324 6712
rect 10318 6672 10324 6684
rect 10376 6672 10382 6724
rect 10686 6672 10692 6724
rect 10744 6672 10750 6724
rect 12452 6712 12480 6743
rect 13538 6740 13544 6752
rect 13596 6740 13602 6792
rect 13725 6783 13783 6789
rect 13725 6749 13737 6783
rect 13771 6780 13783 6783
rect 15304 6780 15332 6820
rect 16022 6808 16028 6820
rect 16080 6808 16086 6860
rect 18141 6851 18199 6857
rect 18141 6848 18153 6851
rect 17236 6820 18153 6848
rect 13771 6752 15332 6780
rect 13771 6749 13783 6752
rect 13725 6743 13783 6749
rect 15930 6740 15936 6792
rect 15988 6780 15994 6792
rect 16301 6783 16359 6789
rect 16301 6780 16313 6783
rect 15988 6752 16313 6780
rect 15988 6740 15994 6752
rect 16301 6749 16313 6752
rect 16347 6749 16359 6783
rect 16301 6743 16359 6749
rect 16390 6740 16396 6792
rect 16448 6780 16454 6792
rect 16448 6752 16493 6780
rect 16448 6740 16454 6752
rect 17126 6740 17132 6792
rect 17184 6780 17190 6792
rect 17236 6789 17264 6820
rect 18141 6817 18153 6820
rect 18187 6817 18199 6851
rect 18141 6811 18199 6817
rect 17221 6783 17279 6789
rect 17221 6780 17233 6783
rect 17184 6752 17233 6780
rect 17184 6740 17190 6752
rect 17221 6749 17233 6752
rect 17267 6749 17279 6783
rect 17221 6743 17279 6749
rect 17405 6783 17463 6789
rect 17405 6749 17417 6783
rect 17451 6780 17463 6783
rect 17865 6783 17923 6789
rect 17865 6780 17877 6783
rect 17451 6752 17877 6780
rect 17451 6749 17463 6752
rect 17405 6743 17463 6749
rect 17865 6749 17877 6752
rect 17911 6749 17923 6783
rect 17865 6743 17923 6749
rect 17957 6783 18015 6789
rect 17957 6749 17969 6783
rect 18003 6749 18015 6783
rect 17957 6743 18015 6749
rect 13446 6712 13452 6724
rect 11164 6684 12480 6712
rect 13407 6684 13452 6712
rect 1765 6647 1823 6653
rect 1765 6613 1777 6647
rect 1811 6644 1823 6647
rect 3694 6644 3700 6656
rect 1811 6616 3700 6644
rect 1811 6613 1823 6616
rect 1765 6607 1823 6613
rect 3694 6604 3700 6616
rect 3752 6604 3758 6656
rect 7650 6644 7656 6656
rect 7611 6616 7656 6644
rect 7650 6604 7656 6616
rect 7708 6604 7714 6656
rect 8573 6647 8631 6653
rect 8573 6613 8585 6647
rect 8619 6644 8631 6647
rect 8662 6644 8668 6656
rect 8619 6616 8668 6644
rect 8619 6613 8631 6616
rect 8573 6607 8631 6613
rect 8662 6604 8668 6616
rect 8720 6604 8726 6656
rect 9217 6647 9275 6653
rect 9217 6613 9229 6647
rect 9263 6644 9275 6647
rect 9398 6644 9404 6656
rect 9263 6616 9404 6644
rect 9263 6613 9275 6616
rect 9217 6607 9275 6613
rect 9398 6604 9404 6616
rect 9456 6604 9462 6656
rect 11164 6653 11192 6684
rect 13446 6672 13452 6684
rect 13504 6672 13510 6724
rect 14522 6715 14580 6721
rect 14522 6712 14534 6715
rect 13740 6684 14534 6712
rect 11149 6647 11207 6653
rect 11149 6613 11161 6647
rect 11195 6613 11207 6647
rect 11149 6607 11207 6613
rect 12897 6647 12955 6653
rect 12897 6613 12909 6647
rect 12943 6644 12955 6647
rect 13078 6644 13084 6656
rect 12943 6616 13084 6644
rect 12943 6613 12955 6616
rect 12897 6607 12955 6613
rect 13078 6604 13084 6616
rect 13136 6604 13142 6656
rect 13740 6653 13768 6684
rect 14522 6681 14534 6684
rect 14568 6681 14580 6715
rect 14522 6675 14580 6681
rect 14642 6672 14648 6724
rect 14700 6712 14706 6724
rect 16117 6715 16175 6721
rect 16117 6712 16129 6715
rect 14700 6684 16129 6712
rect 14700 6672 14706 6684
rect 16117 6681 16129 6684
rect 16163 6681 16175 6715
rect 17420 6712 17448 6743
rect 17972 6712 18000 6743
rect 16117 6675 16175 6681
rect 16592 6684 17448 6712
rect 17880 6684 18000 6712
rect 13725 6647 13783 6653
rect 13725 6613 13737 6647
rect 13771 6613 13783 6647
rect 15654 6644 15660 6656
rect 15615 6616 15660 6644
rect 13725 6607 13783 6613
rect 15654 6604 15660 6616
rect 15712 6604 15718 6656
rect 16592 6653 16620 6684
rect 16577 6647 16635 6653
rect 16577 6613 16589 6647
rect 16623 6613 16635 6647
rect 17034 6644 17040 6656
rect 16995 6616 17040 6644
rect 16577 6607 16635 6613
rect 17034 6604 17040 6616
rect 17092 6604 17098 6656
rect 17218 6604 17224 6656
rect 17276 6644 17282 6656
rect 17880 6644 17908 6684
rect 17276 6616 17908 6644
rect 17276 6604 17282 6616
rect 1104 6554 19019 6576
rect 1104 6502 5388 6554
rect 5440 6502 5452 6554
rect 5504 6502 5516 6554
rect 5568 6502 5580 6554
rect 5632 6502 5644 6554
rect 5696 6502 9827 6554
rect 9879 6502 9891 6554
rect 9943 6502 9955 6554
rect 10007 6502 10019 6554
rect 10071 6502 10083 6554
rect 10135 6502 14266 6554
rect 14318 6502 14330 6554
rect 14382 6502 14394 6554
rect 14446 6502 14458 6554
rect 14510 6502 14522 6554
rect 14574 6502 18705 6554
rect 18757 6502 18769 6554
rect 18821 6502 18833 6554
rect 18885 6502 18897 6554
rect 18949 6502 18961 6554
rect 19013 6502 19019 6554
rect 1104 6480 19019 6502
rect 2958 6440 2964 6452
rect 2792 6412 2964 6440
rect 2792 6381 2820 6412
rect 2958 6400 2964 6412
rect 3016 6400 3022 6452
rect 7190 6400 7196 6452
rect 7248 6440 7254 6452
rect 10502 6440 10508 6452
rect 7248 6412 10508 6440
rect 7248 6400 7254 6412
rect 10502 6400 10508 6412
rect 10560 6440 10566 6452
rect 10965 6443 11023 6449
rect 10965 6440 10977 6443
rect 10560 6412 10977 6440
rect 10560 6400 10566 6412
rect 10965 6409 10977 6412
rect 11011 6409 11023 6443
rect 10965 6403 11023 6409
rect 11793 6443 11851 6449
rect 11793 6409 11805 6443
rect 11839 6440 11851 6443
rect 12713 6443 12771 6449
rect 12713 6440 12725 6443
rect 11839 6412 12725 6440
rect 11839 6409 11851 6412
rect 11793 6403 11851 6409
rect 12713 6409 12725 6412
rect 12759 6409 12771 6443
rect 12713 6403 12771 6409
rect 15473 6443 15531 6449
rect 15473 6409 15485 6443
rect 15519 6440 15531 6443
rect 16114 6440 16120 6452
rect 15519 6412 16120 6440
rect 15519 6409 15531 6412
rect 15473 6403 15531 6409
rect 16114 6400 16120 6412
rect 16172 6400 16178 6452
rect 17037 6443 17095 6449
rect 17037 6409 17049 6443
rect 17083 6440 17095 6443
rect 17770 6440 17776 6452
rect 17083 6412 17776 6440
rect 17083 6409 17095 6412
rect 17037 6403 17095 6409
rect 17770 6400 17776 6412
rect 17828 6400 17834 6452
rect 18046 6440 18052 6452
rect 18007 6412 18052 6440
rect 18046 6400 18052 6412
rect 18104 6400 18110 6452
rect 2777 6375 2835 6381
rect 2777 6341 2789 6375
rect 2823 6341 2835 6375
rect 5074 6372 5080 6384
rect 2777 6335 2835 6341
rect 4172 6344 5080 6372
rect 2961 6307 3019 6313
rect 2961 6273 2973 6307
rect 3007 6273 3019 6307
rect 2961 6267 3019 6273
rect 2866 6196 2872 6248
rect 2924 6236 2930 6248
rect 2976 6236 3004 6267
rect 3050 6264 3056 6316
rect 3108 6304 3114 6316
rect 3970 6304 3976 6316
rect 3108 6276 3153 6304
rect 3931 6276 3976 6304
rect 3108 6264 3114 6276
rect 3970 6264 3976 6276
rect 4028 6264 4034 6316
rect 4172 6313 4200 6344
rect 5074 6332 5080 6344
rect 5132 6332 5138 6384
rect 7837 6375 7895 6381
rect 7837 6341 7849 6375
rect 7883 6372 7895 6375
rect 8018 6372 8024 6384
rect 7883 6344 8024 6372
rect 7883 6341 7895 6344
rect 7837 6335 7895 6341
rect 8018 6332 8024 6344
rect 8076 6332 8082 6384
rect 8386 6332 8392 6384
rect 8444 6332 8450 6384
rect 9030 6332 9036 6384
rect 9088 6372 9094 6384
rect 10045 6375 10103 6381
rect 10045 6372 10057 6375
rect 9088 6344 10057 6372
rect 9088 6332 9094 6344
rect 10045 6341 10057 6344
rect 10091 6341 10103 6375
rect 10045 6335 10103 6341
rect 10413 6375 10471 6381
rect 10413 6341 10425 6375
rect 10459 6372 10471 6375
rect 10686 6372 10692 6384
rect 10459 6344 10692 6372
rect 10459 6341 10471 6344
rect 10413 6335 10471 6341
rect 4157 6307 4215 6313
rect 4157 6273 4169 6307
rect 4203 6273 4215 6307
rect 4614 6304 4620 6316
rect 4575 6276 4620 6304
rect 4157 6267 4215 6273
rect 4614 6264 4620 6276
rect 4672 6264 4678 6316
rect 4884 6307 4942 6313
rect 4884 6273 4896 6307
rect 4930 6304 4942 6307
rect 5166 6304 5172 6316
rect 4930 6276 5172 6304
rect 4930 6273 4942 6276
rect 4884 6267 4942 6273
rect 5166 6264 5172 6276
rect 5224 6264 5230 6316
rect 6730 6304 6736 6316
rect 6691 6276 6736 6304
rect 6730 6264 6736 6276
rect 6788 6264 6794 6316
rect 7650 6304 7656 6316
rect 7611 6276 7656 6304
rect 7650 6264 7656 6276
rect 7708 6264 7714 6316
rect 8113 6307 8171 6313
rect 8113 6273 8125 6307
rect 8159 6304 8171 6307
rect 8202 6304 8208 6316
rect 8159 6276 8208 6304
rect 8159 6273 8171 6276
rect 8113 6267 8171 6273
rect 8202 6264 8208 6276
rect 8260 6264 8266 6316
rect 8297 6307 8355 6313
rect 8297 6273 8309 6307
rect 8343 6304 8355 6307
rect 8404 6304 8432 6332
rect 9217 6307 9275 6313
rect 9217 6304 9229 6307
rect 8343 6276 9229 6304
rect 8343 6273 8355 6276
rect 8297 6267 8355 6273
rect 9217 6273 9229 6276
rect 9263 6273 9275 6307
rect 9398 6304 9404 6316
rect 9359 6276 9404 6304
rect 9217 6267 9275 6273
rect 9398 6264 9404 6276
rect 9456 6264 9462 6316
rect 10060 6304 10088 6335
rect 10686 6332 10692 6344
rect 10744 6332 10750 6384
rect 17218 6372 17224 6384
rect 16868 6344 17224 6372
rect 16868 6316 16896 6344
rect 17218 6332 17224 6344
rect 17276 6372 17282 6384
rect 17681 6375 17739 6381
rect 17681 6372 17693 6375
rect 17276 6344 17693 6372
rect 17276 6332 17282 6344
rect 17681 6341 17693 6344
rect 17727 6341 17739 6375
rect 17681 6335 17739 6341
rect 10873 6307 10931 6313
rect 10873 6304 10885 6307
rect 10060 6276 10885 6304
rect 10873 6273 10885 6276
rect 10919 6273 10931 6307
rect 11698 6304 11704 6316
rect 11659 6276 11704 6304
rect 10873 6267 10931 6273
rect 11698 6264 11704 6276
rect 11756 6264 11762 6316
rect 11882 6264 11888 6316
rect 11940 6304 11946 6316
rect 11977 6307 12035 6313
rect 11977 6304 11989 6307
rect 11940 6276 11989 6304
rect 11940 6264 11946 6276
rect 11977 6273 11989 6276
rect 12023 6273 12035 6307
rect 11977 6267 12035 6273
rect 12713 6307 12771 6313
rect 12713 6273 12725 6307
rect 12759 6304 12771 6307
rect 12802 6304 12808 6316
rect 12759 6276 12808 6304
rect 12759 6273 12771 6276
rect 12713 6267 12771 6273
rect 12802 6264 12808 6276
rect 12860 6264 12866 6316
rect 12897 6307 12955 6313
rect 12897 6273 12909 6307
rect 12943 6304 12955 6307
rect 13262 6304 13268 6316
rect 12943 6276 13268 6304
rect 12943 6273 12955 6276
rect 12897 6267 12955 6273
rect 13262 6264 13268 6276
rect 13320 6264 13326 6316
rect 16850 6304 16856 6316
rect 16811 6276 16856 6304
rect 16850 6264 16856 6276
rect 16908 6264 16914 6316
rect 17034 6304 17040 6316
rect 16995 6276 17040 6304
rect 17034 6264 17040 6276
rect 17092 6304 17098 6316
rect 17497 6307 17555 6313
rect 17497 6304 17509 6307
rect 17092 6276 17509 6304
rect 17092 6264 17098 6276
rect 17497 6273 17509 6276
rect 17543 6273 17555 6307
rect 17497 6267 17555 6273
rect 17773 6307 17831 6313
rect 17773 6273 17785 6307
rect 17819 6273 17831 6307
rect 17773 6267 17831 6273
rect 3234 6236 3240 6248
rect 2924 6208 3240 6236
rect 2924 6196 2930 6208
rect 3234 6196 3240 6208
rect 3292 6236 3298 6248
rect 3988 6236 4016 6264
rect 3292 6208 4016 6236
rect 3292 6196 3298 6208
rect 2222 6128 2228 6180
rect 2280 6168 2286 6180
rect 2777 6171 2835 6177
rect 2777 6168 2789 6171
rect 2280 6140 2789 6168
rect 2280 6128 2286 6140
rect 2777 6137 2789 6140
rect 2823 6137 2835 6171
rect 2777 6131 2835 6137
rect 5997 6171 6055 6177
rect 5997 6137 6009 6171
rect 6043 6168 6055 6171
rect 6914 6168 6920 6180
rect 6043 6140 6920 6168
rect 6043 6137 6055 6140
rect 5997 6131 6055 6137
rect 6914 6128 6920 6140
rect 6972 6128 6978 6180
rect 8220 6168 8248 6264
rect 8481 6239 8539 6245
rect 8481 6205 8493 6239
rect 8527 6236 8539 6239
rect 8754 6236 8760 6248
rect 8527 6208 8760 6236
rect 8527 6205 8539 6208
rect 8481 6199 8539 6205
rect 8754 6196 8760 6208
rect 8812 6236 8818 6248
rect 9125 6239 9183 6245
rect 9125 6236 9137 6239
rect 8812 6208 9137 6236
rect 8812 6196 8818 6208
rect 9125 6205 9137 6208
rect 9171 6205 9183 6239
rect 9125 6199 9183 6205
rect 9309 6239 9367 6245
rect 9309 6205 9321 6239
rect 9355 6205 9367 6239
rect 9309 6199 9367 6205
rect 9324 6168 9352 6199
rect 10318 6196 10324 6248
rect 10376 6236 10382 6248
rect 13446 6236 13452 6248
rect 10376 6208 13452 6236
rect 10376 6196 10382 6208
rect 13446 6196 13452 6208
rect 13504 6196 13510 6248
rect 13538 6196 13544 6248
rect 13596 6236 13602 6248
rect 15013 6239 15071 6245
rect 15013 6236 15025 6239
rect 13596 6208 15025 6236
rect 13596 6196 13602 6208
rect 15013 6205 15025 6208
rect 15059 6236 15071 6239
rect 15746 6236 15752 6248
rect 15059 6208 15752 6236
rect 15059 6205 15071 6208
rect 15013 6199 15071 6205
rect 15746 6196 15752 6208
rect 15804 6196 15810 6248
rect 16942 6196 16948 6248
rect 17000 6236 17006 6248
rect 17788 6236 17816 6267
rect 17862 6264 17868 6316
rect 17920 6304 17926 6316
rect 17920 6276 17965 6304
rect 17920 6264 17926 6276
rect 17000 6208 17816 6236
rect 17000 6196 17006 6208
rect 8220 6140 9352 6168
rect 11422 6128 11428 6180
rect 11480 6168 11486 6180
rect 13722 6168 13728 6180
rect 11480 6140 13728 6168
rect 11480 6128 11486 6140
rect 13722 6128 13728 6140
rect 13780 6128 13786 6180
rect 15381 6171 15439 6177
rect 15381 6137 15393 6171
rect 15427 6168 15439 6171
rect 15654 6168 15660 6180
rect 15427 6140 15660 6168
rect 15427 6137 15439 6140
rect 15381 6131 15439 6137
rect 15654 6128 15660 6140
rect 15712 6168 15718 6180
rect 17402 6168 17408 6180
rect 15712 6140 17408 6168
rect 15712 6128 15718 6140
rect 17402 6128 17408 6140
rect 17460 6128 17466 6180
rect 4154 6100 4160 6112
rect 4115 6072 4160 6100
rect 4154 6060 4160 6072
rect 4212 6060 4218 6112
rect 5258 6060 5264 6112
rect 5316 6100 5322 6112
rect 6549 6103 6607 6109
rect 6549 6100 6561 6103
rect 5316 6072 6561 6100
rect 5316 6060 5322 6072
rect 6549 6069 6561 6072
rect 6595 6069 6607 6103
rect 6549 6063 6607 6069
rect 8478 6060 8484 6112
rect 8536 6100 8542 6112
rect 8941 6103 8999 6109
rect 8941 6100 8953 6103
rect 8536 6072 8953 6100
rect 8536 6060 8542 6072
rect 8941 6069 8953 6072
rect 8987 6069 8999 6103
rect 8941 6063 8999 6069
rect 11790 6060 11796 6112
rect 11848 6100 11854 6112
rect 11977 6103 12035 6109
rect 11977 6100 11989 6103
rect 11848 6072 11989 6100
rect 11848 6060 11854 6072
rect 11977 6069 11989 6072
rect 12023 6069 12035 6103
rect 13446 6100 13452 6112
rect 13359 6072 13452 6100
rect 11977 6063 12035 6069
rect 13446 6060 13452 6072
rect 13504 6100 13510 6112
rect 16206 6100 16212 6112
rect 13504 6072 16212 6100
rect 13504 6060 13510 6072
rect 16206 6060 16212 6072
rect 16264 6060 16270 6112
rect 1104 6010 18860 6032
rect 1104 5958 3169 6010
rect 3221 5958 3233 6010
rect 3285 5958 3297 6010
rect 3349 5958 3361 6010
rect 3413 5958 3425 6010
rect 3477 5958 7608 6010
rect 7660 5958 7672 6010
rect 7724 5958 7736 6010
rect 7788 5958 7800 6010
rect 7852 5958 7864 6010
rect 7916 5958 12047 6010
rect 12099 5958 12111 6010
rect 12163 5958 12175 6010
rect 12227 5958 12239 6010
rect 12291 5958 12303 6010
rect 12355 5958 16486 6010
rect 16538 5958 16550 6010
rect 16602 5958 16614 6010
rect 16666 5958 16678 6010
rect 16730 5958 16742 6010
rect 16794 5958 18860 6010
rect 1104 5936 18860 5958
rect 3694 5856 3700 5908
rect 3752 5896 3758 5908
rect 3973 5899 4031 5905
rect 3973 5896 3985 5899
rect 3752 5868 3985 5896
rect 3752 5856 3758 5868
rect 3973 5865 3985 5868
rect 4019 5896 4031 5899
rect 4062 5896 4068 5908
rect 4019 5868 4068 5896
rect 4019 5865 4031 5868
rect 3973 5859 4031 5865
rect 4062 5856 4068 5868
rect 4120 5856 4126 5908
rect 6086 5896 6092 5908
rect 4448 5868 6092 5896
rect 3050 5828 3056 5840
rect 3011 5800 3056 5828
rect 3050 5788 3056 5800
rect 3108 5788 3114 5840
rect 4448 5828 4476 5868
rect 6086 5856 6092 5868
rect 6144 5856 6150 5908
rect 7653 5899 7711 5905
rect 7653 5896 7665 5899
rect 6380 5868 7665 5896
rect 5902 5828 5908 5840
rect 3896 5800 4476 5828
rect 4540 5800 5908 5828
rect 2317 5763 2375 5769
rect 2317 5729 2329 5763
rect 2363 5760 2375 5763
rect 3896 5760 3924 5800
rect 2363 5732 3924 5760
rect 2363 5729 2375 5732
rect 2317 5723 2375 5729
rect 2777 5695 2835 5701
rect 2777 5661 2789 5695
rect 2823 5692 2835 5695
rect 2958 5692 2964 5704
rect 2823 5664 2964 5692
rect 2823 5661 2835 5664
rect 2777 5655 2835 5661
rect 2958 5652 2964 5664
rect 3016 5652 3022 5704
rect 3068 5701 3096 5732
rect 4062 5720 4068 5772
rect 4120 5760 4126 5772
rect 4540 5769 4568 5800
rect 5902 5788 5908 5800
rect 5960 5788 5966 5840
rect 4525 5763 4583 5769
rect 4525 5760 4537 5763
rect 4120 5732 4537 5760
rect 4120 5720 4126 5732
rect 4525 5729 4537 5732
rect 4571 5729 4583 5763
rect 4525 5723 4583 5729
rect 4614 5720 4620 5772
rect 4672 5760 4678 5772
rect 5261 5763 5319 5769
rect 5261 5760 5273 5763
rect 4672 5732 5273 5760
rect 4672 5720 4678 5732
rect 5261 5729 5273 5732
rect 5307 5729 5319 5763
rect 5261 5723 5319 5729
rect 6380 5704 6408 5868
rect 7653 5865 7665 5868
rect 7699 5865 7711 5899
rect 11422 5896 11428 5908
rect 11383 5868 11428 5896
rect 7653 5859 7711 5865
rect 11422 5856 11428 5868
rect 11480 5856 11486 5908
rect 11882 5856 11888 5908
rect 11940 5896 11946 5908
rect 12069 5899 12127 5905
rect 12069 5896 12081 5899
rect 11940 5868 12081 5896
rect 11940 5856 11946 5868
rect 12069 5865 12081 5868
rect 12115 5865 12127 5899
rect 12069 5859 12127 5865
rect 13725 5899 13783 5905
rect 13725 5865 13737 5899
rect 13771 5896 13783 5899
rect 14642 5896 14648 5908
rect 13771 5868 14648 5896
rect 13771 5865 13783 5868
rect 13725 5859 13783 5865
rect 14642 5856 14648 5868
rect 14700 5856 14706 5908
rect 15930 5896 15936 5908
rect 15891 5868 15936 5896
rect 15930 5856 15936 5868
rect 15988 5856 15994 5908
rect 17310 5896 17316 5908
rect 16040 5868 17316 5896
rect 7926 5788 7932 5840
rect 7984 5828 7990 5840
rect 8297 5831 8355 5837
rect 8297 5828 8309 5831
rect 7984 5800 8309 5828
rect 7984 5788 7990 5800
rect 8297 5797 8309 5800
rect 8343 5797 8355 5831
rect 10410 5828 10416 5840
rect 8297 5791 8355 5797
rect 9692 5800 10416 5828
rect 7282 5720 7288 5772
rect 7340 5760 7346 5772
rect 7745 5763 7803 5769
rect 7745 5760 7757 5763
rect 7340 5732 7757 5760
rect 7340 5720 7346 5732
rect 7745 5729 7757 5732
rect 7791 5760 7803 5763
rect 8110 5760 8116 5772
rect 7791 5732 8116 5760
rect 7791 5729 7803 5732
rect 7745 5723 7803 5729
rect 8110 5720 8116 5732
rect 8168 5760 8174 5772
rect 8168 5732 8340 5760
rect 8168 5720 8174 5732
rect 3053 5695 3111 5701
rect 3053 5661 3065 5695
rect 3099 5661 3111 5695
rect 3053 5655 3111 5661
rect 4709 5695 4767 5701
rect 4709 5661 4721 5695
rect 4755 5661 4767 5695
rect 4709 5655 4767 5661
rect 4801 5695 4859 5701
rect 4801 5661 4813 5695
rect 4847 5692 4859 5695
rect 6362 5692 6368 5704
rect 4847 5664 6368 5692
rect 4847 5661 4859 5664
rect 4801 5655 4859 5661
rect 2866 5624 2872 5636
rect 2827 5596 2872 5624
rect 2866 5584 2872 5596
rect 2924 5584 2930 5636
rect 4724 5624 4752 5655
rect 6362 5652 6368 5664
rect 6420 5652 6426 5704
rect 7006 5692 7012 5704
rect 6967 5664 7012 5692
rect 7006 5652 7012 5664
rect 7064 5652 7070 5704
rect 7837 5695 7895 5701
rect 7837 5661 7849 5695
rect 7883 5692 7895 5695
rect 8202 5692 8208 5704
rect 7883 5664 8208 5692
rect 7883 5661 7895 5664
rect 7837 5655 7895 5661
rect 8202 5652 8208 5664
rect 8260 5652 8266 5704
rect 8312 5701 8340 5732
rect 8297 5695 8355 5701
rect 8297 5661 8309 5695
rect 8343 5661 8355 5695
rect 8478 5692 8484 5704
rect 8439 5664 8484 5692
rect 8297 5655 8355 5661
rect 8478 5652 8484 5664
rect 8536 5652 8542 5704
rect 8570 5652 8576 5704
rect 8628 5692 8634 5704
rect 9493 5695 9551 5701
rect 8628 5664 8673 5692
rect 8628 5652 8634 5664
rect 9493 5661 9505 5695
rect 9539 5692 9551 5695
rect 9692 5692 9720 5800
rect 10410 5788 10416 5800
rect 10468 5788 10474 5840
rect 10612 5800 12940 5828
rect 10318 5760 10324 5772
rect 9784 5732 10324 5760
rect 9784 5701 9812 5732
rect 10318 5720 10324 5732
rect 10376 5760 10382 5772
rect 10612 5760 10640 5800
rect 10376 5732 10640 5760
rect 10376 5720 10382 5732
rect 9539 5664 9720 5692
rect 9769 5695 9827 5701
rect 9539 5661 9551 5664
rect 9493 5655 9551 5661
rect 9769 5661 9781 5695
rect 9815 5661 9827 5695
rect 10410 5692 10416 5704
rect 10371 5664 10416 5692
rect 9769 5655 9827 5661
rect 10410 5652 10416 5664
rect 10468 5652 10474 5704
rect 10612 5701 10640 5732
rect 10686 5720 10692 5772
rect 10744 5760 10750 5772
rect 12802 5760 12808 5772
rect 10744 5732 12296 5760
rect 10744 5720 10750 5732
rect 10597 5695 10655 5701
rect 10597 5661 10609 5695
rect 10643 5661 10655 5695
rect 10597 5655 10655 5661
rect 10781 5695 10839 5701
rect 10781 5661 10793 5695
rect 10827 5692 10839 5695
rect 11146 5692 11152 5704
rect 10827 5664 11152 5692
rect 10827 5661 10839 5664
rect 10781 5655 10839 5661
rect 11146 5652 11152 5664
rect 11204 5652 11210 5704
rect 12268 5701 12296 5732
rect 12452 5732 12808 5760
rect 12253 5695 12311 5701
rect 12253 5661 12265 5695
rect 12299 5661 12311 5695
rect 12253 5655 12311 5661
rect 6546 5624 6552 5636
rect 4724 5596 6552 5624
rect 6546 5584 6552 5596
rect 6604 5584 6610 5636
rect 9585 5627 9643 5633
rect 9585 5593 9597 5627
rect 9631 5624 9643 5627
rect 10689 5627 10747 5633
rect 9631 5596 10548 5624
rect 9631 5593 9643 5596
rect 9585 5587 9643 5593
rect 4801 5559 4859 5565
rect 4801 5525 4813 5559
rect 4847 5556 4859 5559
rect 6178 5556 6184 5568
rect 4847 5528 6184 5556
rect 4847 5525 4859 5528
rect 4801 5519 4859 5525
rect 6178 5516 6184 5528
rect 6236 5516 6242 5568
rect 7466 5556 7472 5568
rect 7427 5528 7472 5556
rect 7466 5516 7472 5528
rect 7524 5516 7530 5568
rect 9953 5559 10011 5565
rect 9953 5525 9965 5559
rect 9999 5556 10011 5559
rect 10226 5556 10232 5568
rect 9999 5528 10232 5556
rect 9999 5525 10011 5528
rect 9953 5519 10011 5525
rect 10226 5516 10232 5528
rect 10284 5516 10290 5568
rect 10520 5556 10548 5596
rect 10689 5593 10701 5627
rect 10735 5624 10747 5627
rect 12452 5624 12480 5732
rect 12802 5720 12808 5732
rect 12860 5720 12866 5772
rect 12529 5695 12587 5701
rect 12529 5661 12541 5695
rect 12575 5661 12587 5695
rect 12529 5655 12587 5661
rect 10735 5596 12480 5624
rect 12544 5624 12572 5655
rect 12912 5624 12940 5800
rect 16040 5760 16068 5868
rect 17310 5856 17316 5868
rect 17368 5896 17374 5908
rect 17589 5899 17647 5905
rect 17589 5896 17601 5899
rect 17368 5868 17601 5896
rect 17368 5856 17374 5868
rect 17589 5865 17601 5868
rect 17635 5865 17647 5899
rect 17589 5859 17647 5865
rect 17773 5899 17831 5905
rect 17773 5865 17785 5899
rect 17819 5896 17831 5899
rect 17862 5896 17868 5908
rect 17819 5868 17868 5896
rect 17819 5865 17831 5868
rect 17773 5859 17831 5865
rect 17862 5856 17868 5868
rect 17920 5856 17926 5908
rect 17954 5856 17960 5908
rect 18012 5896 18018 5908
rect 18233 5899 18291 5905
rect 18233 5896 18245 5899
rect 18012 5868 18245 5896
rect 18012 5856 18018 5868
rect 18233 5865 18245 5868
rect 18279 5865 18291 5899
rect 18233 5859 18291 5865
rect 16669 5831 16727 5837
rect 16669 5797 16681 5831
rect 16715 5797 16727 5831
rect 16669 5791 16727 5797
rect 15488 5732 16068 5760
rect 16684 5760 16712 5791
rect 17586 5760 17592 5772
rect 16684 5732 17592 5760
rect 13078 5692 13084 5704
rect 13039 5664 13084 5692
rect 13078 5652 13084 5664
rect 13136 5652 13142 5704
rect 13262 5692 13268 5704
rect 13223 5664 13268 5692
rect 13262 5652 13268 5664
rect 13320 5652 13326 5704
rect 13538 5692 13544 5704
rect 13499 5664 13544 5692
rect 13538 5652 13544 5664
rect 13596 5652 13602 5704
rect 14642 5652 14648 5704
rect 14700 5692 14706 5704
rect 15488 5701 15516 5732
rect 17586 5720 17592 5732
rect 17644 5720 17650 5772
rect 15289 5695 15347 5701
rect 15289 5692 15301 5695
rect 14700 5664 15301 5692
rect 14700 5652 14706 5664
rect 15289 5661 15301 5664
rect 15335 5661 15347 5695
rect 15289 5655 15347 5661
rect 15473 5695 15531 5701
rect 15473 5661 15485 5695
rect 15519 5661 15531 5695
rect 15746 5692 15752 5704
rect 15659 5664 15752 5692
rect 15473 5655 15531 5661
rect 15746 5652 15752 5664
rect 15804 5692 15810 5704
rect 16945 5695 17003 5701
rect 16945 5692 16957 5695
rect 15804 5664 16957 5692
rect 15804 5652 15810 5664
rect 16945 5661 16957 5664
rect 16991 5692 17003 5695
rect 17678 5692 17684 5704
rect 16991 5664 17684 5692
rect 16991 5661 17003 5664
rect 16945 5655 17003 5661
rect 17678 5652 17684 5664
rect 17736 5652 17742 5704
rect 16022 5624 16028 5636
rect 12544 5596 16028 5624
rect 10735 5593 10747 5596
rect 10689 5587 10747 5593
rect 10704 5556 10732 5587
rect 16022 5584 16028 5596
rect 16080 5584 16086 5636
rect 17402 5624 17408 5636
rect 17363 5596 17408 5624
rect 17402 5584 17408 5596
rect 17460 5584 17466 5636
rect 10520 5528 10732 5556
rect 10778 5516 10784 5568
rect 10836 5556 10842 5568
rect 10965 5559 11023 5565
rect 10965 5556 10977 5559
rect 10836 5528 10977 5556
rect 10836 5516 10842 5528
rect 10965 5525 10977 5528
rect 11011 5525 11023 5559
rect 10965 5519 11023 5525
rect 12437 5559 12495 5565
rect 12437 5525 12449 5559
rect 12483 5556 12495 5559
rect 14182 5556 14188 5568
rect 12483 5528 14188 5556
rect 12483 5525 12495 5528
rect 12437 5519 12495 5525
rect 14182 5516 14188 5528
rect 14240 5516 14246 5568
rect 14829 5559 14887 5565
rect 14829 5525 14841 5559
rect 14875 5556 14887 5559
rect 16206 5556 16212 5568
rect 14875 5528 16212 5556
rect 14875 5525 14887 5528
rect 14829 5519 14887 5525
rect 16206 5516 16212 5528
rect 16264 5516 16270 5568
rect 16298 5516 16304 5568
rect 16356 5556 16362 5568
rect 16485 5559 16543 5565
rect 16485 5556 16497 5559
rect 16356 5528 16497 5556
rect 16356 5516 16362 5528
rect 16485 5525 16497 5528
rect 16531 5556 16543 5559
rect 17605 5559 17663 5565
rect 17605 5556 17617 5559
rect 16531 5528 17617 5556
rect 16531 5525 16543 5528
rect 16485 5519 16543 5525
rect 17605 5525 17617 5528
rect 17651 5525 17663 5559
rect 17605 5519 17663 5525
rect 1104 5466 19019 5488
rect 1104 5414 5388 5466
rect 5440 5414 5452 5466
rect 5504 5414 5516 5466
rect 5568 5414 5580 5466
rect 5632 5414 5644 5466
rect 5696 5414 9827 5466
rect 9879 5414 9891 5466
rect 9943 5414 9955 5466
rect 10007 5414 10019 5466
rect 10071 5414 10083 5466
rect 10135 5414 14266 5466
rect 14318 5414 14330 5466
rect 14382 5414 14394 5466
rect 14446 5414 14458 5466
rect 14510 5414 14522 5466
rect 14574 5414 18705 5466
rect 18757 5414 18769 5466
rect 18821 5414 18833 5466
rect 18885 5414 18897 5466
rect 18949 5414 18961 5466
rect 19013 5414 19019 5466
rect 1104 5392 19019 5414
rect 2225 5355 2283 5361
rect 2225 5321 2237 5355
rect 2271 5352 2283 5355
rect 2958 5352 2964 5364
rect 2271 5324 2964 5352
rect 2271 5321 2283 5324
rect 2225 5315 2283 5321
rect 2958 5312 2964 5324
rect 3016 5312 3022 5364
rect 3970 5312 3976 5364
rect 4028 5352 4034 5364
rect 5445 5355 5503 5361
rect 5445 5352 5457 5355
rect 4028 5324 5457 5352
rect 4028 5312 4034 5324
rect 5445 5321 5457 5324
rect 5491 5321 5503 5355
rect 5902 5352 5908 5364
rect 5863 5324 5908 5352
rect 5445 5315 5503 5321
rect 5902 5312 5908 5324
rect 5960 5312 5966 5364
rect 6914 5352 6920 5364
rect 6875 5324 6920 5352
rect 6914 5312 6920 5324
rect 6972 5312 6978 5364
rect 10597 5355 10655 5361
rect 10597 5321 10609 5355
rect 10643 5352 10655 5355
rect 11054 5352 11060 5364
rect 10643 5324 11060 5352
rect 10643 5321 10655 5324
rect 10597 5315 10655 5321
rect 11054 5312 11060 5324
rect 11112 5352 11118 5364
rect 11698 5352 11704 5364
rect 11112 5324 11704 5352
rect 11112 5312 11118 5324
rect 11698 5312 11704 5324
rect 11756 5312 11762 5364
rect 14182 5312 14188 5364
rect 14240 5312 14246 5364
rect 15289 5355 15347 5361
rect 15289 5321 15301 5355
rect 15335 5352 15347 5355
rect 17034 5352 17040 5364
rect 15335 5324 17040 5352
rect 15335 5321 15347 5324
rect 15289 5315 15347 5321
rect 17034 5312 17040 5324
rect 17092 5312 17098 5364
rect 17954 5352 17960 5364
rect 17236 5324 17960 5352
rect 4614 5284 4620 5296
rect 4080 5256 4620 5284
rect 3349 5219 3407 5225
rect 3349 5185 3361 5219
rect 3395 5216 3407 5219
rect 3510 5216 3516 5228
rect 3395 5188 3516 5216
rect 3395 5185 3407 5188
rect 3349 5179 3407 5185
rect 3510 5176 3516 5188
rect 3568 5176 3574 5228
rect 4080 5225 4108 5256
rect 4614 5244 4620 5256
rect 4672 5244 4678 5296
rect 7006 5244 7012 5296
rect 7064 5284 7070 5296
rect 7837 5287 7895 5293
rect 7837 5284 7849 5287
rect 7064 5256 7849 5284
rect 7064 5244 7070 5256
rect 7837 5253 7849 5256
rect 7883 5253 7895 5287
rect 7837 5247 7895 5253
rect 9585 5287 9643 5293
rect 9585 5253 9597 5287
rect 9631 5284 9643 5287
rect 9674 5284 9680 5296
rect 9631 5256 9680 5284
rect 9631 5253 9643 5256
rect 9585 5247 9643 5253
rect 9674 5244 9680 5256
rect 9732 5284 9738 5296
rect 14200 5284 14228 5312
rect 16117 5287 16175 5293
rect 16117 5284 16129 5287
rect 9732 5256 12434 5284
rect 14200 5256 16129 5284
rect 9732 5244 9738 5256
rect 3605 5219 3663 5225
rect 3605 5185 3617 5219
rect 3651 5216 3663 5219
rect 4065 5219 4123 5225
rect 4065 5216 4077 5219
rect 3651 5188 4077 5216
rect 3651 5185 3663 5188
rect 3605 5179 3663 5185
rect 4065 5185 4077 5188
rect 4111 5185 4123 5219
rect 4065 5179 4123 5185
rect 4154 5176 4160 5228
rect 4212 5216 4218 5228
rect 4321 5219 4379 5225
rect 4321 5216 4333 5219
rect 4212 5188 4333 5216
rect 4212 5176 4218 5188
rect 4321 5185 4333 5188
rect 4367 5185 4379 5219
rect 4321 5179 4379 5185
rect 6825 5219 6883 5225
rect 6825 5185 6837 5219
rect 6871 5216 6883 5219
rect 7098 5216 7104 5228
rect 6871 5188 7104 5216
rect 6871 5185 6883 5188
rect 6825 5179 6883 5185
rect 7098 5176 7104 5188
rect 7156 5176 7162 5228
rect 11146 5216 11152 5228
rect 11107 5188 11152 5216
rect 11146 5176 11152 5188
rect 11204 5176 11210 5228
rect 11900 5225 11928 5256
rect 11885 5219 11943 5225
rect 11885 5185 11897 5219
rect 11931 5185 11943 5219
rect 12141 5219 12199 5225
rect 12141 5216 12153 5219
rect 11885 5179 11943 5185
rect 11992 5188 12153 5216
rect 6733 5151 6791 5157
rect 6733 5117 6745 5151
rect 6779 5148 6791 5151
rect 8662 5148 8668 5160
rect 6779 5120 8668 5148
rect 6779 5117 6791 5120
rect 6733 5111 6791 5117
rect 8662 5108 8668 5120
rect 8720 5108 8726 5160
rect 9950 5108 9956 5160
rect 10008 5148 10014 5160
rect 10873 5151 10931 5157
rect 10873 5148 10885 5151
rect 10008 5120 10885 5148
rect 10008 5108 10014 5120
rect 10873 5117 10885 5120
rect 10919 5117 10931 5151
rect 10873 5111 10931 5117
rect 11790 5108 11796 5160
rect 11848 5148 11854 5160
rect 11992 5148 12020 5188
rect 12141 5185 12153 5188
rect 12187 5185 12199 5219
rect 12406 5216 12434 5256
rect 16117 5253 16129 5256
rect 16163 5253 16175 5287
rect 16117 5247 16175 5253
rect 16301 5287 16359 5293
rect 16301 5253 16313 5287
rect 16347 5284 16359 5287
rect 17126 5284 17132 5296
rect 16347 5256 17132 5284
rect 16347 5253 16359 5256
rect 16301 5247 16359 5253
rect 13909 5219 13967 5225
rect 13909 5216 13921 5219
rect 12406 5188 13921 5216
rect 12141 5179 12199 5185
rect 13909 5185 13921 5188
rect 13955 5216 13967 5219
rect 13998 5216 14004 5228
rect 13955 5188 14004 5216
rect 13955 5185 13967 5188
rect 13909 5179 13967 5185
rect 13998 5176 14004 5188
rect 14056 5176 14062 5228
rect 14176 5219 14234 5225
rect 14176 5185 14188 5219
rect 14222 5216 14234 5219
rect 15838 5216 15844 5228
rect 14222 5188 15844 5216
rect 14222 5185 14234 5188
rect 14176 5179 14234 5185
rect 15838 5176 15844 5188
rect 15896 5176 15902 5228
rect 16022 5216 16028 5228
rect 15983 5188 16028 5216
rect 16022 5176 16028 5188
rect 16080 5176 16086 5228
rect 16132 5216 16160 5247
rect 17126 5244 17132 5256
rect 17184 5244 17190 5296
rect 16942 5216 16948 5228
rect 16132 5188 16948 5216
rect 16942 5176 16948 5188
rect 17000 5176 17006 5228
rect 17034 5176 17040 5228
rect 17092 5216 17098 5228
rect 17236 5225 17264 5324
rect 17954 5312 17960 5324
rect 18012 5352 18018 5364
rect 18233 5355 18291 5361
rect 18233 5352 18245 5355
rect 18012 5324 18245 5352
rect 18012 5312 18018 5324
rect 18233 5321 18245 5324
rect 18279 5321 18291 5355
rect 18233 5315 18291 5321
rect 17586 5284 17592 5296
rect 17547 5256 17592 5284
rect 17586 5244 17592 5256
rect 17644 5244 17650 5296
rect 17221 5219 17279 5225
rect 17221 5216 17233 5219
rect 17092 5188 17233 5216
rect 17092 5176 17098 5188
rect 17221 5185 17233 5188
rect 17267 5185 17279 5219
rect 17221 5179 17279 5185
rect 11848 5120 12020 5148
rect 11848 5108 11854 5120
rect 6362 4972 6368 5024
rect 6420 5012 6426 5024
rect 7098 5012 7104 5024
rect 6420 4984 7104 5012
rect 6420 4972 6426 4984
rect 7098 4972 7104 4984
rect 7156 5012 7162 5024
rect 7285 5015 7343 5021
rect 7285 5012 7297 5015
rect 7156 4984 7297 5012
rect 7156 4972 7162 4984
rect 7285 4981 7297 4984
rect 7331 4981 7343 5015
rect 7285 4975 7343 4981
rect 10965 5015 11023 5021
rect 10965 4981 10977 5015
rect 11011 5012 11023 5015
rect 11422 5012 11428 5024
rect 11011 4984 11428 5012
rect 11011 4981 11023 4984
rect 10965 4975 11023 4981
rect 11422 4972 11428 4984
rect 11480 4972 11486 5024
rect 13262 5012 13268 5024
rect 13223 4984 13268 5012
rect 13262 4972 13268 4984
rect 13320 4972 13326 5024
rect 15930 4972 15936 5024
rect 15988 5012 15994 5024
rect 16301 5015 16359 5021
rect 16301 5012 16313 5015
rect 15988 4984 16313 5012
rect 15988 4972 15994 4984
rect 16301 4981 16313 4984
rect 16347 4981 16359 5015
rect 16301 4975 16359 4981
rect 17402 4972 17408 5024
rect 17460 5012 17466 5024
rect 17589 5015 17647 5021
rect 17589 5012 17601 5015
rect 17460 4984 17601 5012
rect 17460 4972 17466 4984
rect 17589 4981 17601 4984
rect 17635 4981 17647 5015
rect 17770 5012 17776 5024
rect 17731 4984 17776 5012
rect 17589 4975 17647 4981
rect 17770 4972 17776 4984
rect 17828 4972 17834 5024
rect 1104 4922 18860 4944
rect 1104 4870 3169 4922
rect 3221 4870 3233 4922
rect 3285 4870 3297 4922
rect 3349 4870 3361 4922
rect 3413 4870 3425 4922
rect 3477 4870 7608 4922
rect 7660 4870 7672 4922
rect 7724 4870 7736 4922
rect 7788 4870 7800 4922
rect 7852 4870 7864 4922
rect 7916 4870 12047 4922
rect 12099 4870 12111 4922
rect 12163 4870 12175 4922
rect 12227 4870 12239 4922
rect 12291 4870 12303 4922
rect 12355 4870 16486 4922
rect 16538 4870 16550 4922
rect 16602 4870 16614 4922
rect 16666 4870 16678 4922
rect 16730 4870 16742 4922
rect 16794 4870 18860 4922
rect 1104 4848 18860 4870
rect 2958 4808 2964 4820
rect 2919 4780 2964 4808
rect 2958 4768 2964 4780
rect 3016 4768 3022 4820
rect 3329 4811 3387 4817
rect 3329 4777 3341 4811
rect 3375 4808 3387 4811
rect 3510 4808 3516 4820
rect 3375 4780 3516 4808
rect 3375 4777 3387 4780
rect 3329 4771 3387 4777
rect 3510 4768 3516 4780
rect 3568 4768 3574 4820
rect 4341 4811 4399 4817
rect 4341 4777 4353 4811
rect 4387 4808 4399 4811
rect 5074 4808 5080 4820
rect 4387 4780 5080 4808
rect 4387 4777 4399 4780
rect 4341 4771 4399 4777
rect 5074 4768 5080 4780
rect 5132 4808 5138 4820
rect 5261 4811 5319 4817
rect 5261 4808 5273 4811
rect 5132 4780 5273 4808
rect 5132 4768 5138 4780
rect 5261 4777 5273 4780
rect 5307 4777 5319 4811
rect 6730 4808 6736 4820
rect 6691 4780 6736 4808
rect 5261 4771 5319 4777
rect 6730 4768 6736 4780
rect 6788 4768 6794 4820
rect 8573 4811 8631 4817
rect 8573 4777 8585 4811
rect 8619 4808 8631 4811
rect 9122 4808 9128 4820
rect 8619 4780 9128 4808
rect 8619 4777 8631 4780
rect 8573 4771 8631 4777
rect 9122 4768 9128 4780
rect 9180 4768 9186 4820
rect 9953 4811 10011 4817
rect 9953 4777 9965 4811
rect 9999 4808 10011 4811
rect 10226 4808 10232 4820
rect 9999 4780 10232 4808
rect 9999 4777 10011 4780
rect 9953 4771 10011 4777
rect 10226 4768 10232 4780
rect 10284 4768 10290 4820
rect 10778 4808 10784 4820
rect 10739 4780 10784 4808
rect 10778 4768 10784 4780
rect 10836 4768 10842 4820
rect 14182 4768 14188 4820
rect 14240 4808 14246 4820
rect 14277 4811 14335 4817
rect 14277 4808 14289 4811
rect 14240 4780 14289 4808
rect 14240 4768 14246 4780
rect 14277 4777 14289 4780
rect 14323 4777 14335 4811
rect 15838 4808 15844 4820
rect 15799 4780 15844 4808
rect 14277 4771 14335 4777
rect 15838 4768 15844 4780
rect 15896 4768 15902 4820
rect 16669 4811 16727 4817
rect 16669 4777 16681 4811
rect 16715 4808 16727 4811
rect 16942 4808 16948 4820
rect 16715 4780 16948 4808
rect 16715 4777 16727 4780
rect 16669 4771 16727 4777
rect 16942 4768 16948 4780
rect 17000 4808 17006 4820
rect 18138 4808 18144 4820
rect 17000 4780 18000 4808
rect 18099 4780 18144 4808
rect 17000 4768 17006 4780
rect 10965 4743 11023 4749
rect 10965 4709 10977 4743
rect 11011 4709 11023 4743
rect 13722 4740 13728 4752
rect 13635 4712 13728 4740
rect 10965 4703 11023 4709
rect 2866 4672 2872 4684
rect 2827 4644 2872 4672
rect 2866 4632 2872 4644
rect 2924 4632 2930 4684
rect 4614 4632 4620 4684
rect 4672 4672 4678 4684
rect 5258 4672 5264 4684
rect 4672 4644 5264 4672
rect 4672 4632 4678 4644
rect 5258 4632 5264 4644
rect 5316 4672 5322 4684
rect 7190 4672 7196 4684
rect 5316 4644 7196 4672
rect 5316 4632 5322 4644
rect 7190 4632 7196 4644
rect 7248 4632 7254 4684
rect 10318 4672 10324 4684
rect 9140 4644 10324 4672
rect 3050 4564 3056 4616
rect 3108 4604 3114 4616
rect 3145 4607 3203 4613
rect 3145 4604 3157 4607
rect 3108 4576 3157 4604
rect 3108 4564 3114 4576
rect 3145 4573 3157 4576
rect 3191 4573 3203 4607
rect 3145 4567 3203 4573
rect 5537 4607 5595 4613
rect 5537 4573 5549 4607
rect 5583 4604 5595 4607
rect 5902 4604 5908 4616
rect 5583 4576 5908 4604
rect 5583 4573 5595 4576
rect 5537 4567 5595 4573
rect 5902 4564 5908 4576
rect 5960 4564 5966 4616
rect 6362 4604 6368 4616
rect 6323 4576 6368 4604
rect 6362 4564 6368 4576
rect 6420 4564 6426 4616
rect 6549 4607 6607 4613
rect 6549 4573 6561 4607
rect 6595 4604 6607 4607
rect 7282 4604 7288 4616
rect 6595 4576 7288 4604
rect 6595 4573 6607 4576
rect 6549 4567 6607 4573
rect 7282 4564 7288 4576
rect 7340 4564 7346 4616
rect 7460 4607 7518 4613
rect 7460 4573 7472 4607
rect 7506 4604 7518 4607
rect 7926 4604 7932 4616
rect 7506 4576 7932 4604
rect 7506 4573 7518 4576
rect 7460 4567 7518 4573
rect 7576 4548 7604 4576
rect 7926 4564 7932 4576
rect 7984 4564 7990 4616
rect 9140 4613 9168 4644
rect 10318 4632 10324 4644
rect 10376 4632 10382 4684
rect 9125 4607 9183 4613
rect 9125 4573 9137 4607
rect 9171 4573 9183 4607
rect 9125 4567 9183 4573
rect 9309 4607 9367 4613
rect 9309 4573 9321 4607
rect 9355 4604 9367 4607
rect 10410 4604 10416 4616
rect 9355 4576 10416 4604
rect 9355 4573 9367 4576
rect 9309 4567 9367 4573
rect 10410 4564 10416 4576
rect 10468 4564 10474 4616
rect 10980 4604 11008 4703
rect 13722 4700 13728 4712
rect 13780 4740 13786 4752
rect 15930 4740 15936 4752
rect 13780 4712 14964 4740
rect 15891 4712 15936 4740
rect 13780 4700 13786 4712
rect 13262 4632 13268 4684
rect 13320 4672 13326 4684
rect 14436 4675 14494 4681
rect 14436 4672 14448 4675
rect 13320 4644 14448 4672
rect 13320 4632 13326 4644
rect 14436 4641 14448 4644
rect 14482 4641 14494 4675
rect 14436 4635 14494 4641
rect 14553 4675 14611 4681
rect 14553 4641 14565 4675
rect 14599 4672 14611 4675
rect 14642 4672 14648 4684
rect 14599 4644 14648 4672
rect 14599 4641 14611 4644
rect 14553 4635 14611 4641
rect 14642 4632 14648 4644
rect 14700 4632 14706 4684
rect 14936 4681 14964 4712
rect 15930 4700 15936 4712
rect 15988 4700 15994 4752
rect 16022 4700 16028 4752
rect 16080 4740 16086 4752
rect 16080 4712 16712 4740
rect 16080 4700 16086 4712
rect 14921 4675 14979 4681
rect 14921 4641 14933 4675
rect 14967 4672 14979 4675
rect 14967 4644 16620 4672
rect 14967 4641 14979 4644
rect 14921 4635 14979 4641
rect 11425 4607 11483 4613
rect 11425 4604 11437 4607
rect 10980 4576 11437 4604
rect 11425 4573 11437 4576
rect 11471 4573 11483 4607
rect 11425 4567 11483 4573
rect 16025 4607 16083 4613
rect 16025 4573 16037 4607
rect 16071 4604 16083 4607
rect 16071 4576 16528 4604
rect 16071 4573 16083 4576
rect 16025 4567 16083 4573
rect 7558 4496 7564 4548
rect 7616 4496 7622 4548
rect 9950 4545 9956 4548
rect 9217 4539 9275 4545
rect 9217 4505 9229 4539
rect 9263 4536 9275 4539
rect 9937 4539 9956 4545
rect 9937 4536 9949 4539
rect 9263 4508 9949 4536
rect 9263 4505 9275 4508
rect 9217 4499 9275 4505
rect 9937 4505 9949 4508
rect 9937 4499 9956 4505
rect 9950 4496 9956 4499
rect 10008 4496 10014 4548
rect 10137 4539 10195 4545
rect 10137 4505 10149 4539
rect 10183 4536 10195 4539
rect 10502 4536 10508 4548
rect 10183 4508 10508 4536
rect 10183 4505 10195 4508
rect 10137 4499 10195 4505
rect 10502 4496 10508 4508
rect 10560 4536 10566 4548
rect 10597 4539 10655 4545
rect 10597 4536 10609 4539
rect 10560 4508 10609 4536
rect 10560 4496 10566 4508
rect 10597 4505 10609 4508
rect 10643 4505 10655 4539
rect 10597 4499 10655 4505
rect 10813 4539 10871 4545
rect 10813 4505 10825 4539
rect 10859 4536 10871 4539
rect 11054 4536 11060 4548
rect 10859 4508 11060 4536
rect 10859 4505 10871 4508
rect 10813 4499 10871 4505
rect 11054 4496 11060 4508
rect 11112 4496 11118 4548
rect 13078 4536 13084 4548
rect 11164 4508 13084 4536
rect 9674 4428 9680 4480
rect 9732 4468 9738 4480
rect 9769 4471 9827 4477
rect 9769 4468 9781 4471
rect 9732 4440 9781 4468
rect 9732 4428 9738 4440
rect 9769 4437 9781 4440
rect 9815 4437 9827 4471
rect 9769 4431 9827 4437
rect 10410 4428 10416 4480
rect 10468 4468 10474 4480
rect 10686 4468 10692 4480
rect 10468 4440 10692 4468
rect 10468 4428 10474 4440
rect 10686 4428 10692 4440
rect 10744 4468 10750 4480
rect 11164 4468 11192 4508
rect 13078 4496 13084 4508
rect 13136 4536 13142 4548
rect 14645 4539 14703 4545
rect 14645 4536 14657 4539
rect 13136 4508 14657 4536
rect 13136 4496 13142 4508
rect 14645 4505 14657 4508
rect 14691 4505 14703 4539
rect 14645 4499 14703 4505
rect 15749 4539 15807 4545
rect 15749 4505 15761 4539
rect 15795 4536 15807 4539
rect 16206 4536 16212 4548
rect 15795 4508 16212 4536
rect 15795 4505 15807 4508
rect 15749 4499 15807 4505
rect 16206 4496 16212 4508
rect 16264 4536 16270 4548
rect 16390 4536 16396 4548
rect 16264 4508 16396 4536
rect 16264 4496 16270 4508
rect 16390 4496 16396 4508
rect 16448 4496 16454 4548
rect 16500 4480 16528 4576
rect 11606 4468 11612 4480
rect 10744 4440 11192 4468
rect 11567 4440 11612 4468
rect 10744 4428 10750 4440
rect 11606 4428 11612 4440
rect 11664 4428 11670 4480
rect 16482 4468 16488 4480
rect 16443 4440 16488 4468
rect 16482 4428 16488 4440
rect 16540 4428 16546 4480
rect 16592 4468 16620 4644
rect 16684 4545 16712 4712
rect 17770 4700 17776 4752
rect 17828 4740 17834 4752
rect 17828 4712 17908 4740
rect 17828 4700 17834 4712
rect 17218 4564 17224 4616
rect 17276 4604 17282 4616
rect 17880 4613 17908 4712
rect 17972 4613 18000 4780
rect 18138 4768 18144 4780
rect 18196 4768 18202 4820
rect 17737 4607 17795 4613
rect 17737 4604 17749 4607
rect 17276 4576 17749 4604
rect 17276 4564 17282 4576
rect 17737 4573 17749 4576
rect 17783 4573 17795 4607
rect 17737 4567 17795 4573
rect 17845 4607 17908 4613
rect 17845 4573 17857 4607
rect 17891 4576 17908 4607
rect 17957 4607 18015 4613
rect 17891 4573 17903 4576
rect 17845 4567 17903 4573
rect 17957 4573 17969 4607
rect 18003 4573 18015 4607
rect 17957 4567 18015 4573
rect 16653 4539 16712 4545
rect 16653 4505 16665 4539
rect 16699 4508 16712 4539
rect 16853 4539 16911 4545
rect 16699 4505 16711 4508
rect 16653 4499 16711 4505
rect 16853 4505 16865 4539
rect 16899 4536 16911 4539
rect 17126 4536 17132 4548
rect 16899 4508 17132 4536
rect 16899 4505 16911 4508
rect 16853 4499 16911 4505
rect 17126 4496 17132 4508
rect 17184 4496 17190 4548
rect 17034 4468 17040 4480
rect 16592 4440 17040 4468
rect 17034 4428 17040 4440
rect 17092 4428 17098 4480
rect 1104 4378 19019 4400
rect 1104 4326 5388 4378
rect 5440 4326 5452 4378
rect 5504 4326 5516 4378
rect 5568 4326 5580 4378
rect 5632 4326 5644 4378
rect 5696 4326 9827 4378
rect 9879 4326 9891 4378
rect 9943 4326 9955 4378
rect 10007 4326 10019 4378
rect 10071 4326 10083 4378
rect 10135 4326 14266 4378
rect 14318 4326 14330 4378
rect 14382 4326 14394 4378
rect 14446 4326 14458 4378
rect 14510 4326 14522 4378
rect 14574 4326 18705 4378
rect 18757 4326 18769 4378
rect 18821 4326 18833 4378
rect 18885 4326 18897 4378
rect 18949 4326 18961 4378
rect 19013 4326 19019 4378
rect 1104 4304 19019 4326
rect 5166 4224 5172 4276
rect 5224 4264 5230 4276
rect 5224 4236 5396 4264
rect 5224 4224 5230 4236
rect 5368 4205 5396 4236
rect 8478 4224 8484 4276
rect 8536 4264 8542 4276
rect 8665 4267 8723 4273
rect 8665 4264 8677 4267
rect 8536 4236 8677 4264
rect 8536 4224 8542 4236
rect 8665 4233 8677 4236
rect 8711 4233 8723 4267
rect 10686 4264 10692 4276
rect 10647 4236 10692 4264
rect 8665 4227 8723 4233
rect 10686 4224 10692 4236
rect 10744 4224 10750 4276
rect 11146 4224 11152 4276
rect 11204 4264 11210 4276
rect 13081 4267 13139 4273
rect 13081 4264 13093 4267
rect 11204 4236 13093 4264
rect 11204 4224 11210 4236
rect 13081 4233 13093 4236
rect 13127 4264 13139 4267
rect 14642 4264 14648 4276
rect 13127 4236 14648 4264
rect 13127 4233 13139 4236
rect 13081 4227 13139 4233
rect 14642 4224 14648 4236
rect 14700 4224 14706 4276
rect 16942 4224 16948 4276
rect 17000 4264 17006 4276
rect 17221 4267 17279 4273
rect 17221 4264 17233 4267
rect 17000 4236 17233 4264
rect 17000 4224 17006 4236
rect 17221 4233 17233 4236
rect 17267 4264 17279 4267
rect 17586 4264 17592 4276
rect 17267 4236 17592 4264
rect 17267 4233 17279 4236
rect 17221 4227 17279 4233
rect 17586 4224 17592 4236
rect 17644 4224 17650 4276
rect 5353 4199 5411 4205
rect 5353 4165 5365 4199
rect 5399 4165 5411 4199
rect 5353 4159 5411 4165
rect 5537 4199 5595 4205
rect 5537 4165 5549 4199
rect 5583 4196 5595 4199
rect 5583 4168 7972 4196
rect 5583 4165 5595 4168
rect 5537 4159 5595 4165
rect 4525 4131 4583 4137
rect 4525 4097 4537 4131
rect 4571 4128 4583 4131
rect 5169 4131 5227 4137
rect 5169 4128 5181 4131
rect 4571 4100 5181 4128
rect 4571 4097 4583 4100
rect 4525 4091 4583 4097
rect 5169 4097 5181 4100
rect 5215 4097 5227 4131
rect 5368 4128 5396 4159
rect 5368 4100 6684 4128
rect 5169 4091 5227 4097
rect 6546 4060 6552 4072
rect 6507 4032 6552 4060
rect 6546 4020 6552 4032
rect 6604 4020 6610 4072
rect 6656 4060 6684 4100
rect 7374 4088 7380 4140
rect 7432 4128 7438 4140
rect 7469 4131 7527 4137
rect 7469 4128 7481 4131
rect 7432 4100 7481 4128
rect 7432 4088 7438 4100
rect 7469 4097 7481 4100
rect 7515 4128 7527 4131
rect 7558 4128 7564 4140
rect 7515 4100 7564 4128
rect 7515 4097 7527 4100
rect 7469 4091 7527 4097
rect 7558 4088 7564 4100
rect 7616 4088 7622 4140
rect 7944 4072 7972 4168
rect 11606 4156 11612 4208
rect 11664 4196 11670 4208
rect 11946 4199 12004 4205
rect 11946 4196 11958 4199
rect 11664 4168 11958 4196
rect 11664 4156 11670 4168
rect 11946 4165 11958 4168
rect 11992 4165 12004 4199
rect 16853 4199 16911 4205
rect 16853 4196 16865 4199
rect 11946 4159 12004 4165
rect 15488 4168 16865 4196
rect 8389 4131 8447 4137
rect 8389 4097 8401 4131
rect 8435 4097 8447 4131
rect 8389 4091 8447 4097
rect 7926 4060 7932 4072
rect 6656 4032 7512 4060
rect 7839 4032 7932 4060
rect 6730 3952 6736 4004
rect 6788 3992 6794 4004
rect 6917 3995 6975 4001
rect 6917 3992 6929 3995
rect 6788 3964 6929 3992
rect 6788 3952 6794 3964
rect 6917 3961 6929 3964
rect 6963 3992 6975 3995
rect 7374 3992 7380 4004
rect 6963 3964 7380 3992
rect 6963 3961 6975 3964
rect 6917 3955 6975 3961
rect 7374 3952 7380 3964
rect 7432 3952 7438 4004
rect 7484 3992 7512 4032
rect 7926 4020 7932 4032
rect 7984 4020 7990 4072
rect 8404 4060 8432 4091
rect 8662 4088 8668 4140
rect 8720 4128 8726 4140
rect 9582 4137 9588 4140
rect 8757 4131 8815 4137
rect 8757 4128 8769 4131
rect 8720 4100 8769 4128
rect 8720 4088 8726 4100
rect 8757 4097 8769 4100
rect 8803 4097 8815 4131
rect 8757 4091 8815 4097
rect 9576 4091 9588 4137
rect 9640 4128 9646 4140
rect 13909 4131 13967 4137
rect 9640 4100 9676 4128
rect 9582 4088 9588 4091
rect 9640 4088 9646 4100
rect 13909 4097 13921 4131
rect 13955 4128 13967 4131
rect 13998 4128 14004 4140
rect 13955 4100 14004 4128
rect 13955 4097 13967 4100
rect 13909 4091 13967 4097
rect 13998 4088 14004 4100
rect 14056 4088 14062 4140
rect 14176 4131 14234 4137
rect 14176 4097 14188 4131
rect 14222 4128 14234 4131
rect 15488 4128 15516 4168
rect 16853 4165 16865 4168
rect 16899 4165 16911 4199
rect 16853 4159 16911 4165
rect 17126 4156 17132 4208
rect 17184 4196 17190 4208
rect 17313 4199 17371 4205
rect 17313 4196 17325 4199
rect 17184 4168 17325 4196
rect 17184 4156 17190 4168
rect 17313 4165 17325 4168
rect 17359 4165 17371 4199
rect 17313 4159 17371 4165
rect 14222 4100 15516 4128
rect 16117 4131 16175 4137
rect 14222 4097 14234 4100
rect 14176 4091 14234 4097
rect 16117 4097 16129 4131
rect 16163 4097 16175 4131
rect 16298 4128 16304 4140
rect 16259 4100 16304 4128
rect 16117 4091 16175 4097
rect 8036 4032 8432 4060
rect 8573 4063 8631 4069
rect 8036 3992 8064 4032
rect 8573 4029 8585 4063
rect 8619 4029 8631 4063
rect 9306 4060 9312 4072
rect 9267 4032 9312 4060
rect 8573 4023 8631 4029
rect 8588 3992 8616 4023
rect 9306 4020 9312 4032
rect 9364 4020 9370 4072
rect 11698 4060 11704 4072
rect 11659 4032 11704 4060
rect 11698 4020 11704 4032
rect 11756 4020 11762 4072
rect 16132 4060 16160 4091
rect 16298 4088 16304 4100
rect 16356 4088 16362 4140
rect 16574 4128 16580 4140
rect 16408 4100 16580 4128
rect 16408 4060 16436 4100
rect 16574 4088 16580 4100
rect 16632 4128 16638 4140
rect 17144 4128 17172 4156
rect 16632 4100 17172 4128
rect 16632 4088 16638 4100
rect 16132 4032 16436 4060
rect 16482 4020 16488 4072
rect 16540 4060 16546 4072
rect 16945 4063 17003 4069
rect 16945 4060 16957 4063
rect 16540 4032 16957 4060
rect 16540 4020 16546 4032
rect 16945 4029 16957 4032
rect 16991 4060 17003 4063
rect 16991 4032 17908 4060
rect 16991 4029 17003 4032
rect 16945 4023 17003 4029
rect 7484 3964 8064 3992
rect 8312 3964 8616 3992
rect 16117 3995 16175 4001
rect 4706 3924 4712 3936
rect 4667 3896 4712 3924
rect 4706 3884 4712 3896
rect 4764 3884 4770 3936
rect 7006 3924 7012 3936
rect 6967 3896 7012 3924
rect 7006 3884 7012 3896
rect 7064 3884 7070 3936
rect 7282 3884 7288 3936
rect 7340 3924 7346 3936
rect 7561 3927 7619 3933
rect 7561 3924 7573 3927
rect 7340 3896 7573 3924
rect 7340 3884 7346 3896
rect 7561 3893 7573 3896
rect 7607 3924 7619 3927
rect 8312 3924 8340 3964
rect 16117 3961 16129 3995
rect 16163 3992 16175 3995
rect 17037 3995 17095 4001
rect 17037 3992 17049 3995
rect 16163 3964 17049 3992
rect 16163 3961 16175 3964
rect 16117 3955 16175 3961
rect 17037 3961 17049 3964
rect 17083 3961 17095 3995
rect 17037 3955 17095 3961
rect 17880 3936 17908 4032
rect 7607 3896 8340 3924
rect 7607 3893 7619 3896
rect 7561 3887 7619 3893
rect 8386 3884 8392 3936
rect 8444 3924 8450 3936
rect 15289 3927 15347 3933
rect 8444 3896 8489 3924
rect 8444 3884 8450 3896
rect 15289 3893 15301 3927
rect 15335 3924 15347 3927
rect 16942 3924 16948 3936
rect 15335 3896 16948 3924
rect 15335 3893 15347 3896
rect 15289 3887 15347 3893
rect 16942 3884 16948 3896
rect 17000 3884 17006 3936
rect 17862 3924 17868 3936
rect 17823 3896 17868 3924
rect 17862 3884 17868 3896
rect 17920 3884 17926 3936
rect 1104 3834 18860 3856
rect 1104 3782 3169 3834
rect 3221 3782 3233 3834
rect 3285 3782 3297 3834
rect 3349 3782 3361 3834
rect 3413 3782 3425 3834
rect 3477 3782 7608 3834
rect 7660 3782 7672 3834
rect 7724 3782 7736 3834
rect 7788 3782 7800 3834
rect 7852 3782 7864 3834
rect 7916 3782 12047 3834
rect 12099 3782 12111 3834
rect 12163 3782 12175 3834
rect 12227 3782 12239 3834
rect 12291 3782 12303 3834
rect 12355 3782 16486 3834
rect 16538 3782 16550 3834
rect 16602 3782 16614 3834
rect 16666 3782 16678 3834
rect 16730 3782 16742 3834
rect 16794 3782 18860 3834
rect 1104 3760 18860 3782
rect 8294 3680 8300 3732
rect 8352 3720 8358 3732
rect 8481 3723 8539 3729
rect 8481 3720 8493 3723
rect 8352 3692 8493 3720
rect 8352 3680 8358 3692
rect 8481 3689 8493 3692
rect 8527 3689 8539 3723
rect 8481 3683 8539 3689
rect 9493 3723 9551 3729
rect 9493 3689 9505 3723
rect 9539 3720 9551 3723
rect 9582 3720 9588 3732
rect 9539 3692 9588 3720
rect 9539 3689 9551 3692
rect 9493 3683 9551 3689
rect 9582 3680 9588 3692
rect 9640 3680 9646 3732
rect 13262 3680 13268 3732
rect 13320 3720 13326 3732
rect 15102 3720 15108 3732
rect 13320 3692 15108 3720
rect 13320 3680 13326 3692
rect 15102 3680 15108 3692
rect 15160 3680 15166 3732
rect 16574 3680 16580 3732
rect 16632 3720 16638 3732
rect 16850 3720 16856 3732
rect 16632 3692 16856 3720
rect 16632 3680 16638 3692
rect 16850 3680 16856 3692
rect 16908 3720 16914 3732
rect 17129 3723 17187 3729
rect 17129 3720 17141 3723
rect 16908 3692 17141 3720
rect 16908 3680 16914 3692
rect 17129 3689 17141 3692
rect 17175 3689 17187 3723
rect 17129 3683 17187 3689
rect 6546 3612 6552 3664
rect 6604 3652 6610 3664
rect 7282 3652 7288 3664
rect 6604 3624 7288 3652
rect 6604 3612 6610 3624
rect 7006 3584 7012 3596
rect 6288 3556 7012 3584
rect 5258 3476 5264 3528
rect 5316 3516 5322 3528
rect 5353 3519 5411 3525
rect 5353 3516 5365 3519
rect 5316 3488 5365 3516
rect 5316 3476 5322 3488
rect 5353 3485 5365 3488
rect 5399 3485 5411 3519
rect 6178 3516 6184 3528
rect 6139 3488 6184 3516
rect 5353 3479 5411 3485
rect 6178 3476 6184 3488
rect 6236 3476 6242 3528
rect 6288 3525 6316 3556
rect 7006 3544 7012 3556
rect 7064 3544 7070 3596
rect 7208 3593 7236 3624
rect 7282 3612 7288 3624
rect 7340 3612 7346 3664
rect 7374 3612 7380 3664
rect 7432 3612 7438 3664
rect 8386 3612 8392 3664
rect 8444 3652 8450 3664
rect 9030 3652 9036 3664
rect 8444 3624 9036 3652
rect 8444 3612 8450 3624
rect 9030 3612 9036 3624
rect 9088 3612 9094 3664
rect 12986 3612 12992 3664
rect 13044 3652 13050 3664
rect 16485 3655 16543 3661
rect 13044 3624 13308 3652
rect 13044 3612 13050 3624
rect 7193 3587 7251 3593
rect 7193 3553 7205 3587
rect 7239 3553 7251 3587
rect 7392 3584 7420 3612
rect 7653 3587 7711 3593
rect 7653 3584 7665 3587
rect 7392 3556 7665 3584
rect 7193 3547 7251 3553
rect 7653 3553 7665 3556
rect 7699 3553 7711 3587
rect 7653 3547 7711 3553
rect 7926 3544 7932 3596
rect 7984 3584 7990 3596
rect 7984 3556 9996 3584
rect 7984 3544 7990 3556
rect 6273 3519 6331 3525
rect 6273 3485 6285 3519
rect 6319 3485 6331 3519
rect 6454 3516 6460 3528
rect 6415 3488 6460 3516
rect 6273 3479 6331 3485
rect 6454 3476 6460 3488
rect 6512 3476 6518 3528
rect 6549 3519 6607 3525
rect 6549 3485 6561 3519
rect 6595 3516 6607 3519
rect 6822 3516 6828 3528
rect 6595 3488 6828 3516
rect 6595 3485 6607 3488
rect 6549 3479 6607 3485
rect 6822 3476 6828 3488
rect 6880 3516 6886 3528
rect 7466 3516 7472 3528
rect 6880 3488 7472 3516
rect 6880 3476 6886 3488
rect 7466 3476 7472 3488
rect 7524 3476 7530 3528
rect 7561 3519 7619 3525
rect 7561 3485 7573 3519
rect 7607 3485 7619 3519
rect 8386 3516 8392 3528
rect 8347 3488 8392 3516
rect 7561 3479 7619 3485
rect 5108 3451 5166 3457
rect 5108 3417 5120 3451
rect 5154 3448 5166 3451
rect 6362 3448 6368 3460
rect 5154 3420 6368 3448
rect 5154 3417 5166 3420
rect 5108 3411 5166 3417
rect 6362 3408 6368 3420
rect 6420 3408 6426 3460
rect 7098 3408 7104 3460
rect 7156 3448 7162 3460
rect 7576 3448 7604 3479
rect 8386 3476 8392 3488
rect 8444 3476 8450 3528
rect 8478 3476 8484 3528
rect 8536 3516 8542 3528
rect 8573 3519 8631 3525
rect 8573 3516 8585 3519
rect 8536 3488 8585 3516
rect 8536 3476 8542 3488
rect 8573 3485 8585 3488
rect 8619 3485 8631 3519
rect 8573 3479 8631 3485
rect 9309 3519 9367 3525
rect 9309 3485 9321 3519
rect 9355 3516 9367 3519
rect 9674 3516 9680 3528
rect 9355 3488 9680 3516
rect 9355 3485 9367 3488
rect 9309 3479 9367 3485
rect 9674 3476 9680 3488
rect 9732 3476 9738 3528
rect 9968 3525 9996 3556
rect 11790 3544 11796 3596
rect 11848 3584 11854 3596
rect 13280 3584 13308 3624
rect 16485 3621 16497 3655
rect 16531 3652 16543 3655
rect 18138 3652 18144 3664
rect 16531 3624 18144 3652
rect 16531 3621 16543 3624
rect 16485 3615 16543 3621
rect 18138 3612 18144 3624
rect 18196 3612 18202 3664
rect 13722 3584 13728 3596
rect 11848 3556 13216 3584
rect 13280 3556 13728 3584
rect 11848 3544 11854 3556
rect 9953 3519 10011 3525
rect 9953 3485 9965 3519
rect 9999 3485 10011 3519
rect 9953 3479 10011 3485
rect 10137 3519 10195 3525
rect 10137 3485 10149 3519
rect 10183 3485 10195 3519
rect 11238 3516 11244 3528
rect 11199 3488 11244 3516
rect 10137 3479 10195 3485
rect 7156 3420 7604 3448
rect 7837 3451 7895 3457
rect 7156 3408 7162 3420
rect 7837 3417 7849 3451
rect 7883 3448 7895 3451
rect 7926 3448 7932 3460
rect 7883 3420 7932 3448
rect 7883 3417 7895 3420
rect 7837 3411 7895 3417
rect 7926 3408 7932 3420
rect 7984 3448 7990 3460
rect 10152 3448 10180 3479
rect 11238 3476 11244 3488
rect 11296 3476 11302 3528
rect 12802 3476 12808 3528
rect 12860 3516 12866 3528
rect 12897 3519 12955 3525
rect 12897 3516 12909 3519
rect 12860 3488 12909 3516
rect 12860 3476 12866 3488
rect 12897 3485 12909 3488
rect 12943 3485 12955 3519
rect 12897 3479 12955 3485
rect 12986 3476 12992 3528
rect 13044 3516 13050 3528
rect 13188 3525 13216 3556
rect 13722 3544 13728 3556
rect 13780 3584 13786 3596
rect 13780 3556 18092 3584
rect 13780 3544 13786 3556
rect 13173 3519 13231 3525
rect 13044 3488 13089 3516
rect 13044 3476 13050 3488
rect 13173 3485 13185 3519
rect 13219 3485 13231 3519
rect 13173 3479 13231 3485
rect 13262 3476 13268 3528
rect 13320 3516 13326 3528
rect 13320 3488 13365 3516
rect 13320 3476 13326 3488
rect 13446 3476 13452 3528
rect 13504 3516 13510 3528
rect 18064 3525 18092 3556
rect 14277 3519 14335 3525
rect 14277 3516 14289 3519
rect 13504 3488 14289 3516
rect 13504 3476 13510 3488
rect 14277 3485 14289 3488
rect 14323 3485 14335 3519
rect 14277 3479 14335 3485
rect 15473 3519 15531 3525
rect 15473 3485 15485 3519
rect 15519 3485 15531 3519
rect 15473 3479 15531 3485
rect 16209 3519 16267 3525
rect 16209 3485 16221 3519
rect 16255 3516 16267 3519
rect 18049 3519 18107 3525
rect 16255 3488 17172 3516
rect 16255 3485 16267 3488
rect 16209 3479 16267 3485
rect 7984 3420 10180 3448
rect 7984 3408 7990 3420
rect 11330 3408 11336 3460
rect 11388 3448 11394 3460
rect 15488 3448 15516 3479
rect 17144 3460 17172 3488
rect 18049 3485 18061 3519
rect 18095 3485 18107 3519
rect 18049 3479 18107 3485
rect 11388 3420 15516 3448
rect 16485 3451 16543 3457
rect 11388 3408 11394 3420
rect 16485 3417 16497 3451
rect 16531 3448 16543 3451
rect 16574 3448 16580 3460
rect 16531 3420 16580 3448
rect 16531 3417 16543 3420
rect 16485 3411 16543 3417
rect 16574 3408 16580 3420
rect 16632 3408 16638 3460
rect 16942 3448 16948 3460
rect 16903 3420 16948 3448
rect 16942 3408 16948 3420
rect 17000 3408 17006 3460
rect 17126 3408 17132 3460
rect 17184 3457 17190 3460
rect 17184 3451 17203 3457
rect 17191 3417 17203 3451
rect 17184 3411 17203 3417
rect 17184 3408 17190 3411
rect 3970 3380 3976 3392
rect 3931 3352 3976 3380
rect 3970 3340 3976 3352
rect 4028 3340 4034 3392
rect 6733 3383 6791 3389
rect 6733 3349 6745 3383
rect 6779 3380 6791 3383
rect 6914 3380 6920 3392
rect 6779 3352 6920 3380
rect 6779 3349 6791 3352
rect 6733 3343 6791 3349
rect 6914 3340 6920 3352
rect 6972 3340 6978 3392
rect 10045 3383 10103 3389
rect 10045 3349 10057 3383
rect 10091 3380 10103 3383
rect 10318 3380 10324 3392
rect 10091 3352 10324 3380
rect 10091 3349 10103 3352
rect 10045 3343 10103 3349
rect 10318 3340 10324 3352
rect 10376 3340 10382 3392
rect 11146 3340 11152 3392
rect 11204 3380 11210 3392
rect 11425 3383 11483 3389
rect 11425 3380 11437 3383
rect 11204 3352 11437 3380
rect 11204 3340 11210 3352
rect 11425 3349 11437 3352
rect 11471 3349 11483 3383
rect 11425 3343 11483 3349
rect 11790 3340 11796 3392
rect 11848 3380 11854 3392
rect 12161 3383 12219 3389
rect 12161 3380 12173 3383
rect 11848 3352 12173 3380
rect 11848 3340 11854 3352
rect 12161 3349 12173 3352
rect 12207 3349 12219 3383
rect 12710 3380 12716 3392
rect 12671 3352 12716 3380
rect 12161 3343 12219 3349
rect 12710 3340 12716 3352
rect 12768 3340 12774 3392
rect 13630 3340 13636 3392
rect 13688 3380 13694 3392
rect 14461 3383 14519 3389
rect 14461 3380 14473 3383
rect 13688 3352 14473 3380
rect 13688 3340 13694 3352
rect 14461 3349 14473 3352
rect 14507 3349 14519 3383
rect 14461 3343 14519 3349
rect 15657 3383 15715 3389
rect 15657 3349 15669 3383
rect 15703 3380 15715 3383
rect 16114 3380 16120 3392
rect 15703 3352 16120 3380
rect 15703 3349 15715 3352
rect 15657 3343 15715 3349
rect 16114 3340 16120 3352
rect 16172 3340 16178 3392
rect 16301 3383 16359 3389
rect 16301 3349 16313 3383
rect 16347 3380 16359 3383
rect 16960 3380 16988 3408
rect 16347 3352 16988 3380
rect 17313 3383 17371 3389
rect 16347 3349 16359 3352
rect 16301 3343 16359 3349
rect 17313 3349 17325 3383
rect 17359 3380 17371 3383
rect 17402 3380 17408 3392
rect 17359 3352 17408 3380
rect 17359 3349 17371 3352
rect 17313 3343 17371 3349
rect 17402 3340 17408 3352
rect 17460 3340 17466 3392
rect 18233 3383 18291 3389
rect 18233 3349 18245 3383
rect 18279 3380 18291 3383
rect 18598 3380 18604 3392
rect 18279 3352 18604 3380
rect 18279 3349 18291 3352
rect 18233 3343 18291 3349
rect 18598 3340 18604 3352
rect 18656 3340 18662 3392
rect 1104 3290 19019 3312
rect 1104 3238 5388 3290
rect 5440 3238 5452 3290
rect 5504 3238 5516 3290
rect 5568 3238 5580 3290
rect 5632 3238 5644 3290
rect 5696 3238 9827 3290
rect 9879 3238 9891 3290
rect 9943 3238 9955 3290
rect 10007 3238 10019 3290
rect 10071 3238 10083 3290
rect 10135 3238 14266 3290
rect 14318 3238 14330 3290
rect 14382 3238 14394 3290
rect 14446 3238 14458 3290
rect 14510 3238 14522 3290
rect 14574 3238 18705 3290
rect 18757 3238 18769 3290
rect 18821 3238 18833 3290
rect 18885 3238 18897 3290
rect 18949 3238 18961 3290
rect 19013 3238 19019 3290
rect 1104 3216 19019 3238
rect 6362 3136 6368 3188
rect 6420 3176 6426 3188
rect 6549 3179 6607 3185
rect 6549 3176 6561 3179
rect 6420 3148 6561 3176
rect 6420 3136 6426 3148
rect 6549 3145 6561 3148
rect 6595 3145 6607 3179
rect 7098 3176 7104 3188
rect 6549 3139 6607 3145
rect 6748 3148 7104 3176
rect 5258 3108 5264 3120
rect 2792 3080 5264 3108
rect 2792 3049 2820 3080
rect 2777 3043 2835 3049
rect 2777 3009 2789 3043
rect 2823 3009 2835 3043
rect 2777 3003 2835 3009
rect 3044 3043 3102 3049
rect 3044 3009 3056 3043
rect 3090 3040 3102 3043
rect 4522 3040 4528 3052
rect 3090 3012 4528 3040
rect 3090 3009 3102 3012
rect 3044 3003 3102 3009
rect 4522 3000 4528 3012
rect 4580 3000 4586 3052
rect 4632 3049 4660 3080
rect 5258 3068 5264 3080
rect 5316 3068 5322 3120
rect 4617 3043 4675 3049
rect 4617 3009 4629 3043
rect 4663 3009 4675 3043
rect 4617 3003 4675 3009
rect 4706 3000 4712 3052
rect 4764 3040 4770 3052
rect 6748 3049 6776 3148
rect 7098 3136 7104 3148
rect 7156 3176 7162 3188
rect 7374 3176 7380 3188
rect 7156 3148 7380 3176
rect 7156 3136 7162 3148
rect 7374 3136 7380 3148
rect 7432 3136 7438 3188
rect 11149 3179 11207 3185
rect 11149 3145 11161 3179
rect 11195 3176 11207 3179
rect 11330 3176 11336 3188
rect 11195 3148 11336 3176
rect 11195 3145 11207 3148
rect 11149 3139 11207 3145
rect 11330 3136 11336 3148
rect 11388 3136 11394 3188
rect 13081 3179 13139 3185
rect 13081 3145 13093 3179
rect 13127 3176 13139 3179
rect 13446 3176 13452 3188
rect 13127 3148 13452 3176
rect 13127 3145 13139 3148
rect 13081 3139 13139 3145
rect 13446 3136 13452 3148
rect 13504 3136 13510 3188
rect 15381 3179 15439 3185
rect 15381 3145 15393 3179
rect 15427 3176 15439 3179
rect 17218 3176 17224 3188
rect 15427 3148 16712 3176
rect 17179 3148 17224 3176
rect 15427 3145 15439 3148
rect 15381 3139 15439 3145
rect 6914 3068 6920 3120
rect 6972 3108 6978 3120
rect 7990 3111 8048 3117
rect 7990 3108 8002 3111
rect 6972 3080 8002 3108
rect 6972 3068 6978 3080
rect 7990 3077 8002 3080
rect 8036 3077 8048 3111
rect 16301 3111 16359 3117
rect 7990 3071 8048 3077
rect 9784 3080 10640 3108
rect 4873 3043 4931 3049
rect 4873 3040 4885 3043
rect 4764 3012 4885 3040
rect 4764 3000 4770 3012
rect 4873 3009 4885 3012
rect 4919 3009 4931 3043
rect 4873 3003 4931 3009
rect 6733 3043 6791 3049
rect 6733 3009 6745 3043
rect 6779 3009 6791 3043
rect 6733 3003 6791 3009
rect 6825 3043 6883 3049
rect 6825 3009 6837 3043
rect 6871 3009 6883 3043
rect 7006 3040 7012 3052
rect 6967 3012 7012 3040
rect 6825 3003 6883 3009
rect 6546 2932 6552 2984
rect 6604 2972 6610 2984
rect 6840 2972 6868 3003
rect 7006 3000 7012 3012
rect 7064 3000 7070 3052
rect 7101 3043 7159 3049
rect 7101 3009 7113 3043
rect 7147 3009 7159 3043
rect 7101 3003 7159 3009
rect 6604 2944 6868 2972
rect 6604 2932 6610 2944
rect 4157 2839 4215 2845
rect 4157 2805 4169 2839
rect 4203 2836 4215 2839
rect 4246 2836 4252 2848
rect 4203 2808 4252 2836
rect 4203 2805 4215 2808
rect 4157 2799 4215 2805
rect 4246 2796 4252 2808
rect 4304 2796 4310 2848
rect 5994 2836 6000 2848
rect 5955 2808 6000 2836
rect 5994 2796 6000 2808
rect 6052 2796 6058 2848
rect 6178 2796 6184 2848
rect 6236 2836 6242 2848
rect 7116 2836 7144 3003
rect 7190 3000 7196 3052
rect 7248 3040 7254 3052
rect 7745 3043 7803 3049
rect 7745 3040 7757 3043
rect 7248 3012 7757 3040
rect 7248 3000 7254 3012
rect 7745 3009 7757 3012
rect 7791 3009 7803 3043
rect 7745 3003 7803 3009
rect 9306 3000 9312 3052
rect 9364 3040 9370 3052
rect 9784 3049 9812 3080
rect 9769 3043 9827 3049
rect 9769 3040 9781 3043
rect 9364 3012 9781 3040
rect 9364 3000 9370 3012
rect 9769 3009 9781 3012
rect 9815 3009 9827 3043
rect 9769 3003 9827 3009
rect 10036 3043 10094 3049
rect 10036 3009 10048 3043
rect 10082 3040 10094 3043
rect 10318 3040 10324 3052
rect 10082 3012 10324 3040
rect 10082 3009 10094 3012
rect 10036 3003 10094 3009
rect 10318 3000 10324 3012
rect 10376 3000 10382 3052
rect 10612 3040 10640 3080
rect 16301 3077 16313 3111
rect 16347 3108 16359 3111
rect 16574 3108 16580 3120
rect 16347 3080 16580 3108
rect 16347 3077 16359 3080
rect 16301 3071 16359 3077
rect 16574 3068 16580 3080
rect 16632 3068 16638 3120
rect 16684 3108 16712 3148
rect 17218 3136 17224 3148
rect 17276 3136 17282 3188
rect 17310 3108 17316 3120
rect 16684 3080 17316 3108
rect 17310 3068 17316 3080
rect 17368 3068 17374 3120
rect 17862 3068 17868 3120
rect 17920 3108 17926 3120
rect 18325 3111 18383 3117
rect 18325 3108 18337 3111
rect 17920 3080 18337 3108
rect 17920 3068 17926 3080
rect 18325 3077 18337 3080
rect 18371 3077 18383 3111
rect 18325 3071 18383 3077
rect 11698 3040 11704 3052
rect 10612 3012 11704 3040
rect 11698 3000 11704 3012
rect 11756 3000 11762 3052
rect 11957 3043 12015 3049
rect 11957 3040 11969 3043
rect 11808 3012 11969 3040
rect 11054 2932 11060 2984
rect 11112 2972 11118 2984
rect 11808 2972 11836 3012
rect 11957 3009 11969 3012
rect 12003 3009 12015 3043
rect 13998 3040 14004 3052
rect 13959 3012 14004 3040
rect 11957 3003 12015 3009
rect 13998 3000 14004 3012
rect 14056 3000 14062 3052
rect 14268 3043 14326 3049
rect 14268 3009 14280 3043
rect 14314 3040 14326 3043
rect 15746 3040 15752 3052
rect 14314 3012 15752 3040
rect 14314 3009 14326 3012
rect 14268 3003 14326 3009
rect 15746 3000 15752 3012
rect 15804 3000 15810 3052
rect 15930 3040 15936 3052
rect 15891 3012 15936 3040
rect 15930 3000 15936 3012
rect 15988 3000 15994 3052
rect 16117 3043 16175 3049
rect 16117 3009 16129 3043
rect 16163 3040 16175 3043
rect 17034 3040 17040 3052
rect 16163 3012 17040 3040
rect 16163 3009 16175 3012
rect 16117 3003 16175 3009
rect 17034 3000 17040 3012
rect 17092 3000 17098 3052
rect 18049 3043 18107 3049
rect 18049 3040 18061 3043
rect 17420 3012 18061 3040
rect 17420 2984 17448 3012
rect 18049 3009 18061 3012
rect 18095 3009 18107 3043
rect 18049 3003 18107 3009
rect 18138 3000 18144 3052
rect 18196 3040 18202 3052
rect 18196 3012 18241 3040
rect 18196 3000 18202 3012
rect 11112 2944 11836 2972
rect 11112 2932 11118 2944
rect 17402 2932 17408 2984
rect 17460 2972 17466 2984
rect 17460 2944 17505 2972
rect 17460 2932 17466 2944
rect 6236 2808 7144 2836
rect 6236 2796 6242 2808
rect 8662 2796 8668 2848
rect 8720 2836 8726 2848
rect 9125 2839 9183 2845
rect 9125 2836 9137 2839
rect 8720 2808 9137 2836
rect 8720 2796 8726 2808
rect 9125 2805 9137 2808
rect 9171 2805 9183 2839
rect 16850 2836 16856 2848
rect 16811 2808 16856 2836
rect 9125 2799 9183 2805
rect 16850 2796 16856 2808
rect 16908 2796 16914 2848
rect 18046 2836 18052 2848
rect 18007 2808 18052 2836
rect 18046 2796 18052 2808
rect 18104 2796 18110 2848
rect 1104 2746 18860 2768
rect 1104 2694 3169 2746
rect 3221 2694 3233 2746
rect 3285 2694 3297 2746
rect 3349 2694 3361 2746
rect 3413 2694 3425 2746
rect 3477 2694 7608 2746
rect 7660 2694 7672 2746
rect 7724 2694 7736 2746
rect 7788 2694 7800 2746
rect 7852 2694 7864 2746
rect 7916 2694 12047 2746
rect 12099 2694 12111 2746
rect 12163 2694 12175 2746
rect 12227 2694 12239 2746
rect 12291 2694 12303 2746
rect 12355 2694 16486 2746
rect 16538 2694 16550 2746
rect 16602 2694 16614 2746
rect 16666 2694 16678 2746
rect 16730 2694 16742 2746
rect 16794 2694 18860 2746
rect 1104 2672 18860 2694
rect 4522 2592 4528 2644
rect 4580 2632 4586 2644
rect 5169 2635 5227 2641
rect 5169 2632 5181 2635
rect 4580 2604 5181 2632
rect 4580 2592 4586 2604
rect 5169 2601 5181 2604
rect 5215 2601 5227 2635
rect 5169 2595 5227 2601
rect 7561 2635 7619 2641
rect 7561 2601 7573 2635
rect 7607 2632 7619 2635
rect 10505 2635 10563 2641
rect 7607 2604 10088 2632
rect 7607 2601 7619 2604
rect 7561 2595 7619 2601
rect 6454 2564 6460 2576
rect 5092 2536 6460 2564
rect 1857 2431 1915 2437
rect 1857 2397 1869 2431
rect 1903 2428 1915 2431
rect 3970 2428 3976 2440
rect 1903 2400 3976 2428
rect 1903 2397 1915 2400
rect 1857 2391 1915 2397
rect 3970 2388 3976 2400
rect 4028 2388 4034 2440
rect 4246 2428 4252 2440
rect 4207 2400 4252 2428
rect 4246 2388 4252 2400
rect 4304 2388 4310 2440
rect 5092 2437 5120 2536
rect 6454 2524 6460 2536
rect 6512 2564 6518 2576
rect 6733 2567 6791 2573
rect 6733 2564 6745 2567
rect 6512 2536 6745 2564
rect 6512 2524 6518 2536
rect 6733 2533 6745 2536
rect 6779 2533 6791 2567
rect 10060 2564 10088 2604
rect 10505 2601 10517 2635
rect 10551 2632 10563 2635
rect 11238 2632 11244 2644
rect 10551 2604 11244 2632
rect 10551 2601 10563 2604
rect 10505 2595 10563 2601
rect 11238 2592 11244 2604
rect 11296 2592 11302 2644
rect 11790 2632 11796 2644
rect 11751 2604 11796 2632
rect 11790 2592 11796 2604
rect 11848 2632 11854 2644
rect 13633 2635 13691 2641
rect 11848 2604 13584 2632
rect 11848 2592 11854 2604
rect 11054 2564 11060 2576
rect 10060 2536 11060 2564
rect 6733 2527 6791 2533
rect 11054 2524 11060 2536
rect 11112 2524 11118 2576
rect 13556 2564 13584 2604
rect 13633 2601 13645 2635
rect 13679 2632 13691 2635
rect 13722 2632 13728 2644
rect 13679 2604 13728 2632
rect 13679 2601 13691 2604
rect 13633 2595 13691 2601
rect 13722 2592 13728 2604
rect 13780 2592 13786 2644
rect 15657 2635 15715 2641
rect 14292 2604 15332 2632
rect 14292 2564 14320 2604
rect 13556 2536 14320 2564
rect 6914 2496 6920 2508
rect 5276 2468 6920 2496
rect 5276 2437 5304 2468
rect 6914 2456 6920 2468
rect 6972 2496 6978 2508
rect 13998 2496 14004 2508
rect 6972 2468 7512 2496
rect 6972 2456 6978 2468
rect 5077 2431 5135 2437
rect 5077 2397 5089 2431
rect 5123 2397 5135 2431
rect 5077 2391 5135 2397
rect 5261 2431 5319 2437
rect 5261 2397 5273 2431
rect 5307 2397 5319 2431
rect 5994 2428 6000 2440
rect 5955 2400 6000 2428
rect 5261 2391 5319 2397
rect 5994 2388 6000 2400
rect 6052 2388 6058 2440
rect 6546 2428 6552 2440
rect 6507 2400 6552 2428
rect 6546 2388 6552 2400
rect 6604 2388 6610 2440
rect 6730 2388 6736 2440
rect 6788 2428 6794 2440
rect 7484 2437 7512 2468
rect 13832 2468 14004 2496
rect 7009 2431 7067 2437
rect 7009 2428 7021 2431
rect 6788 2400 7021 2428
rect 6788 2388 6794 2400
rect 7009 2397 7021 2400
rect 7055 2397 7067 2431
rect 7009 2391 7067 2397
rect 7469 2431 7527 2437
rect 7469 2397 7481 2431
rect 7515 2397 7527 2431
rect 7469 2391 7527 2397
rect 7653 2431 7711 2437
rect 7653 2397 7665 2431
rect 7699 2428 7711 2431
rect 7926 2428 7932 2440
rect 7699 2400 7932 2428
rect 7699 2397 7711 2400
rect 7653 2391 7711 2397
rect 7926 2388 7932 2400
rect 7984 2388 7990 2440
rect 8573 2431 8631 2437
rect 8573 2397 8585 2431
rect 8619 2428 8631 2431
rect 8662 2428 8668 2440
rect 8619 2400 8668 2428
rect 8619 2397 8631 2400
rect 8573 2391 8631 2397
rect 8662 2388 8668 2400
rect 8720 2388 8726 2440
rect 9125 2431 9183 2437
rect 9125 2397 9137 2431
rect 9171 2428 9183 2431
rect 9214 2428 9220 2440
rect 9171 2400 9220 2428
rect 9171 2397 9183 2400
rect 9125 2391 9183 2397
rect 9214 2388 9220 2400
rect 9272 2388 9278 2440
rect 11698 2388 11704 2440
rect 11756 2428 11762 2440
rect 12253 2431 12311 2437
rect 12253 2428 12265 2431
rect 11756 2400 12265 2428
rect 11756 2388 11762 2400
rect 12253 2397 12265 2400
rect 12299 2428 12311 2431
rect 13832 2428 13860 2468
rect 13998 2456 14004 2468
rect 14056 2496 14062 2508
rect 14277 2499 14335 2505
rect 14277 2496 14289 2499
rect 14056 2468 14289 2496
rect 14056 2456 14062 2468
rect 14277 2465 14289 2468
rect 14323 2465 14335 2499
rect 14277 2459 14335 2465
rect 12299 2400 13860 2428
rect 15304 2428 15332 2604
rect 15657 2601 15669 2635
rect 15703 2632 15715 2635
rect 15930 2632 15936 2644
rect 15703 2604 15936 2632
rect 15703 2601 15715 2604
rect 15657 2595 15715 2601
rect 15930 2592 15936 2604
rect 15988 2592 15994 2644
rect 16942 2592 16948 2644
rect 17000 2632 17006 2644
rect 17313 2635 17371 2641
rect 17313 2632 17325 2635
rect 17000 2604 17325 2632
rect 17000 2592 17006 2604
rect 17313 2601 17325 2604
rect 17359 2632 17371 2635
rect 18141 2635 18199 2641
rect 18141 2632 18153 2635
rect 17359 2604 18153 2632
rect 17359 2601 17371 2604
rect 17313 2595 17371 2601
rect 18141 2601 18153 2604
rect 18187 2601 18199 2635
rect 18141 2595 18199 2601
rect 17218 2524 17224 2576
rect 17276 2564 17282 2576
rect 17681 2567 17739 2573
rect 17681 2564 17693 2567
rect 17276 2536 17693 2564
rect 17276 2524 17282 2536
rect 17681 2533 17693 2536
rect 17727 2533 17739 2567
rect 17681 2527 17739 2533
rect 15746 2456 15752 2508
rect 15804 2496 15810 2508
rect 16209 2499 16267 2505
rect 16209 2496 16221 2499
rect 15804 2468 16221 2496
rect 15804 2456 15810 2468
rect 16209 2465 16221 2468
rect 16255 2465 16267 2499
rect 16209 2459 16267 2465
rect 16117 2431 16175 2437
rect 16117 2428 16129 2431
rect 15304 2400 16129 2428
rect 12299 2397 12311 2400
rect 12253 2391 12311 2397
rect 16117 2397 16129 2400
rect 16163 2397 16175 2431
rect 16117 2391 16175 2397
rect 16301 2431 16359 2437
rect 16301 2397 16313 2431
rect 16347 2428 16359 2431
rect 16850 2428 16856 2440
rect 16347 2400 16856 2428
rect 16347 2397 16359 2400
rect 16301 2391 16359 2397
rect 16850 2388 16856 2400
rect 16908 2388 16914 2440
rect 17221 2431 17279 2437
rect 17221 2397 17233 2431
rect 17267 2428 17279 2431
rect 17310 2428 17316 2440
rect 17267 2400 17316 2428
rect 17267 2397 17279 2400
rect 17221 2391 17279 2397
rect 17310 2388 17316 2400
rect 17368 2388 17374 2440
rect 6917 2363 6975 2369
rect 6917 2329 6929 2363
rect 6963 2360 6975 2363
rect 7374 2360 7380 2372
rect 6963 2332 7380 2360
rect 6963 2329 6975 2332
rect 6917 2323 6975 2329
rect 7374 2320 7380 2332
rect 7432 2320 7438 2372
rect 9030 2320 9036 2372
rect 9088 2360 9094 2372
rect 9370 2363 9428 2369
rect 9370 2360 9382 2363
rect 9088 2332 9382 2360
rect 9088 2320 9094 2332
rect 9370 2329 9382 2332
rect 9416 2329 9428 2363
rect 9370 2323 9428 2329
rect 12520 2363 12578 2369
rect 12520 2329 12532 2363
rect 12566 2360 12578 2363
rect 12710 2360 12716 2372
rect 12566 2332 12716 2360
rect 12566 2329 12578 2332
rect 12520 2323 12578 2329
rect 12710 2320 12716 2332
rect 12768 2320 12774 2372
rect 14544 2363 14602 2369
rect 14544 2329 14556 2363
rect 14590 2360 14602 2363
rect 18046 2360 18052 2372
rect 14590 2332 18052 2360
rect 14590 2329 14602 2332
rect 14544 2323 14602 2329
rect 18046 2320 18052 2332
rect 18104 2320 18110 2372
rect 1210 2252 1216 2304
rect 1268 2292 1274 2304
rect 1673 2295 1731 2301
rect 1673 2292 1685 2295
rect 1268 2264 1685 2292
rect 1268 2252 1274 2264
rect 1673 2261 1685 2264
rect 1719 2261 1731 2295
rect 1673 2255 1731 2261
rect 3694 2252 3700 2304
rect 3752 2292 3758 2304
rect 4065 2295 4123 2301
rect 4065 2292 4077 2295
rect 3752 2264 4077 2292
rect 3752 2252 3758 2264
rect 4065 2261 4077 2264
rect 4111 2261 4123 2295
rect 4065 2255 4123 2261
rect 5813 2295 5871 2301
rect 5813 2261 5825 2295
rect 5859 2292 5871 2295
rect 6178 2292 6184 2304
rect 5859 2264 6184 2292
rect 5859 2261 5871 2264
rect 5813 2255 5871 2261
rect 6178 2252 6184 2264
rect 6236 2252 6242 2304
rect 8389 2295 8447 2301
rect 8389 2261 8401 2295
rect 8435 2292 8447 2295
rect 8662 2292 8668 2304
rect 8435 2264 8668 2292
rect 8435 2261 8447 2264
rect 8389 2255 8447 2261
rect 8662 2252 8668 2264
rect 8720 2252 8726 2304
rect 1104 2202 19019 2224
rect 1104 2150 5388 2202
rect 5440 2150 5452 2202
rect 5504 2150 5516 2202
rect 5568 2150 5580 2202
rect 5632 2150 5644 2202
rect 5696 2150 9827 2202
rect 9879 2150 9891 2202
rect 9943 2150 9955 2202
rect 10007 2150 10019 2202
rect 10071 2150 10083 2202
rect 10135 2150 14266 2202
rect 14318 2150 14330 2202
rect 14382 2150 14394 2202
rect 14446 2150 14458 2202
rect 14510 2150 14522 2202
rect 14574 2150 18705 2202
rect 18757 2150 18769 2202
rect 18821 2150 18833 2202
rect 18885 2150 18897 2202
rect 18949 2150 18961 2202
rect 19013 2150 19019 2202
rect 1104 2128 19019 2150
<< via1 >>
rect 5388 17382 5440 17434
rect 5452 17382 5504 17434
rect 5516 17382 5568 17434
rect 5580 17382 5632 17434
rect 5644 17382 5696 17434
rect 9827 17382 9879 17434
rect 9891 17382 9943 17434
rect 9955 17382 10007 17434
rect 10019 17382 10071 17434
rect 10083 17382 10135 17434
rect 14266 17382 14318 17434
rect 14330 17382 14382 17434
rect 14394 17382 14446 17434
rect 14458 17382 14510 17434
rect 14522 17382 14574 17434
rect 18705 17382 18757 17434
rect 18769 17382 18821 17434
rect 18833 17382 18885 17434
rect 18897 17382 18949 17434
rect 18961 17382 19013 17434
rect 16580 17280 16632 17332
rect 2780 17144 2832 17196
rect 6552 17144 6604 17196
rect 7196 17144 7248 17196
rect 9312 17187 9364 17196
rect 9312 17153 9321 17187
rect 9321 17153 9355 17187
rect 9355 17153 9364 17187
rect 9312 17144 9364 17153
rect 10140 17144 10192 17196
rect 5356 17119 5408 17128
rect 5356 17085 5365 17119
rect 5365 17085 5399 17119
rect 5399 17085 5408 17119
rect 5356 17076 5408 17085
rect 7104 17076 7156 17128
rect 10324 17144 10376 17196
rect 12624 17144 12676 17196
rect 4252 17008 4304 17060
rect 9864 17008 9916 17060
rect 3976 16983 4028 16992
rect 3976 16949 3985 16983
rect 3985 16949 4019 16983
rect 4019 16949 4028 16983
rect 3976 16940 4028 16949
rect 6000 16940 6052 16992
rect 7380 16983 7432 16992
rect 7380 16949 7389 16983
rect 7389 16949 7423 16983
rect 7423 16949 7432 16983
rect 7380 16940 7432 16949
rect 8944 16940 8996 16992
rect 10508 16940 10560 16992
rect 10600 16940 10652 16992
rect 16948 17076 17000 17128
rect 12808 16940 12860 16992
rect 3169 16838 3221 16890
rect 3233 16838 3285 16890
rect 3297 16838 3349 16890
rect 3361 16838 3413 16890
rect 3425 16838 3477 16890
rect 7608 16838 7660 16890
rect 7672 16838 7724 16890
rect 7736 16838 7788 16890
rect 7800 16838 7852 16890
rect 7864 16838 7916 16890
rect 12047 16838 12099 16890
rect 12111 16838 12163 16890
rect 12175 16838 12227 16890
rect 12239 16838 12291 16890
rect 12303 16838 12355 16890
rect 16486 16838 16538 16890
rect 16550 16838 16602 16890
rect 16614 16838 16666 16890
rect 16678 16838 16730 16890
rect 16742 16838 16794 16890
rect 2780 16779 2832 16788
rect 2780 16745 2789 16779
rect 2789 16745 2823 16779
rect 2823 16745 2832 16779
rect 7196 16779 7248 16788
rect 2780 16736 2832 16745
rect 7196 16745 7205 16779
rect 7205 16745 7239 16779
rect 7239 16745 7248 16779
rect 7196 16736 7248 16745
rect 10324 16736 10376 16788
rect 12624 16779 12676 16788
rect 12624 16745 12633 16779
rect 12633 16745 12667 16779
rect 12667 16745 12676 16779
rect 12624 16736 12676 16745
rect 3976 16532 4028 16584
rect 4988 16532 5040 16584
rect 5356 16575 5408 16584
rect 5356 16541 5365 16575
rect 5365 16541 5399 16575
rect 5399 16541 5408 16575
rect 5356 16532 5408 16541
rect 8576 16575 8628 16584
rect 8576 16541 8585 16575
rect 8585 16541 8619 16575
rect 8619 16541 8628 16575
rect 8576 16532 8628 16541
rect 5816 16464 5868 16516
rect 9864 16507 9916 16516
rect 3700 16396 3752 16448
rect 6920 16396 6972 16448
rect 9864 16473 9873 16507
rect 9873 16473 9907 16507
rect 9907 16473 9916 16507
rect 9864 16464 9916 16473
rect 10692 16507 10744 16516
rect 10692 16473 10726 16507
rect 10726 16473 10744 16507
rect 10692 16464 10744 16473
rect 10600 16396 10652 16448
rect 12808 16464 12860 16516
rect 5388 16294 5440 16346
rect 5452 16294 5504 16346
rect 5516 16294 5568 16346
rect 5580 16294 5632 16346
rect 5644 16294 5696 16346
rect 9827 16294 9879 16346
rect 9891 16294 9943 16346
rect 9955 16294 10007 16346
rect 10019 16294 10071 16346
rect 10083 16294 10135 16346
rect 14266 16294 14318 16346
rect 14330 16294 14382 16346
rect 14394 16294 14446 16346
rect 14458 16294 14510 16346
rect 14522 16294 14574 16346
rect 18705 16294 18757 16346
rect 18769 16294 18821 16346
rect 18833 16294 18885 16346
rect 18897 16294 18949 16346
rect 18961 16294 19013 16346
rect 5816 16235 5868 16244
rect 5816 16201 5825 16235
rect 5825 16201 5859 16235
rect 5859 16201 5868 16235
rect 5816 16192 5868 16201
rect 6552 16235 6604 16244
rect 6552 16201 6561 16235
rect 6561 16201 6595 16235
rect 6595 16201 6604 16235
rect 6552 16192 6604 16201
rect 4252 16167 4304 16176
rect 7380 16192 7432 16244
rect 9312 16192 9364 16244
rect 10232 16192 10284 16244
rect 10692 16235 10744 16244
rect 10692 16201 10701 16235
rect 10701 16201 10735 16235
rect 10735 16201 10744 16235
rect 10692 16192 10744 16201
rect 4252 16133 4270 16167
rect 4270 16133 4304 16167
rect 4252 16124 4304 16133
rect 3700 16056 3752 16108
rect 6920 16167 6972 16176
rect 6920 16133 6929 16167
rect 6929 16133 6963 16167
rect 6963 16133 6972 16167
rect 6920 16124 6972 16133
rect 8576 16124 8628 16176
rect 6000 16099 6052 16108
rect 6000 16065 6009 16099
rect 6009 16065 6043 16099
rect 6043 16065 6052 16099
rect 6000 16056 6052 16065
rect 8024 16099 8076 16108
rect 8024 16065 8033 16099
rect 8033 16065 8067 16099
rect 8067 16065 8076 16099
rect 8024 16056 8076 16065
rect 9128 16124 9180 16176
rect 8944 16099 8996 16108
rect 8944 16065 8978 16099
rect 8978 16065 8996 16099
rect 8944 16056 8996 16065
rect 10508 16099 10560 16108
rect 10508 16065 10517 16099
rect 10517 16065 10551 16099
rect 10551 16065 10560 16099
rect 10508 16056 10560 16065
rect 11704 16056 11756 16108
rect 12440 16192 12492 16244
rect 4988 15988 5040 16040
rect 7104 15988 7156 16040
rect 12256 16099 12308 16108
rect 12256 16065 12265 16099
rect 12265 16065 12299 16099
rect 12299 16065 12308 16099
rect 12256 16056 12308 16065
rect 11796 15920 11848 15972
rect 12256 15920 12308 15972
rect 13728 16031 13780 16040
rect 13728 15997 13737 16031
rect 13737 15997 13771 16031
rect 13771 15997 13780 16031
rect 13728 15988 13780 15997
rect 3056 15852 3108 15904
rect 3516 15852 3568 15904
rect 8668 15852 8720 15904
rect 17132 15852 17184 15904
rect 3169 15750 3221 15802
rect 3233 15750 3285 15802
rect 3297 15750 3349 15802
rect 3361 15750 3413 15802
rect 3425 15750 3477 15802
rect 7608 15750 7660 15802
rect 7672 15750 7724 15802
rect 7736 15750 7788 15802
rect 7800 15750 7852 15802
rect 7864 15750 7916 15802
rect 12047 15750 12099 15802
rect 12111 15750 12163 15802
rect 12175 15750 12227 15802
rect 12239 15750 12291 15802
rect 12303 15750 12355 15802
rect 16486 15750 16538 15802
rect 16550 15750 16602 15802
rect 16614 15750 16666 15802
rect 16678 15750 16730 15802
rect 16742 15750 16794 15802
rect 12440 15648 12492 15700
rect 3056 15444 3108 15496
rect 4160 15487 4212 15496
rect 4160 15453 4169 15487
rect 4169 15453 4203 15487
rect 4203 15453 4212 15487
rect 4160 15444 4212 15453
rect 4252 15487 4304 15496
rect 4252 15453 4261 15487
rect 4261 15453 4295 15487
rect 4295 15453 4304 15487
rect 4252 15444 4304 15453
rect 4988 15444 5040 15496
rect 9128 15444 9180 15496
rect 11428 15444 11480 15496
rect 6460 15376 6512 15428
rect 7472 15376 7524 15428
rect 13268 15444 13320 15496
rect 2780 15308 2832 15360
rect 3976 15351 4028 15360
rect 3976 15317 3985 15351
rect 3985 15317 4019 15351
rect 4019 15317 4028 15351
rect 3976 15308 4028 15317
rect 6828 15308 6880 15360
rect 8024 15308 8076 15360
rect 9680 15308 9732 15360
rect 15844 15376 15896 15428
rect 10876 15351 10928 15360
rect 10876 15317 10885 15351
rect 10885 15317 10919 15351
rect 10919 15317 10928 15351
rect 10876 15308 10928 15317
rect 14648 15308 14700 15360
rect 15752 15351 15804 15360
rect 15752 15317 15761 15351
rect 15761 15317 15795 15351
rect 15795 15317 15804 15351
rect 15752 15308 15804 15317
rect 5388 15206 5440 15258
rect 5452 15206 5504 15258
rect 5516 15206 5568 15258
rect 5580 15206 5632 15258
rect 5644 15206 5696 15258
rect 9827 15206 9879 15258
rect 9891 15206 9943 15258
rect 9955 15206 10007 15258
rect 10019 15206 10071 15258
rect 10083 15206 10135 15258
rect 14266 15206 14318 15258
rect 14330 15206 14382 15258
rect 14394 15206 14446 15258
rect 14458 15206 14510 15258
rect 14522 15206 14574 15258
rect 18705 15206 18757 15258
rect 18769 15206 18821 15258
rect 18833 15206 18885 15258
rect 18897 15206 18949 15258
rect 18961 15206 19013 15258
rect 4160 15104 4212 15156
rect 7472 15147 7524 15156
rect 7472 15113 7481 15147
rect 7481 15113 7515 15147
rect 7515 15113 7524 15147
rect 7472 15104 7524 15113
rect 9680 15104 9732 15156
rect 15844 15147 15896 15156
rect 4988 15036 5040 15088
rect 15844 15113 15853 15147
rect 15853 15113 15887 15147
rect 15887 15113 15896 15147
rect 15844 15104 15896 15113
rect 3056 14968 3108 15020
rect 4252 14968 4304 15020
rect 6828 15011 6880 15020
rect 6828 14977 6837 15011
rect 6837 14977 6871 15011
rect 6871 14977 6880 15011
rect 6828 14968 6880 14977
rect 9680 14968 9732 15020
rect 10232 14968 10284 15020
rect 10876 15011 10928 15020
rect 10876 14977 10885 15011
rect 10885 14977 10919 15011
rect 10919 14977 10928 15011
rect 10876 14968 10928 14977
rect 7104 14900 7156 14952
rect 9128 14900 9180 14952
rect 13820 15036 13872 15088
rect 12532 14968 12584 15020
rect 14924 14968 14976 15020
rect 13820 14943 13872 14952
rect 13820 14909 13829 14943
rect 13829 14909 13863 14943
rect 13863 14909 13872 14943
rect 13820 14900 13872 14909
rect 16212 14968 16264 15020
rect 16948 15011 17000 15020
rect 16948 14977 16957 15011
rect 16957 14977 16991 15011
rect 16991 14977 17000 15011
rect 16948 14968 17000 14977
rect 17132 15079 17184 15088
rect 17132 15045 17141 15079
rect 17141 15045 17175 15079
rect 17175 15045 17184 15079
rect 17132 15036 17184 15045
rect 17316 14968 17368 15020
rect 17684 14900 17736 14952
rect 5816 14764 5868 14816
rect 8392 14764 8444 14816
rect 10784 14807 10836 14816
rect 10784 14773 10793 14807
rect 10793 14773 10827 14807
rect 10827 14773 10836 14807
rect 10784 14764 10836 14773
rect 13268 14764 13320 14816
rect 16948 14764 17000 14816
rect 3169 14662 3221 14714
rect 3233 14662 3285 14714
rect 3297 14662 3349 14714
rect 3361 14662 3413 14714
rect 3425 14662 3477 14714
rect 7608 14662 7660 14714
rect 7672 14662 7724 14714
rect 7736 14662 7788 14714
rect 7800 14662 7852 14714
rect 7864 14662 7916 14714
rect 12047 14662 12099 14714
rect 12111 14662 12163 14714
rect 12175 14662 12227 14714
rect 12239 14662 12291 14714
rect 12303 14662 12355 14714
rect 16486 14662 16538 14714
rect 16550 14662 16602 14714
rect 16614 14662 16666 14714
rect 16678 14662 16730 14714
rect 16742 14662 16794 14714
rect 6460 14603 6512 14612
rect 6460 14569 6469 14603
rect 6469 14569 6503 14603
rect 6503 14569 6512 14603
rect 6460 14560 6512 14569
rect 7104 14560 7156 14612
rect 11704 14560 11756 14612
rect 12532 14560 12584 14612
rect 16856 14560 16908 14612
rect 5724 14492 5776 14544
rect 3976 14356 4028 14408
rect 4988 14356 5040 14408
rect 6000 14399 6052 14408
rect 6000 14365 6009 14399
rect 6009 14365 6043 14399
rect 6043 14365 6052 14399
rect 6000 14356 6052 14365
rect 6276 14399 6328 14408
rect 6276 14365 6285 14399
rect 6285 14365 6319 14399
rect 6319 14365 6328 14399
rect 6276 14356 6328 14365
rect 8300 14356 8352 14408
rect 9128 14399 9180 14408
rect 9128 14365 9137 14399
rect 9137 14365 9171 14399
rect 9171 14365 9180 14399
rect 9128 14356 9180 14365
rect 15384 14492 15436 14544
rect 11704 14399 11756 14408
rect 11704 14365 11713 14399
rect 11713 14365 11747 14399
rect 11747 14365 11756 14399
rect 11704 14356 11756 14365
rect 12624 14424 12676 14476
rect 16212 14467 16264 14476
rect 16212 14433 16221 14467
rect 16221 14433 16255 14467
rect 16255 14433 16264 14467
rect 16212 14424 16264 14433
rect 16396 14467 16448 14476
rect 16396 14433 16405 14467
rect 16405 14433 16439 14467
rect 16439 14433 16448 14467
rect 16396 14424 16448 14433
rect 16948 14424 17000 14476
rect 17408 14424 17460 14476
rect 13268 14399 13320 14408
rect 7012 14288 7064 14340
rect 9220 14288 9272 14340
rect 10416 14288 10468 14340
rect 7932 14220 7984 14272
rect 10508 14263 10560 14272
rect 10508 14229 10517 14263
rect 10517 14229 10551 14263
rect 10551 14229 10560 14263
rect 10508 14220 10560 14229
rect 13268 14365 13277 14399
rect 13277 14365 13311 14399
rect 13311 14365 13320 14399
rect 13268 14356 13320 14365
rect 14648 14399 14700 14408
rect 14648 14365 14657 14399
rect 14657 14365 14691 14399
rect 14691 14365 14700 14399
rect 14648 14356 14700 14365
rect 15844 14356 15896 14408
rect 17316 14331 17368 14340
rect 14096 14220 14148 14272
rect 14832 14263 14884 14272
rect 14832 14229 14841 14263
rect 14841 14229 14875 14263
rect 14875 14229 14884 14263
rect 14832 14220 14884 14229
rect 17316 14297 17325 14331
rect 17325 14297 17359 14331
rect 17359 14297 17368 14331
rect 17316 14288 17368 14297
rect 15844 14220 15896 14272
rect 16948 14263 17000 14272
rect 16948 14229 16957 14263
rect 16957 14229 16991 14263
rect 16991 14229 17000 14263
rect 16948 14220 17000 14229
rect 17040 14220 17092 14272
rect 17132 14220 17184 14272
rect 5388 14118 5440 14170
rect 5452 14118 5504 14170
rect 5516 14118 5568 14170
rect 5580 14118 5632 14170
rect 5644 14118 5696 14170
rect 9827 14118 9879 14170
rect 9891 14118 9943 14170
rect 9955 14118 10007 14170
rect 10019 14118 10071 14170
rect 10083 14118 10135 14170
rect 14266 14118 14318 14170
rect 14330 14118 14382 14170
rect 14394 14118 14446 14170
rect 14458 14118 14510 14170
rect 14522 14118 14574 14170
rect 18705 14118 18757 14170
rect 18769 14118 18821 14170
rect 18833 14118 18885 14170
rect 18897 14118 18949 14170
rect 18961 14118 19013 14170
rect 6276 14016 6328 14068
rect 7012 14059 7064 14068
rect 7012 14025 7021 14059
rect 7021 14025 7055 14059
rect 7055 14025 7064 14059
rect 7012 14016 7064 14025
rect 9220 14059 9272 14068
rect 9220 14025 9229 14059
rect 9229 14025 9263 14059
rect 9263 14025 9272 14059
rect 9220 14016 9272 14025
rect 9680 14016 9732 14068
rect 12624 14059 12676 14068
rect 12624 14025 12633 14059
rect 12633 14025 12667 14059
rect 12667 14025 12676 14059
rect 12624 14016 12676 14025
rect 14924 14059 14976 14068
rect 14924 14025 14933 14059
rect 14933 14025 14967 14059
rect 14967 14025 14976 14059
rect 14924 14016 14976 14025
rect 15476 14016 15528 14068
rect 17132 14016 17184 14068
rect 17960 14016 18012 14068
rect 2320 13923 2372 13932
rect 2320 13889 2329 13923
rect 2329 13889 2363 13923
rect 2363 13889 2372 13923
rect 2320 13880 2372 13889
rect 2688 13880 2740 13932
rect 2596 13855 2648 13864
rect 2596 13821 2605 13855
rect 2605 13821 2639 13855
rect 2639 13821 2648 13855
rect 6000 13948 6052 14000
rect 7104 13948 7156 14000
rect 4160 13923 4212 13932
rect 4160 13889 4178 13923
rect 4178 13889 4212 13923
rect 4160 13880 4212 13889
rect 4344 13880 4396 13932
rect 2596 13812 2648 13821
rect 4988 13812 5040 13864
rect 5724 13880 5776 13932
rect 7196 13880 7248 13932
rect 5816 13812 5868 13864
rect 7472 13923 7524 13932
rect 7472 13889 7481 13923
rect 7481 13889 7515 13923
rect 7515 13889 7524 13923
rect 7472 13880 7524 13889
rect 8760 13923 8812 13932
rect 8760 13889 8769 13923
rect 8769 13889 8803 13923
rect 8803 13889 8812 13923
rect 8760 13880 8812 13889
rect 9036 13923 9088 13932
rect 9036 13889 9045 13923
rect 9045 13889 9079 13923
rect 9079 13889 9088 13923
rect 9036 13880 9088 13889
rect 9312 13948 9364 14000
rect 10324 13948 10376 14000
rect 13268 13948 13320 14000
rect 9956 13812 10008 13864
rect 10784 13880 10836 13932
rect 10324 13855 10376 13864
rect 3056 13744 3108 13796
rect 7288 13744 7340 13796
rect 10324 13821 10333 13855
rect 10333 13821 10367 13855
rect 10367 13821 10376 13855
rect 10324 13812 10376 13821
rect 10876 13812 10928 13864
rect 8392 13676 8444 13728
rect 9588 13676 9640 13728
rect 14188 13923 14240 13932
rect 14188 13889 14197 13923
rect 14197 13889 14231 13923
rect 14231 13889 14240 13923
rect 14188 13880 14240 13889
rect 14648 13880 14700 13932
rect 14832 13923 14884 13932
rect 14832 13889 14841 13923
rect 14841 13889 14875 13923
rect 14875 13889 14884 13923
rect 14832 13880 14884 13889
rect 16856 13948 16908 14000
rect 17776 13948 17828 14000
rect 17408 13923 17460 13932
rect 15752 13812 15804 13864
rect 17408 13889 17417 13923
rect 17417 13889 17451 13923
rect 17451 13889 17460 13923
rect 17408 13880 17460 13889
rect 18052 13812 18104 13864
rect 12440 13744 12492 13796
rect 12992 13719 13044 13728
rect 12992 13685 13001 13719
rect 13001 13685 13035 13719
rect 13035 13685 13044 13719
rect 12992 13676 13044 13685
rect 14372 13719 14424 13728
rect 14372 13685 14381 13719
rect 14381 13685 14415 13719
rect 14415 13685 14424 13719
rect 14372 13676 14424 13685
rect 16396 13676 16448 13728
rect 17040 13719 17092 13728
rect 17040 13685 17049 13719
rect 17049 13685 17083 13719
rect 17083 13685 17092 13719
rect 17040 13676 17092 13685
rect 3169 13574 3221 13626
rect 3233 13574 3285 13626
rect 3297 13574 3349 13626
rect 3361 13574 3413 13626
rect 3425 13574 3477 13626
rect 7608 13574 7660 13626
rect 7672 13574 7724 13626
rect 7736 13574 7788 13626
rect 7800 13574 7852 13626
rect 7864 13574 7916 13626
rect 12047 13574 12099 13626
rect 12111 13574 12163 13626
rect 12175 13574 12227 13626
rect 12239 13574 12291 13626
rect 12303 13574 12355 13626
rect 16486 13574 16538 13626
rect 16550 13574 16602 13626
rect 16614 13574 16666 13626
rect 16678 13574 16730 13626
rect 16742 13574 16794 13626
rect 2320 13472 2372 13524
rect 4344 13472 4396 13524
rect 7472 13472 7524 13524
rect 7196 13404 7248 13456
rect 8208 13404 8260 13456
rect 10232 13472 10284 13524
rect 18052 13515 18104 13524
rect 18052 13481 18061 13515
rect 18061 13481 18095 13515
rect 18095 13481 18104 13515
rect 18052 13472 18104 13481
rect 9588 13404 9640 13456
rect 2228 13268 2280 13320
rect 2688 13311 2740 13320
rect 2688 13277 2697 13311
rect 2697 13277 2731 13311
rect 2731 13277 2740 13311
rect 2688 13268 2740 13277
rect 4988 13268 5040 13320
rect 7288 13268 7340 13320
rect 7932 13268 7984 13320
rect 8392 13311 8444 13320
rect 8392 13277 8401 13311
rect 8401 13277 8435 13311
rect 8435 13277 8444 13311
rect 8392 13268 8444 13277
rect 2596 13243 2648 13252
rect 2596 13209 2605 13243
rect 2605 13209 2639 13243
rect 2639 13209 2648 13243
rect 2596 13200 2648 13209
rect 5908 13243 5960 13252
rect 5908 13209 5942 13243
rect 5942 13209 5960 13243
rect 5908 13200 5960 13209
rect 8944 13200 8996 13252
rect 9404 13311 9456 13320
rect 9404 13277 9413 13311
rect 9413 13277 9447 13311
rect 9447 13277 9456 13311
rect 10324 13404 10376 13456
rect 10784 13404 10836 13456
rect 12256 13379 12308 13388
rect 12256 13345 12265 13379
rect 12265 13345 12299 13379
rect 12299 13345 12308 13379
rect 12256 13336 12308 13345
rect 17040 13336 17092 13388
rect 9404 13268 9456 13277
rect 10508 13268 10560 13320
rect 10600 13268 10652 13320
rect 12164 13311 12216 13320
rect 12164 13277 12173 13311
rect 12173 13277 12207 13311
rect 12207 13277 12216 13311
rect 12164 13268 12216 13277
rect 13820 13268 13872 13320
rect 14372 13268 14424 13320
rect 16856 13268 16908 13320
rect 17408 13268 17460 13320
rect 17960 13268 18012 13320
rect 9956 13200 10008 13252
rect 16580 13243 16632 13252
rect 16580 13209 16589 13243
rect 16589 13209 16623 13243
rect 16623 13209 16632 13243
rect 16580 13200 16632 13209
rect 7012 13175 7064 13184
rect 7012 13141 7021 13175
rect 7021 13141 7055 13175
rect 7055 13141 7064 13175
rect 7012 13132 7064 13141
rect 10968 13132 11020 13184
rect 11428 13132 11480 13184
rect 12716 13132 12768 13184
rect 15660 13175 15712 13184
rect 15660 13141 15669 13175
rect 15669 13141 15703 13175
rect 15703 13141 15712 13175
rect 17132 13200 17184 13252
rect 17500 13175 17552 13184
rect 15660 13132 15712 13141
rect 17500 13141 17509 13175
rect 17509 13141 17543 13175
rect 17543 13141 17552 13175
rect 17500 13132 17552 13141
rect 5388 13030 5440 13082
rect 5452 13030 5504 13082
rect 5516 13030 5568 13082
rect 5580 13030 5632 13082
rect 5644 13030 5696 13082
rect 9827 13030 9879 13082
rect 9891 13030 9943 13082
rect 9955 13030 10007 13082
rect 10019 13030 10071 13082
rect 10083 13030 10135 13082
rect 14266 13030 14318 13082
rect 14330 13030 14382 13082
rect 14394 13030 14446 13082
rect 14458 13030 14510 13082
rect 14522 13030 14574 13082
rect 18705 13030 18757 13082
rect 18769 13030 18821 13082
rect 18833 13030 18885 13082
rect 18897 13030 18949 13082
rect 18961 13030 19013 13082
rect 4160 12928 4212 12980
rect 5908 12928 5960 12980
rect 8300 12971 8352 12980
rect 8300 12937 8309 12971
rect 8309 12937 8343 12971
rect 8343 12937 8352 12971
rect 8300 12928 8352 12937
rect 10600 12971 10652 12980
rect 10600 12937 10609 12971
rect 10609 12937 10643 12971
rect 10643 12937 10652 12971
rect 10600 12928 10652 12937
rect 14188 12971 14240 12980
rect 14188 12937 14197 12971
rect 14197 12937 14231 12971
rect 14231 12937 14240 12971
rect 14188 12928 14240 12937
rect 14648 12928 14700 12980
rect 2412 12860 2464 12912
rect 2596 12860 2648 12912
rect 9496 12860 9548 12912
rect 2504 12835 2556 12844
rect 2504 12801 2513 12835
rect 2513 12801 2547 12835
rect 2547 12801 2556 12835
rect 2504 12792 2556 12801
rect 4252 12792 4304 12844
rect 6000 12835 6052 12844
rect 6000 12801 6009 12835
rect 6009 12801 6043 12835
rect 6043 12801 6052 12835
rect 6000 12792 6052 12801
rect 7196 12835 7248 12844
rect 7196 12801 7205 12835
rect 7205 12801 7239 12835
rect 7239 12801 7248 12835
rect 7196 12792 7248 12801
rect 9680 12792 9732 12844
rect 10324 12835 10376 12844
rect 10324 12801 10333 12835
rect 10333 12801 10367 12835
rect 10367 12801 10376 12835
rect 10324 12792 10376 12801
rect 4988 12767 5040 12776
rect 4988 12733 4997 12767
rect 4997 12733 5031 12767
rect 5031 12733 5040 12767
rect 7012 12767 7064 12776
rect 4988 12724 5040 12733
rect 7012 12733 7021 12767
rect 7021 12733 7055 12767
rect 7055 12733 7064 12767
rect 11612 12792 11664 12844
rect 12440 12860 12492 12912
rect 13084 12860 13136 12912
rect 14096 12860 14148 12912
rect 15292 12860 15344 12912
rect 12164 12792 12216 12844
rect 15660 12792 15712 12844
rect 15936 12835 15988 12844
rect 15936 12801 15945 12835
rect 15945 12801 15979 12835
rect 15979 12801 15988 12835
rect 15936 12792 15988 12801
rect 16120 12835 16172 12844
rect 16120 12801 16129 12835
rect 16129 12801 16163 12835
rect 16163 12801 16172 12835
rect 16120 12792 16172 12801
rect 16948 12792 17000 12844
rect 7012 12724 7064 12733
rect 2596 12656 2648 12708
rect 4620 12588 4672 12640
rect 8208 12656 8260 12708
rect 12256 12724 12308 12776
rect 12808 12656 12860 12708
rect 15384 12767 15436 12776
rect 15384 12733 15393 12767
rect 15393 12733 15427 12767
rect 15427 12733 15436 12767
rect 15384 12724 15436 12733
rect 16028 12724 16080 12776
rect 16580 12724 16632 12776
rect 17224 12724 17276 12776
rect 7380 12631 7432 12640
rect 7380 12597 7389 12631
rect 7389 12597 7423 12631
rect 7423 12597 7432 12631
rect 7380 12588 7432 12597
rect 10508 12588 10560 12640
rect 10784 12588 10836 12640
rect 11060 12631 11112 12640
rect 11060 12597 11069 12631
rect 11069 12597 11103 12631
rect 11103 12597 11112 12631
rect 11060 12588 11112 12597
rect 11152 12588 11204 12640
rect 15752 12588 15804 12640
rect 3169 12486 3221 12538
rect 3233 12486 3285 12538
rect 3297 12486 3349 12538
rect 3361 12486 3413 12538
rect 3425 12486 3477 12538
rect 7608 12486 7660 12538
rect 7672 12486 7724 12538
rect 7736 12486 7788 12538
rect 7800 12486 7852 12538
rect 7864 12486 7916 12538
rect 12047 12486 12099 12538
rect 12111 12486 12163 12538
rect 12175 12486 12227 12538
rect 12239 12486 12291 12538
rect 12303 12486 12355 12538
rect 16486 12486 16538 12538
rect 16550 12486 16602 12538
rect 16614 12486 16666 12538
rect 16678 12486 16730 12538
rect 16742 12486 16794 12538
rect 2504 12384 2556 12436
rect 4252 12427 4304 12436
rect 4252 12393 4261 12427
rect 4261 12393 4295 12427
rect 4295 12393 4304 12427
rect 4252 12384 4304 12393
rect 6000 12384 6052 12436
rect 9036 12384 9088 12436
rect 8208 12316 8260 12368
rect 9496 12384 9548 12436
rect 10048 12384 10100 12436
rect 10692 12384 10744 12436
rect 11060 12384 11112 12436
rect 11520 12427 11572 12436
rect 11520 12393 11529 12427
rect 11529 12393 11563 12427
rect 11563 12393 11572 12427
rect 11520 12384 11572 12393
rect 6828 12248 6880 12300
rect 9312 12291 9364 12300
rect 9312 12257 9321 12291
rect 9321 12257 9355 12291
rect 9355 12257 9364 12291
rect 9312 12248 9364 12257
rect 2228 12223 2280 12232
rect 2228 12189 2237 12223
rect 2237 12189 2271 12223
rect 2271 12189 2280 12223
rect 2228 12180 2280 12189
rect 2412 12223 2464 12232
rect 2412 12189 2421 12223
rect 2421 12189 2455 12223
rect 2455 12189 2464 12223
rect 2412 12180 2464 12189
rect 2596 12180 2648 12232
rect 2872 12180 2924 12232
rect 3976 12180 4028 12232
rect 6368 12223 6420 12232
rect 6368 12189 6377 12223
rect 6377 12189 6411 12223
rect 6411 12189 6420 12223
rect 6368 12180 6420 12189
rect 7196 12180 7248 12232
rect 7380 12180 7432 12232
rect 7932 12223 7984 12232
rect 7932 12189 7941 12223
rect 7941 12189 7975 12223
rect 7975 12189 7984 12223
rect 7932 12180 7984 12189
rect 8116 12180 8168 12232
rect 8392 12223 8444 12232
rect 8392 12189 8401 12223
rect 8401 12189 8435 12223
rect 8435 12189 8444 12223
rect 9220 12223 9272 12232
rect 8392 12180 8444 12189
rect 9220 12189 9229 12223
rect 9229 12189 9263 12223
rect 9263 12189 9272 12223
rect 9220 12180 9272 12189
rect 10324 12180 10376 12232
rect 10876 12248 10928 12300
rect 10968 12248 11020 12300
rect 11244 12248 11296 12300
rect 11152 12180 11204 12232
rect 11704 12180 11756 12232
rect 7012 12155 7064 12164
rect 7012 12121 7021 12155
rect 7021 12121 7055 12155
rect 7055 12121 7064 12155
rect 7012 12112 7064 12121
rect 3056 12044 3108 12096
rect 7104 12044 7156 12096
rect 7288 12044 7340 12096
rect 8024 12087 8076 12096
rect 8024 12053 8033 12087
rect 8033 12053 8067 12087
rect 8067 12053 8076 12087
rect 8024 12044 8076 12053
rect 10508 12112 10560 12164
rect 12808 12180 12860 12232
rect 16120 12384 16172 12436
rect 17776 12427 17828 12436
rect 17776 12393 17785 12427
rect 17785 12393 17819 12427
rect 17819 12393 17828 12427
rect 17776 12384 17828 12393
rect 14004 12180 14056 12232
rect 16672 12223 16724 12232
rect 16672 12189 16681 12223
rect 16681 12189 16715 12223
rect 16715 12189 16724 12223
rect 16672 12180 16724 12189
rect 8392 12044 8444 12096
rect 10048 12044 10100 12096
rect 10232 12087 10284 12096
rect 10232 12053 10241 12087
rect 10241 12053 10275 12087
rect 10275 12053 10284 12087
rect 10232 12044 10284 12053
rect 10416 12044 10468 12096
rect 14648 12112 14700 12164
rect 12532 12087 12584 12096
rect 12532 12053 12541 12087
rect 12541 12053 12575 12087
rect 12575 12053 12584 12087
rect 12532 12044 12584 12053
rect 12624 12044 12676 12096
rect 15936 12112 15988 12164
rect 16672 12044 16724 12096
rect 16856 12155 16908 12164
rect 16856 12121 16865 12155
rect 16865 12121 16899 12155
rect 16899 12121 16908 12155
rect 17132 12180 17184 12232
rect 16856 12112 16908 12121
rect 17224 12112 17276 12164
rect 17040 12044 17092 12096
rect 17960 12087 18012 12096
rect 17960 12053 17969 12087
rect 17969 12053 18003 12087
rect 18003 12053 18012 12087
rect 17960 12044 18012 12053
rect 5388 11942 5440 11994
rect 5452 11942 5504 11994
rect 5516 11942 5568 11994
rect 5580 11942 5632 11994
rect 5644 11942 5696 11994
rect 9827 11942 9879 11994
rect 9891 11942 9943 11994
rect 9955 11942 10007 11994
rect 10019 11942 10071 11994
rect 10083 11942 10135 11994
rect 14266 11942 14318 11994
rect 14330 11942 14382 11994
rect 14394 11942 14446 11994
rect 14458 11942 14510 11994
rect 14522 11942 14574 11994
rect 18705 11942 18757 11994
rect 18769 11942 18821 11994
rect 18833 11942 18885 11994
rect 18897 11942 18949 11994
rect 18961 11942 19013 11994
rect 7932 11840 7984 11892
rect 8760 11840 8812 11892
rect 9220 11840 9272 11892
rect 10416 11883 10468 11892
rect 10416 11849 10425 11883
rect 10425 11849 10459 11883
rect 10459 11849 10468 11883
rect 10416 11840 10468 11849
rect 12532 11840 12584 11892
rect 14648 11840 14700 11892
rect 15292 11840 15344 11892
rect 15936 11840 15988 11892
rect 4620 11772 4672 11824
rect 3056 11747 3108 11756
rect 3056 11713 3090 11747
rect 3090 11713 3108 11747
rect 3056 11704 3108 11713
rect 3792 11704 3844 11756
rect 6092 11704 6144 11756
rect 7104 11772 7156 11824
rect 7288 11772 7340 11824
rect 11060 11815 11112 11824
rect 7012 11704 7064 11756
rect 8208 11747 8260 11756
rect 8208 11713 8217 11747
rect 8217 11713 8251 11747
rect 8251 11713 8260 11747
rect 8208 11704 8260 11713
rect 8576 11704 8628 11756
rect 9220 11747 9272 11756
rect 9220 11713 9229 11747
rect 9229 11713 9263 11747
rect 9263 11713 9272 11747
rect 9220 11704 9272 11713
rect 9312 11704 9364 11756
rect 11060 11781 11069 11815
rect 11069 11781 11103 11815
rect 11103 11781 11112 11815
rect 11060 11772 11112 11781
rect 10508 11747 10560 11756
rect 10508 11713 10517 11747
rect 10517 11713 10551 11747
rect 10551 11713 10560 11747
rect 10508 11704 10560 11713
rect 4620 11679 4672 11688
rect 4620 11645 4629 11679
rect 4629 11645 4663 11679
rect 4663 11645 4672 11679
rect 4620 11636 4672 11645
rect 8116 11636 8168 11688
rect 9404 11568 9456 11620
rect 11612 11704 11664 11756
rect 12624 11747 12676 11756
rect 12624 11713 12633 11747
rect 12633 11713 12667 11747
rect 12667 11713 12676 11747
rect 12808 11747 12860 11756
rect 12624 11704 12676 11713
rect 12808 11713 12817 11747
rect 12817 11713 12851 11747
rect 12851 11713 12860 11747
rect 12808 11704 12860 11713
rect 4160 11543 4212 11552
rect 4160 11509 4169 11543
rect 4169 11509 4203 11543
rect 4203 11509 4212 11543
rect 4160 11500 4212 11509
rect 6184 11500 6236 11552
rect 7012 11500 7064 11552
rect 8576 11500 8628 11552
rect 8944 11500 8996 11552
rect 11704 11543 11756 11552
rect 11704 11509 11713 11543
rect 11713 11509 11747 11543
rect 11747 11509 11756 11543
rect 11704 11500 11756 11509
rect 11888 11568 11940 11620
rect 12440 11568 12492 11620
rect 13360 11543 13412 11552
rect 13360 11509 13369 11543
rect 13369 11509 13403 11543
rect 13403 11509 13412 11543
rect 13360 11500 13412 11509
rect 14188 11500 14240 11552
rect 14832 11500 14884 11552
rect 15752 11747 15804 11756
rect 15752 11713 15761 11747
rect 15761 11713 15795 11747
rect 15795 11713 15804 11747
rect 15752 11704 15804 11713
rect 16396 11704 16448 11756
rect 16672 11704 16724 11756
rect 17592 11704 17644 11756
rect 17960 11704 18012 11756
rect 16028 11636 16080 11688
rect 15752 11568 15804 11620
rect 16212 11500 16264 11552
rect 17500 11500 17552 11552
rect 17684 11543 17736 11552
rect 17684 11509 17693 11543
rect 17693 11509 17727 11543
rect 17727 11509 17736 11543
rect 17684 11500 17736 11509
rect 3169 11398 3221 11450
rect 3233 11398 3285 11450
rect 3297 11398 3349 11450
rect 3361 11398 3413 11450
rect 3425 11398 3477 11450
rect 7608 11398 7660 11450
rect 7672 11398 7724 11450
rect 7736 11398 7788 11450
rect 7800 11398 7852 11450
rect 7864 11398 7916 11450
rect 12047 11398 12099 11450
rect 12111 11398 12163 11450
rect 12175 11398 12227 11450
rect 12239 11398 12291 11450
rect 12303 11398 12355 11450
rect 16486 11398 16538 11450
rect 16550 11398 16602 11450
rect 16614 11398 16666 11450
rect 16678 11398 16730 11450
rect 16742 11398 16794 11450
rect 2872 11339 2924 11348
rect 2872 11305 2881 11339
rect 2881 11305 2915 11339
rect 2915 11305 2924 11339
rect 2872 11296 2924 11305
rect 3976 11339 4028 11348
rect 3976 11305 3985 11339
rect 3985 11305 4019 11339
rect 4019 11305 4028 11339
rect 3976 11296 4028 11305
rect 6092 11339 6144 11348
rect 6092 11305 6101 11339
rect 6101 11305 6135 11339
rect 6135 11305 6144 11339
rect 6092 11296 6144 11305
rect 7012 11339 7064 11348
rect 7012 11305 7021 11339
rect 7021 11305 7055 11339
rect 7055 11305 7064 11339
rect 7012 11296 7064 11305
rect 7196 11296 7248 11348
rect 10508 11296 10560 11348
rect 13176 11296 13228 11348
rect 16948 11296 17000 11348
rect 17684 11339 17736 11348
rect 17684 11305 17693 11339
rect 17693 11305 17727 11339
rect 17727 11305 17736 11339
rect 17684 11296 17736 11305
rect 2412 11160 2464 11212
rect 4344 11203 4396 11212
rect 3240 11092 3292 11144
rect 3792 11092 3844 11144
rect 4344 11169 4353 11203
rect 4353 11169 4387 11203
rect 4387 11169 4396 11203
rect 4344 11160 4396 11169
rect 8208 11228 8260 11280
rect 8944 11160 8996 11212
rect 4160 11135 4212 11144
rect 4160 11101 4169 11135
rect 4169 11101 4203 11135
rect 4203 11101 4212 11135
rect 4160 11092 4212 11101
rect 6184 11092 6236 11144
rect 6368 11135 6420 11144
rect 6368 11101 6377 11135
rect 6377 11101 6411 11135
rect 6411 11101 6420 11135
rect 6368 11092 6420 11101
rect 7288 11092 7340 11144
rect 11704 11228 11756 11280
rect 11888 11160 11940 11212
rect 12900 11228 12952 11280
rect 6828 11024 6880 11076
rect 4160 10956 4212 11008
rect 5816 10956 5868 11008
rect 6092 10956 6144 11008
rect 8208 11024 8260 11076
rect 8300 11024 8352 11076
rect 9404 11135 9456 11144
rect 9404 11101 9413 11135
rect 9413 11101 9447 11135
rect 9447 11101 9456 11135
rect 9404 11092 9456 11101
rect 10784 11092 10836 11144
rect 12532 11135 12584 11144
rect 12532 11101 12541 11135
rect 12541 11101 12575 11135
rect 12575 11101 12584 11135
rect 12716 11135 12768 11144
rect 12532 11092 12584 11101
rect 12716 11101 12725 11135
rect 12725 11101 12759 11135
rect 12759 11101 12768 11135
rect 12716 11092 12768 11101
rect 12992 11160 13044 11212
rect 14832 11160 14884 11212
rect 14740 11135 14792 11144
rect 8484 10956 8536 11008
rect 9312 10956 9364 11008
rect 11888 11024 11940 11076
rect 12440 11024 12492 11076
rect 12624 11024 12676 11076
rect 14740 11101 14749 11135
rect 14749 11101 14783 11135
rect 14783 11101 14792 11135
rect 14740 11092 14792 11101
rect 15200 11092 15252 11144
rect 17316 11228 17368 11280
rect 16856 11160 16908 11212
rect 17408 11160 17460 11212
rect 17960 11160 18012 11212
rect 13268 11067 13320 11076
rect 13268 11033 13277 11067
rect 13277 11033 13311 11067
rect 13311 11033 13320 11067
rect 13268 11024 13320 11033
rect 16120 11024 16172 11076
rect 16396 11135 16448 11144
rect 16396 11101 16405 11135
rect 16405 11101 16439 11135
rect 16439 11101 16448 11135
rect 16672 11135 16724 11144
rect 16396 11092 16448 11101
rect 16672 11101 16681 11135
rect 16681 11101 16715 11135
rect 16715 11101 16724 11135
rect 16672 11092 16724 11101
rect 17040 11092 17092 11144
rect 17592 11135 17644 11144
rect 17592 11101 17601 11135
rect 17601 11101 17635 11135
rect 17635 11101 17644 11135
rect 17592 11092 17644 11101
rect 12808 10956 12860 11008
rect 13728 10999 13780 11008
rect 13728 10965 13737 10999
rect 13737 10965 13771 10999
rect 13771 10965 13780 10999
rect 13728 10956 13780 10965
rect 14648 10999 14700 11008
rect 14648 10965 14657 10999
rect 14657 10965 14691 10999
rect 14691 10965 14700 10999
rect 14648 10956 14700 10965
rect 15568 10999 15620 11008
rect 15568 10965 15577 10999
rect 15577 10965 15611 10999
rect 15611 10965 15620 10999
rect 15568 10956 15620 10965
rect 17132 11024 17184 11076
rect 17500 11024 17552 11076
rect 17224 10956 17276 11008
rect 5388 10854 5440 10906
rect 5452 10854 5504 10906
rect 5516 10854 5568 10906
rect 5580 10854 5632 10906
rect 5644 10854 5696 10906
rect 9827 10854 9879 10906
rect 9891 10854 9943 10906
rect 9955 10854 10007 10906
rect 10019 10854 10071 10906
rect 10083 10854 10135 10906
rect 14266 10854 14318 10906
rect 14330 10854 14382 10906
rect 14394 10854 14446 10906
rect 14458 10854 14510 10906
rect 14522 10854 14574 10906
rect 18705 10854 18757 10906
rect 18769 10854 18821 10906
rect 18833 10854 18885 10906
rect 18897 10854 18949 10906
rect 18961 10854 19013 10906
rect 2780 10616 2832 10668
rect 3240 10659 3292 10668
rect 3240 10625 3249 10659
rect 3249 10625 3283 10659
rect 3283 10625 3292 10659
rect 3240 10616 3292 10625
rect 9312 10752 9364 10804
rect 11520 10752 11572 10804
rect 11796 10795 11848 10804
rect 11796 10761 11805 10795
rect 11805 10761 11839 10795
rect 11839 10761 11848 10795
rect 11796 10752 11848 10761
rect 12624 10752 12676 10804
rect 12900 10752 12952 10804
rect 15384 10795 15436 10804
rect 4252 10616 4304 10668
rect 8024 10684 8076 10736
rect 8484 10684 8536 10736
rect 4436 10548 4488 10600
rect 7380 10616 7432 10668
rect 8208 10616 8260 10668
rect 8576 10659 8628 10668
rect 6092 10548 6144 10600
rect 6552 10591 6604 10600
rect 6552 10557 6561 10591
rect 6561 10557 6595 10591
rect 6595 10557 6604 10591
rect 6552 10548 6604 10557
rect 8576 10625 8585 10659
rect 8585 10625 8619 10659
rect 8619 10625 8628 10659
rect 8576 10616 8628 10625
rect 9220 10684 9272 10736
rect 14648 10684 14700 10736
rect 15384 10761 15393 10795
rect 15393 10761 15427 10795
rect 15427 10761 15436 10795
rect 15384 10752 15436 10761
rect 17132 10752 17184 10804
rect 17408 10795 17460 10804
rect 17408 10761 17417 10795
rect 17417 10761 17451 10795
rect 17451 10761 17460 10795
rect 17408 10752 17460 10761
rect 16396 10684 16448 10736
rect 17500 10684 17552 10736
rect 9312 10659 9364 10668
rect 9312 10625 9321 10659
rect 9321 10625 9355 10659
rect 9355 10625 9364 10659
rect 9312 10616 9364 10625
rect 9496 10616 9548 10668
rect 10324 10616 10376 10668
rect 11704 10659 11756 10668
rect 11704 10625 11713 10659
rect 11713 10625 11747 10659
rect 11747 10625 11756 10659
rect 11704 10616 11756 10625
rect 12532 10616 12584 10668
rect 12808 10659 12860 10668
rect 12808 10625 12817 10659
rect 12817 10625 12851 10659
rect 12851 10625 12860 10659
rect 12808 10616 12860 10625
rect 12992 10659 13044 10668
rect 12992 10625 13001 10659
rect 13001 10625 13035 10659
rect 13035 10625 13044 10659
rect 12992 10616 13044 10625
rect 14004 10659 14056 10668
rect 14004 10625 14013 10659
rect 14013 10625 14047 10659
rect 14047 10625 14056 10659
rect 14004 10616 14056 10625
rect 15844 10659 15896 10668
rect 8484 10480 8536 10532
rect 12900 10591 12952 10600
rect 12900 10557 12909 10591
rect 12909 10557 12943 10591
rect 12943 10557 12952 10591
rect 12900 10548 12952 10557
rect 15844 10625 15853 10659
rect 15853 10625 15887 10659
rect 15887 10625 15896 10659
rect 15844 10616 15896 10625
rect 15936 10616 15988 10668
rect 16580 10616 16632 10668
rect 17592 10616 17644 10668
rect 17040 10591 17092 10600
rect 2780 10455 2832 10464
rect 2780 10421 2789 10455
rect 2789 10421 2823 10455
rect 2823 10421 2832 10455
rect 4804 10455 4856 10464
rect 2780 10412 2832 10421
rect 4804 10421 4813 10455
rect 4813 10421 4847 10455
rect 4847 10421 4856 10455
rect 4804 10412 4856 10421
rect 7472 10412 7524 10464
rect 7932 10412 7984 10464
rect 9128 10455 9180 10464
rect 9128 10421 9137 10455
rect 9137 10421 9171 10455
rect 9171 10421 9180 10455
rect 9128 10412 9180 10421
rect 12808 10480 12860 10532
rect 17040 10557 17049 10591
rect 17049 10557 17083 10591
rect 17083 10557 17092 10591
rect 17040 10548 17092 10557
rect 17224 10548 17276 10600
rect 18052 10548 18104 10600
rect 13268 10412 13320 10464
rect 16028 10455 16080 10464
rect 16028 10421 16037 10455
rect 16037 10421 16071 10455
rect 16071 10421 16080 10455
rect 16028 10412 16080 10421
rect 16856 10455 16908 10464
rect 16856 10421 16865 10455
rect 16865 10421 16899 10455
rect 16899 10421 16908 10455
rect 16856 10412 16908 10421
rect 17684 10412 17736 10464
rect 18144 10412 18196 10464
rect 3169 10310 3221 10362
rect 3233 10310 3285 10362
rect 3297 10310 3349 10362
rect 3361 10310 3413 10362
rect 3425 10310 3477 10362
rect 7608 10310 7660 10362
rect 7672 10310 7724 10362
rect 7736 10310 7788 10362
rect 7800 10310 7852 10362
rect 7864 10310 7916 10362
rect 12047 10310 12099 10362
rect 12111 10310 12163 10362
rect 12175 10310 12227 10362
rect 12239 10310 12291 10362
rect 12303 10310 12355 10362
rect 16486 10310 16538 10362
rect 16550 10310 16602 10362
rect 16614 10310 16666 10362
rect 16678 10310 16730 10362
rect 16742 10310 16794 10362
rect 3700 10208 3752 10260
rect 6552 10208 6604 10260
rect 7380 10208 7432 10260
rect 8668 10208 8720 10260
rect 9680 10208 9732 10260
rect 11704 10208 11756 10260
rect 7288 10140 7340 10192
rect 11520 10140 11572 10192
rect 13176 10183 13228 10192
rect 10508 10072 10560 10124
rect 13176 10149 13185 10183
rect 13185 10149 13219 10183
rect 13219 10149 13228 10183
rect 13176 10140 13228 10149
rect 14740 10208 14792 10260
rect 15568 10208 15620 10260
rect 17500 10208 17552 10260
rect 17776 10251 17828 10260
rect 17776 10217 17785 10251
rect 17785 10217 17819 10251
rect 17819 10217 17828 10251
rect 17776 10208 17828 10217
rect 17868 10208 17920 10260
rect 15476 10140 15528 10192
rect 2504 9979 2556 9988
rect 2504 9945 2513 9979
rect 2513 9945 2547 9979
rect 2547 9945 2556 9979
rect 2504 9936 2556 9945
rect 7012 10047 7064 10056
rect 7012 10013 7021 10047
rect 7021 10013 7055 10047
rect 7055 10013 7064 10047
rect 7012 10004 7064 10013
rect 7472 10004 7524 10056
rect 8116 10004 8168 10056
rect 8668 10004 8720 10056
rect 11336 10047 11388 10056
rect 11336 10013 11345 10047
rect 11345 10013 11379 10047
rect 11379 10013 11388 10047
rect 11336 10004 11388 10013
rect 15936 10072 15988 10124
rect 12808 10047 12860 10056
rect 12808 10013 12817 10047
rect 12817 10013 12851 10047
rect 12851 10013 12860 10047
rect 12808 10004 12860 10013
rect 15384 10004 15436 10056
rect 15752 10047 15804 10056
rect 15752 10013 15761 10047
rect 15761 10013 15795 10047
rect 15795 10013 15804 10047
rect 15752 10004 15804 10013
rect 17684 10072 17736 10124
rect 3700 9936 3752 9988
rect 8576 9936 8628 9988
rect 9496 9936 9548 9988
rect 17132 10004 17184 10056
rect 17500 10004 17552 10056
rect 17592 10004 17644 10056
rect 18052 10047 18104 10056
rect 18052 10013 18061 10047
rect 18061 10013 18095 10047
rect 18095 10013 18104 10047
rect 18052 10004 18104 10013
rect 17316 9936 17368 9988
rect 3608 9868 3660 9920
rect 11428 9911 11480 9920
rect 11428 9877 11437 9911
rect 11437 9877 11471 9911
rect 11471 9877 11480 9911
rect 11428 9868 11480 9877
rect 11612 9868 11664 9920
rect 13820 9868 13872 9920
rect 14832 9868 14884 9920
rect 15384 9868 15436 9920
rect 17408 9868 17460 9920
rect 17592 9911 17644 9920
rect 17592 9877 17601 9911
rect 17601 9877 17635 9911
rect 17635 9877 17644 9911
rect 17592 9868 17644 9877
rect 5388 9766 5440 9818
rect 5452 9766 5504 9818
rect 5516 9766 5568 9818
rect 5580 9766 5632 9818
rect 5644 9766 5696 9818
rect 9827 9766 9879 9818
rect 9891 9766 9943 9818
rect 9955 9766 10007 9818
rect 10019 9766 10071 9818
rect 10083 9766 10135 9818
rect 14266 9766 14318 9818
rect 14330 9766 14382 9818
rect 14394 9766 14446 9818
rect 14458 9766 14510 9818
rect 14522 9766 14574 9818
rect 18705 9766 18757 9818
rect 18769 9766 18821 9818
rect 18833 9766 18885 9818
rect 18897 9766 18949 9818
rect 18961 9766 19013 9818
rect 2780 9596 2832 9648
rect 4620 9596 4672 9648
rect 6552 9596 6604 9648
rect 10324 9664 10376 9716
rect 11428 9664 11480 9716
rect 4804 9571 4856 9580
rect 4804 9537 4838 9571
rect 4838 9537 4856 9571
rect 4804 9528 4856 9537
rect 6736 9571 6788 9580
rect 6736 9537 6745 9571
rect 6745 9537 6779 9571
rect 6779 9537 6788 9571
rect 6736 9528 6788 9537
rect 9220 9596 9272 9648
rect 9588 9639 9640 9648
rect 9588 9605 9597 9639
rect 9597 9605 9631 9639
rect 9631 9605 9640 9639
rect 9588 9596 9640 9605
rect 7472 9528 7524 9580
rect 11244 9596 11296 9648
rect 11336 9596 11388 9648
rect 11980 9639 12032 9648
rect 11980 9605 11989 9639
rect 11989 9605 12023 9639
rect 12023 9605 12032 9639
rect 11980 9596 12032 9605
rect 12992 9639 13044 9648
rect 12992 9605 13001 9639
rect 13001 9605 13035 9639
rect 13035 9605 13044 9639
rect 12992 9596 13044 9605
rect 13176 9596 13228 9648
rect 13912 9639 13964 9648
rect 13912 9605 13921 9639
rect 13921 9605 13955 9639
rect 13955 9605 13964 9639
rect 13912 9596 13964 9605
rect 10784 9528 10836 9580
rect 10600 9503 10652 9512
rect 10600 9469 10609 9503
rect 10609 9469 10643 9503
rect 10643 9469 10652 9503
rect 10600 9460 10652 9469
rect 11428 9460 11480 9512
rect 12348 9528 12400 9580
rect 11060 9392 11112 9444
rect 12348 9392 12400 9444
rect 1860 9324 1912 9376
rect 2504 9324 2556 9376
rect 4160 9324 4212 9376
rect 8116 9324 8168 9376
rect 10968 9367 11020 9376
rect 10968 9333 10977 9367
rect 10977 9333 11011 9367
rect 11011 9333 11020 9367
rect 10968 9324 11020 9333
rect 11796 9324 11848 9376
rect 13176 9392 13228 9444
rect 13452 9392 13504 9444
rect 14740 9528 14792 9580
rect 14832 9571 14884 9580
rect 14832 9537 14841 9571
rect 14841 9537 14875 9571
rect 14875 9537 14884 9571
rect 16948 9596 17000 9648
rect 17776 9639 17828 9648
rect 17776 9605 17785 9639
rect 17785 9605 17819 9639
rect 17819 9605 17828 9639
rect 17776 9596 17828 9605
rect 14832 9528 14884 9537
rect 15936 9571 15988 9580
rect 15936 9537 15945 9571
rect 15945 9537 15979 9571
rect 15979 9537 15988 9571
rect 15936 9528 15988 9537
rect 16764 9528 16816 9580
rect 17500 9571 17552 9580
rect 13544 9367 13596 9376
rect 13544 9333 13553 9367
rect 13553 9333 13587 9367
rect 13587 9333 13596 9367
rect 13544 9324 13596 9333
rect 15200 9392 15252 9444
rect 17500 9537 17509 9571
rect 17509 9537 17543 9571
rect 17543 9537 17552 9571
rect 17500 9528 17552 9537
rect 18144 9460 18196 9512
rect 18052 9392 18104 9444
rect 14648 9367 14700 9376
rect 14648 9333 14657 9367
rect 14657 9333 14691 9367
rect 14691 9333 14700 9367
rect 14648 9324 14700 9333
rect 15292 9324 15344 9376
rect 16948 9367 17000 9376
rect 16948 9333 16957 9367
rect 16957 9333 16991 9367
rect 16991 9333 17000 9367
rect 16948 9324 17000 9333
rect 3169 9222 3221 9274
rect 3233 9222 3285 9274
rect 3297 9222 3349 9274
rect 3361 9222 3413 9274
rect 3425 9222 3477 9274
rect 7608 9222 7660 9274
rect 7672 9222 7724 9274
rect 7736 9222 7788 9274
rect 7800 9222 7852 9274
rect 7864 9222 7916 9274
rect 12047 9222 12099 9274
rect 12111 9222 12163 9274
rect 12175 9222 12227 9274
rect 12239 9222 12291 9274
rect 12303 9222 12355 9274
rect 16486 9222 16538 9274
rect 16550 9222 16602 9274
rect 16614 9222 16666 9274
rect 16678 9222 16730 9274
rect 16742 9222 16794 9274
rect 4988 9120 5040 9172
rect 8208 9120 8260 9172
rect 9588 9120 9640 9172
rect 10600 9120 10652 9172
rect 5908 9052 5960 9104
rect 6828 9052 6880 9104
rect 8024 9052 8076 9104
rect 10508 9052 10560 9104
rect 12900 9120 12952 9172
rect 12992 9120 13044 9172
rect 13912 9120 13964 9172
rect 14740 9163 14792 9172
rect 14740 9129 14749 9163
rect 14749 9129 14783 9163
rect 14783 9129 14792 9163
rect 14740 9120 14792 9129
rect 15292 9163 15344 9172
rect 15292 9129 15301 9163
rect 15301 9129 15335 9163
rect 15335 9129 15344 9163
rect 15292 9120 15344 9129
rect 16028 9120 16080 9172
rect 17040 9120 17092 9172
rect 17776 9120 17828 9172
rect 10232 8984 10284 9036
rect 11520 9052 11572 9104
rect 11428 8984 11480 9036
rect 5080 8916 5132 8968
rect 5724 8959 5776 8968
rect 4896 8823 4948 8832
rect 4896 8789 4921 8823
rect 4921 8789 4948 8823
rect 5724 8925 5733 8959
rect 5733 8925 5767 8959
rect 5767 8925 5776 8959
rect 5724 8916 5776 8925
rect 8300 8916 8352 8968
rect 9128 8916 9180 8968
rect 9312 8916 9364 8968
rect 10968 8916 11020 8968
rect 11704 8916 11756 8968
rect 16120 9095 16172 9104
rect 16120 9061 16129 9095
rect 16129 9061 16163 9095
rect 16163 9061 16172 9095
rect 16120 9052 16172 9061
rect 17316 9095 17368 9104
rect 17316 9061 17325 9095
rect 17325 9061 17359 9095
rect 17359 9061 17368 9095
rect 17316 9052 17368 9061
rect 12256 8984 12308 9036
rect 12440 8984 12492 9036
rect 13544 8984 13596 9036
rect 13636 8959 13688 8968
rect 6368 8891 6420 8900
rect 6368 8857 6377 8891
rect 6377 8857 6411 8891
rect 6411 8857 6420 8891
rect 6368 8848 6420 8857
rect 6552 8891 6604 8900
rect 6552 8857 6561 8891
rect 6561 8857 6595 8891
rect 6595 8857 6604 8891
rect 6552 8848 6604 8857
rect 9588 8848 9640 8900
rect 11428 8848 11480 8900
rect 11796 8848 11848 8900
rect 13636 8925 13645 8959
rect 13645 8925 13679 8959
rect 13679 8925 13688 8959
rect 13636 8916 13688 8925
rect 4896 8780 4948 8789
rect 5816 8780 5868 8832
rect 7104 8780 7156 8832
rect 11060 8823 11112 8832
rect 11060 8789 11069 8823
rect 11069 8789 11103 8823
rect 11103 8789 11112 8823
rect 11060 8780 11112 8789
rect 11888 8780 11940 8832
rect 12532 8780 12584 8832
rect 12900 8780 12952 8832
rect 15752 8984 15804 9036
rect 17500 8984 17552 9036
rect 15016 8916 15068 8968
rect 16948 8916 17000 8968
rect 17132 8916 17184 8968
rect 17684 8959 17736 8968
rect 17684 8925 17693 8959
rect 17693 8925 17727 8959
rect 17727 8925 17736 8959
rect 17684 8916 17736 8925
rect 18052 8916 18104 8968
rect 13912 8848 13964 8900
rect 17592 8848 17644 8900
rect 14004 8780 14056 8832
rect 15108 8780 15160 8832
rect 15384 8780 15436 8832
rect 17040 8780 17092 8832
rect 18236 8823 18288 8832
rect 18236 8789 18245 8823
rect 18245 8789 18279 8823
rect 18279 8789 18288 8823
rect 18236 8780 18288 8789
rect 5388 8678 5440 8730
rect 5452 8678 5504 8730
rect 5516 8678 5568 8730
rect 5580 8678 5632 8730
rect 5644 8678 5696 8730
rect 9827 8678 9879 8730
rect 9891 8678 9943 8730
rect 9955 8678 10007 8730
rect 10019 8678 10071 8730
rect 10083 8678 10135 8730
rect 14266 8678 14318 8730
rect 14330 8678 14382 8730
rect 14394 8678 14446 8730
rect 14458 8678 14510 8730
rect 14522 8678 14574 8730
rect 18705 8678 18757 8730
rect 18769 8678 18821 8730
rect 18833 8678 18885 8730
rect 18897 8678 18949 8730
rect 18961 8678 19013 8730
rect 4436 8619 4488 8628
rect 4436 8585 4445 8619
rect 4445 8585 4479 8619
rect 4479 8585 4488 8619
rect 4436 8576 4488 8585
rect 6552 8619 6604 8628
rect 6552 8585 6561 8619
rect 6561 8585 6595 8619
rect 6595 8585 6604 8619
rect 6552 8576 6604 8585
rect 6828 8576 6880 8628
rect 9680 8576 9732 8628
rect 10324 8576 10376 8628
rect 12256 8576 12308 8628
rect 2596 8440 2648 8492
rect 4620 8508 4672 8560
rect 6368 8508 6420 8560
rect 3608 8440 3660 8492
rect 5080 8483 5132 8492
rect 5080 8449 5089 8483
rect 5089 8449 5123 8483
rect 5123 8449 5132 8483
rect 5080 8440 5132 8449
rect 2044 8415 2096 8424
rect 2044 8381 2053 8415
rect 2053 8381 2087 8415
rect 2087 8381 2096 8415
rect 2044 8372 2096 8381
rect 4988 8415 5040 8424
rect 4988 8381 4997 8415
rect 4997 8381 5031 8415
rect 5031 8381 5040 8415
rect 4988 8372 5040 8381
rect 6000 8372 6052 8424
rect 8116 8440 8168 8492
rect 8484 8508 8536 8560
rect 9220 8508 9272 8560
rect 13360 8576 13412 8628
rect 17224 8576 17276 8628
rect 14648 8508 14700 8560
rect 17132 8508 17184 8560
rect 9036 8440 9088 8492
rect 10600 8483 10652 8492
rect 10600 8449 10609 8483
rect 10609 8449 10643 8483
rect 10643 8449 10652 8483
rect 10600 8440 10652 8449
rect 11060 8483 11112 8492
rect 11060 8449 11070 8483
rect 11070 8449 11112 8483
rect 11060 8440 11112 8449
rect 11704 8483 11756 8492
rect 11704 8449 11713 8483
rect 11713 8449 11747 8483
rect 11747 8449 11756 8483
rect 11704 8440 11756 8449
rect 11796 8440 11848 8492
rect 13728 8440 13780 8492
rect 16212 8440 16264 8492
rect 16856 8440 16908 8492
rect 17592 8483 17644 8492
rect 17592 8449 17601 8483
rect 17601 8449 17635 8483
rect 17635 8449 17644 8483
rect 17592 8440 17644 8449
rect 18236 8440 18288 8492
rect 10508 8415 10560 8424
rect 5816 8304 5868 8356
rect 6736 8304 6788 8356
rect 6920 8304 6972 8356
rect 10508 8381 10517 8415
rect 10517 8381 10551 8415
rect 10551 8381 10560 8415
rect 10508 8372 10560 8381
rect 11612 8372 11664 8424
rect 12348 8372 12400 8424
rect 13268 8415 13320 8424
rect 13268 8381 13277 8415
rect 13277 8381 13311 8415
rect 13311 8381 13320 8415
rect 14004 8415 14056 8424
rect 13268 8372 13320 8381
rect 14004 8381 14013 8415
rect 14013 8381 14047 8415
rect 14047 8381 14056 8415
rect 14004 8372 14056 8381
rect 17776 8415 17828 8424
rect 17776 8381 17785 8415
rect 17785 8381 17819 8415
rect 17819 8381 17828 8415
rect 17776 8372 17828 8381
rect 8576 8304 8628 8356
rect 9404 8304 9456 8356
rect 9680 8236 9732 8288
rect 10324 8236 10376 8288
rect 11152 8279 11204 8288
rect 11152 8245 11161 8279
rect 11161 8245 11195 8279
rect 11195 8245 11204 8279
rect 11152 8236 11204 8245
rect 11520 8236 11572 8288
rect 13820 8304 13872 8356
rect 15016 8304 15068 8356
rect 17316 8304 17368 8356
rect 16396 8236 16448 8288
rect 17408 8279 17460 8288
rect 17408 8245 17417 8279
rect 17417 8245 17451 8279
rect 17451 8245 17460 8279
rect 17408 8236 17460 8245
rect 3169 8134 3221 8186
rect 3233 8134 3285 8186
rect 3297 8134 3349 8186
rect 3361 8134 3413 8186
rect 3425 8134 3477 8186
rect 7608 8134 7660 8186
rect 7672 8134 7724 8186
rect 7736 8134 7788 8186
rect 7800 8134 7852 8186
rect 7864 8134 7916 8186
rect 12047 8134 12099 8186
rect 12111 8134 12163 8186
rect 12175 8134 12227 8186
rect 12239 8134 12291 8186
rect 12303 8134 12355 8186
rect 16486 8134 16538 8186
rect 16550 8134 16602 8186
rect 16614 8134 16666 8186
rect 16678 8134 16730 8186
rect 16742 8134 16794 8186
rect 2044 8032 2096 8084
rect 2596 8075 2648 8084
rect 2596 8041 2605 8075
rect 2605 8041 2639 8075
rect 2639 8041 2648 8075
rect 2596 8032 2648 8041
rect 6920 8032 6972 8084
rect 9312 8032 9364 8084
rect 1860 7939 1912 7948
rect 1860 7905 1869 7939
rect 1869 7905 1903 7939
rect 1903 7905 1912 7939
rect 1860 7896 1912 7905
rect 3056 7964 3108 8016
rect 4988 7964 5040 8016
rect 8300 7964 8352 8016
rect 3424 7828 3476 7880
rect 5080 7896 5132 7948
rect 9220 7939 9272 7948
rect 9220 7905 9229 7939
rect 9229 7905 9263 7939
rect 9263 7905 9272 7939
rect 9220 7896 9272 7905
rect 4160 7871 4212 7880
rect 4160 7837 4175 7871
rect 4175 7837 4209 7871
rect 4209 7837 4212 7871
rect 4160 7828 4212 7837
rect 3976 7760 4028 7812
rect 4896 7828 4948 7880
rect 5724 7828 5776 7880
rect 6000 7828 6052 7880
rect 6736 7871 6788 7880
rect 6736 7837 6745 7871
rect 6745 7837 6779 7871
rect 6779 7837 6788 7871
rect 6736 7828 6788 7837
rect 6828 7828 6880 7880
rect 8484 7871 8536 7880
rect 8484 7837 8493 7871
rect 8493 7837 8527 7871
rect 8527 7837 8536 7871
rect 8484 7828 8536 7837
rect 9404 7871 9456 7880
rect 9404 7837 9413 7871
rect 9413 7837 9447 7871
rect 9447 7837 9456 7871
rect 9404 7828 9456 7837
rect 11888 8032 11940 8084
rect 13268 8032 13320 8084
rect 17500 8075 17552 8084
rect 17500 8041 17509 8075
rect 17509 8041 17543 8075
rect 17543 8041 17552 8075
rect 17500 8032 17552 8041
rect 9680 7964 9732 8016
rect 11612 7964 11664 8016
rect 13912 7964 13964 8016
rect 11060 7896 11112 7948
rect 2964 7692 3016 7744
rect 6736 7692 6788 7744
rect 6920 7735 6972 7744
rect 6920 7701 6929 7735
rect 6929 7701 6963 7735
rect 6963 7701 6972 7735
rect 6920 7692 6972 7701
rect 8392 7760 8444 7812
rect 9496 7760 9548 7812
rect 10324 7803 10376 7812
rect 10324 7769 10333 7803
rect 10333 7769 10367 7803
rect 10367 7769 10376 7803
rect 10324 7760 10376 7769
rect 7564 7692 7616 7744
rect 8760 7692 8812 7744
rect 10232 7692 10284 7744
rect 12164 7871 12216 7880
rect 12164 7837 12173 7871
rect 12173 7837 12207 7871
rect 12207 7837 12216 7871
rect 12164 7828 12216 7837
rect 13636 7896 13688 7948
rect 15844 7896 15896 7948
rect 18052 7896 18104 7948
rect 13544 7871 13596 7880
rect 13544 7837 13553 7871
rect 13553 7837 13587 7871
rect 13587 7837 13596 7871
rect 13544 7828 13596 7837
rect 12808 7760 12860 7812
rect 16028 7760 16080 7812
rect 16856 7828 16908 7880
rect 17776 7871 17828 7880
rect 17776 7837 17785 7871
rect 17785 7837 17819 7871
rect 17819 7837 17828 7871
rect 17776 7828 17828 7837
rect 16948 7760 17000 7812
rect 13084 7692 13136 7744
rect 15936 7692 15988 7744
rect 17132 7692 17184 7744
rect 18236 7828 18288 7880
rect 18144 7692 18196 7744
rect 5388 7590 5440 7642
rect 5452 7590 5504 7642
rect 5516 7590 5568 7642
rect 5580 7590 5632 7642
rect 5644 7590 5696 7642
rect 9827 7590 9879 7642
rect 9891 7590 9943 7642
rect 9955 7590 10007 7642
rect 10019 7590 10071 7642
rect 10083 7590 10135 7642
rect 14266 7590 14318 7642
rect 14330 7590 14382 7642
rect 14394 7590 14446 7642
rect 14458 7590 14510 7642
rect 14522 7590 14574 7642
rect 18705 7590 18757 7642
rect 18769 7590 18821 7642
rect 18833 7590 18885 7642
rect 18897 7590 18949 7642
rect 18961 7590 19013 7642
rect 3424 7531 3476 7540
rect 3424 7497 3433 7531
rect 3433 7497 3467 7531
rect 3467 7497 3476 7531
rect 3424 7488 3476 7497
rect 4896 7531 4948 7540
rect 4896 7497 4905 7531
rect 4905 7497 4939 7531
rect 4939 7497 4948 7531
rect 4896 7488 4948 7497
rect 6828 7488 6880 7540
rect 7472 7488 7524 7540
rect 7564 7488 7616 7540
rect 3976 7420 4028 7472
rect 5080 7420 5132 7472
rect 6736 7463 6788 7472
rect 6736 7429 6745 7463
rect 6745 7429 6779 7463
rect 6779 7429 6788 7463
rect 6736 7420 6788 7429
rect 6920 7420 6972 7472
rect 4436 7352 4488 7404
rect 2780 7284 2832 7336
rect 3056 7284 3108 7336
rect 4160 7284 4212 7336
rect 5908 7352 5960 7404
rect 6000 7395 6052 7404
rect 6000 7361 6009 7395
rect 6009 7361 6043 7395
rect 6043 7361 6052 7395
rect 6000 7352 6052 7361
rect 7288 7352 7340 7404
rect 6552 7284 6604 7336
rect 8024 7284 8076 7336
rect 9496 7352 9548 7404
rect 9680 7395 9732 7404
rect 9680 7361 9689 7395
rect 9689 7361 9723 7395
rect 9723 7361 9732 7395
rect 9680 7352 9732 7361
rect 8484 7327 8536 7336
rect 8484 7293 8493 7327
rect 8493 7293 8527 7327
rect 8527 7293 8536 7327
rect 8484 7284 8536 7293
rect 12164 7488 12216 7540
rect 15844 7488 15896 7540
rect 16028 7531 16080 7540
rect 16028 7497 16037 7531
rect 16037 7497 16071 7531
rect 16071 7497 16080 7531
rect 16028 7488 16080 7497
rect 17224 7531 17276 7540
rect 17224 7497 17233 7531
rect 17233 7497 17267 7531
rect 17267 7497 17276 7531
rect 17224 7488 17276 7497
rect 11152 7395 11204 7404
rect 11152 7361 11161 7395
rect 11161 7361 11195 7395
rect 11195 7361 11204 7395
rect 11152 7352 11204 7361
rect 13544 7395 13596 7404
rect 13544 7361 13553 7395
rect 13553 7361 13587 7395
rect 13587 7361 13596 7395
rect 13544 7352 13596 7361
rect 13820 7352 13872 7404
rect 16120 7352 16172 7404
rect 11612 7284 11664 7336
rect 7932 7148 7984 7200
rect 8116 7148 8168 7200
rect 9036 7216 9088 7268
rect 9680 7216 9732 7268
rect 15200 7284 15252 7336
rect 15844 7327 15896 7336
rect 15844 7293 15878 7327
rect 15878 7293 15896 7327
rect 18052 7420 18104 7472
rect 17960 7352 18012 7404
rect 15844 7284 15896 7293
rect 17408 7284 17460 7336
rect 18236 7216 18288 7268
rect 8668 7148 8720 7200
rect 9864 7191 9916 7200
rect 9864 7157 9873 7191
rect 9873 7157 9907 7191
rect 9907 7157 9916 7191
rect 9864 7148 9916 7157
rect 13728 7191 13780 7200
rect 13728 7157 13737 7191
rect 13737 7157 13771 7191
rect 13771 7157 13780 7191
rect 13728 7148 13780 7157
rect 13820 7148 13872 7200
rect 17592 7148 17644 7200
rect 17868 7148 17920 7200
rect 3169 7046 3221 7098
rect 3233 7046 3285 7098
rect 3297 7046 3349 7098
rect 3361 7046 3413 7098
rect 3425 7046 3477 7098
rect 7608 7046 7660 7098
rect 7672 7046 7724 7098
rect 7736 7046 7788 7098
rect 7800 7046 7852 7098
rect 7864 7046 7916 7098
rect 12047 7046 12099 7098
rect 12111 7046 12163 7098
rect 12175 7046 12227 7098
rect 12239 7046 12291 7098
rect 12303 7046 12355 7098
rect 16486 7046 16538 7098
rect 16550 7046 16602 7098
rect 16614 7046 16666 7098
rect 16678 7046 16730 7098
rect 16742 7046 16794 7098
rect 8392 6987 8444 6996
rect 8392 6953 8401 6987
rect 8401 6953 8435 6987
rect 8435 6953 8444 6987
rect 8392 6944 8444 6953
rect 16120 6987 16172 6996
rect 16120 6953 16129 6987
rect 16129 6953 16163 6987
rect 16163 6953 16172 6987
rect 16120 6944 16172 6953
rect 17224 6987 17276 6996
rect 17224 6953 17233 6987
rect 17233 6953 17267 6987
rect 17267 6953 17276 6987
rect 17224 6944 17276 6953
rect 17960 6944 18012 6996
rect 2228 6783 2280 6792
rect 2228 6749 2237 6783
rect 2237 6749 2271 6783
rect 2271 6749 2280 6783
rect 2228 6740 2280 6749
rect 2964 6808 3016 6860
rect 3700 6808 3752 6860
rect 13820 6808 13872 6860
rect 14004 6808 14056 6860
rect 2780 6740 2832 6792
rect 3056 6783 3108 6792
rect 3056 6749 3065 6783
rect 3065 6749 3099 6783
rect 3099 6749 3108 6783
rect 3056 6740 3108 6749
rect 3240 6783 3292 6792
rect 3240 6749 3249 6783
rect 3249 6749 3283 6783
rect 3283 6749 3292 6783
rect 3240 6740 3292 6749
rect 4620 6740 4672 6792
rect 6552 6783 6604 6792
rect 6552 6749 6586 6783
rect 6586 6749 6604 6783
rect 6552 6740 6604 6749
rect 9128 6783 9180 6792
rect 6092 6672 6144 6724
rect 8300 6672 8352 6724
rect 8760 6672 8812 6724
rect 9128 6749 9137 6783
rect 9137 6749 9171 6783
rect 9171 6749 9180 6783
rect 9128 6740 9180 6749
rect 9680 6740 9732 6792
rect 9864 6740 9916 6792
rect 10324 6672 10376 6724
rect 10692 6672 10744 6724
rect 13544 6740 13596 6792
rect 16028 6808 16080 6860
rect 15936 6740 15988 6792
rect 16396 6783 16448 6792
rect 16396 6749 16405 6783
rect 16405 6749 16439 6783
rect 16439 6749 16448 6783
rect 16396 6740 16448 6749
rect 17132 6740 17184 6792
rect 13452 6715 13504 6724
rect 3700 6604 3752 6656
rect 7656 6647 7708 6656
rect 7656 6613 7665 6647
rect 7665 6613 7699 6647
rect 7699 6613 7708 6647
rect 7656 6604 7708 6613
rect 8668 6604 8720 6656
rect 9404 6604 9456 6656
rect 13452 6681 13461 6715
rect 13461 6681 13495 6715
rect 13495 6681 13504 6715
rect 13452 6672 13504 6681
rect 13084 6604 13136 6656
rect 14648 6672 14700 6724
rect 15660 6647 15712 6656
rect 15660 6613 15669 6647
rect 15669 6613 15703 6647
rect 15703 6613 15712 6647
rect 15660 6604 15712 6613
rect 17040 6647 17092 6656
rect 17040 6613 17049 6647
rect 17049 6613 17083 6647
rect 17083 6613 17092 6647
rect 17040 6604 17092 6613
rect 17224 6604 17276 6656
rect 5388 6502 5440 6554
rect 5452 6502 5504 6554
rect 5516 6502 5568 6554
rect 5580 6502 5632 6554
rect 5644 6502 5696 6554
rect 9827 6502 9879 6554
rect 9891 6502 9943 6554
rect 9955 6502 10007 6554
rect 10019 6502 10071 6554
rect 10083 6502 10135 6554
rect 14266 6502 14318 6554
rect 14330 6502 14382 6554
rect 14394 6502 14446 6554
rect 14458 6502 14510 6554
rect 14522 6502 14574 6554
rect 18705 6502 18757 6554
rect 18769 6502 18821 6554
rect 18833 6502 18885 6554
rect 18897 6502 18949 6554
rect 18961 6502 19013 6554
rect 2964 6400 3016 6452
rect 7196 6400 7248 6452
rect 10508 6400 10560 6452
rect 16120 6400 16172 6452
rect 17776 6400 17828 6452
rect 18052 6443 18104 6452
rect 18052 6409 18061 6443
rect 18061 6409 18095 6443
rect 18095 6409 18104 6443
rect 18052 6400 18104 6409
rect 2872 6196 2924 6248
rect 3056 6307 3108 6316
rect 3056 6273 3065 6307
rect 3065 6273 3099 6307
rect 3099 6273 3108 6307
rect 3976 6307 4028 6316
rect 3056 6264 3108 6273
rect 3976 6273 3985 6307
rect 3985 6273 4019 6307
rect 4019 6273 4028 6307
rect 3976 6264 4028 6273
rect 5080 6332 5132 6384
rect 8024 6332 8076 6384
rect 8392 6332 8444 6384
rect 9036 6332 9088 6384
rect 4620 6307 4672 6316
rect 4620 6273 4629 6307
rect 4629 6273 4663 6307
rect 4663 6273 4672 6307
rect 4620 6264 4672 6273
rect 5172 6264 5224 6316
rect 6736 6307 6788 6316
rect 6736 6273 6745 6307
rect 6745 6273 6779 6307
rect 6779 6273 6788 6307
rect 6736 6264 6788 6273
rect 7656 6307 7708 6316
rect 7656 6273 7665 6307
rect 7665 6273 7699 6307
rect 7699 6273 7708 6307
rect 7656 6264 7708 6273
rect 8208 6264 8260 6316
rect 9404 6307 9456 6316
rect 9404 6273 9413 6307
rect 9413 6273 9447 6307
rect 9447 6273 9456 6307
rect 9404 6264 9456 6273
rect 10692 6332 10744 6384
rect 17224 6332 17276 6384
rect 11704 6307 11756 6316
rect 11704 6273 11713 6307
rect 11713 6273 11747 6307
rect 11747 6273 11756 6307
rect 11704 6264 11756 6273
rect 11888 6264 11940 6316
rect 12808 6264 12860 6316
rect 13268 6264 13320 6316
rect 16856 6307 16908 6316
rect 16856 6273 16865 6307
rect 16865 6273 16899 6307
rect 16899 6273 16908 6307
rect 16856 6264 16908 6273
rect 17040 6307 17092 6316
rect 17040 6273 17049 6307
rect 17049 6273 17083 6307
rect 17083 6273 17092 6307
rect 17040 6264 17092 6273
rect 3240 6196 3292 6248
rect 2228 6128 2280 6180
rect 6920 6128 6972 6180
rect 8760 6196 8812 6248
rect 10324 6196 10376 6248
rect 13452 6196 13504 6248
rect 13544 6196 13596 6248
rect 15752 6196 15804 6248
rect 16948 6196 17000 6248
rect 17868 6307 17920 6316
rect 17868 6273 17877 6307
rect 17877 6273 17911 6307
rect 17911 6273 17920 6307
rect 17868 6264 17920 6273
rect 11428 6128 11480 6180
rect 13728 6128 13780 6180
rect 15660 6128 15712 6180
rect 17408 6128 17460 6180
rect 4160 6103 4212 6112
rect 4160 6069 4169 6103
rect 4169 6069 4203 6103
rect 4203 6069 4212 6103
rect 4160 6060 4212 6069
rect 5264 6060 5316 6112
rect 8484 6060 8536 6112
rect 11796 6060 11848 6112
rect 13452 6103 13504 6112
rect 13452 6069 13461 6103
rect 13461 6069 13495 6103
rect 13495 6069 13504 6103
rect 16212 6103 16264 6112
rect 13452 6060 13504 6069
rect 16212 6069 16221 6103
rect 16221 6069 16255 6103
rect 16255 6069 16264 6103
rect 16212 6060 16264 6069
rect 3169 5958 3221 6010
rect 3233 5958 3285 6010
rect 3297 5958 3349 6010
rect 3361 5958 3413 6010
rect 3425 5958 3477 6010
rect 7608 5958 7660 6010
rect 7672 5958 7724 6010
rect 7736 5958 7788 6010
rect 7800 5958 7852 6010
rect 7864 5958 7916 6010
rect 12047 5958 12099 6010
rect 12111 5958 12163 6010
rect 12175 5958 12227 6010
rect 12239 5958 12291 6010
rect 12303 5958 12355 6010
rect 16486 5958 16538 6010
rect 16550 5958 16602 6010
rect 16614 5958 16666 6010
rect 16678 5958 16730 6010
rect 16742 5958 16794 6010
rect 3700 5856 3752 5908
rect 4068 5856 4120 5908
rect 3056 5831 3108 5840
rect 3056 5797 3065 5831
rect 3065 5797 3099 5831
rect 3099 5797 3108 5831
rect 3056 5788 3108 5797
rect 6092 5856 6144 5908
rect 2964 5652 3016 5704
rect 4068 5720 4120 5772
rect 5908 5788 5960 5840
rect 4620 5720 4672 5772
rect 11428 5899 11480 5908
rect 11428 5865 11437 5899
rect 11437 5865 11471 5899
rect 11471 5865 11480 5899
rect 11428 5856 11480 5865
rect 11888 5856 11940 5908
rect 14648 5856 14700 5908
rect 15936 5899 15988 5908
rect 15936 5865 15945 5899
rect 15945 5865 15979 5899
rect 15979 5865 15988 5899
rect 15936 5856 15988 5865
rect 7932 5788 7984 5840
rect 7288 5720 7340 5772
rect 8116 5720 8168 5772
rect 2872 5627 2924 5636
rect 2872 5593 2881 5627
rect 2881 5593 2915 5627
rect 2915 5593 2924 5627
rect 2872 5584 2924 5593
rect 6368 5652 6420 5704
rect 7012 5695 7064 5704
rect 7012 5661 7021 5695
rect 7021 5661 7055 5695
rect 7055 5661 7064 5695
rect 7012 5652 7064 5661
rect 8208 5652 8260 5704
rect 8484 5695 8536 5704
rect 8484 5661 8493 5695
rect 8493 5661 8527 5695
rect 8527 5661 8536 5695
rect 8484 5652 8536 5661
rect 8576 5695 8628 5704
rect 8576 5661 8585 5695
rect 8585 5661 8619 5695
rect 8619 5661 8628 5695
rect 8576 5652 8628 5661
rect 10416 5788 10468 5840
rect 10324 5720 10376 5772
rect 10416 5695 10468 5704
rect 10416 5661 10425 5695
rect 10425 5661 10459 5695
rect 10459 5661 10468 5695
rect 10416 5652 10468 5661
rect 10692 5720 10744 5772
rect 11152 5652 11204 5704
rect 6552 5584 6604 5636
rect 6184 5516 6236 5568
rect 7472 5559 7524 5568
rect 7472 5525 7481 5559
rect 7481 5525 7515 5559
rect 7515 5525 7524 5559
rect 7472 5516 7524 5525
rect 10232 5516 10284 5568
rect 12808 5720 12860 5772
rect 17316 5856 17368 5908
rect 17868 5856 17920 5908
rect 17960 5856 18012 5908
rect 13084 5695 13136 5704
rect 13084 5661 13093 5695
rect 13093 5661 13127 5695
rect 13127 5661 13136 5695
rect 13084 5652 13136 5661
rect 13268 5695 13320 5704
rect 13268 5661 13277 5695
rect 13277 5661 13311 5695
rect 13311 5661 13320 5695
rect 13268 5652 13320 5661
rect 13544 5695 13596 5704
rect 13544 5661 13553 5695
rect 13553 5661 13587 5695
rect 13587 5661 13596 5695
rect 13544 5652 13596 5661
rect 14648 5652 14700 5704
rect 17592 5720 17644 5772
rect 15752 5695 15804 5704
rect 15752 5661 15761 5695
rect 15761 5661 15795 5695
rect 15795 5661 15804 5695
rect 15752 5652 15804 5661
rect 17684 5652 17736 5704
rect 16028 5584 16080 5636
rect 17408 5627 17460 5636
rect 17408 5593 17417 5627
rect 17417 5593 17451 5627
rect 17451 5593 17460 5627
rect 17408 5584 17460 5593
rect 10784 5516 10836 5568
rect 14188 5516 14240 5568
rect 16212 5516 16264 5568
rect 16304 5516 16356 5568
rect 5388 5414 5440 5466
rect 5452 5414 5504 5466
rect 5516 5414 5568 5466
rect 5580 5414 5632 5466
rect 5644 5414 5696 5466
rect 9827 5414 9879 5466
rect 9891 5414 9943 5466
rect 9955 5414 10007 5466
rect 10019 5414 10071 5466
rect 10083 5414 10135 5466
rect 14266 5414 14318 5466
rect 14330 5414 14382 5466
rect 14394 5414 14446 5466
rect 14458 5414 14510 5466
rect 14522 5414 14574 5466
rect 18705 5414 18757 5466
rect 18769 5414 18821 5466
rect 18833 5414 18885 5466
rect 18897 5414 18949 5466
rect 18961 5414 19013 5466
rect 2964 5312 3016 5364
rect 3976 5312 4028 5364
rect 5908 5355 5960 5364
rect 5908 5321 5917 5355
rect 5917 5321 5951 5355
rect 5951 5321 5960 5355
rect 5908 5312 5960 5321
rect 6920 5355 6972 5364
rect 6920 5321 6929 5355
rect 6929 5321 6963 5355
rect 6963 5321 6972 5355
rect 6920 5312 6972 5321
rect 11060 5312 11112 5364
rect 11704 5312 11756 5364
rect 14188 5312 14240 5364
rect 17040 5312 17092 5364
rect 3516 5176 3568 5228
rect 4620 5244 4672 5296
rect 7012 5244 7064 5296
rect 9680 5244 9732 5296
rect 4160 5176 4212 5228
rect 7104 5176 7156 5228
rect 11152 5219 11204 5228
rect 11152 5185 11161 5219
rect 11161 5185 11195 5219
rect 11195 5185 11204 5219
rect 11152 5176 11204 5185
rect 8668 5108 8720 5160
rect 9956 5108 10008 5160
rect 11796 5108 11848 5160
rect 14004 5176 14056 5228
rect 15844 5176 15896 5228
rect 16028 5219 16080 5228
rect 16028 5185 16037 5219
rect 16037 5185 16071 5219
rect 16071 5185 16080 5219
rect 16028 5176 16080 5185
rect 17132 5244 17184 5296
rect 16948 5176 17000 5228
rect 17040 5176 17092 5228
rect 17960 5312 18012 5364
rect 17592 5287 17644 5296
rect 17592 5253 17601 5287
rect 17601 5253 17635 5287
rect 17635 5253 17644 5287
rect 17592 5244 17644 5253
rect 6368 4972 6420 5024
rect 7104 4972 7156 5024
rect 11428 4972 11480 5024
rect 13268 5015 13320 5024
rect 13268 4981 13277 5015
rect 13277 4981 13311 5015
rect 13311 4981 13320 5015
rect 13268 4972 13320 4981
rect 15936 4972 15988 5024
rect 17408 4972 17460 5024
rect 17776 5015 17828 5024
rect 17776 4981 17785 5015
rect 17785 4981 17819 5015
rect 17819 4981 17828 5015
rect 17776 4972 17828 4981
rect 3169 4870 3221 4922
rect 3233 4870 3285 4922
rect 3297 4870 3349 4922
rect 3361 4870 3413 4922
rect 3425 4870 3477 4922
rect 7608 4870 7660 4922
rect 7672 4870 7724 4922
rect 7736 4870 7788 4922
rect 7800 4870 7852 4922
rect 7864 4870 7916 4922
rect 12047 4870 12099 4922
rect 12111 4870 12163 4922
rect 12175 4870 12227 4922
rect 12239 4870 12291 4922
rect 12303 4870 12355 4922
rect 16486 4870 16538 4922
rect 16550 4870 16602 4922
rect 16614 4870 16666 4922
rect 16678 4870 16730 4922
rect 16742 4870 16794 4922
rect 2964 4811 3016 4820
rect 2964 4777 2973 4811
rect 2973 4777 3007 4811
rect 3007 4777 3016 4811
rect 2964 4768 3016 4777
rect 3516 4768 3568 4820
rect 5080 4768 5132 4820
rect 6736 4811 6788 4820
rect 6736 4777 6745 4811
rect 6745 4777 6779 4811
rect 6779 4777 6788 4811
rect 6736 4768 6788 4777
rect 9128 4768 9180 4820
rect 10232 4768 10284 4820
rect 10784 4811 10836 4820
rect 10784 4777 10793 4811
rect 10793 4777 10827 4811
rect 10827 4777 10836 4811
rect 10784 4768 10836 4777
rect 14188 4768 14240 4820
rect 15844 4811 15896 4820
rect 15844 4777 15853 4811
rect 15853 4777 15887 4811
rect 15887 4777 15896 4811
rect 15844 4768 15896 4777
rect 16948 4768 17000 4820
rect 18144 4811 18196 4820
rect 13728 4743 13780 4752
rect 2872 4675 2924 4684
rect 2872 4641 2881 4675
rect 2881 4641 2915 4675
rect 2915 4641 2924 4675
rect 2872 4632 2924 4641
rect 4620 4632 4672 4684
rect 5264 4632 5316 4684
rect 7196 4675 7248 4684
rect 7196 4641 7205 4675
rect 7205 4641 7239 4675
rect 7239 4641 7248 4675
rect 7196 4632 7248 4641
rect 3056 4564 3108 4616
rect 5908 4564 5960 4616
rect 6368 4607 6420 4616
rect 6368 4573 6377 4607
rect 6377 4573 6411 4607
rect 6411 4573 6420 4607
rect 6368 4564 6420 4573
rect 7288 4564 7340 4616
rect 7932 4564 7984 4616
rect 10324 4632 10376 4684
rect 10416 4564 10468 4616
rect 13728 4709 13737 4743
rect 13737 4709 13771 4743
rect 13771 4709 13780 4743
rect 15936 4743 15988 4752
rect 13728 4700 13780 4709
rect 13268 4632 13320 4684
rect 14648 4632 14700 4684
rect 15936 4709 15945 4743
rect 15945 4709 15979 4743
rect 15979 4709 15988 4743
rect 15936 4700 15988 4709
rect 16028 4700 16080 4752
rect 7564 4496 7616 4548
rect 9956 4539 10008 4548
rect 9956 4505 9983 4539
rect 9983 4505 10008 4539
rect 9956 4496 10008 4505
rect 10508 4496 10560 4548
rect 11060 4496 11112 4548
rect 9680 4428 9732 4480
rect 10416 4428 10468 4480
rect 10692 4428 10744 4480
rect 13084 4496 13136 4548
rect 16212 4496 16264 4548
rect 16396 4496 16448 4548
rect 11612 4471 11664 4480
rect 11612 4437 11621 4471
rect 11621 4437 11655 4471
rect 11655 4437 11664 4471
rect 11612 4428 11664 4437
rect 16488 4471 16540 4480
rect 16488 4437 16497 4471
rect 16497 4437 16531 4471
rect 16531 4437 16540 4471
rect 16488 4428 16540 4437
rect 17776 4700 17828 4752
rect 17224 4564 17276 4616
rect 18144 4777 18153 4811
rect 18153 4777 18187 4811
rect 18187 4777 18196 4811
rect 18144 4768 18196 4777
rect 17132 4496 17184 4548
rect 17040 4428 17092 4480
rect 5388 4326 5440 4378
rect 5452 4326 5504 4378
rect 5516 4326 5568 4378
rect 5580 4326 5632 4378
rect 5644 4326 5696 4378
rect 9827 4326 9879 4378
rect 9891 4326 9943 4378
rect 9955 4326 10007 4378
rect 10019 4326 10071 4378
rect 10083 4326 10135 4378
rect 14266 4326 14318 4378
rect 14330 4326 14382 4378
rect 14394 4326 14446 4378
rect 14458 4326 14510 4378
rect 14522 4326 14574 4378
rect 18705 4326 18757 4378
rect 18769 4326 18821 4378
rect 18833 4326 18885 4378
rect 18897 4326 18949 4378
rect 18961 4326 19013 4378
rect 5172 4224 5224 4276
rect 8484 4224 8536 4276
rect 10692 4267 10744 4276
rect 10692 4233 10701 4267
rect 10701 4233 10735 4267
rect 10735 4233 10744 4267
rect 10692 4224 10744 4233
rect 11152 4224 11204 4276
rect 14648 4224 14700 4276
rect 16948 4224 17000 4276
rect 17592 4224 17644 4276
rect 6552 4063 6604 4072
rect 6552 4029 6561 4063
rect 6561 4029 6595 4063
rect 6595 4029 6604 4063
rect 6552 4020 6604 4029
rect 7380 4088 7432 4140
rect 7564 4088 7616 4140
rect 11612 4156 11664 4208
rect 7932 4063 7984 4072
rect 6736 3952 6788 4004
rect 7380 3952 7432 4004
rect 7932 4029 7941 4063
rect 7941 4029 7975 4063
rect 7975 4029 7984 4063
rect 7932 4020 7984 4029
rect 8668 4088 8720 4140
rect 9588 4131 9640 4140
rect 9588 4097 9622 4131
rect 9622 4097 9640 4131
rect 9588 4088 9640 4097
rect 14004 4088 14056 4140
rect 17132 4156 17184 4208
rect 16304 4131 16356 4140
rect 9312 4063 9364 4072
rect 9312 4029 9321 4063
rect 9321 4029 9355 4063
rect 9355 4029 9364 4063
rect 9312 4020 9364 4029
rect 11704 4063 11756 4072
rect 11704 4029 11713 4063
rect 11713 4029 11747 4063
rect 11747 4029 11756 4063
rect 11704 4020 11756 4029
rect 16304 4097 16313 4131
rect 16313 4097 16347 4131
rect 16347 4097 16356 4131
rect 16304 4088 16356 4097
rect 16580 4088 16632 4140
rect 16488 4020 16540 4072
rect 4712 3927 4764 3936
rect 4712 3893 4721 3927
rect 4721 3893 4755 3927
rect 4755 3893 4764 3927
rect 4712 3884 4764 3893
rect 7012 3927 7064 3936
rect 7012 3893 7021 3927
rect 7021 3893 7055 3927
rect 7055 3893 7064 3927
rect 7012 3884 7064 3893
rect 7288 3884 7340 3936
rect 8392 3927 8444 3936
rect 8392 3893 8401 3927
rect 8401 3893 8435 3927
rect 8435 3893 8444 3927
rect 8392 3884 8444 3893
rect 16948 3884 17000 3936
rect 17868 3927 17920 3936
rect 17868 3893 17877 3927
rect 17877 3893 17911 3927
rect 17911 3893 17920 3927
rect 17868 3884 17920 3893
rect 3169 3782 3221 3834
rect 3233 3782 3285 3834
rect 3297 3782 3349 3834
rect 3361 3782 3413 3834
rect 3425 3782 3477 3834
rect 7608 3782 7660 3834
rect 7672 3782 7724 3834
rect 7736 3782 7788 3834
rect 7800 3782 7852 3834
rect 7864 3782 7916 3834
rect 12047 3782 12099 3834
rect 12111 3782 12163 3834
rect 12175 3782 12227 3834
rect 12239 3782 12291 3834
rect 12303 3782 12355 3834
rect 16486 3782 16538 3834
rect 16550 3782 16602 3834
rect 16614 3782 16666 3834
rect 16678 3782 16730 3834
rect 16742 3782 16794 3834
rect 8300 3680 8352 3732
rect 9588 3680 9640 3732
rect 13268 3680 13320 3732
rect 15108 3680 15160 3732
rect 16580 3680 16632 3732
rect 16856 3680 16908 3732
rect 6552 3612 6604 3664
rect 5264 3476 5316 3528
rect 6184 3519 6236 3528
rect 6184 3485 6193 3519
rect 6193 3485 6227 3519
rect 6227 3485 6236 3519
rect 6184 3476 6236 3485
rect 7012 3544 7064 3596
rect 7288 3612 7340 3664
rect 7380 3612 7432 3664
rect 8392 3612 8444 3664
rect 9036 3612 9088 3664
rect 12992 3612 13044 3664
rect 7932 3544 7984 3596
rect 6460 3519 6512 3528
rect 6460 3485 6469 3519
rect 6469 3485 6503 3519
rect 6503 3485 6512 3519
rect 6460 3476 6512 3485
rect 6828 3476 6880 3528
rect 7472 3476 7524 3528
rect 8392 3519 8444 3528
rect 6368 3408 6420 3460
rect 7104 3408 7156 3460
rect 8392 3485 8401 3519
rect 8401 3485 8435 3519
rect 8435 3485 8444 3519
rect 8392 3476 8444 3485
rect 8484 3476 8536 3528
rect 9680 3476 9732 3528
rect 11796 3544 11848 3596
rect 18144 3612 18196 3664
rect 11244 3519 11296 3528
rect 7932 3408 7984 3460
rect 11244 3485 11253 3519
rect 11253 3485 11287 3519
rect 11287 3485 11296 3519
rect 11244 3476 11296 3485
rect 12808 3476 12860 3528
rect 12992 3519 13044 3528
rect 12992 3485 13001 3519
rect 13001 3485 13035 3519
rect 13035 3485 13044 3519
rect 13728 3544 13780 3596
rect 12992 3476 13044 3485
rect 13268 3519 13320 3528
rect 13268 3485 13277 3519
rect 13277 3485 13311 3519
rect 13311 3485 13320 3519
rect 13268 3476 13320 3485
rect 13452 3476 13504 3528
rect 11336 3408 11388 3460
rect 16580 3408 16632 3460
rect 16948 3451 17000 3460
rect 16948 3417 16957 3451
rect 16957 3417 16991 3451
rect 16991 3417 17000 3451
rect 16948 3408 17000 3417
rect 17132 3451 17184 3460
rect 17132 3417 17157 3451
rect 17157 3417 17184 3451
rect 17132 3408 17184 3417
rect 3976 3383 4028 3392
rect 3976 3349 3985 3383
rect 3985 3349 4019 3383
rect 4019 3349 4028 3383
rect 3976 3340 4028 3349
rect 6920 3340 6972 3392
rect 10324 3340 10376 3392
rect 11152 3340 11204 3392
rect 11796 3340 11848 3392
rect 12716 3383 12768 3392
rect 12716 3349 12725 3383
rect 12725 3349 12759 3383
rect 12759 3349 12768 3383
rect 12716 3340 12768 3349
rect 13636 3340 13688 3392
rect 16120 3340 16172 3392
rect 17408 3340 17460 3392
rect 18604 3340 18656 3392
rect 5388 3238 5440 3290
rect 5452 3238 5504 3290
rect 5516 3238 5568 3290
rect 5580 3238 5632 3290
rect 5644 3238 5696 3290
rect 9827 3238 9879 3290
rect 9891 3238 9943 3290
rect 9955 3238 10007 3290
rect 10019 3238 10071 3290
rect 10083 3238 10135 3290
rect 14266 3238 14318 3290
rect 14330 3238 14382 3290
rect 14394 3238 14446 3290
rect 14458 3238 14510 3290
rect 14522 3238 14574 3290
rect 18705 3238 18757 3290
rect 18769 3238 18821 3290
rect 18833 3238 18885 3290
rect 18897 3238 18949 3290
rect 18961 3238 19013 3290
rect 6368 3136 6420 3188
rect 4528 3000 4580 3052
rect 5264 3068 5316 3120
rect 4712 3000 4764 3052
rect 7104 3136 7156 3188
rect 7380 3136 7432 3188
rect 11336 3136 11388 3188
rect 13452 3136 13504 3188
rect 17224 3179 17276 3188
rect 6920 3068 6972 3120
rect 7012 3043 7064 3052
rect 6552 2932 6604 2984
rect 7012 3009 7021 3043
rect 7021 3009 7055 3043
rect 7055 3009 7064 3043
rect 7012 3000 7064 3009
rect 4252 2796 4304 2848
rect 6000 2839 6052 2848
rect 6000 2805 6009 2839
rect 6009 2805 6043 2839
rect 6043 2805 6052 2839
rect 6000 2796 6052 2805
rect 6184 2796 6236 2848
rect 7196 3000 7248 3052
rect 9312 3000 9364 3052
rect 10324 3000 10376 3052
rect 16580 3068 16632 3120
rect 17224 3145 17233 3179
rect 17233 3145 17267 3179
rect 17267 3145 17276 3179
rect 17224 3136 17276 3145
rect 17316 3111 17368 3120
rect 17316 3077 17325 3111
rect 17325 3077 17359 3111
rect 17359 3077 17368 3111
rect 17316 3068 17368 3077
rect 17868 3068 17920 3120
rect 11704 3043 11756 3052
rect 11704 3009 11713 3043
rect 11713 3009 11747 3043
rect 11747 3009 11756 3043
rect 11704 3000 11756 3009
rect 11060 2932 11112 2984
rect 14004 3043 14056 3052
rect 14004 3009 14013 3043
rect 14013 3009 14047 3043
rect 14047 3009 14056 3043
rect 14004 3000 14056 3009
rect 15752 3000 15804 3052
rect 15936 3043 15988 3052
rect 15936 3009 15945 3043
rect 15945 3009 15979 3043
rect 15979 3009 15988 3043
rect 15936 3000 15988 3009
rect 17040 3000 17092 3052
rect 18144 3043 18196 3052
rect 18144 3009 18153 3043
rect 18153 3009 18187 3043
rect 18187 3009 18196 3043
rect 18144 3000 18196 3009
rect 17408 2975 17460 2984
rect 17408 2941 17417 2975
rect 17417 2941 17451 2975
rect 17451 2941 17460 2975
rect 17408 2932 17460 2941
rect 8668 2796 8720 2848
rect 16856 2839 16908 2848
rect 16856 2805 16865 2839
rect 16865 2805 16899 2839
rect 16899 2805 16908 2839
rect 16856 2796 16908 2805
rect 18052 2839 18104 2848
rect 18052 2805 18061 2839
rect 18061 2805 18095 2839
rect 18095 2805 18104 2839
rect 18052 2796 18104 2805
rect 3169 2694 3221 2746
rect 3233 2694 3285 2746
rect 3297 2694 3349 2746
rect 3361 2694 3413 2746
rect 3425 2694 3477 2746
rect 7608 2694 7660 2746
rect 7672 2694 7724 2746
rect 7736 2694 7788 2746
rect 7800 2694 7852 2746
rect 7864 2694 7916 2746
rect 12047 2694 12099 2746
rect 12111 2694 12163 2746
rect 12175 2694 12227 2746
rect 12239 2694 12291 2746
rect 12303 2694 12355 2746
rect 16486 2694 16538 2746
rect 16550 2694 16602 2746
rect 16614 2694 16666 2746
rect 16678 2694 16730 2746
rect 16742 2694 16794 2746
rect 4528 2592 4580 2644
rect 3976 2388 4028 2440
rect 4252 2431 4304 2440
rect 4252 2397 4261 2431
rect 4261 2397 4295 2431
rect 4295 2397 4304 2431
rect 4252 2388 4304 2397
rect 6460 2524 6512 2576
rect 11244 2592 11296 2644
rect 11796 2635 11848 2644
rect 11796 2601 11805 2635
rect 11805 2601 11839 2635
rect 11839 2601 11848 2635
rect 11796 2592 11848 2601
rect 11060 2524 11112 2576
rect 13728 2592 13780 2644
rect 6920 2456 6972 2508
rect 6000 2431 6052 2440
rect 6000 2397 6009 2431
rect 6009 2397 6043 2431
rect 6043 2397 6052 2431
rect 6000 2388 6052 2397
rect 6552 2431 6604 2440
rect 6552 2397 6561 2431
rect 6561 2397 6595 2431
rect 6595 2397 6604 2431
rect 6552 2388 6604 2397
rect 6736 2388 6788 2440
rect 7932 2388 7984 2440
rect 8668 2388 8720 2440
rect 9220 2388 9272 2440
rect 11704 2388 11756 2440
rect 14004 2456 14056 2508
rect 15936 2592 15988 2644
rect 16948 2592 17000 2644
rect 17224 2524 17276 2576
rect 15752 2456 15804 2508
rect 16856 2388 16908 2440
rect 17316 2388 17368 2440
rect 7380 2320 7432 2372
rect 9036 2320 9088 2372
rect 12716 2320 12768 2372
rect 18052 2320 18104 2372
rect 1216 2252 1268 2304
rect 3700 2252 3752 2304
rect 6184 2252 6236 2304
rect 8668 2252 8720 2304
rect 5388 2150 5440 2202
rect 5452 2150 5504 2202
rect 5516 2150 5568 2202
rect 5580 2150 5632 2202
rect 5644 2150 5696 2202
rect 9827 2150 9879 2202
rect 9891 2150 9943 2202
rect 9955 2150 10007 2202
rect 10019 2150 10071 2202
rect 10083 2150 10135 2202
rect 14266 2150 14318 2202
rect 14330 2150 14382 2202
rect 14394 2150 14446 2202
rect 14458 2150 14510 2202
rect 14522 2150 14574 2202
rect 18705 2150 18757 2202
rect 18769 2150 18821 2202
rect 18833 2150 18885 2202
rect 18897 2150 18949 2202
rect 18961 2150 19013 2202
<< metal2 >>
rect 3330 19200 3386 20000
rect 9954 19200 10010 20000
rect 10060 19230 10364 19258
rect 2780 17196 2832 17202
rect 2780 17138 2832 17144
rect 2792 16794 2820 17138
rect 3344 16980 3372 19200
rect 9968 19122 9996 19200
rect 10060 19122 10088 19230
rect 9968 19094 10088 19122
rect 5388 17436 5696 17445
rect 5388 17434 5394 17436
rect 5450 17434 5474 17436
rect 5530 17434 5554 17436
rect 5610 17434 5634 17436
rect 5690 17434 5696 17436
rect 5450 17382 5452 17434
rect 5632 17382 5634 17434
rect 5388 17380 5394 17382
rect 5450 17380 5474 17382
rect 5530 17380 5554 17382
rect 5610 17380 5634 17382
rect 5690 17380 5696 17382
rect 5388 17371 5696 17380
rect 9827 17436 10135 17445
rect 9827 17434 9833 17436
rect 9889 17434 9913 17436
rect 9969 17434 9993 17436
rect 10049 17434 10073 17436
rect 10129 17434 10135 17436
rect 9889 17382 9891 17434
rect 10071 17382 10073 17434
rect 9827 17380 9833 17382
rect 9889 17380 9913 17382
rect 9969 17380 9993 17382
rect 10049 17380 10073 17382
rect 10129 17380 10135 17382
rect 9827 17371 10135 17380
rect 10336 17202 10364 19230
rect 16578 19200 16634 20000
rect 14266 17436 14574 17445
rect 14266 17434 14272 17436
rect 14328 17434 14352 17436
rect 14408 17434 14432 17436
rect 14488 17434 14512 17436
rect 14568 17434 14574 17436
rect 14328 17382 14330 17434
rect 14510 17382 14512 17434
rect 14266 17380 14272 17382
rect 14328 17380 14352 17382
rect 14408 17380 14432 17382
rect 14488 17380 14512 17382
rect 14568 17380 14574 17382
rect 14266 17371 14574 17380
rect 16592 17338 16620 19200
rect 18705 17436 19013 17445
rect 18705 17434 18711 17436
rect 18767 17434 18791 17436
rect 18847 17434 18871 17436
rect 18927 17434 18951 17436
rect 19007 17434 19013 17436
rect 18767 17382 18769 17434
rect 18949 17382 18951 17434
rect 18705 17380 18711 17382
rect 18767 17380 18791 17382
rect 18847 17380 18871 17382
rect 18927 17380 18951 17382
rect 19007 17380 19013 17382
rect 18705 17371 19013 17380
rect 16580 17332 16632 17338
rect 16580 17274 16632 17280
rect 6552 17196 6604 17202
rect 6552 17138 6604 17144
rect 7196 17196 7248 17202
rect 7196 17138 7248 17144
rect 9312 17196 9364 17202
rect 9312 17138 9364 17144
rect 10140 17196 10192 17202
rect 10324 17196 10376 17202
rect 10192 17156 10272 17184
rect 10140 17138 10192 17144
rect 5356 17128 5408 17134
rect 5356 17070 5408 17076
rect 4252 17060 4304 17066
rect 4252 17002 4304 17008
rect 3976 16992 4028 16998
rect 3344 16952 3556 16980
rect 3169 16892 3477 16901
rect 3169 16890 3175 16892
rect 3231 16890 3255 16892
rect 3311 16890 3335 16892
rect 3391 16890 3415 16892
rect 3471 16890 3477 16892
rect 3231 16838 3233 16890
rect 3413 16838 3415 16890
rect 3169 16836 3175 16838
rect 3231 16836 3255 16838
rect 3311 16836 3335 16838
rect 3391 16836 3415 16838
rect 3471 16836 3477 16838
rect 3169 16827 3477 16836
rect 2780 16788 2832 16794
rect 2780 16730 2832 16736
rect 3528 15910 3556 16952
rect 3976 16934 4028 16940
rect 3988 16590 4016 16934
rect 3976 16584 4028 16590
rect 3976 16526 4028 16532
rect 3700 16448 3752 16454
rect 3700 16390 3752 16396
rect 3712 16114 3740 16390
rect 4264 16182 4292 17002
rect 5368 16590 5396 17070
rect 6000 16992 6052 16998
rect 6000 16934 6052 16940
rect 4988 16584 5040 16590
rect 4988 16526 5040 16532
rect 5356 16584 5408 16590
rect 5356 16526 5408 16532
rect 4252 16176 4304 16182
rect 4252 16118 4304 16124
rect 3700 16108 3752 16114
rect 3700 16050 3752 16056
rect 3056 15904 3108 15910
rect 3056 15846 3108 15852
rect 3516 15904 3568 15910
rect 3516 15846 3568 15852
rect 3068 15502 3096 15846
rect 3169 15804 3477 15813
rect 3169 15802 3175 15804
rect 3231 15802 3255 15804
rect 3311 15802 3335 15804
rect 3391 15802 3415 15804
rect 3471 15802 3477 15804
rect 3231 15750 3233 15802
rect 3413 15750 3415 15802
rect 3169 15748 3175 15750
rect 3231 15748 3255 15750
rect 3311 15748 3335 15750
rect 3391 15748 3415 15750
rect 3471 15748 3477 15750
rect 3169 15739 3477 15748
rect 3056 15496 3108 15502
rect 3056 15438 3108 15444
rect 2780 15360 2832 15366
rect 2780 15302 2832 15308
rect 2320 13932 2372 13938
rect 2320 13874 2372 13880
rect 2688 13932 2740 13938
rect 2688 13874 2740 13880
rect 2332 13530 2360 13874
rect 2596 13864 2648 13870
rect 2596 13806 2648 13812
rect 2320 13524 2372 13530
rect 2320 13466 2372 13472
rect 2228 13320 2280 13326
rect 2228 13262 2280 13268
rect 2240 12238 2268 13262
rect 2608 13258 2636 13806
rect 2700 13326 2728 13874
rect 2688 13320 2740 13326
rect 2688 13262 2740 13268
rect 2596 13252 2648 13258
rect 2596 13194 2648 13200
rect 2608 12918 2636 13194
rect 2412 12912 2464 12918
rect 2412 12854 2464 12860
rect 2596 12912 2648 12918
rect 2596 12854 2648 12860
rect 2424 12238 2452 12854
rect 2504 12844 2556 12850
rect 2504 12786 2556 12792
rect 2516 12442 2544 12786
rect 2596 12708 2648 12714
rect 2596 12650 2648 12656
rect 2504 12436 2556 12442
rect 2504 12378 2556 12384
rect 2608 12238 2636 12650
rect 2228 12232 2280 12238
rect 2228 12174 2280 12180
rect 2412 12232 2464 12238
rect 2412 12174 2464 12180
rect 2596 12232 2648 12238
rect 2596 12174 2648 12180
rect 2424 11218 2452 12174
rect 2412 11212 2464 11218
rect 2412 11154 2464 11160
rect 2792 10674 2820 15302
rect 3056 15020 3108 15026
rect 3056 14962 3108 14968
rect 3068 13802 3096 14962
rect 3169 14716 3477 14725
rect 3169 14714 3175 14716
rect 3231 14714 3255 14716
rect 3311 14714 3335 14716
rect 3391 14714 3415 14716
rect 3471 14714 3477 14716
rect 3231 14662 3233 14714
rect 3413 14662 3415 14714
rect 3169 14660 3175 14662
rect 3231 14660 3255 14662
rect 3311 14660 3335 14662
rect 3391 14660 3415 14662
rect 3471 14660 3477 14662
rect 3169 14651 3477 14660
rect 3056 13796 3108 13802
rect 3056 13738 3108 13744
rect 3169 13628 3477 13637
rect 3169 13626 3175 13628
rect 3231 13626 3255 13628
rect 3311 13626 3335 13628
rect 3391 13626 3415 13628
rect 3471 13626 3477 13628
rect 3231 13574 3233 13626
rect 3413 13574 3415 13626
rect 3169 13572 3175 13574
rect 3231 13572 3255 13574
rect 3311 13572 3335 13574
rect 3391 13572 3415 13574
rect 3471 13572 3477 13574
rect 3169 13563 3477 13572
rect 3169 12540 3477 12549
rect 3169 12538 3175 12540
rect 3231 12538 3255 12540
rect 3311 12538 3335 12540
rect 3391 12538 3415 12540
rect 3471 12538 3477 12540
rect 3231 12486 3233 12538
rect 3413 12486 3415 12538
rect 3169 12484 3175 12486
rect 3231 12484 3255 12486
rect 3311 12484 3335 12486
rect 3391 12484 3415 12486
rect 3471 12484 3477 12486
rect 3169 12475 3477 12484
rect 2872 12232 2924 12238
rect 2872 12174 2924 12180
rect 2884 11354 2912 12174
rect 3056 12096 3108 12102
rect 3056 12038 3108 12044
rect 3068 11762 3096 12038
rect 3056 11756 3108 11762
rect 3056 11698 3108 11704
rect 3169 11452 3477 11461
rect 3169 11450 3175 11452
rect 3231 11450 3255 11452
rect 3311 11450 3335 11452
rect 3391 11450 3415 11452
rect 3471 11450 3477 11452
rect 3231 11398 3233 11450
rect 3413 11398 3415 11450
rect 3169 11396 3175 11398
rect 3231 11396 3255 11398
rect 3311 11396 3335 11398
rect 3391 11396 3415 11398
rect 3471 11396 3477 11398
rect 3169 11387 3477 11396
rect 2872 11348 2924 11354
rect 2872 11290 2924 11296
rect 3240 11144 3292 11150
rect 3240 11086 3292 11092
rect 3252 10674 3280 11086
rect 2780 10668 2832 10674
rect 2780 10610 2832 10616
rect 3240 10668 3292 10674
rect 3240 10610 3292 10616
rect 2780 10464 2832 10470
rect 2780 10406 2832 10412
rect 2504 9988 2556 9994
rect 2504 9930 2556 9936
rect 2516 9382 2544 9930
rect 2792 9654 2820 10406
rect 3169 10364 3477 10373
rect 3169 10362 3175 10364
rect 3231 10362 3255 10364
rect 3311 10362 3335 10364
rect 3391 10362 3415 10364
rect 3471 10362 3477 10364
rect 3231 10310 3233 10362
rect 3413 10310 3415 10362
rect 3169 10308 3175 10310
rect 3231 10308 3255 10310
rect 3311 10308 3335 10310
rect 3391 10308 3415 10310
rect 3471 10308 3477 10310
rect 3169 10299 3477 10308
rect 3712 10266 3740 16050
rect 5000 16046 5028 16526
rect 5816 16516 5868 16522
rect 5816 16458 5868 16464
rect 5388 16348 5696 16357
rect 5388 16346 5394 16348
rect 5450 16346 5474 16348
rect 5530 16346 5554 16348
rect 5610 16346 5634 16348
rect 5690 16346 5696 16348
rect 5450 16294 5452 16346
rect 5632 16294 5634 16346
rect 5388 16292 5394 16294
rect 5450 16292 5474 16294
rect 5530 16292 5554 16294
rect 5610 16292 5634 16294
rect 5690 16292 5696 16294
rect 5388 16283 5696 16292
rect 5828 16250 5856 16458
rect 5816 16244 5868 16250
rect 5816 16186 5868 16192
rect 6012 16114 6040 16934
rect 6564 16250 6592 17138
rect 7104 17128 7156 17134
rect 7104 17070 7156 17076
rect 6920 16448 6972 16454
rect 6920 16390 6972 16396
rect 6552 16244 6604 16250
rect 6552 16186 6604 16192
rect 6932 16182 6960 16390
rect 6920 16176 6972 16182
rect 6920 16118 6972 16124
rect 6000 16108 6052 16114
rect 6000 16050 6052 16056
rect 7116 16046 7144 17070
rect 7208 16794 7236 17138
rect 7380 16992 7432 16998
rect 7380 16934 7432 16940
rect 8944 16992 8996 16998
rect 8944 16934 8996 16940
rect 7196 16788 7248 16794
rect 7196 16730 7248 16736
rect 7392 16250 7420 16934
rect 7608 16892 7916 16901
rect 7608 16890 7614 16892
rect 7670 16890 7694 16892
rect 7750 16890 7774 16892
rect 7830 16890 7854 16892
rect 7910 16890 7916 16892
rect 7670 16838 7672 16890
rect 7852 16838 7854 16890
rect 7608 16836 7614 16838
rect 7670 16836 7694 16838
rect 7750 16836 7774 16838
rect 7830 16836 7854 16838
rect 7910 16836 7916 16838
rect 7608 16827 7916 16836
rect 8576 16584 8628 16590
rect 8576 16526 8628 16532
rect 7380 16244 7432 16250
rect 7380 16186 7432 16192
rect 8588 16182 8616 16526
rect 8576 16176 8628 16182
rect 8576 16118 8628 16124
rect 8956 16114 8984 16934
rect 9324 16250 9352 17138
rect 9864 17060 9916 17066
rect 9864 17002 9916 17008
rect 9876 16522 9904 17002
rect 9864 16516 9916 16522
rect 9864 16458 9916 16464
rect 9827 16348 10135 16357
rect 9827 16346 9833 16348
rect 9889 16346 9913 16348
rect 9969 16346 9993 16348
rect 10049 16346 10073 16348
rect 10129 16346 10135 16348
rect 9889 16294 9891 16346
rect 10071 16294 10073 16346
rect 9827 16292 9833 16294
rect 9889 16292 9913 16294
rect 9969 16292 9993 16294
rect 10049 16292 10073 16294
rect 10129 16292 10135 16294
rect 9827 16283 10135 16292
rect 10244 16250 10272 17156
rect 10324 17138 10376 17144
rect 12624 17196 12676 17202
rect 12624 17138 12676 17144
rect 10508 16992 10560 16998
rect 10508 16934 10560 16940
rect 10600 16992 10652 16998
rect 10600 16934 10652 16940
rect 10324 16788 10376 16794
rect 10324 16730 10376 16736
rect 9312 16244 9364 16250
rect 9312 16186 9364 16192
rect 10232 16244 10284 16250
rect 10232 16186 10284 16192
rect 9128 16176 9180 16182
rect 9128 16118 9180 16124
rect 8024 16108 8076 16114
rect 8024 16050 8076 16056
rect 8944 16108 8996 16114
rect 8944 16050 8996 16056
rect 4988 16040 5040 16046
rect 4988 15982 5040 15988
rect 7104 16040 7156 16046
rect 7104 15982 7156 15988
rect 5000 15502 5028 15982
rect 4160 15496 4212 15502
rect 4160 15438 4212 15444
rect 4252 15496 4304 15502
rect 4252 15438 4304 15444
rect 4988 15496 5040 15502
rect 4988 15438 5040 15444
rect 3976 15360 4028 15366
rect 3976 15302 4028 15308
rect 3988 14414 4016 15302
rect 4172 15162 4200 15438
rect 4160 15156 4212 15162
rect 4160 15098 4212 15104
rect 4264 15026 4292 15438
rect 5000 15094 5028 15438
rect 6460 15428 6512 15434
rect 6460 15370 6512 15376
rect 5388 15260 5696 15269
rect 5388 15258 5394 15260
rect 5450 15258 5474 15260
rect 5530 15258 5554 15260
rect 5610 15258 5634 15260
rect 5690 15258 5696 15260
rect 5450 15206 5452 15258
rect 5632 15206 5634 15258
rect 5388 15204 5394 15206
rect 5450 15204 5474 15206
rect 5530 15204 5554 15206
rect 5610 15204 5634 15206
rect 5690 15204 5696 15206
rect 5388 15195 5696 15204
rect 4988 15088 5040 15094
rect 4988 15030 5040 15036
rect 4252 15020 4304 15026
rect 4252 14962 4304 14968
rect 3976 14408 4028 14414
rect 3976 14350 4028 14356
rect 4160 13932 4212 13938
rect 4160 13874 4212 13880
rect 4172 12986 4200 13874
rect 4264 13410 4292 14962
rect 5000 14414 5028 15030
rect 5816 14816 5868 14822
rect 5816 14758 5868 14764
rect 5724 14544 5776 14550
rect 5724 14486 5776 14492
rect 4988 14408 5040 14414
rect 4988 14350 5040 14356
rect 4344 13932 4396 13938
rect 4344 13874 4396 13880
rect 4356 13530 4384 13874
rect 5000 13870 5028 14350
rect 5388 14172 5696 14181
rect 5388 14170 5394 14172
rect 5450 14170 5474 14172
rect 5530 14170 5554 14172
rect 5610 14170 5634 14172
rect 5690 14170 5696 14172
rect 5450 14118 5452 14170
rect 5632 14118 5634 14170
rect 5388 14116 5394 14118
rect 5450 14116 5474 14118
rect 5530 14116 5554 14118
rect 5610 14116 5634 14118
rect 5690 14116 5696 14118
rect 5388 14107 5696 14116
rect 5736 13938 5764 14486
rect 5724 13932 5776 13938
rect 5724 13874 5776 13880
rect 5828 13870 5856 14758
rect 6472 14618 6500 15370
rect 6828 15360 6880 15366
rect 6828 15302 6880 15308
rect 6840 15026 6868 15302
rect 6828 15020 6880 15026
rect 6828 14962 6880 14968
rect 7116 14958 7144 15982
rect 7608 15804 7916 15813
rect 7608 15802 7614 15804
rect 7670 15802 7694 15804
rect 7750 15802 7774 15804
rect 7830 15802 7854 15804
rect 7910 15802 7916 15804
rect 7670 15750 7672 15802
rect 7852 15750 7854 15802
rect 7608 15748 7614 15750
rect 7670 15748 7694 15750
rect 7750 15748 7774 15750
rect 7830 15748 7854 15750
rect 7910 15748 7916 15750
rect 7608 15739 7916 15748
rect 7472 15428 7524 15434
rect 7472 15370 7524 15376
rect 7484 15162 7512 15370
rect 8036 15366 8064 16050
rect 8668 15904 8720 15910
rect 8668 15846 8720 15852
rect 8024 15360 8076 15366
rect 8024 15302 8076 15308
rect 7472 15156 7524 15162
rect 7472 15098 7524 15104
rect 7104 14952 7156 14958
rect 7104 14894 7156 14900
rect 7116 14618 7144 14894
rect 8392 14816 8444 14822
rect 8392 14758 8444 14764
rect 7608 14716 7916 14725
rect 7608 14714 7614 14716
rect 7670 14714 7694 14716
rect 7750 14714 7774 14716
rect 7830 14714 7854 14716
rect 7910 14714 7916 14716
rect 7670 14662 7672 14714
rect 7852 14662 7854 14714
rect 7608 14660 7614 14662
rect 7670 14660 7694 14662
rect 7750 14660 7774 14662
rect 7830 14660 7854 14662
rect 7910 14660 7916 14662
rect 7608 14651 7916 14660
rect 6460 14612 6512 14618
rect 6460 14554 6512 14560
rect 7104 14612 7156 14618
rect 7104 14554 7156 14560
rect 6000 14408 6052 14414
rect 6000 14350 6052 14356
rect 6276 14408 6328 14414
rect 6276 14350 6328 14356
rect 6012 14006 6040 14350
rect 6288 14074 6316 14350
rect 7012 14340 7064 14346
rect 7012 14282 7064 14288
rect 7024 14074 7052 14282
rect 6276 14068 6328 14074
rect 6276 14010 6328 14016
rect 7012 14068 7064 14074
rect 7012 14010 7064 14016
rect 7116 14006 7144 14554
rect 8300 14408 8352 14414
rect 8300 14350 8352 14356
rect 7932 14272 7984 14278
rect 7932 14214 7984 14220
rect 6000 14000 6052 14006
rect 6000 13942 6052 13948
rect 7104 14000 7156 14006
rect 7104 13942 7156 13948
rect 7196 13932 7248 13938
rect 7196 13874 7248 13880
rect 7472 13932 7524 13938
rect 7472 13874 7524 13880
rect 4988 13864 5040 13870
rect 4988 13806 5040 13812
rect 5816 13864 5868 13870
rect 5816 13806 5868 13812
rect 4344 13524 4396 13530
rect 4344 13466 4396 13472
rect 4264 13382 4384 13410
rect 4160 12980 4212 12986
rect 4160 12922 4212 12928
rect 4252 12844 4304 12850
rect 4252 12786 4304 12792
rect 4264 12442 4292 12786
rect 4252 12436 4304 12442
rect 4252 12378 4304 12384
rect 3976 12232 4028 12238
rect 3976 12174 4028 12180
rect 3792 11756 3844 11762
rect 3792 11698 3844 11704
rect 3804 11150 3832 11698
rect 3988 11354 4016 12174
rect 4160 11552 4212 11558
rect 4160 11494 4212 11500
rect 3976 11348 4028 11354
rect 3976 11290 4028 11296
rect 4172 11150 4200 11494
rect 4356 11218 4384 13382
rect 5000 13326 5028 13806
rect 4988 13320 5040 13326
rect 4988 13262 5040 13268
rect 5000 12782 5028 13262
rect 5388 13084 5696 13093
rect 5388 13082 5394 13084
rect 5450 13082 5474 13084
rect 5530 13082 5554 13084
rect 5610 13082 5634 13084
rect 5690 13082 5696 13084
rect 5450 13030 5452 13082
rect 5632 13030 5634 13082
rect 5388 13028 5394 13030
rect 5450 13028 5474 13030
rect 5530 13028 5554 13030
rect 5610 13028 5634 13030
rect 5690 13028 5696 13030
rect 5388 13019 5696 13028
rect 4988 12776 5040 12782
rect 4988 12718 5040 12724
rect 4620 12640 4672 12646
rect 4620 12582 4672 12588
rect 4632 11830 4660 12582
rect 5388 11996 5696 12005
rect 5388 11994 5394 11996
rect 5450 11994 5474 11996
rect 5530 11994 5554 11996
rect 5610 11994 5634 11996
rect 5690 11994 5696 11996
rect 5450 11942 5452 11994
rect 5632 11942 5634 11994
rect 5388 11940 5394 11942
rect 5450 11940 5474 11942
rect 5530 11940 5554 11942
rect 5610 11940 5634 11942
rect 5690 11940 5696 11942
rect 5388 11931 5696 11940
rect 4620 11824 4672 11830
rect 4620 11766 4672 11772
rect 4632 11694 4660 11766
rect 4620 11688 4672 11694
rect 4620 11630 4672 11636
rect 4344 11212 4396 11218
rect 4344 11154 4396 11160
rect 3792 11144 3844 11150
rect 3792 11086 3844 11092
rect 4160 11144 4212 11150
rect 4160 11086 4212 11092
rect 4160 11008 4212 11014
rect 4160 10950 4212 10956
rect 3700 10260 3752 10266
rect 3700 10202 3752 10208
rect 3712 9994 3740 10202
rect 3700 9988 3752 9994
rect 3700 9930 3752 9936
rect 3608 9920 3660 9926
rect 3608 9862 3660 9868
rect 2780 9648 2832 9654
rect 2780 9590 2832 9596
rect 1860 9376 1912 9382
rect 1860 9318 1912 9324
rect 2504 9376 2556 9382
rect 2504 9318 2556 9324
rect 1872 7954 1900 9318
rect 3169 9276 3477 9285
rect 3169 9274 3175 9276
rect 3231 9274 3255 9276
rect 3311 9274 3335 9276
rect 3391 9274 3415 9276
rect 3471 9274 3477 9276
rect 3231 9222 3233 9274
rect 3413 9222 3415 9274
rect 3169 9220 3175 9222
rect 3231 9220 3255 9222
rect 3311 9220 3335 9222
rect 3391 9220 3415 9222
rect 3471 9220 3477 9222
rect 3169 9211 3477 9220
rect 3620 8498 3648 9862
rect 2596 8492 2648 8498
rect 2596 8434 2648 8440
rect 3608 8492 3660 8498
rect 3608 8434 3660 8440
rect 2044 8424 2096 8430
rect 2044 8366 2096 8372
rect 2056 8090 2084 8366
rect 2608 8090 2636 8434
rect 3169 8188 3477 8197
rect 3169 8186 3175 8188
rect 3231 8186 3255 8188
rect 3311 8186 3335 8188
rect 3391 8186 3415 8188
rect 3471 8186 3477 8188
rect 3231 8134 3233 8186
rect 3413 8134 3415 8186
rect 3169 8132 3175 8134
rect 3231 8132 3255 8134
rect 3311 8132 3335 8134
rect 3391 8132 3415 8134
rect 3471 8132 3477 8134
rect 3169 8123 3477 8132
rect 2044 8084 2096 8090
rect 2044 8026 2096 8032
rect 2596 8084 2648 8090
rect 2596 8026 2648 8032
rect 3056 8016 3108 8022
rect 3056 7958 3108 7964
rect 1860 7948 1912 7954
rect 1860 7890 1912 7896
rect 2964 7744 3016 7750
rect 2964 7686 3016 7692
rect 2780 7336 2832 7342
rect 2780 7278 2832 7284
rect 2792 6798 2820 7278
rect 2976 6866 3004 7686
rect 3068 7342 3096 7958
rect 3424 7880 3476 7886
rect 3424 7822 3476 7828
rect 3436 7546 3464 7822
rect 3424 7540 3476 7546
rect 3424 7482 3476 7488
rect 3056 7336 3108 7342
rect 3056 7278 3108 7284
rect 3169 7100 3477 7109
rect 3169 7098 3175 7100
rect 3231 7098 3255 7100
rect 3311 7098 3335 7100
rect 3391 7098 3415 7100
rect 3471 7098 3477 7100
rect 3231 7046 3233 7098
rect 3413 7046 3415 7098
rect 3169 7044 3175 7046
rect 3231 7044 3255 7046
rect 3311 7044 3335 7046
rect 3391 7044 3415 7046
rect 3471 7044 3477 7046
rect 3169 7035 3477 7044
rect 3712 6866 3740 9930
rect 4172 9382 4200 10950
rect 4252 10668 4304 10674
rect 4356 10656 4384 11154
rect 4304 10628 4384 10656
rect 4252 10610 4304 10616
rect 4436 10600 4488 10606
rect 4436 10542 4488 10548
rect 4160 9376 4212 9382
rect 4160 9318 4212 9324
rect 4172 7886 4200 9318
rect 4448 8634 4476 10542
rect 4632 9654 4660 11630
rect 5828 11014 5856 13806
rect 7208 13462 7236 13874
rect 7288 13796 7340 13802
rect 7288 13738 7340 13744
rect 7196 13456 7248 13462
rect 7196 13398 7248 13404
rect 5908 13252 5960 13258
rect 5908 13194 5960 13200
rect 5920 12986 5948 13194
rect 7012 13184 7064 13190
rect 7012 13126 7064 13132
rect 5908 12980 5960 12986
rect 5908 12922 5960 12928
rect 6000 12844 6052 12850
rect 6000 12786 6052 12792
rect 6012 12442 6040 12786
rect 7024 12782 7052 13126
rect 7208 12850 7236 13398
rect 7300 13326 7328 13738
rect 7484 13530 7512 13874
rect 7608 13628 7916 13637
rect 7608 13626 7614 13628
rect 7670 13626 7694 13628
rect 7750 13626 7774 13628
rect 7830 13626 7854 13628
rect 7910 13626 7916 13628
rect 7670 13574 7672 13626
rect 7852 13574 7854 13626
rect 7608 13572 7614 13574
rect 7670 13572 7694 13574
rect 7750 13572 7774 13574
rect 7830 13572 7854 13574
rect 7910 13572 7916 13574
rect 7608 13563 7916 13572
rect 7472 13524 7524 13530
rect 7472 13466 7524 13472
rect 7944 13326 7972 14214
rect 8208 13456 8260 13462
rect 8208 13398 8260 13404
rect 7288 13320 7340 13326
rect 7288 13262 7340 13268
rect 7932 13320 7984 13326
rect 7932 13262 7984 13268
rect 7196 12844 7248 12850
rect 7196 12786 7248 12792
rect 7012 12776 7064 12782
rect 7012 12718 7064 12724
rect 6000 12436 6052 12442
rect 6000 12378 6052 12384
rect 7010 12336 7066 12345
rect 6828 12300 6880 12306
rect 7010 12271 7066 12280
rect 6828 12242 6880 12248
rect 6368 12232 6420 12238
rect 6368 12174 6420 12180
rect 6092 11756 6144 11762
rect 6092 11698 6144 11704
rect 6104 11354 6132 11698
rect 6184 11552 6236 11558
rect 6184 11494 6236 11500
rect 6092 11348 6144 11354
rect 6092 11290 6144 11296
rect 6196 11150 6224 11494
rect 6380 11150 6408 12174
rect 6184 11144 6236 11150
rect 6184 11086 6236 11092
rect 6368 11144 6420 11150
rect 6368 11086 6420 11092
rect 6840 11082 6868 12242
rect 7024 12170 7052 12271
rect 7196 12232 7248 12238
rect 7196 12174 7248 12180
rect 7012 12164 7064 12170
rect 7012 12106 7064 12112
rect 7104 12096 7156 12102
rect 7104 12038 7156 12044
rect 7116 11830 7144 12038
rect 7104 11824 7156 11830
rect 7104 11766 7156 11772
rect 7012 11756 7064 11762
rect 7012 11698 7064 11704
rect 7024 11642 7052 11698
rect 7024 11614 7144 11642
rect 7012 11552 7064 11558
rect 7012 11494 7064 11500
rect 7024 11354 7052 11494
rect 7012 11348 7064 11354
rect 7012 11290 7064 11296
rect 6828 11076 6880 11082
rect 6828 11018 6880 11024
rect 5816 11008 5868 11014
rect 5816 10950 5868 10956
rect 6092 11008 6144 11014
rect 6092 10950 6144 10956
rect 5388 10908 5696 10917
rect 5388 10906 5394 10908
rect 5450 10906 5474 10908
rect 5530 10906 5554 10908
rect 5610 10906 5634 10908
rect 5690 10906 5696 10908
rect 5450 10854 5452 10906
rect 5632 10854 5634 10906
rect 5388 10852 5394 10854
rect 5450 10852 5474 10854
rect 5530 10852 5554 10854
rect 5610 10852 5634 10854
rect 5690 10852 5696 10854
rect 5388 10843 5696 10852
rect 6104 10606 6132 10950
rect 6092 10600 6144 10606
rect 6092 10542 6144 10548
rect 6552 10600 6604 10606
rect 6552 10542 6604 10548
rect 4804 10464 4856 10470
rect 4804 10406 4856 10412
rect 4620 9648 4672 9654
rect 4620 9590 4672 9596
rect 4816 9586 4844 10406
rect 5388 9820 5696 9829
rect 5388 9818 5394 9820
rect 5450 9818 5474 9820
rect 5530 9818 5554 9820
rect 5610 9818 5634 9820
rect 5690 9818 5696 9820
rect 5450 9766 5452 9818
rect 5632 9766 5634 9818
rect 5388 9764 5394 9766
rect 5450 9764 5474 9766
rect 5530 9764 5554 9766
rect 5610 9764 5634 9766
rect 5690 9764 5696 9766
rect 5388 9755 5696 9764
rect 4804 9580 4856 9586
rect 4804 9522 4856 9528
rect 4988 9172 5040 9178
rect 4988 9114 5040 9120
rect 4896 8832 4948 8838
rect 4896 8774 4948 8780
rect 4436 8628 4488 8634
rect 4436 8570 4488 8576
rect 4160 7880 4212 7886
rect 4160 7822 4212 7828
rect 3976 7812 4028 7818
rect 3976 7754 4028 7760
rect 3988 7478 4016 7754
rect 3976 7472 4028 7478
rect 3976 7414 4028 7420
rect 2964 6860 3016 6866
rect 2964 6802 3016 6808
rect 3700 6860 3752 6866
rect 3700 6802 3752 6808
rect 2228 6792 2280 6798
rect 2228 6734 2280 6740
rect 2780 6792 2832 6798
rect 2780 6734 2832 6740
rect 2240 6186 2268 6734
rect 2976 6458 3004 6802
rect 3056 6792 3108 6798
rect 3056 6734 3108 6740
rect 3240 6792 3292 6798
rect 3240 6734 3292 6740
rect 2964 6452 3016 6458
rect 2964 6394 3016 6400
rect 3068 6322 3096 6734
rect 3056 6316 3108 6322
rect 2976 6276 3056 6304
rect 2872 6248 2924 6254
rect 2872 6190 2924 6196
rect 2228 6180 2280 6186
rect 2228 6122 2280 6128
rect 2884 5642 2912 6190
rect 2976 5710 3004 6276
rect 3056 6258 3108 6264
rect 3252 6254 3280 6734
rect 3712 6662 3740 6802
rect 3700 6656 3752 6662
rect 3700 6598 3752 6604
rect 3240 6248 3292 6254
rect 3240 6190 3292 6196
rect 3169 6012 3477 6021
rect 3169 6010 3175 6012
rect 3231 6010 3255 6012
rect 3311 6010 3335 6012
rect 3391 6010 3415 6012
rect 3471 6010 3477 6012
rect 3231 5958 3233 6010
rect 3413 5958 3415 6010
rect 3169 5956 3175 5958
rect 3231 5956 3255 5958
rect 3311 5956 3335 5958
rect 3391 5956 3415 5958
rect 3471 5956 3477 5958
rect 3169 5947 3477 5956
rect 3712 5914 3740 6598
rect 3988 6322 4016 7414
rect 4172 7342 4200 7822
rect 4448 7410 4476 8570
rect 4620 8560 4672 8566
rect 4620 8502 4672 8508
rect 4436 7404 4488 7410
rect 4436 7346 4488 7352
rect 4160 7336 4212 7342
rect 4160 7278 4212 7284
rect 4632 6798 4660 8502
rect 4908 7886 4936 8774
rect 5000 8430 5028 9114
rect 5908 9104 5960 9110
rect 5908 9046 5960 9052
rect 5080 8968 5132 8974
rect 5080 8910 5132 8916
rect 5724 8968 5776 8974
rect 5724 8910 5776 8916
rect 5092 8498 5120 8910
rect 5388 8732 5696 8741
rect 5388 8730 5394 8732
rect 5450 8730 5474 8732
rect 5530 8730 5554 8732
rect 5610 8730 5634 8732
rect 5690 8730 5696 8732
rect 5450 8678 5452 8730
rect 5632 8678 5634 8730
rect 5388 8676 5394 8678
rect 5450 8676 5474 8678
rect 5530 8676 5554 8678
rect 5610 8676 5634 8678
rect 5690 8676 5696 8678
rect 5388 8667 5696 8676
rect 5080 8492 5132 8498
rect 5080 8434 5132 8440
rect 4988 8424 5040 8430
rect 4988 8366 5040 8372
rect 5000 8022 5028 8366
rect 4988 8016 5040 8022
rect 4988 7958 5040 7964
rect 5092 7954 5120 8434
rect 5080 7948 5132 7954
rect 5080 7890 5132 7896
rect 5736 7886 5764 8910
rect 5816 8832 5868 8838
rect 5816 8774 5868 8780
rect 5828 8362 5856 8774
rect 5816 8356 5868 8362
rect 5816 8298 5868 8304
rect 4896 7880 4948 7886
rect 4896 7822 4948 7828
rect 5724 7880 5776 7886
rect 5724 7822 5776 7828
rect 4908 7546 4936 7822
rect 5388 7644 5696 7653
rect 5388 7642 5394 7644
rect 5450 7642 5474 7644
rect 5530 7642 5554 7644
rect 5610 7642 5634 7644
rect 5690 7642 5696 7644
rect 5450 7590 5452 7642
rect 5632 7590 5634 7642
rect 5388 7588 5394 7590
rect 5450 7588 5474 7590
rect 5530 7588 5554 7590
rect 5610 7588 5634 7590
rect 5690 7588 5696 7590
rect 5388 7579 5696 7588
rect 4896 7540 4948 7546
rect 4896 7482 4948 7488
rect 5080 7472 5132 7478
rect 5080 7414 5132 7420
rect 4620 6792 4672 6798
rect 4620 6734 4672 6740
rect 4632 6322 4660 6734
rect 5092 6390 5120 7414
rect 5920 7410 5948 9046
rect 6000 8424 6052 8430
rect 6000 8366 6052 8372
rect 6012 7886 6040 8366
rect 6000 7880 6052 7886
rect 6000 7822 6052 7828
rect 6012 7410 6040 7822
rect 5908 7404 5960 7410
rect 5908 7346 5960 7352
rect 6000 7404 6052 7410
rect 6000 7346 6052 7352
rect 6104 6730 6132 10542
rect 6564 10266 6592 10542
rect 6552 10260 6604 10266
rect 6552 10202 6604 10208
rect 6564 9654 6592 10202
rect 7012 10056 7064 10062
rect 7012 9998 7064 10004
rect 6552 9648 6604 9654
rect 6552 9590 6604 9596
rect 6736 9580 6788 9586
rect 6736 9522 6788 9528
rect 6368 8900 6420 8906
rect 6368 8842 6420 8848
rect 6552 8900 6604 8906
rect 6552 8842 6604 8848
rect 6380 8566 6408 8842
rect 6564 8634 6592 8842
rect 6552 8628 6604 8634
rect 6552 8570 6604 8576
rect 6368 8560 6420 8566
rect 6368 8502 6420 8508
rect 6748 8480 6776 9522
rect 6828 9104 6880 9110
rect 6828 9046 6880 9052
rect 6840 8634 6868 9046
rect 6828 8628 6880 8634
rect 6828 8570 6880 8576
rect 6748 8452 6868 8480
rect 6736 8356 6788 8362
rect 6736 8298 6788 8304
rect 6748 7886 6776 8298
rect 6840 7886 6868 8452
rect 6920 8356 6972 8362
rect 6920 8298 6972 8304
rect 6932 8090 6960 8298
rect 6920 8084 6972 8090
rect 6920 8026 6972 8032
rect 6736 7880 6788 7886
rect 6736 7822 6788 7828
rect 6828 7880 6880 7886
rect 6828 7822 6880 7828
rect 6736 7744 6788 7750
rect 6736 7686 6788 7692
rect 6748 7478 6776 7686
rect 6840 7546 6868 7822
rect 6920 7744 6972 7750
rect 6920 7686 6972 7692
rect 6828 7540 6880 7546
rect 6828 7482 6880 7488
rect 6932 7478 6960 7686
rect 6736 7472 6788 7478
rect 6736 7414 6788 7420
rect 6920 7472 6972 7478
rect 6920 7414 6972 7420
rect 6552 7336 6604 7342
rect 6552 7278 6604 7284
rect 6564 6798 6592 7278
rect 6552 6792 6604 6798
rect 6552 6734 6604 6740
rect 6092 6724 6144 6730
rect 6092 6666 6144 6672
rect 5388 6556 5696 6565
rect 5388 6554 5394 6556
rect 5450 6554 5474 6556
rect 5530 6554 5554 6556
rect 5610 6554 5634 6556
rect 5690 6554 5696 6556
rect 5450 6502 5452 6554
rect 5632 6502 5634 6554
rect 5388 6500 5394 6502
rect 5450 6500 5474 6502
rect 5530 6500 5554 6502
rect 5610 6500 5634 6502
rect 5690 6500 5696 6502
rect 5388 6491 5696 6500
rect 5080 6384 5132 6390
rect 5080 6326 5132 6332
rect 3976 6316 4028 6322
rect 3976 6258 4028 6264
rect 4620 6316 4672 6322
rect 4620 6258 4672 6264
rect 3700 5908 3752 5914
rect 3700 5850 3752 5856
rect 3056 5840 3108 5846
rect 3056 5782 3108 5788
rect 2964 5704 3016 5710
rect 2964 5646 3016 5652
rect 2872 5636 2924 5642
rect 2872 5578 2924 5584
rect 2884 4690 2912 5578
rect 2976 5370 3004 5646
rect 2964 5364 3016 5370
rect 2964 5306 3016 5312
rect 2976 4826 3004 5306
rect 2964 4820 3016 4826
rect 2964 4762 3016 4768
rect 2872 4684 2924 4690
rect 2872 4626 2924 4632
rect 3068 4622 3096 5782
rect 3988 5370 4016 6258
rect 4160 6112 4212 6118
rect 4160 6054 4212 6060
rect 4068 5908 4120 5914
rect 4068 5850 4120 5856
rect 4080 5778 4108 5850
rect 4068 5772 4120 5778
rect 4068 5714 4120 5720
rect 3976 5364 4028 5370
rect 3976 5306 4028 5312
rect 4172 5234 4200 6054
rect 4632 5778 4660 6258
rect 4620 5772 4672 5778
rect 4620 5714 4672 5720
rect 4632 5302 4660 5714
rect 4620 5296 4672 5302
rect 4620 5238 4672 5244
rect 3516 5228 3568 5234
rect 3516 5170 3568 5176
rect 4160 5228 4212 5234
rect 4160 5170 4212 5176
rect 3169 4924 3477 4933
rect 3169 4922 3175 4924
rect 3231 4922 3255 4924
rect 3311 4922 3335 4924
rect 3391 4922 3415 4924
rect 3471 4922 3477 4924
rect 3231 4870 3233 4922
rect 3413 4870 3415 4922
rect 3169 4868 3175 4870
rect 3231 4868 3255 4870
rect 3311 4868 3335 4870
rect 3391 4868 3415 4870
rect 3471 4868 3477 4870
rect 3169 4859 3477 4868
rect 3528 4826 3556 5170
rect 3516 4820 3568 4826
rect 3516 4762 3568 4768
rect 4632 4690 4660 5238
rect 5092 4826 5120 6326
rect 5172 6316 5224 6322
rect 5172 6258 5224 6264
rect 5184 6066 5212 6258
rect 5264 6112 5316 6118
rect 5184 6060 5264 6066
rect 5184 6054 5316 6060
rect 5184 6038 5304 6054
rect 5080 4820 5132 4826
rect 5080 4762 5132 4768
rect 4620 4684 4672 4690
rect 4620 4626 4672 4632
rect 3056 4616 3108 4622
rect 3056 4558 3108 4564
rect 5184 4282 5212 6038
rect 6104 5914 6132 6666
rect 6092 5908 6144 5914
rect 6092 5850 6144 5856
rect 5908 5840 5960 5846
rect 5908 5782 5960 5788
rect 5388 5468 5696 5477
rect 5388 5466 5394 5468
rect 5450 5466 5474 5468
rect 5530 5466 5554 5468
rect 5610 5466 5634 5468
rect 5690 5466 5696 5468
rect 5450 5414 5452 5466
rect 5632 5414 5634 5466
rect 5388 5412 5394 5414
rect 5450 5412 5474 5414
rect 5530 5412 5554 5414
rect 5610 5412 5634 5414
rect 5690 5412 5696 5414
rect 5388 5403 5696 5412
rect 5920 5370 5948 5782
rect 6368 5704 6420 5710
rect 6368 5646 6420 5652
rect 6184 5568 6236 5574
rect 6184 5510 6236 5516
rect 5908 5364 5960 5370
rect 5908 5306 5960 5312
rect 5264 4684 5316 4690
rect 5264 4626 5316 4632
rect 5172 4276 5224 4282
rect 5172 4218 5224 4224
rect 4712 3936 4764 3942
rect 4712 3878 4764 3884
rect 3169 3836 3477 3845
rect 3169 3834 3175 3836
rect 3231 3834 3255 3836
rect 3311 3834 3335 3836
rect 3391 3834 3415 3836
rect 3471 3834 3477 3836
rect 3231 3782 3233 3834
rect 3413 3782 3415 3834
rect 3169 3780 3175 3782
rect 3231 3780 3255 3782
rect 3311 3780 3335 3782
rect 3391 3780 3415 3782
rect 3471 3780 3477 3782
rect 3169 3771 3477 3780
rect 3976 3392 4028 3398
rect 3976 3334 4028 3340
rect 3169 2748 3477 2757
rect 3169 2746 3175 2748
rect 3231 2746 3255 2748
rect 3311 2746 3335 2748
rect 3391 2746 3415 2748
rect 3471 2746 3477 2748
rect 3231 2694 3233 2746
rect 3413 2694 3415 2746
rect 3169 2692 3175 2694
rect 3231 2692 3255 2694
rect 3311 2692 3335 2694
rect 3391 2692 3415 2694
rect 3471 2692 3477 2694
rect 3169 2683 3477 2692
rect 3988 2446 4016 3334
rect 4724 3058 4752 3878
rect 5276 3534 5304 4626
rect 5920 4622 5948 5306
rect 5908 4616 5960 4622
rect 5908 4558 5960 4564
rect 5388 4380 5696 4389
rect 5388 4378 5394 4380
rect 5450 4378 5474 4380
rect 5530 4378 5554 4380
rect 5610 4378 5634 4380
rect 5690 4378 5696 4380
rect 5450 4326 5452 4378
rect 5632 4326 5634 4378
rect 5388 4324 5394 4326
rect 5450 4324 5474 4326
rect 5530 4324 5554 4326
rect 5610 4324 5634 4326
rect 5690 4324 5696 4326
rect 5388 4315 5696 4324
rect 6196 3534 6224 5510
rect 6380 5030 6408 5646
rect 6564 5642 6592 6734
rect 6736 6316 6788 6322
rect 6736 6258 6788 6264
rect 6552 5636 6604 5642
rect 6552 5578 6604 5584
rect 6368 5024 6420 5030
rect 6368 4966 6420 4972
rect 6380 4622 6408 4966
rect 6368 4616 6420 4622
rect 6368 4558 6420 4564
rect 6564 4078 6592 5578
rect 6748 4826 6776 6258
rect 6920 6180 6972 6186
rect 6920 6122 6972 6128
rect 6932 5370 6960 6122
rect 7024 5710 7052 9998
rect 7116 8922 7144 11614
rect 7208 11354 7236 12174
rect 7300 12102 7328 13262
rect 8220 12714 8248 13398
rect 8312 12986 8340 14350
rect 8404 13734 8432 14758
rect 8392 13728 8444 13734
rect 8392 13670 8444 13676
rect 8404 13326 8432 13670
rect 8392 13320 8444 13326
rect 8392 13262 8444 13268
rect 8300 12980 8352 12986
rect 8300 12922 8352 12928
rect 8208 12708 8260 12714
rect 8208 12650 8260 12656
rect 7380 12640 7432 12646
rect 7380 12582 7432 12588
rect 7392 12238 7420 12582
rect 7608 12540 7916 12549
rect 7608 12538 7614 12540
rect 7670 12538 7694 12540
rect 7750 12538 7774 12540
rect 7830 12538 7854 12540
rect 7910 12538 7916 12540
rect 7670 12486 7672 12538
rect 7852 12486 7854 12538
rect 7608 12484 7614 12486
rect 7670 12484 7694 12486
rect 7750 12484 7774 12486
rect 7830 12484 7854 12486
rect 7910 12484 7916 12486
rect 7608 12475 7916 12484
rect 8208 12368 8260 12374
rect 8208 12310 8260 12316
rect 7380 12232 7432 12238
rect 7380 12174 7432 12180
rect 7932 12232 7984 12238
rect 7932 12174 7984 12180
rect 8116 12232 8168 12238
rect 8116 12174 8168 12180
rect 7288 12096 7340 12102
rect 7288 12038 7340 12044
rect 7944 11898 7972 12174
rect 8024 12096 8076 12102
rect 8024 12038 8076 12044
rect 7932 11892 7984 11898
rect 7932 11834 7984 11840
rect 7288 11824 7340 11830
rect 7288 11766 7340 11772
rect 7196 11348 7248 11354
rect 7196 11290 7248 11296
rect 7300 11150 7328 11766
rect 7608 11452 7916 11461
rect 7608 11450 7614 11452
rect 7670 11450 7694 11452
rect 7750 11450 7774 11452
rect 7830 11450 7854 11452
rect 7910 11450 7916 11452
rect 7670 11398 7672 11450
rect 7852 11398 7854 11450
rect 7608 11396 7614 11398
rect 7670 11396 7694 11398
rect 7750 11396 7774 11398
rect 7830 11396 7854 11398
rect 7910 11396 7916 11398
rect 7608 11387 7916 11396
rect 7288 11144 7340 11150
rect 7288 11086 7340 11092
rect 7300 10198 7328 11086
rect 8036 10742 8064 12038
rect 8128 11694 8156 12174
rect 8220 11762 8248 12310
rect 8392 12232 8444 12238
rect 8392 12174 8444 12180
rect 8404 12102 8432 12174
rect 8392 12096 8444 12102
rect 8392 12038 8444 12044
rect 8208 11756 8260 11762
rect 8208 11698 8260 11704
rect 8576 11756 8628 11762
rect 8576 11698 8628 11704
rect 8116 11688 8168 11694
rect 8116 11630 8168 11636
rect 8220 11286 8248 11698
rect 8588 11558 8616 11698
rect 8576 11552 8628 11558
rect 8576 11494 8628 11500
rect 8208 11280 8260 11286
rect 8128 11228 8208 11234
rect 8128 11222 8260 11228
rect 8128 11206 8248 11222
rect 8024 10736 8076 10742
rect 8024 10678 8076 10684
rect 7380 10668 7432 10674
rect 7380 10610 7432 10616
rect 7392 10266 7420 10610
rect 7472 10464 7524 10470
rect 7472 10406 7524 10412
rect 7932 10464 7984 10470
rect 7932 10406 7984 10412
rect 7380 10260 7432 10266
rect 7380 10202 7432 10208
rect 7288 10192 7340 10198
rect 7288 10134 7340 10140
rect 7116 8894 7236 8922
rect 7104 8832 7156 8838
rect 7104 8774 7156 8780
rect 7012 5704 7064 5710
rect 7012 5646 7064 5652
rect 6920 5364 6972 5370
rect 6920 5306 6972 5312
rect 7024 5302 7052 5646
rect 7012 5296 7064 5302
rect 7012 5238 7064 5244
rect 7116 5234 7144 8774
rect 7208 6458 7236 8894
rect 7300 7410 7328 10134
rect 7484 10062 7512 10406
rect 7608 10364 7916 10373
rect 7608 10362 7614 10364
rect 7670 10362 7694 10364
rect 7750 10362 7774 10364
rect 7830 10362 7854 10364
rect 7910 10362 7916 10364
rect 7670 10310 7672 10362
rect 7852 10310 7854 10362
rect 7608 10308 7614 10310
rect 7670 10308 7694 10310
rect 7750 10308 7774 10310
rect 7830 10308 7854 10310
rect 7910 10308 7916 10310
rect 7608 10299 7916 10308
rect 7472 10056 7524 10062
rect 7472 9998 7524 10004
rect 7472 9580 7524 9586
rect 7472 9522 7524 9528
rect 7484 7546 7512 9522
rect 7608 9276 7916 9285
rect 7608 9274 7614 9276
rect 7670 9274 7694 9276
rect 7750 9274 7774 9276
rect 7830 9274 7854 9276
rect 7910 9274 7916 9276
rect 7670 9222 7672 9274
rect 7852 9222 7854 9274
rect 7608 9220 7614 9222
rect 7670 9220 7694 9222
rect 7750 9220 7774 9222
rect 7830 9220 7854 9222
rect 7910 9220 7916 9222
rect 7608 9211 7916 9220
rect 7608 8188 7916 8197
rect 7608 8186 7614 8188
rect 7670 8186 7694 8188
rect 7750 8186 7774 8188
rect 7830 8186 7854 8188
rect 7910 8186 7916 8188
rect 7670 8134 7672 8186
rect 7852 8134 7854 8186
rect 7608 8132 7614 8134
rect 7670 8132 7694 8134
rect 7750 8132 7774 8134
rect 7830 8132 7854 8134
rect 7910 8132 7916 8134
rect 7608 8123 7916 8132
rect 7564 7744 7616 7750
rect 7564 7686 7616 7692
rect 7576 7546 7604 7686
rect 7472 7540 7524 7546
rect 7472 7482 7524 7488
rect 7564 7540 7616 7546
rect 7564 7482 7616 7488
rect 7288 7404 7340 7410
rect 7288 7346 7340 7352
rect 7944 7206 7972 10406
rect 8036 9110 8064 10678
rect 8128 10062 8156 11206
rect 8208 11076 8260 11082
rect 8208 11018 8260 11024
rect 8300 11076 8352 11082
rect 8300 11018 8352 11024
rect 8220 10674 8248 11018
rect 8208 10668 8260 10674
rect 8208 10610 8260 10616
rect 8116 10056 8168 10062
rect 8168 10016 8248 10044
rect 8116 9998 8168 10004
rect 8116 9376 8168 9382
rect 8116 9318 8168 9324
rect 8024 9104 8076 9110
rect 8024 9046 8076 9052
rect 8128 8498 8156 9318
rect 8220 9178 8248 10016
rect 8208 9172 8260 9178
rect 8208 9114 8260 9120
rect 8312 8974 8340 11018
rect 8484 11008 8536 11014
rect 8484 10950 8536 10956
rect 8496 10742 8524 10950
rect 8484 10736 8536 10742
rect 8484 10678 8536 10684
rect 8496 10538 8524 10678
rect 8588 10674 8616 11494
rect 8576 10668 8628 10674
rect 8576 10610 8628 10616
rect 8484 10532 8536 10538
rect 8484 10474 8536 10480
rect 8300 8968 8352 8974
rect 8300 8910 8352 8916
rect 8496 8566 8524 10474
rect 8588 9994 8616 10610
rect 8680 10266 8708 15846
rect 9140 15502 9168 16118
rect 9128 15496 9180 15502
rect 9128 15438 9180 15444
rect 9140 14958 9168 15438
rect 9680 15360 9732 15366
rect 9680 15302 9732 15308
rect 9692 15162 9720 15302
rect 9827 15260 10135 15269
rect 9827 15258 9833 15260
rect 9889 15258 9913 15260
rect 9969 15258 9993 15260
rect 10049 15258 10073 15260
rect 10129 15258 10135 15260
rect 9889 15206 9891 15258
rect 10071 15206 10073 15258
rect 9827 15204 9833 15206
rect 9889 15204 9913 15206
rect 9969 15204 9993 15206
rect 10049 15204 10073 15206
rect 10129 15204 10135 15206
rect 9827 15195 10135 15204
rect 9680 15156 9732 15162
rect 9680 15098 9732 15104
rect 9680 15020 9732 15026
rect 9680 14962 9732 14968
rect 10232 15020 10284 15026
rect 10232 14962 10284 14968
rect 9128 14952 9180 14958
rect 9128 14894 9180 14900
rect 9140 14414 9168 14894
rect 9128 14408 9180 14414
rect 9128 14350 9180 14356
rect 9220 14340 9272 14346
rect 9220 14282 9272 14288
rect 9232 14074 9260 14282
rect 9692 14074 9720 14962
rect 9827 14172 10135 14181
rect 9827 14170 9833 14172
rect 9889 14170 9913 14172
rect 9969 14170 9993 14172
rect 10049 14170 10073 14172
rect 10129 14170 10135 14172
rect 9889 14118 9891 14170
rect 10071 14118 10073 14170
rect 9827 14116 9833 14118
rect 9889 14116 9913 14118
rect 9969 14116 9993 14118
rect 10049 14116 10073 14118
rect 10129 14116 10135 14118
rect 9827 14107 10135 14116
rect 9220 14068 9272 14074
rect 9220 14010 9272 14016
rect 9680 14068 9732 14074
rect 9680 14010 9732 14016
rect 9312 14000 9364 14006
rect 9312 13942 9364 13948
rect 8760 13932 8812 13938
rect 8760 13874 8812 13880
rect 9036 13932 9088 13938
rect 9036 13874 9088 13880
rect 8772 11898 8800 13874
rect 8944 13252 8996 13258
rect 8944 13194 8996 13200
rect 8760 11892 8812 11898
rect 8760 11834 8812 11840
rect 8956 11558 8984 13194
rect 9048 12442 9076 13874
rect 9036 12436 9088 12442
rect 9324 12434 9352 13942
rect 9956 13864 10008 13870
rect 9956 13806 10008 13812
rect 9588 13728 9640 13734
rect 9588 13670 9640 13676
rect 9600 13462 9628 13670
rect 9588 13456 9640 13462
rect 9588 13398 9640 13404
rect 9404 13320 9456 13326
rect 9404 13262 9456 13268
rect 9036 12378 9088 12384
rect 9232 12406 9352 12434
rect 9232 12345 9260 12406
rect 9218 12336 9274 12345
rect 9140 12294 9218 12322
rect 8944 11552 8996 11558
rect 8944 11494 8996 11500
rect 8956 11218 8984 11494
rect 8944 11212 8996 11218
rect 8944 11154 8996 11160
rect 9140 10554 9168 12294
rect 9218 12271 9274 12280
rect 9312 12300 9364 12306
rect 9312 12242 9364 12248
rect 9220 12232 9272 12238
rect 9220 12174 9272 12180
rect 9232 11898 9260 12174
rect 9220 11892 9272 11898
rect 9220 11834 9272 11840
rect 9324 11762 9352 12242
rect 9220 11756 9272 11762
rect 9220 11698 9272 11704
rect 9312 11756 9364 11762
rect 9312 11698 9364 11704
rect 9232 10742 9260 11698
rect 9416 11626 9444 13262
rect 9496 12912 9548 12918
rect 9496 12854 9548 12860
rect 9508 12442 9536 12854
rect 9496 12436 9548 12442
rect 9496 12378 9548 12384
rect 9404 11620 9456 11626
rect 9404 11562 9456 11568
rect 9416 11150 9444 11562
rect 9404 11144 9456 11150
rect 9404 11086 9456 11092
rect 9312 11008 9364 11014
rect 9312 10950 9364 10956
rect 9324 10810 9352 10950
rect 9312 10804 9364 10810
rect 9312 10746 9364 10752
rect 9220 10736 9272 10742
rect 9220 10678 9272 10684
rect 9048 10526 9168 10554
rect 8668 10260 8720 10266
rect 8668 10202 8720 10208
rect 8680 10062 8708 10202
rect 8668 10056 8720 10062
rect 8668 9998 8720 10004
rect 8576 9988 8628 9994
rect 8576 9930 8628 9936
rect 8484 8560 8536 8566
rect 8484 8502 8536 8508
rect 9048 8498 9076 10526
rect 9128 10464 9180 10470
rect 9128 10406 9180 10412
rect 9140 8974 9168 10406
rect 9232 9654 9260 10678
rect 9312 10668 9364 10674
rect 9312 10610 9364 10616
rect 9496 10668 9548 10674
rect 9496 10610 9548 10616
rect 9220 9648 9272 9654
rect 9220 9590 9272 9596
rect 9324 8974 9352 10610
rect 9508 9994 9536 10610
rect 9496 9988 9548 9994
rect 9496 9930 9548 9936
rect 9128 8968 9180 8974
rect 9128 8910 9180 8916
rect 9312 8968 9364 8974
rect 9312 8910 9364 8916
rect 9220 8560 9272 8566
rect 9220 8502 9272 8508
rect 8116 8492 8168 8498
rect 8116 8434 8168 8440
rect 9036 8492 9088 8498
rect 9036 8434 9088 8440
rect 8576 8356 8628 8362
rect 8576 8298 8628 8304
rect 8300 8016 8352 8022
rect 8300 7958 8352 7964
rect 8024 7336 8076 7342
rect 8024 7278 8076 7284
rect 7932 7200 7984 7206
rect 7932 7142 7984 7148
rect 7608 7100 7916 7109
rect 7608 7098 7614 7100
rect 7670 7098 7694 7100
rect 7750 7098 7774 7100
rect 7830 7098 7854 7100
rect 7910 7098 7916 7100
rect 7670 7046 7672 7098
rect 7852 7046 7854 7098
rect 7608 7044 7614 7046
rect 7670 7044 7694 7046
rect 7750 7044 7774 7046
rect 7830 7044 7854 7046
rect 7910 7044 7916 7046
rect 7608 7035 7916 7044
rect 7656 6656 7708 6662
rect 7656 6598 7708 6604
rect 7196 6452 7248 6458
rect 7196 6394 7248 6400
rect 7668 6322 7696 6598
rect 8036 6390 8064 7278
rect 8116 7200 8168 7206
rect 8116 7142 8168 7148
rect 8024 6384 8076 6390
rect 8024 6326 8076 6332
rect 7656 6316 7708 6322
rect 7656 6258 7708 6264
rect 7608 6012 7916 6021
rect 7608 6010 7614 6012
rect 7670 6010 7694 6012
rect 7750 6010 7774 6012
rect 7830 6010 7854 6012
rect 7910 6010 7916 6012
rect 7670 5958 7672 6010
rect 7852 5958 7854 6010
rect 7608 5956 7614 5958
rect 7670 5956 7694 5958
rect 7750 5956 7774 5958
rect 7830 5956 7854 5958
rect 7910 5956 7916 5958
rect 7608 5947 7916 5956
rect 7932 5840 7984 5846
rect 7932 5782 7984 5788
rect 7288 5772 7340 5778
rect 7288 5714 7340 5720
rect 7104 5228 7156 5234
rect 7104 5170 7156 5176
rect 7104 5024 7156 5030
rect 7104 4966 7156 4972
rect 6736 4820 6788 4826
rect 6736 4762 6788 4768
rect 6552 4072 6604 4078
rect 6552 4014 6604 4020
rect 6564 3670 6592 4014
rect 6736 4004 6788 4010
rect 6736 3946 6788 3952
rect 6552 3664 6604 3670
rect 6552 3606 6604 3612
rect 5264 3528 5316 3534
rect 5264 3470 5316 3476
rect 6184 3528 6236 3534
rect 6184 3470 6236 3476
rect 6460 3528 6512 3534
rect 6460 3470 6512 3476
rect 5276 3126 5304 3470
rect 5388 3292 5696 3301
rect 5388 3290 5394 3292
rect 5450 3290 5474 3292
rect 5530 3290 5554 3292
rect 5610 3290 5634 3292
rect 5690 3290 5696 3292
rect 5450 3238 5452 3290
rect 5632 3238 5634 3290
rect 5388 3236 5394 3238
rect 5450 3236 5474 3238
rect 5530 3236 5554 3238
rect 5610 3236 5634 3238
rect 5690 3236 5696 3238
rect 5388 3227 5696 3236
rect 5264 3120 5316 3126
rect 5264 3062 5316 3068
rect 4528 3052 4580 3058
rect 4528 2994 4580 3000
rect 4712 3052 4764 3058
rect 4712 2994 4764 3000
rect 4252 2848 4304 2854
rect 4252 2790 4304 2796
rect 4264 2446 4292 2790
rect 4540 2650 4568 2994
rect 6196 2854 6224 3470
rect 6368 3460 6420 3466
rect 6368 3402 6420 3408
rect 6380 3194 6408 3402
rect 6368 3188 6420 3194
rect 6368 3130 6420 3136
rect 6000 2848 6052 2854
rect 6000 2790 6052 2796
rect 6184 2848 6236 2854
rect 6184 2790 6236 2796
rect 4528 2644 4580 2650
rect 4528 2586 4580 2592
rect 6012 2446 6040 2790
rect 6472 2582 6500 3470
rect 6564 2990 6592 3606
rect 6552 2984 6604 2990
rect 6552 2926 6604 2932
rect 6460 2576 6512 2582
rect 6460 2518 6512 2524
rect 6564 2446 6592 2926
rect 6748 2446 6776 3946
rect 7012 3936 7064 3942
rect 7012 3878 7064 3884
rect 7024 3602 7052 3878
rect 7012 3596 7064 3602
rect 7012 3538 7064 3544
rect 6828 3528 6880 3534
rect 6828 3470 6880 3476
rect 6840 2774 6868 3470
rect 6920 3392 6972 3398
rect 6920 3334 6972 3340
rect 6932 3126 6960 3334
rect 6920 3120 6972 3126
rect 6920 3062 6972 3068
rect 7024 3058 7052 3538
rect 7116 3466 7144 4966
rect 7196 4684 7248 4690
rect 7196 4626 7248 4632
rect 7104 3460 7156 3466
rect 7104 3402 7156 3408
rect 7116 3194 7144 3402
rect 7104 3188 7156 3194
rect 7104 3130 7156 3136
rect 7208 3058 7236 4626
rect 7300 4622 7328 5714
rect 7472 5568 7524 5574
rect 7472 5510 7524 5516
rect 7288 4616 7340 4622
rect 7288 4558 7340 4564
rect 7380 4140 7432 4146
rect 7380 4082 7432 4088
rect 7392 4010 7420 4082
rect 7380 4004 7432 4010
rect 7380 3946 7432 3952
rect 7288 3936 7340 3942
rect 7288 3878 7340 3884
rect 7300 3670 7328 3878
rect 7392 3670 7420 3946
rect 7288 3664 7340 3670
rect 7288 3606 7340 3612
rect 7380 3664 7432 3670
rect 7380 3606 7432 3612
rect 7484 3534 7512 5510
rect 7608 4924 7916 4933
rect 7608 4922 7614 4924
rect 7670 4922 7694 4924
rect 7750 4922 7774 4924
rect 7830 4922 7854 4924
rect 7910 4922 7916 4924
rect 7670 4870 7672 4922
rect 7852 4870 7854 4922
rect 7608 4868 7614 4870
rect 7670 4868 7694 4870
rect 7750 4868 7774 4870
rect 7830 4868 7854 4870
rect 7910 4868 7916 4870
rect 7608 4859 7916 4868
rect 7944 4622 7972 5782
rect 8128 5778 8156 7142
rect 8312 6730 8340 7958
rect 8484 7880 8536 7886
rect 8484 7822 8536 7828
rect 8392 7812 8444 7818
rect 8392 7754 8444 7760
rect 8404 7002 8432 7754
rect 8496 7342 8524 7822
rect 8484 7336 8536 7342
rect 8484 7278 8536 7284
rect 8392 6996 8444 7002
rect 8392 6938 8444 6944
rect 8300 6724 8352 6730
rect 8300 6666 8352 6672
rect 8208 6316 8260 6322
rect 8312 6304 8340 6666
rect 8404 6390 8432 6938
rect 8392 6384 8444 6390
rect 8392 6326 8444 6332
rect 8260 6276 8340 6304
rect 8208 6258 8260 6264
rect 8484 6112 8536 6118
rect 8484 6054 8536 6060
rect 8116 5772 8168 5778
rect 8116 5714 8168 5720
rect 8496 5710 8524 6054
rect 8588 5710 8616 8298
rect 8760 7744 8812 7750
rect 8760 7686 8812 7692
rect 8668 7200 8720 7206
rect 8668 7142 8720 7148
rect 8680 6662 8708 7142
rect 8772 6730 8800 7686
rect 9048 7274 9076 8434
rect 9232 7954 9260 8502
rect 9324 8090 9352 8910
rect 9404 8356 9456 8362
rect 9404 8298 9456 8304
rect 9312 8084 9364 8090
rect 9312 8026 9364 8032
rect 9220 7948 9272 7954
rect 9220 7890 9272 7896
rect 9416 7886 9444 8298
rect 9404 7880 9456 7886
rect 9404 7822 9456 7828
rect 9508 7818 9536 9930
rect 9600 9654 9628 13398
rect 9968 13258 9996 13806
rect 10244 13530 10272 14962
rect 10336 14006 10364 16730
rect 10520 16114 10548 16934
rect 10612 16454 10640 16934
rect 12047 16892 12355 16901
rect 12047 16890 12053 16892
rect 12109 16890 12133 16892
rect 12189 16890 12213 16892
rect 12269 16890 12293 16892
rect 12349 16890 12355 16892
rect 12109 16838 12111 16890
rect 12291 16838 12293 16890
rect 12047 16836 12053 16838
rect 12109 16836 12133 16838
rect 12189 16836 12213 16838
rect 12269 16836 12293 16838
rect 12349 16836 12355 16838
rect 12047 16827 12355 16836
rect 12636 16794 12664 17138
rect 16948 17128 17000 17134
rect 16948 17070 17000 17076
rect 12808 16992 12860 16998
rect 12808 16934 12860 16940
rect 12624 16788 12676 16794
rect 12624 16730 12676 16736
rect 12820 16522 12848 16934
rect 16486 16892 16794 16901
rect 16486 16890 16492 16892
rect 16548 16890 16572 16892
rect 16628 16890 16652 16892
rect 16708 16890 16732 16892
rect 16788 16890 16794 16892
rect 16548 16838 16550 16890
rect 16730 16838 16732 16890
rect 16486 16836 16492 16838
rect 16548 16836 16572 16838
rect 16628 16836 16652 16838
rect 16708 16836 16732 16838
rect 16788 16836 16794 16838
rect 16486 16827 16794 16836
rect 10692 16516 10744 16522
rect 10692 16458 10744 16464
rect 12808 16516 12860 16522
rect 12808 16458 12860 16464
rect 10600 16448 10652 16454
rect 10600 16390 10652 16396
rect 10704 16250 10732 16458
rect 10692 16244 10744 16250
rect 10692 16186 10744 16192
rect 12440 16244 12492 16250
rect 12440 16186 12492 16192
rect 10508 16108 10560 16114
rect 10508 16050 10560 16056
rect 11704 16108 11756 16114
rect 11704 16050 11756 16056
rect 12256 16108 12308 16114
rect 12256 16050 12308 16056
rect 11428 15496 11480 15502
rect 11428 15438 11480 15444
rect 10876 15360 10928 15366
rect 10876 15302 10928 15308
rect 10888 15026 10916 15302
rect 10876 15020 10928 15026
rect 10876 14962 10928 14968
rect 10784 14816 10836 14822
rect 10784 14758 10836 14764
rect 10416 14340 10468 14346
rect 10416 14282 10468 14288
rect 10324 14000 10376 14006
rect 10324 13942 10376 13948
rect 10336 13870 10364 13942
rect 10324 13864 10376 13870
rect 10324 13806 10376 13812
rect 10232 13524 10284 13530
rect 10232 13466 10284 13472
rect 10324 13456 10376 13462
rect 10324 13398 10376 13404
rect 9956 13252 10008 13258
rect 9956 13194 10008 13200
rect 9827 13084 10135 13093
rect 9827 13082 9833 13084
rect 9889 13082 9913 13084
rect 9969 13082 9993 13084
rect 10049 13082 10073 13084
rect 10129 13082 10135 13084
rect 9889 13030 9891 13082
rect 10071 13030 10073 13082
rect 9827 13028 9833 13030
rect 9889 13028 9913 13030
rect 9969 13028 9993 13030
rect 10049 13028 10073 13030
rect 10129 13028 10135 13030
rect 9827 13019 10135 13028
rect 10336 12850 10364 13398
rect 9680 12844 9732 12850
rect 9680 12786 9732 12792
rect 10324 12844 10376 12850
rect 10324 12786 10376 12792
rect 9692 10266 9720 12786
rect 10428 12730 10456 14282
rect 10508 14272 10560 14278
rect 10508 14214 10560 14220
rect 10520 13326 10548 14214
rect 10796 13938 10824 14758
rect 10784 13932 10836 13938
rect 10784 13874 10836 13880
rect 10796 13462 10824 13874
rect 10876 13864 10928 13870
rect 10876 13806 10928 13812
rect 10784 13456 10836 13462
rect 10784 13398 10836 13404
rect 10508 13320 10560 13326
rect 10508 13262 10560 13268
rect 10600 13320 10652 13326
rect 10600 13262 10652 13268
rect 10244 12702 10456 12730
rect 10048 12436 10100 12442
rect 10048 12378 10100 12384
rect 10060 12102 10088 12378
rect 10244 12102 10272 12702
rect 10520 12646 10548 13262
rect 10612 12986 10640 13262
rect 10600 12980 10652 12986
rect 10600 12922 10652 12928
rect 10508 12640 10560 12646
rect 10508 12582 10560 12588
rect 10784 12640 10836 12646
rect 10784 12582 10836 12588
rect 10692 12436 10744 12442
rect 10692 12378 10744 12384
rect 10324 12232 10376 12238
rect 10324 12174 10376 12180
rect 10048 12096 10100 12102
rect 10048 12038 10100 12044
rect 10232 12096 10284 12102
rect 10232 12038 10284 12044
rect 9827 11996 10135 12005
rect 9827 11994 9833 11996
rect 9889 11994 9913 11996
rect 9969 11994 9993 11996
rect 10049 11994 10073 11996
rect 10129 11994 10135 11996
rect 9889 11942 9891 11994
rect 10071 11942 10073 11994
rect 9827 11940 9833 11942
rect 9889 11940 9913 11942
rect 9969 11940 9993 11942
rect 10049 11940 10073 11942
rect 10129 11940 10135 11942
rect 9827 11931 10135 11940
rect 9827 10908 10135 10917
rect 9827 10906 9833 10908
rect 9889 10906 9913 10908
rect 9969 10906 9993 10908
rect 10049 10906 10073 10908
rect 10129 10906 10135 10908
rect 9889 10854 9891 10906
rect 10071 10854 10073 10906
rect 9827 10852 9833 10854
rect 9889 10852 9913 10854
rect 9969 10852 9993 10854
rect 10049 10852 10073 10854
rect 10129 10852 10135 10854
rect 9827 10843 10135 10852
rect 9680 10260 9732 10266
rect 9680 10202 9732 10208
rect 9827 9820 10135 9829
rect 9827 9818 9833 9820
rect 9889 9818 9913 9820
rect 9969 9818 9993 9820
rect 10049 9818 10073 9820
rect 10129 9818 10135 9820
rect 9889 9766 9891 9818
rect 10071 9766 10073 9818
rect 9827 9764 9833 9766
rect 9889 9764 9913 9766
rect 9969 9764 9993 9766
rect 10049 9764 10073 9766
rect 10129 9764 10135 9766
rect 9827 9755 10135 9764
rect 9588 9648 9640 9654
rect 9588 9590 9640 9596
rect 10244 9602 10272 12038
rect 10336 10674 10364 12174
rect 10508 12164 10560 12170
rect 10508 12106 10560 12112
rect 10416 12096 10468 12102
rect 10416 12038 10468 12044
rect 10428 11898 10456 12038
rect 10416 11892 10468 11898
rect 10416 11834 10468 11840
rect 10520 11762 10548 12106
rect 10508 11756 10560 11762
rect 10508 11698 10560 11704
rect 10520 11354 10548 11698
rect 10508 11348 10560 11354
rect 10508 11290 10560 11296
rect 10324 10668 10376 10674
rect 10324 10610 10376 10616
rect 10336 9722 10364 10610
rect 10520 10130 10548 11290
rect 10508 10124 10560 10130
rect 10508 10066 10560 10072
rect 10324 9716 10376 9722
rect 10324 9658 10376 9664
rect 9600 9178 9628 9590
rect 10244 9574 10364 9602
rect 9588 9172 9640 9178
rect 9588 9114 9640 9120
rect 9600 8906 9628 9114
rect 10232 9036 10284 9042
rect 10232 8978 10284 8984
rect 9588 8900 9640 8906
rect 9588 8842 9640 8848
rect 9827 8732 10135 8741
rect 9827 8730 9833 8732
rect 9889 8730 9913 8732
rect 9969 8730 9993 8732
rect 10049 8730 10073 8732
rect 10129 8730 10135 8732
rect 9889 8678 9891 8730
rect 10071 8678 10073 8730
rect 9827 8676 9833 8678
rect 9889 8676 9913 8678
rect 9969 8676 9993 8678
rect 10049 8676 10073 8678
rect 10129 8676 10135 8678
rect 9827 8667 10135 8676
rect 9680 8628 9732 8634
rect 9680 8570 9732 8576
rect 9692 8294 9720 8570
rect 9680 8288 9732 8294
rect 9680 8230 9732 8236
rect 9680 8016 9732 8022
rect 9680 7958 9732 7964
rect 9496 7812 9548 7818
rect 9496 7754 9548 7760
rect 9508 7410 9536 7754
rect 9692 7410 9720 7958
rect 10244 7750 10272 8978
rect 10336 8634 10364 9574
rect 10600 9512 10652 9518
rect 10600 9454 10652 9460
rect 10612 9178 10640 9454
rect 10600 9172 10652 9178
rect 10600 9114 10652 9120
rect 10508 9104 10560 9110
rect 10508 9046 10560 9052
rect 10324 8628 10376 8634
rect 10324 8570 10376 8576
rect 10520 8430 10548 9046
rect 10612 8498 10640 9114
rect 10600 8492 10652 8498
rect 10600 8434 10652 8440
rect 10508 8424 10560 8430
rect 10508 8366 10560 8372
rect 10324 8288 10376 8294
rect 10324 8230 10376 8236
rect 10336 7818 10364 8230
rect 10324 7812 10376 7818
rect 10324 7754 10376 7760
rect 10232 7744 10284 7750
rect 10232 7686 10284 7692
rect 9827 7644 10135 7653
rect 9827 7642 9833 7644
rect 9889 7642 9913 7644
rect 9969 7642 9993 7644
rect 10049 7642 10073 7644
rect 10129 7642 10135 7644
rect 9889 7590 9891 7642
rect 10071 7590 10073 7642
rect 9827 7588 9833 7590
rect 9889 7588 9913 7590
rect 9969 7588 9993 7590
rect 10049 7588 10073 7590
rect 10129 7588 10135 7590
rect 9827 7579 10135 7588
rect 9496 7404 9548 7410
rect 9496 7346 9548 7352
rect 9680 7404 9732 7410
rect 9680 7346 9732 7352
rect 9036 7268 9088 7274
rect 9036 7210 9088 7216
rect 9680 7268 9732 7274
rect 9680 7210 9732 7216
rect 8760 6724 8812 6730
rect 8760 6666 8812 6672
rect 8668 6656 8720 6662
rect 8668 6598 8720 6604
rect 8208 5704 8260 5710
rect 8484 5704 8536 5710
rect 8260 5652 8340 5658
rect 8208 5646 8340 5652
rect 8484 5646 8536 5652
rect 8576 5704 8628 5710
rect 8576 5646 8628 5652
rect 8220 5630 8340 5646
rect 7932 4616 7984 4622
rect 7932 4558 7984 4564
rect 7564 4548 7616 4554
rect 7564 4490 7616 4496
rect 7576 4146 7604 4490
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 7932 4072 7984 4078
rect 7932 4014 7984 4020
rect 7608 3836 7916 3845
rect 7608 3834 7614 3836
rect 7670 3834 7694 3836
rect 7750 3834 7774 3836
rect 7830 3834 7854 3836
rect 7910 3834 7916 3836
rect 7670 3782 7672 3834
rect 7852 3782 7854 3834
rect 7608 3780 7614 3782
rect 7670 3780 7694 3782
rect 7750 3780 7774 3782
rect 7830 3780 7854 3782
rect 7910 3780 7916 3782
rect 7608 3771 7916 3780
rect 7944 3602 7972 4014
rect 8312 3738 8340 5630
rect 8496 4282 8524 5646
rect 8484 4276 8536 4282
rect 8484 4218 8536 4224
rect 8392 3936 8444 3942
rect 8392 3878 8444 3884
rect 8300 3732 8352 3738
rect 8300 3674 8352 3680
rect 8404 3670 8432 3878
rect 8392 3664 8444 3670
rect 8392 3606 8444 3612
rect 7932 3596 7984 3602
rect 7932 3538 7984 3544
rect 8496 3534 8524 4218
rect 8588 4162 8616 5646
rect 8680 5166 8708 6598
rect 8772 6254 8800 6666
rect 9048 6390 9076 7210
rect 9692 6798 9720 7210
rect 9864 7200 9916 7206
rect 9864 7142 9916 7148
rect 9876 6798 9904 7142
rect 9128 6792 9180 6798
rect 9128 6734 9180 6740
rect 9680 6792 9732 6798
rect 9680 6734 9732 6740
rect 9864 6792 9916 6798
rect 9864 6734 9916 6740
rect 9036 6384 9088 6390
rect 9036 6326 9088 6332
rect 8760 6248 8812 6254
rect 8760 6190 8812 6196
rect 8668 5160 8720 5166
rect 8668 5102 8720 5108
rect 9140 4826 9168 6734
rect 9404 6656 9456 6662
rect 9404 6598 9456 6604
rect 9416 6322 9444 6598
rect 9404 6316 9456 6322
rect 9404 6258 9456 6264
rect 9692 5302 9720 6734
rect 10336 6730 10364 7754
rect 10704 6730 10732 12378
rect 10796 11150 10824 12582
rect 10888 12306 10916 13806
rect 11440 13190 11468 15438
rect 11716 14618 11744 16050
rect 12268 15978 12296 16050
rect 11796 15972 11848 15978
rect 11796 15914 11848 15920
rect 12256 15972 12308 15978
rect 12256 15914 12308 15920
rect 11704 14612 11756 14618
rect 11704 14554 11756 14560
rect 11716 14414 11744 14554
rect 11704 14408 11756 14414
rect 11704 14350 11756 14356
rect 10968 13184 11020 13190
rect 10968 13126 11020 13132
rect 11428 13184 11480 13190
rect 11428 13126 11480 13132
rect 10980 12306 11008 13126
rect 11060 12640 11112 12646
rect 11060 12582 11112 12588
rect 11152 12640 11204 12646
rect 11152 12582 11204 12588
rect 11072 12442 11100 12582
rect 11060 12436 11112 12442
rect 11060 12378 11112 12384
rect 10876 12300 10928 12306
rect 10876 12242 10928 12248
rect 10968 12300 11020 12306
rect 10968 12242 11020 12248
rect 11164 12238 11192 12582
rect 11244 12300 11296 12306
rect 11244 12242 11296 12248
rect 11152 12232 11204 12238
rect 11152 12174 11204 12180
rect 11060 11824 11112 11830
rect 11060 11766 11112 11772
rect 10784 11144 10836 11150
rect 10784 11086 10836 11092
rect 10796 9586 10824 11086
rect 10784 9580 10836 9586
rect 10784 9522 10836 9528
rect 11072 9450 11100 11766
rect 11256 9654 11284 12242
rect 11336 10056 11388 10062
rect 11440 10044 11468 13126
rect 11612 12844 11664 12850
rect 11612 12786 11664 12792
rect 11520 12436 11572 12442
rect 11520 12378 11572 12384
rect 11532 10810 11560 12378
rect 11624 11762 11652 12786
rect 11704 12232 11756 12238
rect 11704 12174 11756 12180
rect 11612 11756 11664 11762
rect 11612 11698 11664 11704
rect 11716 11558 11744 12174
rect 11704 11552 11756 11558
rect 11704 11494 11756 11500
rect 11716 11286 11744 11494
rect 11704 11280 11756 11286
rect 11704 11222 11756 11228
rect 11808 10810 11836 15914
rect 12047 15804 12355 15813
rect 12047 15802 12053 15804
rect 12109 15802 12133 15804
rect 12189 15802 12213 15804
rect 12269 15802 12293 15804
rect 12349 15802 12355 15804
rect 12109 15750 12111 15802
rect 12291 15750 12293 15802
rect 12047 15748 12053 15750
rect 12109 15748 12133 15750
rect 12189 15748 12213 15750
rect 12269 15748 12293 15750
rect 12349 15748 12355 15750
rect 12047 15739 12355 15748
rect 12452 15706 12480 16186
rect 12440 15700 12492 15706
rect 12440 15642 12492 15648
rect 12532 15020 12584 15026
rect 12532 14962 12584 14968
rect 12047 14716 12355 14725
rect 12047 14714 12053 14716
rect 12109 14714 12133 14716
rect 12189 14714 12213 14716
rect 12269 14714 12293 14716
rect 12349 14714 12355 14716
rect 12109 14662 12111 14714
rect 12291 14662 12293 14714
rect 12047 14660 12053 14662
rect 12109 14660 12133 14662
rect 12189 14660 12213 14662
rect 12269 14660 12293 14662
rect 12349 14660 12355 14662
rect 12047 14651 12355 14660
rect 12544 14618 12572 14962
rect 12532 14612 12584 14618
rect 12532 14554 12584 14560
rect 12624 14476 12676 14482
rect 12624 14418 12676 14424
rect 12636 14074 12664 14418
rect 12624 14068 12676 14074
rect 12624 14010 12676 14016
rect 12440 13796 12492 13802
rect 12440 13738 12492 13744
rect 12047 13628 12355 13637
rect 12047 13626 12053 13628
rect 12109 13626 12133 13628
rect 12189 13626 12213 13628
rect 12269 13626 12293 13628
rect 12349 13626 12355 13628
rect 12109 13574 12111 13626
rect 12291 13574 12293 13626
rect 12047 13572 12053 13574
rect 12109 13572 12133 13574
rect 12189 13572 12213 13574
rect 12269 13572 12293 13574
rect 12349 13572 12355 13574
rect 12047 13563 12355 13572
rect 12256 13388 12308 13394
rect 12256 13330 12308 13336
rect 12164 13320 12216 13326
rect 12164 13262 12216 13268
rect 12176 12850 12204 13262
rect 12164 12844 12216 12850
rect 12164 12786 12216 12792
rect 12268 12782 12296 13330
rect 12452 12918 12480 13738
rect 12716 13184 12768 13190
rect 12716 13126 12768 13132
rect 12440 12912 12492 12918
rect 12440 12854 12492 12860
rect 12256 12776 12308 12782
rect 12256 12718 12308 12724
rect 12047 12540 12355 12549
rect 12047 12538 12053 12540
rect 12109 12538 12133 12540
rect 12189 12538 12213 12540
rect 12269 12538 12293 12540
rect 12349 12538 12355 12540
rect 12109 12486 12111 12538
rect 12291 12486 12293 12538
rect 12047 12484 12053 12486
rect 12109 12484 12133 12486
rect 12189 12484 12213 12486
rect 12269 12484 12293 12486
rect 12349 12484 12355 12486
rect 12047 12475 12355 12484
rect 12532 12096 12584 12102
rect 12532 12038 12584 12044
rect 12624 12096 12676 12102
rect 12624 12038 12676 12044
rect 12544 11898 12572 12038
rect 12532 11892 12584 11898
rect 12532 11834 12584 11840
rect 11888 11620 11940 11626
rect 11888 11562 11940 11568
rect 12440 11620 12492 11626
rect 12440 11562 12492 11568
rect 11900 11218 11928 11562
rect 12047 11452 12355 11461
rect 12047 11450 12053 11452
rect 12109 11450 12133 11452
rect 12189 11450 12213 11452
rect 12269 11450 12293 11452
rect 12349 11450 12355 11452
rect 12109 11398 12111 11450
rect 12291 11398 12293 11450
rect 12047 11396 12053 11398
rect 12109 11396 12133 11398
rect 12189 11396 12213 11398
rect 12269 11396 12293 11398
rect 12349 11396 12355 11398
rect 12047 11387 12355 11396
rect 11888 11212 11940 11218
rect 11888 11154 11940 11160
rect 12452 11082 12480 11562
rect 12544 11150 12572 11834
rect 12636 11762 12664 12038
rect 12624 11756 12676 11762
rect 12624 11698 12676 11704
rect 12728 11150 12756 13126
rect 12820 12714 12848 16458
rect 14266 16348 14574 16357
rect 14266 16346 14272 16348
rect 14328 16346 14352 16348
rect 14408 16346 14432 16348
rect 14488 16346 14512 16348
rect 14568 16346 14574 16348
rect 14328 16294 14330 16346
rect 14510 16294 14512 16346
rect 14266 16292 14272 16294
rect 14328 16292 14352 16294
rect 14408 16292 14432 16294
rect 14488 16292 14512 16294
rect 14568 16292 14574 16294
rect 14266 16283 14574 16292
rect 13728 16040 13780 16046
rect 13728 15982 13780 15988
rect 13268 15496 13320 15502
rect 13268 15438 13320 15444
rect 13280 14822 13308 15438
rect 13740 15178 13768 15982
rect 16486 15804 16794 15813
rect 16486 15802 16492 15804
rect 16548 15802 16572 15804
rect 16628 15802 16652 15804
rect 16708 15802 16732 15804
rect 16788 15802 16794 15804
rect 16548 15750 16550 15802
rect 16730 15750 16732 15802
rect 16486 15748 16492 15750
rect 16548 15748 16572 15750
rect 16628 15748 16652 15750
rect 16708 15748 16732 15750
rect 16788 15748 16794 15750
rect 16486 15739 16794 15748
rect 15844 15428 15896 15434
rect 15844 15370 15896 15376
rect 14648 15360 14700 15366
rect 14648 15302 14700 15308
rect 15752 15360 15804 15366
rect 15752 15302 15804 15308
rect 14266 15260 14574 15269
rect 14266 15258 14272 15260
rect 14328 15258 14352 15260
rect 14408 15258 14432 15260
rect 14488 15258 14512 15260
rect 14568 15258 14574 15260
rect 14328 15206 14330 15258
rect 14510 15206 14512 15258
rect 14266 15204 14272 15206
rect 14328 15204 14352 15206
rect 14408 15204 14432 15206
rect 14488 15204 14512 15206
rect 14568 15204 14574 15206
rect 14266 15195 14574 15204
rect 13740 15150 13860 15178
rect 13832 15094 13860 15150
rect 13820 15088 13872 15094
rect 13820 15030 13872 15036
rect 13832 14958 13860 15030
rect 13820 14952 13872 14958
rect 13820 14894 13872 14900
rect 13268 14816 13320 14822
rect 13268 14758 13320 14764
rect 13280 14414 13308 14758
rect 13268 14408 13320 14414
rect 13268 14350 13320 14356
rect 13280 14006 13308 14350
rect 13268 14000 13320 14006
rect 13268 13942 13320 13948
rect 12992 13728 13044 13734
rect 12992 13670 13044 13676
rect 12808 12708 12860 12714
rect 12808 12650 12860 12656
rect 12808 12232 12860 12238
rect 12808 12174 12860 12180
rect 12820 11762 12848 12174
rect 12808 11756 12860 11762
rect 12808 11698 12860 11704
rect 12900 11280 12952 11286
rect 12900 11222 12952 11228
rect 12532 11144 12584 11150
rect 12532 11086 12584 11092
rect 12716 11144 12768 11150
rect 12716 11086 12768 11092
rect 11888 11076 11940 11082
rect 11888 11018 11940 11024
rect 12440 11076 12492 11082
rect 12440 11018 12492 11024
rect 12624 11076 12676 11082
rect 12624 11018 12676 11024
rect 11520 10804 11572 10810
rect 11520 10746 11572 10752
rect 11796 10804 11848 10810
rect 11796 10746 11848 10752
rect 11532 10198 11560 10746
rect 11704 10668 11756 10674
rect 11704 10610 11756 10616
rect 11716 10266 11744 10610
rect 11704 10260 11756 10266
rect 11704 10202 11756 10208
rect 11520 10192 11572 10198
rect 11520 10134 11572 10140
rect 11440 10016 11560 10044
rect 11336 9998 11388 10004
rect 11348 9654 11376 9998
rect 11428 9920 11480 9926
rect 11428 9862 11480 9868
rect 11440 9722 11468 9862
rect 11428 9716 11480 9722
rect 11428 9658 11480 9664
rect 11244 9648 11296 9654
rect 11244 9590 11296 9596
rect 11336 9648 11388 9654
rect 11336 9590 11388 9596
rect 11440 9518 11468 9658
rect 11428 9512 11480 9518
rect 11428 9454 11480 9460
rect 11060 9444 11112 9450
rect 11060 9386 11112 9392
rect 10968 9376 11020 9382
rect 10968 9318 11020 9324
rect 10980 8974 11008 9318
rect 11440 9042 11468 9454
rect 11532 9110 11560 10016
rect 11612 9920 11664 9926
rect 11612 9862 11664 9868
rect 11520 9104 11572 9110
rect 11520 9046 11572 9052
rect 11428 9036 11480 9042
rect 11428 8978 11480 8984
rect 10968 8968 11020 8974
rect 10968 8910 11020 8916
rect 11428 8900 11480 8906
rect 11428 8842 11480 8848
rect 11060 8832 11112 8838
rect 11060 8774 11112 8780
rect 11072 8498 11100 8774
rect 11060 8492 11112 8498
rect 11060 8434 11112 8440
rect 11072 7954 11100 8434
rect 11152 8288 11204 8294
rect 11152 8230 11204 8236
rect 11060 7948 11112 7954
rect 11060 7890 11112 7896
rect 11164 7410 11192 8230
rect 11152 7404 11204 7410
rect 11152 7346 11204 7352
rect 10324 6724 10376 6730
rect 10324 6666 10376 6672
rect 10692 6724 10744 6730
rect 10692 6666 10744 6672
rect 9827 6556 10135 6565
rect 9827 6554 9833 6556
rect 9889 6554 9913 6556
rect 9969 6554 9993 6556
rect 10049 6554 10073 6556
rect 10129 6554 10135 6556
rect 9889 6502 9891 6554
rect 10071 6502 10073 6554
rect 9827 6500 9833 6502
rect 9889 6500 9913 6502
rect 9969 6500 9993 6502
rect 10049 6500 10073 6502
rect 10129 6500 10135 6502
rect 9827 6491 10135 6500
rect 10336 6254 10364 6666
rect 10508 6452 10560 6458
rect 10508 6394 10560 6400
rect 10324 6248 10376 6254
rect 10324 6190 10376 6196
rect 10416 5840 10468 5846
rect 10416 5782 10468 5788
rect 10324 5772 10376 5778
rect 10324 5714 10376 5720
rect 10232 5568 10284 5574
rect 10232 5510 10284 5516
rect 9827 5468 10135 5477
rect 9827 5466 9833 5468
rect 9889 5466 9913 5468
rect 9969 5466 9993 5468
rect 10049 5466 10073 5468
rect 10129 5466 10135 5468
rect 9889 5414 9891 5466
rect 10071 5414 10073 5466
rect 9827 5412 9833 5414
rect 9889 5412 9913 5414
rect 9969 5412 9993 5414
rect 10049 5412 10073 5414
rect 10129 5412 10135 5414
rect 9827 5403 10135 5412
rect 9680 5296 9732 5302
rect 9680 5238 9732 5244
rect 9956 5160 10008 5166
rect 9956 5102 10008 5108
rect 9128 4820 9180 4826
rect 9128 4762 9180 4768
rect 9968 4554 9996 5102
rect 10244 4826 10272 5510
rect 10232 4820 10284 4826
rect 10232 4762 10284 4768
rect 10336 4690 10364 5714
rect 10428 5710 10456 5782
rect 10416 5704 10468 5710
rect 10416 5646 10468 5652
rect 10324 4684 10376 4690
rect 10324 4626 10376 4632
rect 10428 4622 10456 5646
rect 10416 4616 10468 4622
rect 10416 4558 10468 4564
rect 9956 4548 10008 4554
rect 9956 4490 10008 4496
rect 10428 4486 10456 4558
rect 10520 4554 10548 6394
rect 10704 6390 10732 6666
rect 10692 6384 10744 6390
rect 10692 6326 10744 6332
rect 10704 5778 10732 6326
rect 11440 6186 11468 8842
rect 11532 8294 11560 9046
rect 11624 8430 11652 9862
rect 11796 9376 11848 9382
rect 11796 9318 11848 9324
rect 11704 8968 11756 8974
rect 11704 8910 11756 8916
rect 11716 8498 11744 8910
rect 11808 8906 11836 9318
rect 11900 9024 11928 11018
rect 12636 10810 12664 11018
rect 12808 11008 12860 11014
rect 12808 10950 12860 10956
rect 12624 10804 12676 10810
rect 12624 10746 12676 10752
rect 12820 10674 12848 10950
rect 12912 10810 12940 11222
rect 13004 11218 13032 13670
rect 13832 13326 13860 14894
rect 14660 14414 14688 15302
rect 14924 15020 14976 15026
rect 14924 14962 14976 14968
rect 14648 14408 14700 14414
rect 14648 14350 14700 14356
rect 14096 14272 14148 14278
rect 14096 14214 14148 14220
rect 14832 14272 14884 14278
rect 14832 14214 14884 14220
rect 13820 13320 13872 13326
rect 13820 13262 13872 13268
rect 13084 12912 13136 12918
rect 13084 12854 13136 12860
rect 12992 11212 13044 11218
rect 12992 11154 13044 11160
rect 12900 10804 12952 10810
rect 12900 10746 12952 10752
rect 12532 10668 12584 10674
rect 12532 10610 12584 10616
rect 12808 10668 12860 10674
rect 12808 10610 12860 10616
rect 12047 10364 12355 10373
rect 12047 10362 12053 10364
rect 12109 10362 12133 10364
rect 12189 10362 12213 10364
rect 12269 10362 12293 10364
rect 12349 10362 12355 10364
rect 12109 10310 12111 10362
rect 12291 10310 12293 10362
rect 12047 10308 12053 10310
rect 12109 10308 12133 10310
rect 12189 10308 12213 10310
rect 12269 10308 12293 10310
rect 12349 10308 12355 10310
rect 12047 10299 12355 10308
rect 11980 9648 12032 9654
rect 11978 9616 11980 9625
rect 12032 9616 12034 9625
rect 11978 9551 12034 9560
rect 12348 9580 12400 9586
rect 12348 9522 12400 9528
rect 12360 9450 12388 9522
rect 12348 9444 12400 9450
rect 12348 9386 12400 9392
rect 12047 9276 12355 9285
rect 12047 9274 12053 9276
rect 12109 9274 12133 9276
rect 12189 9274 12213 9276
rect 12269 9274 12293 9276
rect 12349 9274 12355 9276
rect 12109 9222 12111 9274
rect 12291 9222 12293 9274
rect 12047 9220 12053 9222
rect 12109 9220 12133 9222
rect 12189 9220 12213 9222
rect 12269 9220 12293 9222
rect 12349 9220 12355 9222
rect 12047 9211 12355 9220
rect 12360 9042 12480 9058
rect 12256 9036 12308 9042
rect 11900 8996 12256 9024
rect 12256 8978 12308 8984
rect 12360 9036 12492 9042
rect 12360 9030 12440 9036
rect 11796 8900 11848 8906
rect 11796 8842 11848 8848
rect 11808 8498 11836 8842
rect 11888 8832 11940 8838
rect 11888 8774 11940 8780
rect 12254 8800 12310 8809
rect 11704 8492 11756 8498
rect 11704 8434 11756 8440
rect 11796 8492 11848 8498
rect 11796 8434 11848 8440
rect 11612 8424 11664 8430
rect 11612 8366 11664 8372
rect 11520 8288 11572 8294
rect 11520 8230 11572 8236
rect 11900 8090 11928 8774
rect 12254 8735 12310 8744
rect 12268 8634 12296 8735
rect 12256 8628 12308 8634
rect 12256 8570 12308 8576
rect 12360 8430 12388 9030
rect 12440 8978 12492 8984
rect 12544 8838 12572 10610
rect 12912 10606 12940 10746
rect 13004 10674 13032 11154
rect 12992 10668 13044 10674
rect 12992 10610 13044 10616
rect 12900 10600 12952 10606
rect 12900 10542 12952 10548
rect 12808 10532 12860 10538
rect 12808 10474 12860 10480
rect 12820 10062 12848 10474
rect 12808 10056 12860 10062
rect 12808 9998 12860 10004
rect 12912 9330 12940 10542
rect 12992 9648 13044 9654
rect 12992 9590 13044 9596
rect 12820 9302 12940 9330
rect 12532 8832 12584 8838
rect 12532 8774 12584 8780
rect 12348 8424 12400 8430
rect 12348 8366 12400 8372
rect 12047 8188 12355 8197
rect 12047 8186 12053 8188
rect 12109 8186 12133 8188
rect 12189 8186 12213 8188
rect 12269 8186 12293 8188
rect 12349 8186 12355 8188
rect 12109 8134 12111 8186
rect 12291 8134 12293 8186
rect 12047 8132 12053 8134
rect 12109 8132 12133 8134
rect 12189 8132 12213 8134
rect 12269 8132 12293 8134
rect 12349 8132 12355 8134
rect 12047 8123 12355 8132
rect 11888 8084 11940 8090
rect 11888 8026 11940 8032
rect 11612 8016 11664 8022
rect 11612 7958 11664 7964
rect 11624 7342 11652 7958
rect 12164 7880 12216 7886
rect 12164 7822 12216 7828
rect 12176 7546 12204 7822
rect 12820 7818 12848 9302
rect 13004 9178 13032 9590
rect 12900 9172 12952 9178
rect 12900 9114 12952 9120
rect 12992 9172 13044 9178
rect 12992 9114 13044 9120
rect 12912 8838 12940 9114
rect 12900 8832 12952 8838
rect 12900 8774 12952 8780
rect 12808 7812 12860 7818
rect 12808 7754 12860 7760
rect 12164 7540 12216 7546
rect 12164 7482 12216 7488
rect 11612 7336 11664 7342
rect 11612 7278 11664 7284
rect 11428 6180 11480 6186
rect 11428 6122 11480 6128
rect 11440 5914 11468 6122
rect 11428 5908 11480 5914
rect 11428 5850 11480 5856
rect 10692 5772 10744 5778
rect 10692 5714 10744 5720
rect 11152 5704 11204 5710
rect 11152 5646 11204 5652
rect 10784 5568 10836 5574
rect 10784 5510 10836 5516
rect 10796 4826 10824 5510
rect 11060 5364 11112 5370
rect 11060 5306 11112 5312
rect 10784 4820 10836 4826
rect 10784 4762 10836 4768
rect 11072 4554 11100 5306
rect 11164 5234 11192 5646
rect 11152 5228 11204 5234
rect 11152 5170 11204 5176
rect 10508 4548 10560 4554
rect 10508 4490 10560 4496
rect 11060 4548 11112 4554
rect 11060 4490 11112 4496
rect 9680 4480 9732 4486
rect 9680 4422 9732 4428
rect 10416 4480 10468 4486
rect 10416 4422 10468 4428
rect 10692 4480 10744 4486
rect 10692 4422 10744 4428
rect 8588 4146 8708 4162
rect 8588 4140 8720 4146
rect 8588 4134 8668 4140
rect 7472 3528 7524 3534
rect 7472 3470 7524 3476
rect 8392 3528 8444 3534
rect 8392 3470 8444 3476
rect 8484 3528 8536 3534
rect 8484 3470 8536 3476
rect 7932 3460 7984 3466
rect 7932 3402 7984 3408
rect 7380 3188 7432 3194
rect 7380 3130 7432 3136
rect 7012 3052 7064 3058
rect 7012 2994 7064 3000
rect 7196 3052 7248 3058
rect 7196 2994 7248 3000
rect 6840 2746 6960 2774
rect 6932 2514 6960 2746
rect 6920 2508 6972 2514
rect 6920 2450 6972 2456
rect 3976 2440 4028 2446
rect 3976 2382 4028 2388
rect 4252 2440 4304 2446
rect 4252 2382 4304 2388
rect 6000 2440 6052 2446
rect 6000 2382 6052 2388
rect 6552 2440 6604 2446
rect 6552 2382 6604 2388
rect 6736 2440 6788 2446
rect 6736 2382 6788 2388
rect 7392 2378 7420 3130
rect 7608 2748 7916 2757
rect 7608 2746 7614 2748
rect 7670 2746 7694 2748
rect 7750 2746 7774 2748
rect 7830 2746 7854 2748
rect 7910 2746 7916 2748
rect 7670 2694 7672 2746
rect 7852 2694 7854 2746
rect 7608 2692 7614 2694
rect 7670 2692 7694 2694
rect 7750 2692 7774 2694
rect 7830 2692 7854 2694
rect 7910 2692 7916 2694
rect 7608 2683 7916 2692
rect 7944 2446 7972 3402
rect 8404 3380 8432 3470
rect 8588 3380 8616 4134
rect 8668 4082 8720 4088
rect 9588 4140 9640 4146
rect 9588 4082 9640 4088
rect 9312 4072 9364 4078
rect 9312 4014 9364 4020
rect 9036 3664 9088 3670
rect 9036 3606 9088 3612
rect 8404 3352 8616 3380
rect 8668 2848 8720 2854
rect 8668 2790 8720 2796
rect 8680 2446 8708 2790
rect 7932 2440 7984 2446
rect 7932 2382 7984 2388
rect 8668 2440 8720 2446
rect 8668 2382 8720 2388
rect 9048 2378 9076 3606
rect 9324 3058 9352 4014
rect 9600 3738 9628 4082
rect 9588 3732 9640 3738
rect 9588 3674 9640 3680
rect 9692 3534 9720 4422
rect 9827 4380 10135 4389
rect 9827 4378 9833 4380
rect 9889 4378 9913 4380
rect 9969 4378 9993 4380
rect 10049 4378 10073 4380
rect 10129 4378 10135 4380
rect 9889 4326 9891 4378
rect 10071 4326 10073 4378
rect 9827 4324 9833 4326
rect 9889 4324 9913 4326
rect 9969 4324 9993 4326
rect 10049 4324 10073 4326
rect 10129 4324 10135 4326
rect 9827 4315 10135 4324
rect 10704 4282 10732 4422
rect 11164 4282 11192 5170
rect 11440 5030 11468 5850
rect 11428 5024 11480 5030
rect 11428 4966 11480 4972
rect 11624 4978 11652 7278
rect 12047 7100 12355 7109
rect 12047 7098 12053 7100
rect 12109 7098 12133 7100
rect 12189 7098 12213 7100
rect 12269 7098 12293 7100
rect 12349 7098 12355 7100
rect 12109 7046 12111 7098
rect 12291 7046 12293 7098
rect 12047 7044 12053 7046
rect 12109 7044 12133 7046
rect 12189 7044 12213 7046
rect 12269 7044 12293 7046
rect 12349 7044 12355 7046
rect 12047 7035 12355 7044
rect 12820 6322 12848 7754
rect 13096 7750 13124 12854
rect 13832 12434 13860 13262
rect 14108 12918 14136 14214
rect 14266 14172 14574 14181
rect 14266 14170 14272 14172
rect 14328 14170 14352 14172
rect 14408 14170 14432 14172
rect 14488 14170 14512 14172
rect 14568 14170 14574 14172
rect 14328 14118 14330 14170
rect 14510 14118 14512 14170
rect 14266 14116 14272 14118
rect 14328 14116 14352 14118
rect 14408 14116 14432 14118
rect 14488 14116 14512 14118
rect 14568 14116 14574 14118
rect 14266 14107 14574 14116
rect 14844 13938 14872 14214
rect 14936 14074 14964 14962
rect 15384 14544 15436 14550
rect 15384 14486 15436 14492
rect 14924 14068 14976 14074
rect 14924 14010 14976 14016
rect 14188 13932 14240 13938
rect 14188 13874 14240 13880
rect 14648 13932 14700 13938
rect 14648 13874 14700 13880
rect 14832 13932 14884 13938
rect 14832 13874 14884 13880
rect 14200 12986 14228 13874
rect 14372 13728 14424 13734
rect 14372 13670 14424 13676
rect 14384 13326 14412 13670
rect 14372 13320 14424 13326
rect 14372 13262 14424 13268
rect 14266 13084 14574 13093
rect 14266 13082 14272 13084
rect 14328 13082 14352 13084
rect 14408 13082 14432 13084
rect 14488 13082 14512 13084
rect 14568 13082 14574 13084
rect 14328 13030 14330 13082
rect 14510 13030 14512 13082
rect 14266 13028 14272 13030
rect 14328 13028 14352 13030
rect 14408 13028 14432 13030
rect 14488 13028 14512 13030
rect 14568 13028 14574 13030
rect 14266 13019 14574 13028
rect 14660 12986 14688 13874
rect 14188 12980 14240 12986
rect 14188 12922 14240 12928
rect 14648 12980 14700 12986
rect 14648 12922 14700 12928
rect 14096 12912 14148 12918
rect 14096 12854 14148 12860
rect 13832 12406 14044 12434
rect 14016 12238 14044 12406
rect 14004 12232 14056 12238
rect 14004 12174 14056 12180
rect 13360 11552 13412 11558
rect 13360 11494 13412 11500
rect 13176 11348 13228 11354
rect 13176 11290 13228 11296
rect 13188 10198 13216 11290
rect 13268 11076 13320 11082
rect 13268 11018 13320 11024
rect 13280 10470 13308 11018
rect 13268 10464 13320 10470
rect 13268 10406 13320 10412
rect 13176 10192 13228 10198
rect 13176 10134 13228 10140
rect 13176 9648 13228 9654
rect 13176 9590 13228 9596
rect 13188 9450 13216 9590
rect 13176 9444 13228 9450
rect 13176 9386 13228 9392
rect 13372 8634 13400 11494
rect 13728 11008 13780 11014
rect 13728 10950 13780 10956
rect 13464 9450 13676 9466
rect 13452 9444 13676 9450
rect 13504 9438 13676 9444
rect 13452 9386 13504 9392
rect 13544 9376 13596 9382
rect 13544 9318 13596 9324
rect 13556 9042 13584 9318
rect 13544 9036 13596 9042
rect 13544 8978 13596 8984
rect 13360 8628 13412 8634
rect 13360 8570 13412 8576
rect 13268 8424 13320 8430
rect 13268 8366 13320 8372
rect 13280 8090 13308 8366
rect 13268 8084 13320 8090
rect 13268 8026 13320 8032
rect 13556 7886 13584 8978
rect 13648 8974 13676 9438
rect 13636 8968 13688 8974
rect 13636 8910 13688 8916
rect 13648 7954 13676 8910
rect 13740 8498 13768 10950
rect 14016 10674 14044 12174
rect 14200 11558 14228 12922
rect 15292 12912 15344 12918
rect 15292 12854 15344 12860
rect 14648 12164 14700 12170
rect 14648 12106 14700 12112
rect 14266 11996 14574 12005
rect 14266 11994 14272 11996
rect 14328 11994 14352 11996
rect 14408 11994 14432 11996
rect 14488 11994 14512 11996
rect 14568 11994 14574 11996
rect 14328 11942 14330 11994
rect 14510 11942 14512 11994
rect 14266 11940 14272 11942
rect 14328 11940 14352 11942
rect 14408 11940 14432 11942
rect 14488 11940 14512 11942
rect 14568 11940 14574 11942
rect 14266 11931 14574 11940
rect 14660 11898 14688 12106
rect 15304 11898 15332 12854
rect 15396 12782 15424 14486
rect 15476 14068 15528 14074
rect 15476 14010 15528 14016
rect 15384 12776 15436 12782
rect 15384 12718 15436 12724
rect 14648 11892 14700 11898
rect 14648 11834 14700 11840
rect 15292 11892 15344 11898
rect 15292 11834 15344 11840
rect 14188 11552 14240 11558
rect 14188 11494 14240 11500
rect 14832 11552 14884 11558
rect 14832 11494 14884 11500
rect 14844 11218 14872 11494
rect 14832 11212 14884 11218
rect 14832 11154 14884 11160
rect 14740 11144 14792 11150
rect 14740 11086 14792 11092
rect 14648 11008 14700 11014
rect 14648 10950 14700 10956
rect 14266 10908 14574 10917
rect 14266 10906 14272 10908
rect 14328 10906 14352 10908
rect 14408 10906 14432 10908
rect 14488 10906 14512 10908
rect 14568 10906 14574 10908
rect 14328 10854 14330 10906
rect 14510 10854 14512 10906
rect 14266 10852 14272 10854
rect 14328 10852 14352 10854
rect 14408 10852 14432 10854
rect 14488 10852 14512 10854
rect 14568 10852 14574 10854
rect 14266 10843 14574 10852
rect 14660 10742 14688 10950
rect 14648 10736 14700 10742
rect 14648 10678 14700 10684
rect 14004 10668 14056 10674
rect 14004 10610 14056 10616
rect 14752 10266 14780 11086
rect 14740 10260 14792 10266
rect 14740 10202 14792 10208
rect 14844 9926 14872 11154
rect 15200 11144 15252 11150
rect 15200 11086 15252 11092
rect 13820 9920 13872 9926
rect 13820 9862 13872 9868
rect 14832 9920 14884 9926
rect 14832 9862 14884 9868
rect 13832 8786 13860 9862
rect 14266 9820 14574 9829
rect 14266 9818 14272 9820
rect 14328 9818 14352 9820
rect 14408 9818 14432 9820
rect 14488 9818 14512 9820
rect 14568 9818 14574 9820
rect 14328 9766 14330 9818
rect 14510 9766 14512 9818
rect 14266 9764 14272 9766
rect 14328 9764 14352 9766
rect 14408 9764 14432 9766
rect 14488 9764 14512 9766
rect 14568 9764 14574 9766
rect 14266 9755 14574 9764
rect 13912 9648 13964 9654
rect 13912 9590 13964 9596
rect 13924 9178 13952 9590
rect 14844 9586 14872 9862
rect 14740 9580 14792 9586
rect 14740 9522 14792 9528
rect 14832 9580 14884 9586
rect 14832 9522 14884 9528
rect 14648 9376 14700 9382
rect 14648 9318 14700 9324
rect 13912 9172 13964 9178
rect 13912 9114 13964 9120
rect 13924 8906 13952 9114
rect 13912 8900 13964 8906
rect 13912 8842 13964 8848
rect 14004 8832 14056 8838
rect 14002 8800 14004 8809
rect 14056 8800 14058 8809
rect 13832 8758 13952 8786
rect 13728 8492 13780 8498
rect 13728 8434 13780 8440
rect 13820 8356 13872 8362
rect 13820 8298 13872 8304
rect 13636 7948 13688 7954
rect 13636 7890 13688 7896
rect 13544 7880 13596 7886
rect 13544 7822 13596 7828
rect 13084 7744 13136 7750
rect 13084 7686 13136 7692
rect 13096 6662 13124 7686
rect 13832 7410 13860 8298
rect 13924 8022 13952 8758
rect 14002 8735 14058 8744
rect 14266 8732 14574 8741
rect 14266 8730 14272 8732
rect 14328 8730 14352 8732
rect 14408 8730 14432 8732
rect 14488 8730 14512 8732
rect 14568 8730 14574 8732
rect 14328 8678 14330 8730
rect 14510 8678 14512 8730
rect 14266 8676 14272 8678
rect 14328 8676 14352 8678
rect 14408 8676 14432 8678
rect 14488 8676 14512 8678
rect 14568 8676 14574 8678
rect 14266 8667 14574 8676
rect 14660 8566 14688 9318
rect 14752 9178 14780 9522
rect 15212 9450 15240 11086
rect 15384 10804 15436 10810
rect 15384 10746 15436 10752
rect 15396 10062 15424 10746
rect 15488 10198 15516 14010
rect 15764 13870 15792 15302
rect 15856 15162 15884 15370
rect 15844 15156 15896 15162
rect 15844 15098 15896 15104
rect 15856 14414 15884 15098
rect 16960 15026 16988 17070
rect 18705 16348 19013 16357
rect 18705 16346 18711 16348
rect 18767 16346 18791 16348
rect 18847 16346 18871 16348
rect 18927 16346 18951 16348
rect 19007 16346 19013 16348
rect 18767 16294 18769 16346
rect 18949 16294 18951 16346
rect 18705 16292 18711 16294
rect 18767 16292 18791 16294
rect 18847 16292 18871 16294
rect 18927 16292 18951 16294
rect 19007 16292 19013 16294
rect 18705 16283 19013 16292
rect 17132 15904 17184 15910
rect 17132 15846 17184 15852
rect 17144 15094 17172 15846
rect 18705 15260 19013 15269
rect 18705 15258 18711 15260
rect 18767 15258 18791 15260
rect 18847 15258 18871 15260
rect 18927 15258 18951 15260
rect 19007 15258 19013 15260
rect 18767 15206 18769 15258
rect 18949 15206 18951 15258
rect 18705 15204 18711 15206
rect 18767 15204 18791 15206
rect 18847 15204 18871 15206
rect 18927 15204 18951 15206
rect 19007 15204 19013 15206
rect 18705 15195 19013 15204
rect 17132 15088 17184 15094
rect 17132 15030 17184 15036
rect 16212 15020 16264 15026
rect 16212 14962 16264 14968
rect 16948 15020 17000 15026
rect 16948 14962 17000 14968
rect 16224 14482 16252 14962
rect 16960 14822 16988 14962
rect 16948 14816 17000 14822
rect 16948 14758 17000 14764
rect 16486 14716 16794 14725
rect 16486 14714 16492 14716
rect 16548 14714 16572 14716
rect 16628 14714 16652 14716
rect 16708 14714 16732 14716
rect 16788 14714 16794 14716
rect 16548 14662 16550 14714
rect 16730 14662 16732 14714
rect 16486 14660 16492 14662
rect 16548 14660 16572 14662
rect 16628 14660 16652 14662
rect 16708 14660 16732 14662
rect 16788 14660 16794 14662
rect 16486 14651 16794 14660
rect 16856 14612 16908 14618
rect 16856 14554 16908 14560
rect 16212 14476 16264 14482
rect 16212 14418 16264 14424
rect 16396 14476 16448 14482
rect 16396 14418 16448 14424
rect 15844 14408 15896 14414
rect 15844 14350 15896 14356
rect 15844 14272 15896 14278
rect 15844 14214 15896 14220
rect 15752 13864 15804 13870
rect 15752 13806 15804 13812
rect 15660 13184 15712 13190
rect 15660 13126 15712 13132
rect 15672 12850 15700 13126
rect 15660 12844 15712 12850
rect 15660 12786 15712 12792
rect 15752 12640 15804 12646
rect 15752 12582 15804 12588
rect 15764 11762 15792 12582
rect 15752 11756 15804 11762
rect 15752 11698 15804 11704
rect 15752 11620 15804 11626
rect 15752 11562 15804 11568
rect 15568 11008 15620 11014
rect 15568 10950 15620 10956
rect 15580 10266 15608 10950
rect 15568 10260 15620 10266
rect 15568 10202 15620 10208
rect 15476 10192 15528 10198
rect 15476 10134 15528 10140
rect 15764 10062 15792 11562
rect 15856 10674 15884 14214
rect 16408 13734 16436 14418
rect 16868 14006 16896 14554
rect 16960 14482 16988 14758
rect 16948 14476 17000 14482
rect 16948 14418 17000 14424
rect 17144 14278 17172 15030
rect 17316 15020 17368 15026
rect 17316 14962 17368 14968
rect 17328 14346 17356 14962
rect 17684 14952 17736 14958
rect 17684 14894 17736 14900
rect 17408 14476 17460 14482
rect 17408 14418 17460 14424
rect 17316 14340 17368 14346
rect 17316 14282 17368 14288
rect 16948 14272 17000 14278
rect 16948 14214 17000 14220
rect 17040 14272 17092 14278
rect 17040 14214 17092 14220
rect 17132 14272 17184 14278
rect 17132 14214 17184 14220
rect 16856 14000 16908 14006
rect 16856 13942 16908 13948
rect 16396 13728 16448 13734
rect 16396 13670 16448 13676
rect 16486 13628 16794 13637
rect 16486 13626 16492 13628
rect 16548 13626 16572 13628
rect 16628 13626 16652 13628
rect 16708 13626 16732 13628
rect 16788 13626 16794 13628
rect 16548 13574 16550 13626
rect 16730 13574 16732 13626
rect 16486 13572 16492 13574
rect 16548 13572 16572 13574
rect 16628 13572 16652 13574
rect 16708 13572 16732 13574
rect 16788 13572 16794 13574
rect 16486 13563 16794 13572
rect 16868 13326 16896 13942
rect 16856 13320 16908 13326
rect 16856 13262 16908 13268
rect 16580 13252 16632 13258
rect 16580 13194 16632 13200
rect 15936 12844 15988 12850
rect 15936 12786 15988 12792
rect 16120 12844 16172 12850
rect 16120 12786 16172 12792
rect 15948 12170 15976 12786
rect 16028 12776 16080 12782
rect 16028 12718 16080 12724
rect 15936 12164 15988 12170
rect 15936 12106 15988 12112
rect 15948 11898 15976 12106
rect 15936 11892 15988 11898
rect 15936 11834 15988 11840
rect 16040 11694 16068 12718
rect 16132 12442 16160 12786
rect 16592 12782 16620 13194
rect 16960 12850 16988 14214
rect 17052 13734 17080 14214
rect 17144 14074 17172 14214
rect 17132 14068 17184 14074
rect 17132 14010 17184 14016
rect 17420 13938 17448 14418
rect 17408 13932 17460 13938
rect 17408 13874 17460 13880
rect 17040 13728 17092 13734
rect 17040 13670 17092 13676
rect 17052 13394 17080 13670
rect 17040 13388 17092 13394
rect 17040 13330 17092 13336
rect 17420 13326 17448 13874
rect 17408 13320 17460 13326
rect 17408 13262 17460 13268
rect 17132 13252 17184 13258
rect 17132 13194 17184 13200
rect 16948 12844 17000 12850
rect 16948 12786 17000 12792
rect 16580 12776 16632 12782
rect 16580 12718 16632 12724
rect 16486 12540 16794 12549
rect 16486 12538 16492 12540
rect 16548 12538 16572 12540
rect 16628 12538 16652 12540
rect 16708 12538 16732 12540
rect 16788 12538 16794 12540
rect 16548 12486 16550 12538
rect 16730 12486 16732 12538
rect 16486 12484 16492 12486
rect 16548 12484 16572 12486
rect 16628 12484 16652 12486
rect 16708 12484 16732 12486
rect 16788 12484 16794 12486
rect 16486 12475 16794 12484
rect 16120 12436 16172 12442
rect 16960 12434 16988 12786
rect 16120 12378 16172 12384
rect 16868 12406 16988 12434
rect 16672 12232 16724 12238
rect 16672 12174 16724 12180
rect 16684 12102 16712 12174
rect 16868 12170 16896 12406
rect 17144 12238 17172 13194
rect 17500 13184 17552 13190
rect 17500 13126 17552 13132
rect 17224 12776 17276 12782
rect 17224 12718 17276 12724
rect 17132 12232 17184 12238
rect 17132 12174 17184 12180
rect 17236 12170 17264 12718
rect 16856 12164 16908 12170
rect 16856 12106 16908 12112
rect 17224 12164 17276 12170
rect 17224 12106 17276 12112
rect 16672 12096 16724 12102
rect 16672 12038 16724 12044
rect 16684 11762 16712 12038
rect 16396 11756 16448 11762
rect 16396 11698 16448 11704
rect 16672 11756 16724 11762
rect 16672 11698 16724 11704
rect 16028 11688 16080 11694
rect 16028 11630 16080 11636
rect 16212 11552 16264 11558
rect 16212 11494 16264 11500
rect 16120 11076 16172 11082
rect 16120 11018 16172 11024
rect 15844 10668 15896 10674
rect 15844 10610 15896 10616
rect 15936 10668 15988 10674
rect 15936 10610 15988 10616
rect 15948 10130 15976 10610
rect 16028 10464 16080 10470
rect 16028 10406 16080 10412
rect 15936 10124 15988 10130
rect 15936 10066 15988 10072
rect 15384 10056 15436 10062
rect 15384 9998 15436 10004
rect 15752 10056 15804 10062
rect 15752 9998 15804 10004
rect 15384 9920 15436 9926
rect 15384 9862 15436 9868
rect 15200 9444 15252 9450
rect 15200 9386 15252 9392
rect 15292 9376 15344 9382
rect 15292 9318 15344 9324
rect 15304 9178 15332 9318
rect 14740 9172 14792 9178
rect 14740 9114 14792 9120
rect 15292 9172 15344 9178
rect 15292 9114 15344 9120
rect 15016 8968 15068 8974
rect 15016 8910 15068 8916
rect 14648 8560 14700 8566
rect 14648 8502 14700 8508
rect 14004 8424 14056 8430
rect 14004 8366 14056 8372
rect 13912 8016 13964 8022
rect 13912 7958 13964 7964
rect 13544 7404 13596 7410
rect 13544 7346 13596 7352
rect 13820 7404 13872 7410
rect 13820 7346 13872 7352
rect 13556 6798 13584 7346
rect 13728 7200 13780 7206
rect 13728 7142 13780 7148
rect 13820 7200 13872 7206
rect 13820 7142 13872 7148
rect 13544 6792 13596 6798
rect 13544 6734 13596 6740
rect 13452 6724 13504 6730
rect 13452 6666 13504 6672
rect 13084 6656 13136 6662
rect 13084 6598 13136 6604
rect 11704 6316 11756 6322
rect 11704 6258 11756 6264
rect 11888 6316 11940 6322
rect 11888 6258 11940 6264
rect 12808 6316 12860 6322
rect 12808 6258 12860 6264
rect 13268 6316 13320 6322
rect 13268 6258 13320 6264
rect 11716 5370 11744 6258
rect 11796 6112 11848 6118
rect 11796 6054 11848 6060
rect 11704 5364 11756 5370
rect 11704 5306 11756 5312
rect 11808 5166 11836 6054
rect 11900 5914 11928 6258
rect 12047 6012 12355 6021
rect 12047 6010 12053 6012
rect 12109 6010 12133 6012
rect 12189 6010 12213 6012
rect 12269 6010 12293 6012
rect 12349 6010 12355 6012
rect 12109 5958 12111 6010
rect 12291 5958 12293 6010
rect 12047 5956 12053 5958
rect 12109 5956 12133 5958
rect 12189 5956 12213 5958
rect 12269 5956 12293 5958
rect 12349 5956 12355 5958
rect 12047 5947 12355 5956
rect 11888 5908 11940 5914
rect 11888 5850 11940 5856
rect 12820 5778 12848 6258
rect 12808 5772 12860 5778
rect 12808 5714 12860 5720
rect 11796 5160 11848 5166
rect 11796 5102 11848 5108
rect 11624 4950 11836 4978
rect 11612 4480 11664 4486
rect 11612 4422 11664 4428
rect 10692 4276 10744 4282
rect 10692 4218 10744 4224
rect 11152 4276 11204 4282
rect 11152 4218 11204 4224
rect 11624 4214 11652 4422
rect 11612 4208 11664 4214
rect 11612 4150 11664 4156
rect 11704 4072 11756 4078
rect 11704 4014 11756 4020
rect 9680 3528 9732 3534
rect 9680 3470 9732 3476
rect 11244 3528 11296 3534
rect 11244 3470 11296 3476
rect 10324 3392 10376 3398
rect 10324 3334 10376 3340
rect 11152 3392 11204 3398
rect 11152 3334 11204 3340
rect 9827 3292 10135 3301
rect 9827 3290 9833 3292
rect 9889 3290 9913 3292
rect 9969 3290 9993 3292
rect 10049 3290 10073 3292
rect 10129 3290 10135 3292
rect 9889 3238 9891 3290
rect 10071 3238 10073 3290
rect 9827 3236 9833 3238
rect 9889 3236 9913 3238
rect 9969 3236 9993 3238
rect 10049 3236 10073 3238
rect 10129 3236 10135 3238
rect 9827 3227 10135 3236
rect 10336 3058 10364 3334
rect 9312 3052 9364 3058
rect 9312 2994 9364 3000
rect 10324 3052 10376 3058
rect 10324 2994 10376 3000
rect 9220 2440 9272 2446
rect 9324 2428 9352 2994
rect 11060 2984 11112 2990
rect 11060 2926 11112 2932
rect 11072 2582 11100 2926
rect 11060 2576 11112 2582
rect 11060 2518 11112 2524
rect 9272 2400 9352 2428
rect 9220 2382 9272 2388
rect 7380 2372 7432 2378
rect 7380 2314 7432 2320
rect 9036 2372 9088 2378
rect 9036 2314 9088 2320
rect 1216 2304 1268 2310
rect 1216 2246 1268 2252
rect 3700 2304 3752 2310
rect 3700 2246 3752 2252
rect 6184 2304 6236 2310
rect 6184 2246 6236 2252
rect 8668 2304 8720 2310
rect 8668 2246 8720 2252
rect 1228 800 1256 2246
rect 3712 800 3740 2246
rect 5388 2204 5696 2213
rect 5388 2202 5394 2204
rect 5450 2202 5474 2204
rect 5530 2202 5554 2204
rect 5610 2202 5634 2204
rect 5690 2202 5696 2204
rect 5450 2150 5452 2202
rect 5632 2150 5634 2202
rect 5388 2148 5394 2150
rect 5450 2148 5474 2150
rect 5530 2148 5554 2150
rect 5610 2148 5634 2150
rect 5690 2148 5696 2150
rect 5388 2139 5696 2148
rect 6196 800 6224 2246
rect 8680 800 8708 2246
rect 9827 2204 10135 2213
rect 9827 2202 9833 2204
rect 9889 2202 9913 2204
rect 9969 2202 9993 2204
rect 10049 2202 10073 2204
rect 10129 2202 10135 2204
rect 9889 2150 9891 2202
rect 10071 2150 10073 2202
rect 9827 2148 9833 2150
rect 9889 2148 9913 2150
rect 9969 2148 9993 2150
rect 10049 2148 10073 2150
rect 10129 2148 10135 2150
rect 9827 2139 10135 2148
rect 11164 800 11192 3334
rect 11256 2650 11284 3470
rect 11336 3460 11388 3466
rect 11336 3402 11388 3408
rect 11348 3194 11376 3402
rect 11336 3188 11388 3194
rect 11336 3130 11388 3136
rect 11716 3058 11744 4014
rect 11808 3602 11836 4950
rect 12047 4924 12355 4933
rect 12047 4922 12053 4924
rect 12109 4922 12133 4924
rect 12189 4922 12213 4924
rect 12269 4922 12293 4924
rect 12349 4922 12355 4924
rect 12109 4870 12111 4922
rect 12291 4870 12293 4922
rect 12047 4868 12053 4870
rect 12109 4868 12133 4870
rect 12189 4868 12213 4870
rect 12269 4868 12293 4870
rect 12349 4868 12355 4870
rect 12047 4859 12355 4868
rect 12047 3836 12355 3845
rect 12047 3834 12053 3836
rect 12109 3834 12133 3836
rect 12189 3834 12213 3836
rect 12269 3834 12293 3836
rect 12349 3834 12355 3836
rect 12109 3782 12111 3834
rect 12291 3782 12293 3834
rect 12047 3780 12053 3782
rect 12109 3780 12133 3782
rect 12189 3780 12213 3782
rect 12269 3780 12293 3782
rect 12349 3780 12355 3782
rect 12047 3771 12355 3780
rect 11796 3596 11848 3602
rect 11796 3538 11848 3544
rect 11808 3398 11836 3538
rect 12820 3534 12848 5714
rect 13280 5710 13308 6258
rect 13464 6254 13492 6666
rect 13556 6254 13584 6734
rect 13452 6248 13504 6254
rect 13452 6190 13504 6196
rect 13544 6248 13596 6254
rect 13544 6190 13596 6196
rect 13464 6118 13492 6190
rect 13452 6112 13504 6118
rect 13452 6054 13504 6060
rect 13556 5710 13584 6190
rect 13740 6186 13768 7142
rect 13832 6866 13860 7142
rect 14016 6866 14044 8366
rect 15028 8362 15056 8910
rect 15396 8838 15424 9862
rect 15764 9042 15792 9998
rect 15934 9616 15990 9625
rect 15934 9551 15936 9560
rect 15988 9551 15990 9560
rect 15936 9522 15988 9528
rect 16040 9178 16068 10406
rect 16028 9172 16080 9178
rect 16028 9114 16080 9120
rect 16132 9110 16160 11018
rect 16120 9104 16172 9110
rect 16120 9046 16172 9052
rect 15752 9036 15804 9042
rect 15752 8978 15804 8984
rect 15108 8832 15160 8838
rect 15108 8774 15160 8780
rect 15384 8832 15436 8838
rect 15384 8774 15436 8780
rect 15016 8356 15068 8362
rect 15016 8298 15068 8304
rect 14266 7644 14574 7653
rect 14266 7642 14272 7644
rect 14328 7642 14352 7644
rect 14408 7642 14432 7644
rect 14488 7642 14512 7644
rect 14568 7642 14574 7644
rect 14328 7590 14330 7642
rect 14510 7590 14512 7642
rect 14266 7588 14272 7590
rect 14328 7588 14352 7590
rect 14408 7588 14432 7590
rect 14488 7588 14512 7590
rect 14568 7588 14574 7590
rect 14266 7579 14574 7588
rect 15120 7290 15148 8774
rect 16224 8498 16252 11494
rect 16408 11150 16436 11698
rect 16486 11452 16794 11461
rect 16486 11450 16492 11452
rect 16548 11450 16572 11452
rect 16628 11450 16652 11452
rect 16708 11450 16732 11452
rect 16788 11450 16794 11452
rect 16548 11398 16550 11450
rect 16730 11398 16732 11450
rect 16486 11396 16492 11398
rect 16548 11396 16572 11398
rect 16628 11396 16652 11398
rect 16708 11396 16732 11398
rect 16788 11396 16794 11398
rect 16486 11387 16794 11396
rect 16868 11218 16896 12106
rect 17040 12096 17092 12102
rect 17040 12038 17092 12044
rect 16948 11348 17000 11354
rect 16948 11290 17000 11296
rect 16856 11212 16908 11218
rect 16856 11154 16908 11160
rect 16396 11144 16448 11150
rect 16672 11144 16724 11150
rect 16448 11092 16620 11098
rect 16396 11086 16620 11092
rect 16672 11086 16724 11092
rect 16408 11070 16620 11086
rect 16396 10736 16448 10742
rect 16396 10678 16448 10684
rect 16408 10554 16436 10678
rect 16592 10674 16620 11070
rect 16580 10668 16632 10674
rect 16580 10610 16632 10616
rect 16684 10554 16712 11086
rect 16408 10526 16712 10554
rect 16212 8492 16264 8498
rect 16212 8434 16264 8440
rect 16408 8294 16436 10526
rect 16856 10464 16908 10470
rect 16856 10406 16908 10412
rect 16486 10364 16794 10373
rect 16486 10362 16492 10364
rect 16548 10362 16572 10364
rect 16628 10362 16652 10364
rect 16708 10362 16732 10364
rect 16788 10362 16794 10364
rect 16548 10310 16550 10362
rect 16730 10310 16732 10362
rect 16486 10308 16492 10310
rect 16548 10308 16572 10310
rect 16628 10308 16652 10310
rect 16708 10308 16732 10310
rect 16788 10308 16794 10310
rect 16486 10299 16794 10308
rect 16764 9580 16816 9586
rect 16868 9568 16896 10406
rect 16960 9654 16988 11290
rect 17052 11150 17080 12038
rect 17040 11144 17092 11150
rect 17040 11086 17092 11092
rect 17132 11076 17184 11082
rect 17132 11018 17184 11024
rect 17144 10810 17172 11018
rect 17236 11014 17264 12106
rect 17512 11558 17540 13126
rect 17592 11756 17644 11762
rect 17592 11698 17644 11704
rect 17500 11552 17552 11558
rect 17500 11494 17552 11500
rect 17316 11280 17368 11286
rect 17316 11222 17368 11228
rect 17224 11008 17276 11014
rect 17224 10950 17276 10956
rect 17132 10804 17184 10810
rect 17132 10746 17184 10752
rect 17040 10600 17092 10606
rect 17040 10542 17092 10548
rect 16948 9648 17000 9654
rect 16948 9590 17000 9596
rect 16816 9540 16896 9568
rect 16764 9522 16816 9528
rect 16948 9376 17000 9382
rect 16948 9318 17000 9324
rect 16486 9276 16794 9285
rect 16486 9274 16492 9276
rect 16548 9274 16572 9276
rect 16628 9274 16652 9276
rect 16708 9274 16732 9276
rect 16788 9274 16794 9276
rect 16548 9222 16550 9274
rect 16730 9222 16732 9274
rect 16486 9220 16492 9222
rect 16548 9220 16572 9222
rect 16628 9220 16652 9222
rect 16708 9220 16732 9222
rect 16788 9220 16794 9222
rect 16486 9211 16794 9220
rect 16960 8974 16988 9318
rect 17052 9178 17080 10542
rect 17144 10062 17172 10746
rect 17236 10606 17264 10950
rect 17328 10690 17356 11222
rect 17408 11212 17460 11218
rect 17408 11154 17460 11160
rect 17420 10810 17448 11154
rect 17604 11150 17632 11698
rect 17696 11558 17724 14894
rect 18705 14172 19013 14181
rect 18705 14170 18711 14172
rect 18767 14170 18791 14172
rect 18847 14170 18871 14172
rect 18927 14170 18951 14172
rect 19007 14170 19013 14172
rect 18767 14118 18769 14170
rect 18949 14118 18951 14170
rect 18705 14116 18711 14118
rect 18767 14116 18791 14118
rect 18847 14116 18871 14118
rect 18927 14116 18951 14118
rect 19007 14116 19013 14118
rect 18705 14107 19013 14116
rect 17960 14068 18012 14074
rect 17960 14010 18012 14016
rect 17776 14000 17828 14006
rect 17776 13942 17828 13948
rect 17788 12442 17816 13942
rect 17972 13326 18000 14010
rect 18052 13864 18104 13870
rect 18052 13806 18104 13812
rect 18064 13530 18092 13806
rect 18052 13524 18104 13530
rect 18052 13466 18104 13472
rect 17960 13320 18012 13326
rect 17960 13262 18012 13268
rect 18705 13084 19013 13093
rect 18705 13082 18711 13084
rect 18767 13082 18791 13084
rect 18847 13082 18871 13084
rect 18927 13082 18951 13084
rect 19007 13082 19013 13084
rect 18767 13030 18769 13082
rect 18949 13030 18951 13082
rect 18705 13028 18711 13030
rect 18767 13028 18791 13030
rect 18847 13028 18871 13030
rect 18927 13028 18951 13030
rect 19007 13028 19013 13030
rect 18705 13019 19013 13028
rect 17776 12436 17828 12442
rect 17776 12378 17828 12384
rect 17684 11552 17736 11558
rect 17684 11494 17736 11500
rect 17696 11354 17724 11494
rect 17684 11348 17736 11354
rect 17684 11290 17736 11296
rect 17592 11144 17644 11150
rect 17592 11086 17644 11092
rect 17500 11076 17552 11082
rect 17500 11018 17552 11024
rect 17408 10804 17460 10810
rect 17408 10746 17460 10752
rect 17512 10742 17540 11018
rect 17500 10736 17552 10742
rect 17328 10662 17448 10690
rect 17500 10678 17552 10684
rect 17224 10600 17276 10606
rect 17224 10542 17276 10548
rect 17132 10056 17184 10062
rect 17132 9998 17184 10004
rect 17316 9988 17368 9994
rect 17316 9930 17368 9936
rect 17040 9172 17092 9178
rect 17040 9114 17092 9120
rect 17328 9110 17356 9930
rect 17420 9926 17448 10662
rect 17512 10266 17540 10678
rect 17604 10674 17632 11086
rect 17592 10668 17644 10674
rect 17592 10610 17644 10616
rect 17500 10260 17552 10266
rect 17500 10202 17552 10208
rect 17604 10062 17632 10610
rect 17696 10470 17724 11290
rect 17684 10464 17736 10470
rect 17684 10406 17736 10412
rect 17788 10418 17816 12378
rect 17960 12096 18012 12102
rect 17960 12038 18012 12044
rect 17972 11762 18000 12038
rect 18705 11996 19013 12005
rect 18705 11994 18711 11996
rect 18767 11994 18791 11996
rect 18847 11994 18871 11996
rect 18927 11994 18951 11996
rect 19007 11994 19013 11996
rect 18767 11942 18769 11994
rect 18949 11942 18951 11994
rect 18705 11940 18711 11942
rect 18767 11940 18791 11942
rect 18847 11940 18871 11942
rect 18927 11940 18951 11942
rect 19007 11940 19013 11942
rect 18705 11931 19013 11940
rect 17960 11756 18012 11762
rect 17960 11698 18012 11704
rect 17972 11218 18000 11698
rect 17960 11212 18012 11218
rect 17960 11154 18012 11160
rect 17972 10690 18000 11154
rect 18705 10908 19013 10917
rect 18705 10906 18711 10908
rect 18767 10906 18791 10908
rect 18847 10906 18871 10908
rect 18927 10906 18951 10908
rect 19007 10906 19013 10908
rect 18767 10854 18769 10906
rect 18949 10854 18951 10906
rect 18705 10852 18711 10854
rect 18767 10852 18791 10854
rect 18847 10852 18871 10854
rect 18927 10852 18951 10854
rect 19007 10852 19013 10854
rect 18705 10843 19013 10852
rect 17972 10662 18092 10690
rect 18064 10606 18092 10662
rect 18052 10600 18104 10606
rect 18052 10542 18104 10548
rect 17696 10130 17724 10406
rect 17788 10390 17908 10418
rect 17880 10266 17908 10390
rect 17776 10260 17828 10266
rect 17776 10202 17828 10208
rect 17868 10260 17920 10266
rect 17868 10202 17920 10208
rect 17684 10124 17736 10130
rect 17684 10066 17736 10072
rect 17500 10056 17552 10062
rect 17500 9998 17552 10004
rect 17592 10056 17644 10062
rect 17592 9998 17644 10004
rect 17408 9920 17460 9926
rect 17408 9862 17460 9868
rect 17512 9586 17540 9998
rect 17592 9920 17644 9926
rect 17592 9862 17644 9868
rect 17500 9580 17552 9586
rect 17500 9522 17552 9528
rect 17316 9104 17368 9110
rect 17316 9046 17368 9052
rect 16948 8968 17000 8974
rect 16948 8910 17000 8916
rect 17132 8968 17184 8974
rect 17132 8910 17184 8916
rect 17040 8832 17092 8838
rect 17040 8774 17092 8780
rect 16856 8492 16908 8498
rect 16856 8434 16908 8440
rect 16396 8288 16448 8294
rect 16396 8230 16448 8236
rect 16486 8188 16794 8197
rect 16486 8186 16492 8188
rect 16548 8186 16572 8188
rect 16628 8186 16652 8188
rect 16708 8186 16732 8188
rect 16788 8186 16794 8188
rect 16548 8134 16550 8186
rect 16730 8134 16732 8186
rect 16486 8132 16492 8134
rect 16548 8132 16572 8134
rect 16628 8132 16652 8134
rect 16708 8132 16732 8134
rect 16788 8132 16794 8134
rect 16486 8123 16794 8132
rect 15844 7948 15896 7954
rect 15844 7890 15896 7896
rect 15856 7546 15884 7890
rect 16868 7886 16896 8434
rect 16856 7880 16908 7886
rect 16856 7822 16908 7828
rect 16028 7812 16080 7818
rect 16028 7754 16080 7760
rect 16948 7812 17000 7818
rect 16948 7754 17000 7760
rect 15936 7744 15988 7750
rect 15936 7686 15988 7692
rect 15844 7540 15896 7546
rect 15844 7482 15896 7488
rect 15856 7342 15884 7482
rect 15948 7426 15976 7686
rect 16040 7546 16068 7754
rect 16028 7540 16080 7546
rect 16028 7482 16080 7488
rect 15948 7398 16068 7426
rect 15200 7336 15252 7342
rect 15120 7284 15200 7290
rect 15120 7278 15252 7284
rect 15844 7336 15896 7342
rect 15844 7278 15896 7284
rect 15120 7262 15240 7278
rect 13820 6860 13872 6866
rect 13820 6802 13872 6808
rect 14004 6860 14056 6866
rect 14004 6802 14056 6808
rect 13728 6180 13780 6186
rect 13728 6122 13780 6128
rect 13084 5704 13136 5710
rect 13084 5646 13136 5652
rect 13268 5704 13320 5710
rect 13268 5646 13320 5652
rect 13544 5704 13596 5710
rect 13544 5646 13596 5652
rect 13096 4554 13124 5646
rect 13280 5030 13308 5646
rect 13268 5024 13320 5030
rect 13268 4966 13320 4972
rect 13280 4690 13308 4966
rect 13740 4758 13768 6122
rect 14016 5234 14044 6802
rect 14648 6724 14700 6730
rect 14648 6666 14700 6672
rect 14266 6556 14574 6565
rect 14266 6554 14272 6556
rect 14328 6554 14352 6556
rect 14408 6554 14432 6556
rect 14488 6554 14512 6556
rect 14568 6554 14574 6556
rect 14328 6502 14330 6554
rect 14510 6502 14512 6554
rect 14266 6500 14272 6502
rect 14328 6500 14352 6502
rect 14408 6500 14432 6502
rect 14488 6500 14512 6502
rect 14568 6500 14574 6502
rect 14266 6491 14574 6500
rect 14660 5914 14688 6666
rect 14648 5908 14700 5914
rect 14648 5850 14700 5856
rect 14648 5704 14700 5710
rect 14648 5646 14700 5652
rect 14188 5568 14240 5574
rect 14188 5510 14240 5516
rect 14200 5370 14228 5510
rect 14266 5468 14574 5477
rect 14266 5466 14272 5468
rect 14328 5466 14352 5468
rect 14408 5466 14432 5468
rect 14488 5466 14512 5468
rect 14568 5466 14574 5468
rect 14328 5414 14330 5466
rect 14510 5414 14512 5466
rect 14266 5412 14272 5414
rect 14328 5412 14352 5414
rect 14408 5412 14432 5414
rect 14488 5412 14512 5414
rect 14568 5412 14574 5414
rect 14266 5403 14574 5412
rect 14188 5364 14240 5370
rect 14188 5306 14240 5312
rect 14004 5228 14056 5234
rect 14004 5170 14056 5176
rect 13728 4752 13780 4758
rect 13728 4694 13780 4700
rect 13268 4684 13320 4690
rect 13268 4626 13320 4632
rect 13084 4548 13136 4554
rect 13084 4490 13136 4496
rect 14016 4146 14044 5170
rect 14200 4826 14228 5306
rect 14188 4820 14240 4826
rect 14188 4762 14240 4768
rect 14660 4690 14688 5646
rect 14648 4684 14700 4690
rect 14648 4626 14700 4632
rect 14266 4380 14574 4389
rect 14266 4378 14272 4380
rect 14328 4378 14352 4380
rect 14408 4378 14432 4380
rect 14488 4378 14512 4380
rect 14568 4378 14574 4380
rect 14328 4326 14330 4378
rect 14510 4326 14512 4378
rect 14266 4324 14272 4326
rect 14328 4324 14352 4326
rect 14408 4324 14432 4326
rect 14488 4324 14512 4326
rect 14568 4324 14574 4326
rect 14266 4315 14574 4324
rect 14660 4282 14688 4626
rect 14648 4276 14700 4282
rect 14648 4218 14700 4224
rect 14004 4140 14056 4146
rect 14004 4082 14056 4088
rect 13268 3732 13320 3738
rect 13268 3674 13320 3680
rect 12992 3664 13044 3670
rect 12992 3606 13044 3612
rect 13004 3534 13032 3606
rect 13280 3534 13308 3674
rect 13728 3596 13780 3602
rect 13728 3538 13780 3544
rect 12808 3528 12860 3534
rect 12808 3470 12860 3476
rect 12992 3528 13044 3534
rect 12992 3470 13044 3476
rect 13268 3528 13320 3534
rect 13268 3470 13320 3476
rect 13452 3528 13504 3534
rect 13452 3470 13504 3476
rect 11796 3392 11848 3398
rect 11796 3334 11848 3340
rect 12716 3392 12768 3398
rect 12716 3334 12768 3340
rect 11704 3052 11756 3058
rect 11704 2994 11756 3000
rect 11244 2644 11296 2650
rect 11244 2586 11296 2592
rect 11716 2446 11744 2994
rect 11808 2650 11836 3334
rect 12047 2748 12355 2757
rect 12047 2746 12053 2748
rect 12109 2746 12133 2748
rect 12189 2746 12213 2748
rect 12269 2746 12293 2748
rect 12349 2746 12355 2748
rect 12109 2694 12111 2746
rect 12291 2694 12293 2746
rect 12047 2692 12053 2694
rect 12109 2692 12133 2694
rect 12189 2692 12213 2694
rect 12269 2692 12293 2694
rect 12349 2692 12355 2694
rect 12047 2683 12355 2692
rect 11796 2644 11848 2650
rect 11796 2586 11848 2592
rect 11704 2440 11756 2446
rect 11704 2382 11756 2388
rect 12728 2378 12756 3334
rect 13464 3194 13492 3470
rect 13636 3392 13688 3398
rect 13636 3334 13688 3340
rect 13452 3188 13504 3194
rect 13452 3130 13504 3136
rect 12716 2372 12768 2378
rect 12716 2314 12768 2320
rect 13648 800 13676 3334
rect 13740 2650 13768 3538
rect 14016 3058 14044 4082
rect 15120 3738 15148 7262
rect 16040 6866 16068 7398
rect 16120 7404 16172 7410
rect 16120 7346 16172 7352
rect 16132 7002 16160 7346
rect 16486 7100 16794 7109
rect 16486 7098 16492 7100
rect 16548 7098 16572 7100
rect 16628 7098 16652 7100
rect 16708 7098 16732 7100
rect 16788 7098 16794 7100
rect 16548 7046 16550 7098
rect 16730 7046 16732 7098
rect 16486 7044 16492 7046
rect 16548 7044 16572 7046
rect 16628 7044 16652 7046
rect 16708 7044 16732 7046
rect 16788 7044 16794 7046
rect 16486 7035 16794 7044
rect 16120 6996 16172 7002
rect 16120 6938 16172 6944
rect 16028 6860 16080 6866
rect 16028 6802 16080 6808
rect 15936 6792 15988 6798
rect 15936 6734 15988 6740
rect 15660 6656 15712 6662
rect 15660 6598 15712 6604
rect 15672 6186 15700 6598
rect 15752 6248 15804 6254
rect 15752 6190 15804 6196
rect 15660 6180 15712 6186
rect 15660 6122 15712 6128
rect 15764 5710 15792 6190
rect 15948 5914 15976 6734
rect 15936 5908 15988 5914
rect 15936 5850 15988 5856
rect 15752 5704 15804 5710
rect 15752 5646 15804 5652
rect 16040 5642 16068 6802
rect 16132 6458 16160 6938
rect 16396 6792 16448 6798
rect 16396 6734 16448 6740
rect 16120 6452 16172 6458
rect 16120 6394 16172 6400
rect 16212 6112 16264 6118
rect 16212 6054 16264 6060
rect 16028 5636 16080 5642
rect 16028 5578 16080 5584
rect 16040 5234 16068 5578
rect 16224 5574 16252 6054
rect 16408 5658 16436 6734
rect 16960 6474 16988 7754
rect 17052 6662 17080 8774
rect 17144 8566 17172 8910
rect 17224 8628 17276 8634
rect 17224 8570 17276 8576
rect 17132 8560 17184 8566
rect 17132 8502 17184 8508
rect 17132 7744 17184 7750
rect 17132 7686 17184 7692
rect 17144 6798 17172 7686
rect 17236 7546 17264 8570
rect 17328 8362 17356 9046
rect 17500 9036 17552 9042
rect 17500 8978 17552 8984
rect 17316 8356 17368 8362
rect 17316 8298 17368 8304
rect 17408 8288 17460 8294
rect 17408 8230 17460 8236
rect 17224 7540 17276 7546
rect 17224 7482 17276 7488
rect 17420 7342 17448 8230
rect 17512 8090 17540 8978
rect 17604 8906 17632 9862
rect 17788 9654 17816 10202
rect 17776 9648 17828 9654
rect 17776 9590 17828 9596
rect 17776 9172 17828 9178
rect 17776 9114 17828 9120
rect 17684 8968 17736 8974
rect 17684 8910 17736 8916
rect 17592 8900 17644 8906
rect 17592 8842 17644 8848
rect 17604 8498 17632 8842
rect 17592 8492 17644 8498
rect 17592 8434 17644 8440
rect 17696 8106 17724 8910
rect 17788 8430 17816 9114
rect 17776 8424 17828 8430
rect 17776 8366 17828 8372
rect 17500 8084 17552 8090
rect 17500 8026 17552 8032
rect 17604 8078 17724 8106
rect 17408 7336 17460 7342
rect 17408 7278 17460 7284
rect 17604 7206 17632 8078
rect 17880 7970 17908 10202
rect 18064 10062 18092 10542
rect 18144 10464 18196 10470
rect 18144 10406 18196 10412
rect 18052 10056 18104 10062
rect 18052 9998 18104 10004
rect 18156 9518 18184 10406
rect 18705 9820 19013 9829
rect 18705 9818 18711 9820
rect 18767 9818 18791 9820
rect 18847 9818 18871 9820
rect 18927 9818 18951 9820
rect 19007 9818 19013 9820
rect 18767 9766 18769 9818
rect 18949 9766 18951 9818
rect 18705 9764 18711 9766
rect 18767 9764 18791 9766
rect 18847 9764 18871 9766
rect 18927 9764 18951 9766
rect 19007 9764 19013 9766
rect 18705 9755 19013 9764
rect 18144 9512 18196 9518
rect 18144 9454 18196 9460
rect 18052 9444 18104 9450
rect 18052 9386 18104 9392
rect 18064 8974 18092 9386
rect 18052 8968 18104 8974
rect 18052 8910 18104 8916
rect 17696 7942 17908 7970
rect 18064 7954 18092 8910
rect 18052 7948 18104 7954
rect 17592 7200 17644 7206
rect 17592 7142 17644 7148
rect 17224 6996 17276 7002
rect 17224 6938 17276 6944
rect 17132 6792 17184 6798
rect 17132 6734 17184 6740
rect 17040 6656 17092 6662
rect 17040 6598 17092 6604
rect 16960 6446 17080 6474
rect 17052 6322 17080 6446
rect 16856 6316 16908 6322
rect 16856 6258 16908 6264
rect 17040 6316 17092 6322
rect 17040 6258 17092 6264
rect 16486 6012 16794 6021
rect 16486 6010 16492 6012
rect 16548 6010 16572 6012
rect 16628 6010 16652 6012
rect 16708 6010 16732 6012
rect 16788 6010 16794 6012
rect 16548 5958 16550 6010
rect 16730 5958 16732 6010
rect 16486 5956 16492 5958
rect 16548 5956 16572 5958
rect 16628 5956 16652 5958
rect 16708 5956 16732 5958
rect 16788 5956 16794 5958
rect 16486 5947 16794 5956
rect 16316 5630 16436 5658
rect 16316 5574 16344 5630
rect 16212 5568 16264 5574
rect 16212 5510 16264 5516
rect 16304 5568 16356 5574
rect 16304 5510 16356 5516
rect 15844 5228 15896 5234
rect 15844 5170 15896 5176
rect 16028 5228 16080 5234
rect 16028 5170 16080 5176
rect 15856 4826 15884 5170
rect 15936 5024 15988 5030
rect 15936 4966 15988 4972
rect 15844 4820 15896 4826
rect 15844 4762 15896 4768
rect 15948 4758 15976 4966
rect 16040 4758 16068 5170
rect 15936 4752 15988 4758
rect 15936 4694 15988 4700
rect 16028 4752 16080 4758
rect 16028 4694 16080 4700
rect 16224 4554 16252 5510
rect 16212 4548 16264 4554
rect 16212 4490 16264 4496
rect 16316 4146 16344 5510
rect 16486 4924 16794 4933
rect 16486 4922 16492 4924
rect 16548 4922 16572 4924
rect 16628 4922 16652 4924
rect 16708 4922 16732 4924
rect 16788 4922 16794 4924
rect 16548 4870 16550 4922
rect 16730 4870 16732 4922
rect 16486 4868 16492 4870
rect 16548 4868 16572 4870
rect 16628 4868 16652 4870
rect 16708 4868 16732 4870
rect 16788 4868 16794 4870
rect 16486 4859 16794 4868
rect 16396 4548 16448 4554
rect 16396 4490 16448 4496
rect 16408 4298 16436 4490
rect 16488 4480 16540 4486
rect 16540 4428 16620 4434
rect 16488 4422 16620 4428
rect 16500 4406 16620 4422
rect 16408 4270 16528 4298
rect 16304 4140 16356 4146
rect 16304 4082 16356 4088
rect 16500 4078 16528 4270
rect 16592 4146 16620 4406
rect 16580 4140 16632 4146
rect 16580 4082 16632 4088
rect 16488 4072 16540 4078
rect 16488 4014 16540 4020
rect 16486 3836 16794 3845
rect 16486 3834 16492 3836
rect 16548 3834 16572 3836
rect 16628 3834 16652 3836
rect 16708 3834 16732 3836
rect 16788 3834 16794 3836
rect 16548 3782 16550 3834
rect 16730 3782 16732 3834
rect 16486 3780 16492 3782
rect 16548 3780 16572 3782
rect 16628 3780 16652 3782
rect 16708 3780 16732 3782
rect 16788 3780 16794 3782
rect 16486 3771 16794 3780
rect 16868 3738 16896 6258
rect 16948 6248 17000 6254
rect 16948 6190 17000 6196
rect 16960 5234 16988 6190
rect 17052 5370 17080 6258
rect 17040 5364 17092 5370
rect 17040 5306 17092 5312
rect 17144 5302 17172 6734
rect 17236 6662 17264 6938
rect 17224 6656 17276 6662
rect 17224 6598 17276 6604
rect 17236 6390 17264 6598
rect 17224 6384 17276 6390
rect 17224 6326 17276 6332
rect 17408 6180 17460 6186
rect 17408 6122 17460 6128
rect 17316 5908 17368 5914
rect 17316 5850 17368 5856
rect 17132 5296 17184 5302
rect 17132 5238 17184 5244
rect 16948 5228 17000 5234
rect 16948 5170 17000 5176
rect 17040 5228 17092 5234
rect 17040 5170 17092 5176
rect 16960 4826 16988 5170
rect 16948 4820 17000 4826
rect 16948 4762 17000 4768
rect 17052 4486 17080 5170
rect 17144 4554 17172 5238
rect 17224 4616 17276 4622
rect 17224 4558 17276 4564
rect 17132 4548 17184 4554
rect 17132 4490 17184 4496
rect 17040 4480 17092 4486
rect 17040 4422 17092 4428
rect 16948 4276 17000 4282
rect 16948 4218 17000 4224
rect 16960 3942 16988 4218
rect 16948 3936 17000 3942
rect 16948 3878 17000 3884
rect 15108 3732 15160 3738
rect 15108 3674 15160 3680
rect 16580 3732 16632 3738
rect 16580 3674 16632 3680
rect 16856 3732 16908 3738
rect 16856 3674 16908 3680
rect 16592 3466 16620 3674
rect 16960 3466 16988 3878
rect 16580 3460 16632 3466
rect 16580 3402 16632 3408
rect 16948 3460 17000 3466
rect 16948 3402 17000 3408
rect 16120 3392 16172 3398
rect 16120 3334 16172 3340
rect 14266 3292 14574 3301
rect 14266 3290 14272 3292
rect 14328 3290 14352 3292
rect 14408 3290 14432 3292
rect 14488 3290 14512 3292
rect 14568 3290 14574 3292
rect 14328 3238 14330 3290
rect 14510 3238 14512 3290
rect 14266 3236 14272 3238
rect 14328 3236 14352 3238
rect 14408 3236 14432 3238
rect 14488 3236 14512 3238
rect 14568 3236 14574 3238
rect 14266 3227 14574 3236
rect 14004 3052 14056 3058
rect 14004 2994 14056 3000
rect 15752 3052 15804 3058
rect 15752 2994 15804 3000
rect 15936 3052 15988 3058
rect 15936 2994 15988 3000
rect 13728 2644 13780 2650
rect 13728 2586 13780 2592
rect 14016 2514 14044 2994
rect 15764 2514 15792 2994
rect 15948 2650 15976 2994
rect 15936 2644 15988 2650
rect 15936 2586 15988 2592
rect 14004 2508 14056 2514
rect 14004 2450 14056 2456
rect 15752 2508 15804 2514
rect 15752 2450 15804 2456
rect 14266 2204 14574 2213
rect 14266 2202 14272 2204
rect 14328 2202 14352 2204
rect 14408 2202 14432 2204
rect 14488 2202 14512 2204
rect 14568 2202 14574 2204
rect 14328 2150 14330 2202
rect 14510 2150 14512 2202
rect 14266 2148 14272 2150
rect 14328 2148 14352 2150
rect 14408 2148 14432 2150
rect 14488 2148 14512 2150
rect 14568 2148 14574 2150
rect 14266 2139 14574 2148
rect 16132 800 16160 3334
rect 16592 3126 16620 3402
rect 16580 3120 16632 3126
rect 16580 3062 16632 3068
rect 17052 3058 17080 4422
rect 17132 4208 17184 4214
rect 17132 4150 17184 4156
rect 17144 3466 17172 4150
rect 17132 3460 17184 3466
rect 17132 3402 17184 3408
rect 17236 3194 17264 4558
rect 17224 3188 17276 3194
rect 17224 3130 17276 3136
rect 17040 3052 17092 3058
rect 17040 2994 17092 3000
rect 16856 2848 16908 2854
rect 16856 2790 16908 2796
rect 16486 2748 16794 2757
rect 16486 2746 16492 2748
rect 16548 2746 16572 2748
rect 16628 2746 16652 2748
rect 16708 2746 16732 2748
rect 16788 2746 16794 2748
rect 16548 2694 16550 2746
rect 16730 2694 16732 2746
rect 16486 2692 16492 2694
rect 16548 2692 16572 2694
rect 16628 2692 16652 2694
rect 16708 2692 16732 2694
rect 16788 2692 16794 2694
rect 16486 2683 16794 2692
rect 16868 2446 16896 2790
rect 17052 2774 17080 2994
rect 16960 2746 17080 2774
rect 16960 2650 16988 2746
rect 16948 2644 17000 2650
rect 16948 2586 17000 2592
rect 17236 2582 17264 3130
rect 17328 3126 17356 5850
rect 17420 5642 17448 6122
rect 17592 5772 17644 5778
rect 17592 5714 17644 5720
rect 17408 5636 17460 5642
rect 17408 5578 17460 5584
rect 17420 5030 17448 5578
rect 17604 5302 17632 5714
rect 17696 5710 17724 7942
rect 18052 7890 18104 7896
rect 17776 7880 17828 7886
rect 18156 7868 18184 9454
rect 18236 8832 18288 8838
rect 18236 8774 18288 8780
rect 18248 8498 18276 8774
rect 18705 8732 19013 8741
rect 18705 8730 18711 8732
rect 18767 8730 18791 8732
rect 18847 8730 18871 8732
rect 18927 8730 18951 8732
rect 19007 8730 19013 8732
rect 18767 8678 18769 8730
rect 18949 8678 18951 8730
rect 18705 8676 18711 8678
rect 18767 8676 18791 8678
rect 18847 8676 18871 8678
rect 18927 8676 18951 8678
rect 19007 8676 19013 8678
rect 18705 8667 19013 8676
rect 18236 8492 18288 8498
rect 18236 8434 18288 8440
rect 18236 7880 18288 7886
rect 18156 7840 18236 7868
rect 17776 7822 17828 7828
rect 18236 7822 18288 7828
rect 17788 6458 17816 7822
rect 18144 7744 18196 7750
rect 18144 7686 18196 7692
rect 18052 7472 18104 7478
rect 18052 7414 18104 7420
rect 17960 7404 18012 7410
rect 17960 7346 18012 7352
rect 17868 7200 17920 7206
rect 17868 7142 17920 7148
rect 17880 6882 17908 7142
rect 17972 7002 18000 7346
rect 17960 6996 18012 7002
rect 17960 6938 18012 6944
rect 17880 6854 18000 6882
rect 17776 6452 17828 6458
rect 17776 6394 17828 6400
rect 17868 6316 17920 6322
rect 17868 6258 17920 6264
rect 17880 5914 17908 6258
rect 17972 5914 18000 6854
rect 18064 6458 18092 7414
rect 18052 6452 18104 6458
rect 18052 6394 18104 6400
rect 17868 5908 17920 5914
rect 17868 5850 17920 5856
rect 17960 5908 18012 5914
rect 17960 5850 18012 5856
rect 17684 5704 17736 5710
rect 17684 5646 17736 5652
rect 17972 5370 18000 5850
rect 17960 5364 18012 5370
rect 17960 5306 18012 5312
rect 17592 5296 17644 5302
rect 17592 5238 17644 5244
rect 17408 5024 17460 5030
rect 17408 4966 17460 4972
rect 17604 4282 17632 5238
rect 17776 5024 17828 5030
rect 17776 4966 17828 4972
rect 17788 4758 17816 4966
rect 18156 4826 18184 7686
rect 18248 7274 18276 7822
rect 18705 7644 19013 7653
rect 18705 7642 18711 7644
rect 18767 7642 18791 7644
rect 18847 7642 18871 7644
rect 18927 7642 18951 7644
rect 19007 7642 19013 7644
rect 18767 7590 18769 7642
rect 18949 7590 18951 7642
rect 18705 7588 18711 7590
rect 18767 7588 18791 7590
rect 18847 7588 18871 7590
rect 18927 7588 18951 7590
rect 19007 7588 19013 7590
rect 18705 7579 19013 7588
rect 18236 7268 18288 7274
rect 18236 7210 18288 7216
rect 18705 6556 19013 6565
rect 18705 6554 18711 6556
rect 18767 6554 18791 6556
rect 18847 6554 18871 6556
rect 18927 6554 18951 6556
rect 19007 6554 19013 6556
rect 18767 6502 18769 6554
rect 18949 6502 18951 6554
rect 18705 6500 18711 6502
rect 18767 6500 18791 6502
rect 18847 6500 18871 6502
rect 18927 6500 18951 6502
rect 19007 6500 19013 6502
rect 18705 6491 19013 6500
rect 18705 5468 19013 5477
rect 18705 5466 18711 5468
rect 18767 5466 18791 5468
rect 18847 5466 18871 5468
rect 18927 5466 18951 5468
rect 19007 5466 19013 5468
rect 18767 5414 18769 5466
rect 18949 5414 18951 5466
rect 18705 5412 18711 5414
rect 18767 5412 18791 5414
rect 18847 5412 18871 5414
rect 18927 5412 18951 5414
rect 19007 5412 19013 5414
rect 18705 5403 19013 5412
rect 18144 4820 18196 4826
rect 18144 4762 18196 4768
rect 17776 4752 17828 4758
rect 17776 4694 17828 4700
rect 18705 4380 19013 4389
rect 18705 4378 18711 4380
rect 18767 4378 18791 4380
rect 18847 4378 18871 4380
rect 18927 4378 18951 4380
rect 19007 4378 19013 4380
rect 18767 4326 18769 4378
rect 18949 4326 18951 4378
rect 18705 4324 18711 4326
rect 18767 4324 18791 4326
rect 18847 4324 18871 4326
rect 18927 4324 18951 4326
rect 19007 4324 19013 4326
rect 18705 4315 19013 4324
rect 17592 4276 17644 4282
rect 17592 4218 17644 4224
rect 17868 3936 17920 3942
rect 17868 3878 17920 3884
rect 17408 3392 17460 3398
rect 17408 3334 17460 3340
rect 17316 3120 17368 3126
rect 17316 3062 17368 3068
rect 17224 2576 17276 2582
rect 17224 2518 17276 2524
rect 17328 2446 17356 3062
rect 17420 2990 17448 3334
rect 17880 3126 17908 3878
rect 18144 3664 18196 3670
rect 18144 3606 18196 3612
rect 17868 3120 17920 3126
rect 17868 3062 17920 3068
rect 18156 3058 18184 3606
rect 18604 3392 18656 3398
rect 18604 3334 18656 3340
rect 18144 3052 18196 3058
rect 18144 2994 18196 3000
rect 17408 2984 17460 2990
rect 17408 2926 17460 2932
rect 18052 2848 18104 2854
rect 18052 2790 18104 2796
rect 16856 2440 16908 2446
rect 16856 2382 16908 2388
rect 17316 2440 17368 2446
rect 17316 2382 17368 2388
rect 18064 2378 18092 2790
rect 18052 2372 18104 2378
rect 18052 2314 18104 2320
rect 18616 800 18644 3334
rect 18705 3292 19013 3301
rect 18705 3290 18711 3292
rect 18767 3290 18791 3292
rect 18847 3290 18871 3292
rect 18927 3290 18951 3292
rect 19007 3290 19013 3292
rect 18767 3238 18769 3290
rect 18949 3238 18951 3290
rect 18705 3236 18711 3238
rect 18767 3236 18791 3238
rect 18847 3236 18871 3238
rect 18927 3236 18951 3238
rect 19007 3236 19013 3238
rect 18705 3227 19013 3236
rect 18705 2204 19013 2213
rect 18705 2202 18711 2204
rect 18767 2202 18791 2204
rect 18847 2202 18871 2204
rect 18927 2202 18951 2204
rect 19007 2202 19013 2204
rect 18767 2150 18769 2202
rect 18949 2150 18951 2202
rect 18705 2148 18711 2150
rect 18767 2148 18791 2150
rect 18847 2148 18871 2150
rect 18927 2148 18951 2150
rect 19007 2148 19013 2150
rect 18705 2139 19013 2148
rect 1214 0 1270 800
rect 3698 0 3754 800
rect 6182 0 6238 800
rect 8666 0 8722 800
rect 11150 0 11206 800
rect 13634 0 13690 800
rect 16118 0 16174 800
rect 18602 0 18658 800
<< via2 >>
rect 5394 17434 5450 17436
rect 5474 17434 5530 17436
rect 5554 17434 5610 17436
rect 5634 17434 5690 17436
rect 5394 17382 5440 17434
rect 5440 17382 5450 17434
rect 5474 17382 5504 17434
rect 5504 17382 5516 17434
rect 5516 17382 5530 17434
rect 5554 17382 5568 17434
rect 5568 17382 5580 17434
rect 5580 17382 5610 17434
rect 5634 17382 5644 17434
rect 5644 17382 5690 17434
rect 5394 17380 5450 17382
rect 5474 17380 5530 17382
rect 5554 17380 5610 17382
rect 5634 17380 5690 17382
rect 9833 17434 9889 17436
rect 9913 17434 9969 17436
rect 9993 17434 10049 17436
rect 10073 17434 10129 17436
rect 9833 17382 9879 17434
rect 9879 17382 9889 17434
rect 9913 17382 9943 17434
rect 9943 17382 9955 17434
rect 9955 17382 9969 17434
rect 9993 17382 10007 17434
rect 10007 17382 10019 17434
rect 10019 17382 10049 17434
rect 10073 17382 10083 17434
rect 10083 17382 10129 17434
rect 9833 17380 9889 17382
rect 9913 17380 9969 17382
rect 9993 17380 10049 17382
rect 10073 17380 10129 17382
rect 14272 17434 14328 17436
rect 14352 17434 14408 17436
rect 14432 17434 14488 17436
rect 14512 17434 14568 17436
rect 14272 17382 14318 17434
rect 14318 17382 14328 17434
rect 14352 17382 14382 17434
rect 14382 17382 14394 17434
rect 14394 17382 14408 17434
rect 14432 17382 14446 17434
rect 14446 17382 14458 17434
rect 14458 17382 14488 17434
rect 14512 17382 14522 17434
rect 14522 17382 14568 17434
rect 14272 17380 14328 17382
rect 14352 17380 14408 17382
rect 14432 17380 14488 17382
rect 14512 17380 14568 17382
rect 18711 17434 18767 17436
rect 18791 17434 18847 17436
rect 18871 17434 18927 17436
rect 18951 17434 19007 17436
rect 18711 17382 18757 17434
rect 18757 17382 18767 17434
rect 18791 17382 18821 17434
rect 18821 17382 18833 17434
rect 18833 17382 18847 17434
rect 18871 17382 18885 17434
rect 18885 17382 18897 17434
rect 18897 17382 18927 17434
rect 18951 17382 18961 17434
rect 18961 17382 19007 17434
rect 18711 17380 18767 17382
rect 18791 17380 18847 17382
rect 18871 17380 18927 17382
rect 18951 17380 19007 17382
rect 3175 16890 3231 16892
rect 3255 16890 3311 16892
rect 3335 16890 3391 16892
rect 3415 16890 3471 16892
rect 3175 16838 3221 16890
rect 3221 16838 3231 16890
rect 3255 16838 3285 16890
rect 3285 16838 3297 16890
rect 3297 16838 3311 16890
rect 3335 16838 3349 16890
rect 3349 16838 3361 16890
rect 3361 16838 3391 16890
rect 3415 16838 3425 16890
rect 3425 16838 3471 16890
rect 3175 16836 3231 16838
rect 3255 16836 3311 16838
rect 3335 16836 3391 16838
rect 3415 16836 3471 16838
rect 3175 15802 3231 15804
rect 3255 15802 3311 15804
rect 3335 15802 3391 15804
rect 3415 15802 3471 15804
rect 3175 15750 3221 15802
rect 3221 15750 3231 15802
rect 3255 15750 3285 15802
rect 3285 15750 3297 15802
rect 3297 15750 3311 15802
rect 3335 15750 3349 15802
rect 3349 15750 3361 15802
rect 3361 15750 3391 15802
rect 3415 15750 3425 15802
rect 3425 15750 3471 15802
rect 3175 15748 3231 15750
rect 3255 15748 3311 15750
rect 3335 15748 3391 15750
rect 3415 15748 3471 15750
rect 3175 14714 3231 14716
rect 3255 14714 3311 14716
rect 3335 14714 3391 14716
rect 3415 14714 3471 14716
rect 3175 14662 3221 14714
rect 3221 14662 3231 14714
rect 3255 14662 3285 14714
rect 3285 14662 3297 14714
rect 3297 14662 3311 14714
rect 3335 14662 3349 14714
rect 3349 14662 3361 14714
rect 3361 14662 3391 14714
rect 3415 14662 3425 14714
rect 3425 14662 3471 14714
rect 3175 14660 3231 14662
rect 3255 14660 3311 14662
rect 3335 14660 3391 14662
rect 3415 14660 3471 14662
rect 3175 13626 3231 13628
rect 3255 13626 3311 13628
rect 3335 13626 3391 13628
rect 3415 13626 3471 13628
rect 3175 13574 3221 13626
rect 3221 13574 3231 13626
rect 3255 13574 3285 13626
rect 3285 13574 3297 13626
rect 3297 13574 3311 13626
rect 3335 13574 3349 13626
rect 3349 13574 3361 13626
rect 3361 13574 3391 13626
rect 3415 13574 3425 13626
rect 3425 13574 3471 13626
rect 3175 13572 3231 13574
rect 3255 13572 3311 13574
rect 3335 13572 3391 13574
rect 3415 13572 3471 13574
rect 3175 12538 3231 12540
rect 3255 12538 3311 12540
rect 3335 12538 3391 12540
rect 3415 12538 3471 12540
rect 3175 12486 3221 12538
rect 3221 12486 3231 12538
rect 3255 12486 3285 12538
rect 3285 12486 3297 12538
rect 3297 12486 3311 12538
rect 3335 12486 3349 12538
rect 3349 12486 3361 12538
rect 3361 12486 3391 12538
rect 3415 12486 3425 12538
rect 3425 12486 3471 12538
rect 3175 12484 3231 12486
rect 3255 12484 3311 12486
rect 3335 12484 3391 12486
rect 3415 12484 3471 12486
rect 3175 11450 3231 11452
rect 3255 11450 3311 11452
rect 3335 11450 3391 11452
rect 3415 11450 3471 11452
rect 3175 11398 3221 11450
rect 3221 11398 3231 11450
rect 3255 11398 3285 11450
rect 3285 11398 3297 11450
rect 3297 11398 3311 11450
rect 3335 11398 3349 11450
rect 3349 11398 3361 11450
rect 3361 11398 3391 11450
rect 3415 11398 3425 11450
rect 3425 11398 3471 11450
rect 3175 11396 3231 11398
rect 3255 11396 3311 11398
rect 3335 11396 3391 11398
rect 3415 11396 3471 11398
rect 3175 10362 3231 10364
rect 3255 10362 3311 10364
rect 3335 10362 3391 10364
rect 3415 10362 3471 10364
rect 3175 10310 3221 10362
rect 3221 10310 3231 10362
rect 3255 10310 3285 10362
rect 3285 10310 3297 10362
rect 3297 10310 3311 10362
rect 3335 10310 3349 10362
rect 3349 10310 3361 10362
rect 3361 10310 3391 10362
rect 3415 10310 3425 10362
rect 3425 10310 3471 10362
rect 3175 10308 3231 10310
rect 3255 10308 3311 10310
rect 3335 10308 3391 10310
rect 3415 10308 3471 10310
rect 5394 16346 5450 16348
rect 5474 16346 5530 16348
rect 5554 16346 5610 16348
rect 5634 16346 5690 16348
rect 5394 16294 5440 16346
rect 5440 16294 5450 16346
rect 5474 16294 5504 16346
rect 5504 16294 5516 16346
rect 5516 16294 5530 16346
rect 5554 16294 5568 16346
rect 5568 16294 5580 16346
rect 5580 16294 5610 16346
rect 5634 16294 5644 16346
rect 5644 16294 5690 16346
rect 5394 16292 5450 16294
rect 5474 16292 5530 16294
rect 5554 16292 5610 16294
rect 5634 16292 5690 16294
rect 7614 16890 7670 16892
rect 7694 16890 7750 16892
rect 7774 16890 7830 16892
rect 7854 16890 7910 16892
rect 7614 16838 7660 16890
rect 7660 16838 7670 16890
rect 7694 16838 7724 16890
rect 7724 16838 7736 16890
rect 7736 16838 7750 16890
rect 7774 16838 7788 16890
rect 7788 16838 7800 16890
rect 7800 16838 7830 16890
rect 7854 16838 7864 16890
rect 7864 16838 7910 16890
rect 7614 16836 7670 16838
rect 7694 16836 7750 16838
rect 7774 16836 7830 16838
rect 7854 16836 7910 16838
rect 9833 16346 9889 16348
rect 9913 16346 9969 16348
rect 9993 16346 10049 16348
rect 10073 16346 10129 16348
rect 9833 16294 9879 16346
rect 9879 16294 9889 16346
rect 9913 16294 9943 16346
rect 9943 16294 9955 16346
rect 9955 16294 9969 16346
rect 9993 16294 10007 16346
rect 10007 16294 10019 16346
rect 10019 16294 10049 16346
rect 10073 16294 10083 16346
rect 10083 16294 10129 16346
rect 9833 16292 9889 16294
rect 9913 16292 9969 16294
rect 9993 16292 10049 16294
rect 10073 16292 10129 16294
rect 5394 15258 5450 15260
rect 5474 15258 5530 15260
rect 5554 15258 5610 15260
rect 5634 15258 5690 15260
rect 5394 15206 5440 15258
rect 5440 15206 5450 15258
rect 5474 15206 5504 15258
rect 5504 15206 5516 15258
rect 5516 15206 5530 15258
rect 5554 15206 5568 15258
rect 5568 15206 5580 15258
rect 5580 15206 5610 15258
rect 5634 15206 5644 15258
rect 5644 15206 5690 15258
rect 5394 15204 5450 15206
rect 5474 15204 5530 15206
rect 5554 15204 5610 15206
rect 5634 15204 5690 15206
rect 5394 14170 5450 14172
rect 5474 14170 5530 14172
rect 5554 14170 5610 14172
rect 5634 14170 5690 14172
rect 5394 14118 5440 14170
rect 5440 14118 5450 14170
rect 5474 14118 5504 14170
rect 5504 14118 5516 14170
rect 5516 14118 5530 14170
rect 5554 14118 5568 14170
rect 5568 14118 5580 14170
rect 5580 14118 5610 14170
rect 5634 14118 5644 14170
rect 5644 14118 5690 14170
rect 5394 14116 5450 14118
rect 5474 14116 5530 14118
rect 5554 14116 5610 14118
rect 5634 14116 5690 14118
rect 7614 15802 7670 15804
rect 7694 15802 7750 15804
rect 7774 15802 7830 15804
rect 7854 15802 7910 15804
rect 7614 15750 7660 15802
rect 7660 15750 7670 15802
rect 7694 15750 7724 15802
rect 7724 15750 7736 15802
rect 7736 15750 7750 15802
rect 7774 15750 7788 15802
rect 7788 15750 7800 15802
rect 7800 15750 7830 15802
rect 7854 15750 7864 15802
rect 7864 15750 7910 15802
rect 7614 15748 7670 15750
rect 7694 15748 7750 15750
rect 7774 15748 7830 15750
rect 7854 15748 7910 15750
rect 7614 14714 7670 14716
rect 7694 14714 7750 14716
rect 7774 14714 7830 14716
rect 7854 14714 7910 14716
rect 7614 14662 7660 14714
rect 7660 14662 7670 14714
rect 7694 14662 7724 14714
rect 7724 14662 7736 14714
rect 7736 14662 7750 14714
rect 7774 14662 7788 14714
rect 7788 14662 7800 14714
rect 7800 14662 7830 14714
rect 7854 14662 7864 14714
rect 7864 14662 7910 14714
rect 7614 14660 7670 14662
rect 7694 14660 7750 14662
rect 7774 14660 7830 14662
rect 7854 14660 7910 14662
rect 5394 13082 5450 13084
rect 5474 13082 5530 13084
rect 5554 13082 5610 13084
rect 5634 13082 5690 13084
rect 5394 13030 5440 13082
rect 5440 13030 5450 13082
rect 5474 13030 5504 13082
rect 5504 13030 5516 13082
rect 5516 13030 5530 13082
rect 5554 13030 5568 13082
rect 5568 13030 5580 13082
rect 5580 13030 5610 13082
rect 5634 13030 5644 13082
rect 5644 13030 5690 13082
rect 5394 13028 5450 13030
rect 5474 13028 5530 13030
rect 5554 13028 5610 13030
rect 5634 13028 5690 13030
rect 5394 11994 5450 11996
rect 5474 11994 5530 11996
rect 5554 11994 5610 11996
rect 5634 11994 5690 11996
rect 5394 11942 5440 11994
rect 5440 11942 5450 11994
rect 5474 11942 5504 11994
rect 5504 11942 5516 11994
rect 5516 11942 5530 11994
rect 5554 11942 5568 11994
rect 5568 11942 5580 11994
rect 5580 11942 5610 11994
rect 5634 11942 5644 11994
rect 5644 11942 5690 11994
rect 5394 11940 5450 11942
rect 5474 11940 5530 11942
rect 5554 11940 5610 11942
rect 5634 11940 5690 11942
rect 3175 9274 3231 9276
rect 3255 9274 3311 9276
rect 3335 9274 3391 9276
rect 3415 9274 3471 9276
rect 3175 9222 3221 9274
rect 3221 9222 3231 9274
rect 3255 9222 3285 9274
rect 3285 9222 3297 9274
rect 3297 9222 3311 9274
rect 3335 9222 3349 9274
rect 3349 9222 3361 9274
rect 3361 9222 3391 9274
rect 3415 9222 3425 9274
rect 3425 9222 3471 9274
rect 3175 9220 3231 9222
rect 3255 9220 3311 9222
rect 3335 9220 3391 9222
rect 3415 9220 3471 9222
rect 3175 8186 3231 8188
rect 3255 8186 3311 8188
rect 3335 8186 3391 8188
rect 3415 8186 3471 8188
rect 3175 8134 3221 8186
rect 3221 8134 3231 8186
rect 3255 8134 3285 8186
rect 3285 8134 3297 8186
rect 3297 8134 3311 8186
rect 3335 8134 3349 8186
rect 3349 8134 3361 8186
rect 3361 8134 3391 8186
rect 3415 8134 3425 8186
rect 3425 8134 3471 8186
rect 3175 8132 3231 8134
rect 3255 8132 3311 8134
rect 3335 8132 3391 8134
rect 3415 8132 3471 8134
rect 3175 7098 3231 7100
rect 3255 7098 3311 7100
rect 3335 7098 3391 7100
rect 3415 7098 3471 7100
rect 3175 7046 3221 7098
rect 3221 7046 3231 7098
rect 3255 7046 3285 7098
rect 3285 7046 3297 7098
rect 3297 7046 3311 7098
rect 3335 7046 3349 7098
rect 3349 7046 3361 7098
rect 3361 7046 3391 7098
rect 3415 7046 3425 7098
rect 3425 7046 3471 7098
rect 3175 7044 3231 7046
rect 3255 7044 3311 7046
rect 3335 7044 3391 7046
rect 3415 7044 3471 7046
rect 7614 13626 7670 13628
rect 7694 13626 7750 13628
rect 7774 13626 7830 13628
rect 7854 13626 7910 13628
rect 7614 13574 7660 13626
rect 7660 13574 7670 13626
rect 7694 13574 7724 13626
rect 7724 13574 7736 13626
rect 7736 13574 7750 13626
rect 7774 13574 7788 13626
rect 7788 13574 7800 13626
rect 7800 13574 7830 13626
rect 7854 13574 7864 13626
rect 7864 13574 7910 13626
rect 7614 13572 7670 13574
rect 7694 13572 7750 13574
rect 7774 13572 7830 13574
rect 7854 13572 7910 13574
rect 7010 12280 7066 12336
rect 5394 10906 5450 10908
rect 5474 10906 5530 10908
rect 5554 10906 5610 10908
rect 5634 10906 5690 10908
rect 5394 10854 5440 10906
rect 5440 10854 5450 10906
rect 5474 10854 5504 10906
rect 5504 10854 5516 10906
rect 5516 10854 5530 10906
rect 5554 10854 5568 10906
rect 5568 10854 5580 10906
rect 5580 10854 5610 10906
rect 5634 10854 5644 10906
rect 5644 10854 5690 10906
rect 5394 10852 5450 10854
rect 5474 10852 5530 10854
rect 5554 10852 5610 10854
rect 5634 10852 5690 10854
rect 5394 9818 5450 9820
rect 5474 9818 5530 9820
rect 5554 9818 5610 9820
rect 5634 9818 5690 9820
rect 5394 9766 5440 9818
rect 5440 9766 5450 9818
rect 5474 9766 5504 9818
rect 5504 9766 5516 9818
rect 5516 9766 5530 9818
rect 5554 9766 5568 9818
rect 5568 9766 5580 9818
rect 5580 9766 5610 9818
rect 5634 9766 5644 9818
rect 5644 9766 5690 9818
rect 5394 9764 5450 9766
rect 5474 9764 5530 9766
rect 5554 9764 5610 9766
rect 5634 9764 5690 9766
rect 3175 6010 3231 6012
rect 3255 6010 3311 6012
rect 3335 6010 3391 6012
rect 3415 6010 3471 6012
rect 3175 5958 3221 6010
rect 3221 5958 3231 6010
rect 3255 5958 3285 6010
rect 3285 5958 3297 6010
rect 3297 5958 3311 6010
rect 3335 5958 3349 6010
rect 3349 5958 3361 6010
rect 3361 5958 3391 6010
rect 3415 5958 3425 6010
rect 3425 5958 3471 6010
rect 3175 5956 3231 5958
rect 3255 5956 3311 5958
rect 3335 5956 3391 5958
rect 3415 5956 3471 5958
rect 5394 8730 5450 8732
rect 5474 8730 5530 8732
rect 5554 8730 5610 8732
rect 5634 8730 5690 8732
rect 5394 8678 5440 8730
rect 5440 8678 5450 8730
rect 5474 8678 5504 8730
rect 5504 8678 5516 8730
rect 5516 8678 5530 8730
rect 5554 8678 5568 8730
rect 5568 8678 5580 8730
rect 5580 8678 5610 8730
rect 5634 8678 5644 8730
rect 5644 8678 5690 8730
rect 5394 8676 5450 8678
rect 5474 8676 5530 8678
rect 5554 8676 5610 8678
rect 5634 8676 5690 8678
rect 5394 7642 5450 7644
rect 5474 7642 5530 7644
rect 5554 7642 5610 7644
rect 5634 7642 5690 7644
rect 5394 7590 5440 7642
rect 5440 7590 5450 7642
rect 5474 7590 5504 7642
rect 5504 7590 5516 7642
rect 5516 7590 5530 7642
rect 5554 7590 5568 7642
rect 5568 7590 5580 7642
rect 5580 7590 5610 7642
rect 5634 7590 5644 7642
rect 5644 7590 5690 7642
rect 5394 7588 5450 7590
rect 5474 7588 5530 7590
rect 5554 7588 5610 7590
rect 5634 7588 5690 7590
rect 5394 6554 5450 6556
rect 5474 6554 5530 6556
rect 5554 6554 5610 6556
rect 5634 6554 5690 6556
rect 5394 6502 5440 6554
rect 5440 6502 5450 6554
rect 5474 6502 5504 6554
rect 5504 6502 5516 6554
rect 5516 6502 5530 6554
rect 5554 6502 5568 6554
rect 5568 6502 5580 6554
rect 5580 6502 5610 6554
rect 5634 6502 5644 6554
rect 5644 6502 5690 6554
rect 5394 6500 5450 6502
rect 5474 6500 5530 6502
rect 5554 6500 5610 6502
rect 5634 6500 5690 6502
rect 3175 4922 3231 4924
rect 3255 4922 3311 4924
rect 3335 4922 3391 4924
rect 3415 4922 3471 4924
rect 3175 4870 3221 4922
rect 3221 4870 3231 4922
rect 3255 4870 3285 4922
rect 3285 4870 3297 4922
rect 3297 4870 3311 4922
rect 3335 4870 3349 4922
rect 3349 4870 3361 4922
rect 3361 4870 3391 4922
rect 3415 4870 3425 4922
rect 3425 4870 3471 4922
rect 3175 4868 3231 4870
rect 3255 4868 3311 4870
rect 3335 4868 3391 4870
rect 3415 4868 3471 4870
rect 5394 5466 5450 5468
rect 5474 5466 5530 5468
rect 5554 5466 5610 5468
rect 5634 5466 5690 5468
rect 5394 5414 5440 5466
rect 5440 5414 5450 5466
rect 5474 5414 5504 5466
rect 5504 5414 5516 5466
rect 5516 5414 5530 5466
rect 5554 5414 5568 5466
rect 5568 5414 5580 5466
rect 5580 5414 5610 5466
rect 5634 5414 5644 5466
rect 5644 5414 5690 5466
rect 5394 5412 5450 5414
rect 5474 5412 5530 5414
rect 5554 5412 5610 5414
rect 5634 5412 5690 5414
rect 3175 3834 3231 3836
rect 3255 3834 3311 3836
rect 3335 3834 3391 3836
rect 3415 3834 3471 3836
rect 3175 3782 3221 3834
rect 3221 3782 3231 3834
rect 3255 3782 3285 3834
rect 3285 3782 3297 3834
rect 3297 3782 3311 3834
rect 3335 3782 3349 3834
rect 3349 3782 3361 3834
rect 3361 3782 3391 3834
rect 3415 3782 3425 3834
rect 3425 3782 3471 3834
rect 3175 3780 3231 3782
rect 3255 3780 3311 3782
rect 3335 3780 3391 3782
rect 3415 3780 3471 3782
rect 3175 2746 3231 2748
rect 3255 2746 3311 2748
rect 3335 2746 3391 2748
rect 3415 2746 3471 2748
rect 3175 2694 3221 2746
rect 3221 2694 3231 2746
rect 3255 2694 3285 2746
rect 3285 2694 3297 2746
rect 3297 2694 3311 2746
rect 3335 2694 3349 2746
rect 3349 2694 3361 2746
rect 3361 2694 3391 2746
rect 3415 2694 3425 2746
rect 3425 2694 3471 2746
rect 3175 2692 3231 2694
rect 3255 2692 3311 2694
rect 3335 2692 3391 2694
rect 3415 2692 3471 2694
rect 5394 4378 5450 4380
rect 5474 4378 5530 4380
rect 5554 4378 5610 4380
rect 5634 4378 5690 4380
rect 5394 4326 5440 4378
rect 5440 4326 5450 4378
rect 5474 4326 5504 4378
rect 5504 4326 5516 4378
rect 5516 4326 5530 4378
rect 5554 4326 5568 4378
rect 5568 4326 5580 4378
rect 5580 4326 5610 4378
rect 5634 4326 5644 4378
rect 5644 4326 5690 4378
rect 5394 4324 5450 4326
rect 5474 4324 5530 4326
rect 5554 4324 5610 4326
rect 5634 4324 5690 4326
rect 7614 12538 7670 12540
rect 7694 12538 7750 12540
rect 7774 12538 7830 12540
rect 7854 12538 7910 12540
rect 7614 12486 7660 12538
rect 7660 12486 7670 12538
rect 7694 12486 7724 12538
rect 7724 12486 7736 12538
rect 7736 12486 7750 12538
rect 7774 12486 7788 12538
rect 7788 12486 7800 12538
rect 7800 12486 7830 12538
rect 7854 12486 7864 12538
rect 7864 12486 7910 12538
rect 7614 12484 7670 12486
rect 7694 12484 7750 12486
rect 7774 12484 7830 12486
rect 7854 12484 7910 12486
rect 7614 11450 7670 11452
rect 7694 11450 7750 11452
rect 7774 11450 7830 11452
rect 7854 11450 7910 11452
rect 7614 11398 7660 11450
rect 7660 11398 7670 11450
rect 7694 11398 7724 11450
rect 7724 11398 7736 11450
rect 7736 11398 7750 11450
rect 7774 11398 7788 11450
rect 7788 11398 7800 11450
rect 7800 11398 7830 11450
rect 7854 11398 7864 11450
rect 7864 11398 7910 11450
rect 7614 11396 7670 11398
rect 7694 11396 7750 11398
rect 7774 11396 7830 11398
rect 7854 11396 7910 11398
rect 7614 10362 7670 10364
rect 7694 10362 7750 10364
rect 7774 10362 7830 10364
rect 7854 10362 7910 10364
rect 7614 10310 7660 10362
rect 7660 10310 7670 10362
rect 7694 10310 7724 10362
rect 7724 10310 7736 10362
rect 7736 10310 7750 10362
rect 7774 10310 7788 10362
rect 7788 10310 7800 10362
rect 7800 10310 7830 10362
rect 7854 10310 7864 10362
rect 7864 10310 7910 10362
rect 7614 10308 7670 10310
rect 7694 10308 7750 10310
rect 7774 10308 7830 10310
rect 7854 10308 7910 10310
rect 7614 9274 7670 9276
rect 7694 9274 7750 9276
rect 7774 9274 7830 9276
rect 7854 9274 7910 9276
rect 7614 9222 7660 9274
rect 7660 9222 7670 9274
rect 7694 9222 7724 9274
rect 7724 9222 7736 9274
rect 7736 9222 7750 9274
rect 7774 9222 7788 9274
rect 7788 9222 7800 9274
rect 7800 9222 7830 9274
rect 7854 9222 7864 9274
rect 7864 9222 7910 9274
rect 7614 9220 7670 9222
rect 7694 9220 7750 9222
rect 7774 9220 7830 9222
rect 7854 9220 7910 9222
rect 7614 8186 7670 8188
rect 7694 8186 7750 8188
rect 7774 8186 7830 8188
rect 7854 8186 7910 8188
rect 7614 8134 7660 8186
rect 7660 8134 7670 8186
rect 7694 8134 7724 8186
rect 7724 8134 7736 8186
rect 7736 8134 7750 8186
rect 7774 8134 7788 8186
rect 7788 8134 7800 8186
rect 7800 8134 7830 8186
rect 7854 8134 7864 8186
rect 7864 8134 7910 8186
rect 7614 8132 7670 8134
rect 7694 8132 7750 8134
rect 7774 8132 7830 8134
rect 7854 8132 7910 8134
rect 9833 15258 9889 15260
rect 9913 15258 9969 15260
rect 9993 15258 10049 15260
rect 10073 15258 10129 15260
rect 9833 15206 9879 15258
rect 9879 15206 9889 15258
rect 9913 15206 9943 15258
rect 9943 15206 9955 15258
rect 9955 15206 9969 15258
rect 9993 15206 10007 15258
rect 10007 15206 10019 15258
rect 10019 15206 10049 15258
rect 10073 15206 10083 15258
rect 10083 15206 10129 15258
rect 9833 15204 9889 15206
rect 9913 15204 9969 15206
rect 9993 15204 10049 15206
rect 10073 15204 10129 15206
rect 9833 14170 9889 14172
rect 9913 14170 9969 14172
rect 9993 14170 10049 14172
rect 10073 14170 10129 14172
rect 9833 14118 9879 14170
rect 9879 14118 9889 14170
rect 9913 14118 9943 14170
rect 9943 14118 9955 14170
rect 9955 14118 9969 14170
rect 9993 14118 10007 14170
rect 10007 14118 10019 14170
rect 10019 14118 10049 14170
rect 10073 14118 10083 14170
rect 10083 14118 10129 14170
rect 9833 14116 9889 14118
rect 9913 14116 9969 14118
rect 9993 14116 10049 14118
rect 10073 14116 10129 14118
rect 9218 12280 9274 12336
rect 7614 7098 7670 7100
rect 7694 7098 7750 7100
rect 7774 7098 7830 7100
rect 7854 7098 7910 7100
rect 7614 7046 7660 7098
rect 7660 7046 7670 7098
rect 7694 7046 7724 7098
rect 7724 7046 7736 7098
rect 7736 7046 7750 7098
rect 7774 7046 7788 7098
rect 7788 7046 7800 7098
rect 7800 7046 7830 7098
rect 7854 7046 7864 7098
rect 7864 7046 7910 7098
rect 7614 7044 7670 7046
rect 7694 7044 7750 7046
rect 7774 7044 7830 7046
rect 7854 7044 7910 7046
rect 7614 6010 7670 6012
rect 7694 6010 7750 6012
rect 7774 6010 7830 6012
rect 7854 6010 7910 6012
rect 7614 5958 7660 6010
rect 7660 5958 7670 6010
rect 7694 5958 7724 6010
rect 7724 5958 7736 6010
rect 7736 5958 7750 6010
rect 7774 5958 7788 6010
rect 7788 5958 7800 6010
rect 7800 5958 7830 6010
rect 7854 5958 7864 6010
rect 7864 5958 7910 6010
rect 7614 5956 7670 5958
rect 7694 5956 7750 5958
rect 7774 5956 7830 5958
rect 7854 5956 7910 5958
rect 5394 3290 5450 3292
rect 5474 3290 5530 3292
rect 5554 3290 5610 3292
rect 5634 3290 5690 3292
rect 5394 3238 5440 3290
rect 5440 3238 5450 3290
rect 5474 3238 5504 3290
rect 5504 3238 5516 3290
rect 5516 3238 5530 3290
rect 5554 3238 5568 3290
rect 5568 3238 5580 3290
rect 5580 3238 5610 3290
rect 5634 3238 5644 3290
rect 5644 3238 5690 3290
rect 5394 3236 5450 3238
rect 5474 3236 5530 3238
rect 5554 3236 5610 3238
rect 5634 3236 5690 3238
rect 7614 4922 7670 4924
rect 7694 4922 7750 4924
rect 7774 4922 7830 4924
rect 7854 4922 7910 4924
rect 7614 4870 7660 4922
rect 7660 4870 7670 4922
rect 7694 4870 7724 4922
rect 7724 4870 7736 4922
rect 7736 4870 7750 4922
rect 7774 4870 7788 4922
rect 7788 4870 7800 4922
rect 7800 4870 7830 4922
rect 7854 4870 7864 4922
rect 7864 4870 7910 4922
rect 7614 4868 7670 4870
rect 7694 4868 7750 4870
rect 7774 4868 7830 4870
rect 7854 4868 7910 4870
rect 12053 16890 12109 16892
rect 12133 16890 12189 16892
rect 12213 16890 12269 16892
rect 12293 16890 12349 16892
rect 12053 16838 12099 16890
rect 12099 16838 12109 16890
rect 12133 16838 12163 16890
rect 12163 16838 12175 16890
rect 12175 16838 12189 16890
rect 12213 16838 12227 16890
rect 12227 16838 12239 16890
rect 12239 16838 12269 16890
rect 12293 16838 12303 16890
rect 12303 16838 12349 16890
rect 12053 16836 12109 16838
rect 12133 16836 12189 16838
rect 12213 16836 12269 16838
rect 12293 16836 12349 16838
rect 16492 16890 16548 16892
rect 16572 16890 16628 16892
rect 16652 16890 16708 16892
rect 16732 16890 16788 16892
rect 16492 16838 16538 16890
rect 16538 16838 16548 16890
rect 16572 16838 16602 16890
rect 16602 16838 16614 16890
rect 16614 16838 16628 16890
rect 16652 16838 16666 16890
rect 16666 16838 16678 16890
rect 16678 16838 16708 16890
rect 16732 16838 16742 16890
rect 16742 16838 16788 16890
rect 16492 16836 16548 16838
rect 16572 16836 16628 16838
rect 16652 16836 16708 16838
rect 16732 16836 16788 16838
rect 9833 13082 9889 13084
rect 9913 13082 9969 13084
rect 9993 13082 10049 13084
rect 10073 13082 10129 13084
rect 9833 13030 9879 13082
rect 9879 13030 9889 13082
rect 9913 13030 9943 13082
rect 9943 13030 9955 13082
rect 9955 13030 9969 13082
rect 9993 13030 10007 13082
rect 10007 13030 10019 13082
rect 10019 13030 10049 13082
rect 10073 13030 10083 13082
rect 10083 13030 10129 13082
rect 9833 13028 9889 13030
rect 9913 13028 9969 13030
rect 9993 13028 10049 13030
rect 10073 13028 10129 13030
rect 9833 11994 9889 11996
rect 9913 11994 9969 11996
rect 9993 11994 10049 11996
rect 10073 11994 10129 11996
rect 9833 11942 9879 11994
rect 9879 11942 9889 11994
rect 9913 11942 9943 11994
rect 9943 11942 9955 11994
rect 9955 11942 9969 11994
rect 9993 11942 10007 11994
rect 10007 11942 10019 11994
rect 10019 11942 10049 11994
rect 10073 11942 10083 11994
rect 10083 11942 10129 11994
rect 9833 11940 9889 11942
rect 9913 11940 9969 11942
rect 9993 11940 10049 11942
rect 10073 11940 10129 11942
rect 9833 10906 9889 10908
rect 9913 10906 9969 10908
rect 9993 10906 10049 10908
rect 10073 10906 10129 10908
rect 9833 10854 9879 10906
rect 9879 10854 9889 10906
rect 9913 10854 9943 10906
rect 9943 10854 9955 10906
rect 9955 10854 9969 10906
rect 9993 10854 10007 10906
rect 10007 10854 10019 10906
rect 10019 10854 10049 10906
rect 10073 10854 10083 10906
rect 10083 10854 10129 10906
rect 9833 10852 9889 10854
rect 9913 10852 9969 10854
rect 9993 10852 10049 10854
rect 10073 10852 10129 10854
rect 9833 9818 9889 9820
rect 9913 9818 9969 9820
rect 9993 9818 10049 9820
rect 10073 9818 10129 9820
rect 9833 9766 9879 9818
rect 9879 9766 9889 9818
rect 9913 9766 9943 9818
rect 9943 9766 9955 9818
rect 9955 9766 9969 9818
rect 9993 9766 10007 9818
rect 10007 9766 10019 9818
rect 10019 9766 10049 9818
rect 10073 9766 10083 9818
rect 10083 9766 10129 9818
rect 9833 9764 9889 9766
rect 9913 9764 9969 9766
rect 9993 9764 10049 9766
rect 10073 9764 10129 9766
rect 9833 8730 9889 8732
rect 9913 8730 9969 8732
rect 9993 8730 10049 8732
rect 10073 8730 10129 8732
rect 9833 8678 9879 8730
rect 9879 8678 9889 8730
rect 9913 8678 9943 8730
rect 9943 8678 9955 8730
rect 9955 8678 9969 8730
rect 9993 8678 10007 8730
rect 10007 8678 10019 8730
rect 10019 8678 10049 8730
rect 10073 8678 10083 8730
rect 10083 8678 10129 8730
rect 9833 8676 9889 8678
rect 9913 8676 9969 8678
rect 9993 8676 10049 8678
rect 10073 8676 10129 8678
rect 9833 7642 9889 7644
rect 9913 7642 9969 7644
rect 9993 7642 10049 7644
rect 10073 7642 10129 7644
rect 9833 7590 9879 7642
rect 9879 7590 9889 7642
rect 9913 7590 9943 7642
rect 9943 7590 9955 7642
rect 9955 7590 9969 7642
rect 9993 7590 10007 7642
rect 10007 7590 10019 7642
rect 10019 7590 10049 7642
rect 10073 7590 10083 7642
rect 10083 7590 10129 7642
rect 9833 7588 9889 7590
rect 9913 7588 9969 7590
rect 9993 7588 10049 7590
rect 10073 7588 10129 7590
rect 7614 3834 7670 3836
rect 7694 3834 7750 3836
rect 7774 3834 7830 3836
rect 7854 3834 7910 3836
rect 7614 3782 7660 3834
rect 7660 3782 7670 3834
rect 7694 3782 7724 3834
rect 7724 3782 7736 3834
rect 7736 3782 7750 3834
rect 7774 3782 7788 3834
rect 7788 3782 7800 3834
rect 7800 3782 7830 3834
rect 7854 3782 7864 3834
rect 7864 3782 7910 3834
rect 7614 3780 7670 3782
rect 7694 3780 7750 3782
rect 7774 3780 7830 3782
rect 7854 3780 7910 3782
rect 12053 15802 12109 15804
rect 12133 15802 12189 15804
rect 12213 15802 12269 15804
rect 12293 15802 12349 15804
rect 12053 15750 12099 15802
rect 12099 15750 12109 15802
rect 12133 15750 12163 15802
rect 12163 15750 12175 15802
rect 12175 15750 12189 15802
rect 12213 15750 12227 15802
rect 12227 15750 12239 15802
rect 12239 15750 12269 15802
rect 12293 15750 12303 15802
rect 12303 15750 12349 15802
rect 12053 15748 12109 15750
rect 12133 15748 12189 15750
rect 12213 15748 12269 15750
rect 12293 15748 12349 15750
rect 12053 14714 12109 14716
rect 12133 14714 12189 14716
rect 12213 14714 12269 14716
rect 12293 14714 12349 14716
rect 12053 14662 12099 14714
rect 12099 14662 12109 14714
rect 12133 14662 12163 14714
rect 12163 14662 12175 14714
rect 12175 14662 12189 14714
rect 12213 14662 12227 14714
rect 12227 14662 12239 14714
rect 12239 14662 12269 14714
rect 12293 14662 12303 14714
rect 12303 14662 12349 14714
rect 12053 14660 12109 14662
rect 12133 14660 12189 14662
rect 12213 14660 12269 14662
rect 12293 14660 12349 14662
rect 12053 13626 12109 13628
rect 12133 13626 12189 13628
rect 12213 13626 12269 13628
rect 12293 13626 12349 13628
rect 12053 13574 12099 13626
rect 12099 13574 12109 13626
rect 12133 13574 12163 13626
rect 12163 13574 12175 13626
rect 12175 13574 12189 13626
rect 12213 13574 12227 13626
rect 12227 13574 12239 13626
rect 12239 13574 12269 13626
rect 12293 13574 12303 13626
rect 12303 13574 12349 13626
rect 12053 13572 12109 13574
rect 12133 13572 12189 13574
rect 12213 13572 12269 13574
rect 12293 13572 12349 13574
rect 12053 12538 12109 12540
rect 12133 12538 12189 12540
rect 12213 12538 12269 12540
rect 12293 12538 12349 12540
rect 12053 12486 12099 12538
rect 12099 12486 12109 12538
rect 12133 12486 12163 12538
rect 12163 12486 12175 12538
rect 12175 12486 12189 12538
rect 12213 12486 12227 12538
rect 12227 12486 12239 12538
rect 12239 12486 12269 12538
rect 12293 12486 12303 12538
rect 12303 12486 12349 12538
rect 12053 12484 12109 12486
rect 12133 12484 12189 12486
rect 12213 12484 12269 12486
rect 12293 12484 12349 12486
rect 12053 11450 12109 11452
rect 12133 11450 12189 11452
rect 12213 11450 12269 11452
rect 12293 11450 12349 11452
rect 12053 11398 12099 11450
rect 12099 11398 12109 11450
rect 12133 11398 12163 11450
rect 12163 11398 12175 11450
rect 12175 11398 12189 11450
rect 12213 11398 12227 11450
rect 12227 11398 12239 11450
rect 12239 11398 12269 11450
rect 12293 11398 12303 11450
rect 12303 11398 12349 11450
rect 12053 11396 12109 11398
rect 12133 11396 12189 11398
rect 12213 11396 12269 11398
rect 12293 11396 12349 11398
rect 14272 16346 14328 16348
rect 14352 16346 14408 16348
rect 14432 16346 14488 16348
rect 14512 16346 14568 16348
rect 14272 16294 14318 16346
rect 14318 16294 14328 16346
rect 14352 16294 14382 16346
rect 14382 16294 14394 16346
rect 14394 16294 14408 16346
rect 14432 16294 14446 16346
rect 14446 16294 14458 16346
rect 14458 16294 14488 16346
rect 14512 16294 14522 16346
rect 14522 16294 14568 16346
rect 14272 16292 14328 16294
rect 14352 16292 14408 16294
rect 14432 16292 14488 16294
rect 14512 16292 14568 16294
rect 16492 15802 16548 15804
rect 16572 15802 16628 15804
rect 16652 15802 16708 15804
rect 16732 15802 16788 15804
rect 16492 15750 16538 15802
rect 16538 15750 16548 15802
rect 16572 15750 16602 15802
rect 16602 15750 16614 15802
rect 16614 15750 16628 15802
rect 16652 15750 16666 15802
rect 16666 15750 16678 15802
rect 16678 15750 16708 15802
rect 16732 15750 16742 15802
rect 16742 15750 16788 15802
rect 16492 15748 16548 15750
rect 16572 15748 16628 15750
rect 16652 15748 16708 15750
rect 16732 15748 16788 15750
rect 14272 15258 14328 15260
rect 14352 15258 14408 15260
rect 14432 15258 14488 15260
rect 14512 15258 14568 15260
rect 14272 15206 14318 15258
rect 14318 15206 14328 15258
rect 14352 15206 14382 15258
rect 14382 15206 14394 15258
rect 14394 15206 14408 15258
rect 14432 15206 14446 15258
rect 14446 15206 14458 15258
rect 14458 15206 14488 15258
rect 14512 15206 14522 15258
rect 14522 15206 14568 15258
rect 14272 15204 14328 15206
rect 14352 15204 14408 15206
rect 14432 15204 14488 15206
rect 14512 15204 14568 15206
rect 9833 6554 9889 6556
rect 9913 6554 9969 6556
rect 9993 6554 10049 6556
rect 10073 6554 10129 6556
rect 9833 6502 9879 6554
rect 9879 6502 9889 6554
rect 9913 6502 9943 6554
rect 9943 6502 9955 6554
rect 9955 6502 9969 6554
rect 9993 6502 10007 6554
rect 10007 6502 10019 6554
rect 10019 6502 10049 6554
rect 10073 6502 10083 6554
rect 10083 6502 10129 6554
rect 9833 6500 9889 6502
rect 9913 6500 9969 6502
rect 9993 6500 10049 6502
rect 10073 6500 10129 6502
rect 9833 5466 9889 5468
rect 9913 5466 9969 5468
rect 9993 5466 10049 5468
rect 10073 5466 10129 5468
rect 9833 5414 9879 5466
rect 9879 5414 9889 5466
rect 9913 5414 9943 5466
rect 9943 5414 9955 5466
rect 9955 5414 9969 5466
rect 9993 5414 10007 5466
rect 10007 5414 10019 5466
rect 10019 5414 10049 5466
rect 10073 5414 10083 5466
rect 10083 5414 10129 5466
rect 9833 5412 9889 5414
rect 9913 5412 9969 5414
rect 9993 5412 10049 5414
rect 10073 5412 10129 5414
rect 12053 10362 12109 10364
rect 12133 10362 12189 10364
rect 12213 10362 12269 10364
rect 12293 10362 12349 10364
rect 12053 10310 12099 10362
rect 12099 10310 12109 10362
rect 12133 10310 12163 10362
rect 12163 10310 12175 10362
rect 12175 10310 12189 10362
rect 12213 10310 12227 10362
rect 12227 10310 12239 10362
rect 12239 10310 12269 10362
rect 12293 10310 12303 10362
rect 12303 10310 12349 10362
rect 12053 10308 12109 10310
rect 12133 10308 12189 10310
rect 12213 10308 12269 10310
rect 12293 10308 12349 10310
rect 11978 9596 11980 9616
rect 11980 9596 12032 9616
rect 12032 9596 12034 9616
rect 11978 9560 12034 9596
rect 12053 9274 12109 9276
rect 12133 9274 12189 9276
rect 12213 9274 12269 9276
rect 12293 9274 12349 9276
rect 12053 9222 12099 9274
rect 12099 9222 12109 9274
rect 12133 9222 12163 9274
rect 12163 9222 12175 9274
rect 12175 9222 12189 9274
rect 12213 9222 12227 9274
rect 12227 9222 12239 9274
rect 12239 9222 12269 9274
rect 12293 9222 12303 9274
rect 12303 9222 12349 9274
rect 12053 9220 12109 9222
rect 12133 9220 12189 9222
rect 12213 9220 12269 9222
rect 12293 9220 12349 9222
rect 12254 8744 12310 8800
rect 12053 8186 12109 8188
rect 12133 8186 12189 8188
rect 12213 8186 12269 8188
rect 12293 8186 12349 8188
rect 12053 8134 12099 8186
rect 12099 8134 12109 8186
rect 12133 8134 12163 8186
rect 12163 8134 12175 8186
rect 12175 8134 12189 8186
rect 12213 8134 12227 8186
rect 12227 8134 12239 8186
rect 12239 8134 12269 8186
rect 12293 8134 12303 8186
rect 12303 8134 12349 8186
rect 12053 8132 12109 8134
rect 12133 8132 12189 8134
rect 12213 8132 12269 8134
rect 12293 8132 12349 8134
rect 7614 2746 7670 2748
rect 7694 2746 7750 2748
rect 7774 2746 7830 2748
rect 7854 2746 7910 2748
rect 7614 2694 7660 2746
rect 7660 2694 7670 2746
rect 7694 2694 7724 2746
rect 7724 2694 7736 2746
rect 7736 2694 7750 2746
rect 7774 2694 7788 2746
rect 7788 2694 7800 2746
rect 7800 2694 7830 2746
rect 7854 2694 7864 2746
rect 7864 2694 7910 2746
rect 7614 2692 7670 2694
rect 7694 2692 7750 2694
rect 7774 2692 7830 2694
rect 7854 2692 7910 2694
rect 9833 4378 9889 4380
rect 9913 4378 9969 4380
rect 9993 4378 10049 4380
rect 10073 4378 10129 4380
rect 9833 4326 9879 4378
rect 9879 4326 9889 4378
rect 9913 4326 9943 4378
rect 9943 4326 9955 4378
rect 9955 4326 9969 4378
rect 9993 4326 10007 4378
rect 10007 4326 10019 4378
rect 10019 4326 10049 4378
rect 10073 4326 10083 4378
rect 10083 4326 10129 4378
rect 9833 4324 9889 4326
rect 9913 4324 9969 4326
rect 9993 4324 10049 4326
rect 10073 4324 10129 4326
rect 12053 7098 12109 7100
rect 12133 7098 12189 7100
rect 12213 7098 12269 7100
rect 12293 7098 12349 7100
rect 12053 7046 12099 7098
rect 12099 7046 12109 7098
rect 12133 7046 12163 7098
rect 12163 7046 12175 7098
rect 12175 7046 12189 7098
rect 12213 7046 12227 7098
rect 12227 7046 12239 7098
rect 12239 7046 12269 7098
rect 12293 7046 12303 7098
rect 12303 7046 12349 7098
rect 12053 7044 12109 7046
rect 12133 7044 12189 7046
rect 12213 7044 12269 7046
rect 12293 7044 12349 7046
rect 14272 14170 14328 14172
rect 14352 14170 14408 14172
rect 14432 14170 14488 14172
rect 14512 14170 14568 14172
rect 14272 14118 14318 14170
rect 14318 14118 14328 14170
rect 14352 14118 14382 14170
rect 14382 14118 14394 14170
rect 14394 14118 14408 14170
rect 14432 14118 14446 14170
rect 14446 14118 14458 14170
rect 14458 14118 14488 14170
rect 14512 14118 14522 14170
rect 14522 14118 14568 14170
rect 14272 14116 14328 14118
rect 14352 14116 14408 14118
rect 14432 14116 14488 14118
rect 14512 14116 14568 14118
rect 14272 13082 14328 13084
rect 14352 13082 14408 13084
rect 14432 13082 14488 13084
rect 14512 13082 14568 13084
rect 14272 13030 14318 13082
rect 14318 13030 14328 13082
rect 14352 13030 14382 13082
rect 14382 13030 14394 13082
rect 14394 13030 14408 13082
rect 14432 13030 14446 13082
rect 14446 13030 14458 13082
rect 14458 13030 14488 13082
rect 14512 13030 14522 13082
rect 14522 13030 14568 13082
rect 14272 13028 14328 13030
rect 14352 13028 14408 13030
rect 14432 13028 14488 13030
rect 14512 13028 14568 13030
rect 14272 11994 14328 11996
rect 14352 11994 14408 11996
rect 14432 11994 14488 11996
rect 14512 11994 14568 11996
rect 14272 11942 14318 11994
rect 14318 11942 14328 11994
rect 14352 11942 14382 11994
rect 14382 11942 14394 11994
rect 14394 11942 14408 11994
rect 14432 11942 14446 11994
rect 14446 11942 14458 11994
rect 14458 11942 14488 11994
rect 14512 11942 14522 11994
rect 14522 11942 14568 11994
rect 14272 11940 14328 11942
rect 14352 11940 14408 11942
rect 14432 11940 14488 11942
rect 14512 11940 14568 11942
rect 14272 10906 14328 10908
rect 14352 10906 14408 10908
rect 14432 10906 14488 10908
rect 14512 10906 14568 10908
rect 14272 10854 14318 10906
rect 14318 10854 14328 10906
rect 14352 10854 14382 10906
rect 14382 10854 14394 10906
rect 14394 10854 14408 10906
rect 14432 10854 14446 10906
rect 14446 10854 14458 10906
rect 14458 10854 14488 10906
rect 14512 10854 14522 10906
rect 14522 10854 14568 10906
rect 14272 10852 14328 10854
rect 14352 10852 14408 10854
rect 14432 10852 14488 10854
rect 14512 10852 14568 10854
rect 14272 9818 14328 9820
rect 14352 9818 14408 9820
rect 14432 9818 14488 9820
rect 14512 9818 14568 9820
rect 14272 9766 14318 9818
rect 14318 9766 14328 9818
rect 14352 9766 14382 9818
rect 14382 9766 14394 9818
rect 14394 9766 14408 9818
rect 14432 9766 14446 9818
rect 14446 9766 14458 9818
rect 14458 9766 14488 9818
rect 14512 9766 14522 9818
rect 14522 9766 14568 9818
rect 14272 9764 14328 9766
rect 14352 9764 14408 9766
rect 14432 9764 14488 9766
rect 14512 9764 14568 9766
rect 14002 8780 14004 8800
rect 14004 8780 14056 8800
rect 14056 8780 14058 8800
rect 14002 8744 14058 8780
rect 14272 8730 14328 8732
rect 14352 8730 14408 8732
rect 14432 8730 14488 8732
rect 14512 8730 14568 8732
rect 14272 8678 14318 8730
rect 14318 8678 14328 8730
rect 14352 8678 14382 8730
rect 14382 8678 14394 8730
rect 14394 8678 14408 8730
rect 14432 8678 14446 8730
rect 14446 8678 14458 8730
rect 14458 8678 14488 8730
rect 14512 8678 14522 8730
rect 14522 8678 14568 8730
rect 14272 8676 14328 8678
rect 14352 8676 14408 8678
rect 14432 8676 14488 8678
rect 14512 8676 14568 8678
rect 18711 16346 18767 16348
rect 18791 16346 18847 16348
rect 18871 16346 18927 16348
rect 18951 16346 19007 16348
rect 18711 16294 18757 16346
rect 18757 16294 18767 16346
rect 18791 16294 18821 16346
rect 18821 16294 18833 16346
rect 18833 16294 18847 16346
rect 18871 16294 18885 16346
rect 18885 16294 18897 16346
rect 18897 16294 18927 16346
rect 18951 16294 18961 16346
rect 18961 16294 19007 16346
rect 18711 16292 18767 16294
rect 18791 16292 18847 16294
rect 18871 16292 18927 16294
rect 18951 16292 19007 16294
rect 18711 15258 18767 15260
rect 18791 15258 18847 15260
rect 18871 15258 18927 15260
rect 18951 15258 19007 15260
rect 18711 15206 18757 15258
rect 18757 15206 18767 15258
rect 18791 15206 18821 15258
rect 18821 15206 18833 15258
rect 18833 15206 18847 15258
rect 18871 15206 18885 15258
rect 18885 15206 18897 15258
rect 18897 15206 18927 15258
rect 18951 15206 18961 15258
rect 18961 15206 19007 15258
rect 18711 15204 18767 15206
rect 18791 15204 18847 15206
rect 18871 15204 18927 15206
rect 18951 15204 19007 15206
rect 16492 14714 16548 14716
rect 16572 14714 16628 14716
rect 16652 14714 16708 14716
rect 16732 14714 16788 14716
rect 16492 14662 16538 14714
rect 16538 14662 16548 14714
rect 16572 14662 16602 14714
rect 16602 14662 16614 14714
rect 16614 14662 16628 14714
rect 16652 14662 16666 14714
rect 16666 14662 16678 14714
rect 16678 14662 16708 14714
rect 16732 14662 16742 14714
rect 16742 14662 16788 14714
rect 16492 14660 16548 14662
rect 16572 14660 16628 14662
rect 16652 14660 16708 14662
rect 16732 14660 16788 14662
rect 16492 13626 16548 13628
rect 16572 13626 16628 13628
rect 16652 13626 16708 13628
rect 16732 13626 16788 13628
rect 16492 13574 16538 13626
rect 16538 13574 16548 13626
rect 16572 13574 16602 13626
rect 16602 13574 16614 13626
rect 16614 13574 16628 13626
rect 16652 13574 16666 13626
rect 16666 13574 16678 13626
rect 16678 13574 16708 13626
rect 16732 13574 16742 13626
rect 16742 13574 16788 13626
rect 16492 13572 16548 13574
rect 16572 13572 16628 13574
rect 16652 13572 16708 13574
rect 16732 13572 16788 13574
rect 16492 12538 16548 12540
rect 16572 12538 16628 12540
rect 16652 12538 16708 12540
rect 16732 12538 16788 12540
rect 16492 12486 16538 12538
rect 16538 12486 16548 12538
rect 16572 12486 16602 12538
rect 16602 12486 16614 12538
rect 16614 12486 16628 12538
rect 16652 12486 16666 12538
rect 16666 12486 16678 12538
rect 16678 12486 16708 12538
rect 16732 12486 16742 12538
rect 16742 12486 16788 12538
rect 16492 12484 16548 12486
rect 16572 12484 16628 12486
rect 16652 12484 16708 12486
rect 16732 12484 16788 12486
rect 12053 6010 12109 6012
rect 12133 6010 12189 6012
rect 12213 6010 12269 6012
rect 12293 6010 12349 6012
rect 12053 5958 12099 6010
rect 12099 5958 12109 6010
rect 12133 5958 12163 6010
rect 12163 5958 12175 6010
rect 12175 5958 12189 6010
rect 12213 5958 12227 6010
rect 12227 5958 12239 6010
rect 12239 5958 12269 6010
rect 12293 5958 12303 6010
rect 12303 5958 12349 6010
rect 12053 5956 12109 5958
rect 12133 5956 12189 5958
rect 12213 5956 12269 5958
rect 12293 5956 12349 5958
rect 9833 3290 9889 3292
rect 9913 3290 9969 3292
rect 9993 3290 10049 3292
rect 10073 3290 10129 3292
rect 9833 3238 9879 3290
rect 9879 3238 9889 3290
rect 9913 3238 9943 3290
rect 9943 3238 9955 3290
rect 9955 3238 9969 3290
rect 9993 3238 10007 3290
rect 10007 3238 10019 3290
rect 10019 3238 10049 3290
rect 10073 3238 10083 3290
rect 10083 3238 10129 3290
rect 9833 3236 9889 3238
rect 9913 3236 9969 3238
rect 9993 3236 10049 3238
rect 10073 3236 10129 3238
rect 5394 2202 5450 2204
rect 5474 2202 5530 2204
rect 5554 2202 5610 2204
rect 5634 2202 5690 2204
rect 5394 2150 5440 2202
rect 5440 2150 5450 2202
rect 5474 2150 5504 2202
rect 5504 2150 5516 2202
rect 5516 2150 5530 2202
rect 5554 2150 5568 2202
rect 5568 2150 5580 2202
rect 5580 2150 5610 2202
rect 5634 2150 5644 2202
rect 5644 2150 5690 2202
rect 5394 2148 5450 2150
rect 5474 2148 5530 2150
rect 5554 2148 5610 2150
rect 5634 2148 5690 2150
rect 9833 2202 9889 2204
rect 9913 2202 9969 2204
rect 9993 2202 10049 2204
rect 10073 2202 10129 2204
rect 9833 2150 9879 2202
rect 9879 2150 9889 2202
rect 9913 2150 9943 2202
rect 9943 2150 9955 2202
rect 9955 2150 9969 2202
rect 9993 2150 10007 2202
rect 10007 2150 10019 2202
rect 10019 2150 10049 2202
rect 10073 2150 10083 2202
rect 10083 2150 10129 2202
rect 9833 2148 9889 2150
rect 9913 2148 9969 2150
rect 9993 2148 10049 2150
rect 10073 2148 10129 2150
rect 12053 4922 12109 4924
rect 12133 4922 12189 4924
rect 12213 4922 12269 4924
rect 12293 4922 12349 4924
rect 12053 4870 12099 4922
rect 12099 4870 12109 4922
rect 12133 4870 12163 4922
rect 12163 4870 12175 4922
rect 12175 4870 12189 4922
rect 12213 4870 12227 4922
rect 12227 4870 12239 4922
rect 12239 4870 12269 4922
rect 12293 4870 12303 4922
rect 12303 4870 12349 4922
rect 12053 4868 12109 4870
rect 12133 4868 12189 4870
rect 12213 4868 12269 4870
rect 12293 4868 12349 4870
rect 12053 3834 12109 3836
rect 12133 3834 12189 3836
rect 12213 3834 12269 3836
rect 12293 3834 12349 3836
rect 12053 3782 12099 3834
rect 12099 3782 12109 3834
rect 12133 3782 12163 3834
rect 12163 3782 12175 3834
rect 12175 3782 12189 3834
rect 12213 3782 12227 3834
rect 12227 3782 12239 3834
rect 12239 3782 12269 3834
rect 12293 3782 12303 3834
rect 12303 3782 12349 3834
rect 12053 3780 12109 3782
rect 12133 3780 12189 3782
rect 12213 3780 12269 3782
rect 12293 3780 12349 3782
rect 15934 9580 15990 9616
rect 15934 9560 15936 9580
rect 15936 9560 15988 9580
rect 15988 9560 15990 9580
rect 14272 7642 14328 7644
rect 14352 7642 14408 7644
rect 14432 7642 14488 7644
rect 14512 7642 14568 7644
rect 14272 7590 14318 7642
rect 14318 7590 14328 7642
rect 14352 7590 14382 7642
rect 14382 7590 14394 7642
rect 14394 7590 14408 7642
rect 14432 7590 14446 7642
rect 14446 7590 14458 7642
rect 14458 7590 14488 7642
rect 14512 7590 14522 7642
rect 14522 7590 14568 7642
rect 14272 7588 14328 7590
rect 14352 7588 14408 7590
rect 14432 7588 14488 7590
rect 14512 7588 14568 7590
rect 16492 11450 16548 11452
rect 16572 11450 16628 11452
rect 16652 11450 16708 11452
rect 16732 11450 16788 11452
rect 16492 11398 16538 11450
rect 16538 11398 16548 11450
rect 16572 11398 16602 11450
rect 16602 11398 16614 11450
rect 16614 11398 16628 11450
rect 16652 11398 16666 11450
rect 16666 11398 16678 11450
rect 16678 11398 16708 11450
rect 16732 11398 16742 11450
rect 16742 11398 16788 11450
rect 16492 11396 16548 11398
rect 16572 11396 16628 11398
rect 16652 11396 16708 11398
rect 16732 11396 16788 11398
rect 16492 10362 16548 10364
rect 16572 10362 16628 10364
rect 16652 10362 16708 10364
rect 16732 10362 16788 10364
rect 16492 10310 16538 10362
rect 16538 10310 16548 10362
rect 16572 10310 16602 10362
rect 16602 10310 16614 10362
rect 16614 10310 16628 10362
rect 16652 10310 16666 10362
rect 16666 10310 16678 10362
rect 16678 10310 16708 10362
rect 16732 10310 16742 10362
rect 16742 10310 16788 10362
rect 16492 10308 16548 10310
rect 16572 10308 16628 10310
rect 16652 10308 16708 10310
rect 16732 10308 16788 10310
rect 16492 9274 16548 9276
rect 16572 9274 16628 9276
rect 16652 9274 16708 9276
rect 16732 9274 16788 9276
rect 16492 9222 16538 9274
rect 16538 9222 16548 9274
rect 16572 9222 16602 9274
rect 16602 9222 16614 9274
rect 16614 9222 16628 9274
rect 16652 9222 16666 9274
rect 16666 9222 16678 9274
rect 16678 9222 16708 9274
rect 16732 9222 16742 9274
rect 16742 9222 16788 9274
rect 16492 9220 16548 9222
rect 16572 9220 16628 9222
rect 16652 9220 16708 9222
rect 16732 9220 16788 9222
rect 18711 14170 18767 14172
rect 18791 14170 18847 14172
rect 18871 14170 18927 14172
rect 18951 14170 19007 14172
rect 18711 14118 18757 14170
rect 18757 14118 18767 14170
rect 18791 14118 18821 14170
rect 18821 14118 18833 14170
rect 18833 14118 18847 14170
rect 18871 14118 18885 14170
rect 18885 14118 18897 14170
rect 18897 14118 18927 14170
rect 18951 14118 18961 14170
rect 18961 14118 19007 14170
rect 18711 14116 18767 14118
rect 18791 14116 18847 14118
rect 18871 14116 18927 14118
rect 18951 14116 19007 14118
rect 18711 13082 18767 13084
rect 18791 13082 18847 13084
rect 18871 13082 18927 13084
rect 18951 13082 19007 13084
rect 18711 13030 18757 13082
rect 18757 13030 18767 13082
rect 18791 13030 18821 13082
rect 18821 13030 18833 13082
rect 18833 13030 18847 13082
rect 18871 13030 18885 13082
rect 18885 13030 18897 13082
rect 18897 13030 18927 13082
rect 18951 13030 18961 13082
rect 18961 13030 19007 13082
rect 18711 13028 18767 13030
rect 18791 13028 18847 13030
rect 18871 13028 18927 13030
rect 18951 13028 19007 13030
rect 18711 11994 18767 11996
rect 18791 11994 18847 11996
rect 18871 11994 18927 11996
rect 18951 11994 19007 11996
rect 18711 11942 18757 11994
rect 18757 11942 18767 11994
rect 18791 11942 18821 11994
rect 18821 11942 18833 11994
rect 18833 11942 18847 11994
rect 18871 11942 18885 11994
rect 18885 11942 18897 11994
rect 18897 11942 18927 11994
rect 18951 11942 18961 11994
rect 18961 11942 19007 11994
rect 18711 11940 18767 11942
rect 18791 11940 18847 11942
rect 18871 11940 18927 11942
rect 18951 11940 19007 11942
rect 18711 10906 18767 10908
rect 18791 10906 18847 10908
rect 18871 10906 18927 10908
rect 18951 10906 19007 10908
rect 18711 10854 18757 10906
rect 18757 10854 18767 10906
rect 18791 10854 18821 10906
rect 18821 10854 18833 10906
rect 18833 10854 18847 10906
rect 18871 10854 18885 10906
rect 18885 10854 18897 10906
rect 18897 10854 18927 10906
rect 18951 10854 18961 10906
rect 18961 10854 19007 10906
rect 18711 10852 18767 10854
rect 18791 10852 18847 10854
rect 18871 10852 18927 10854
rect 18951 10852 19007 10854
rect 16492 8186 16548 8188
rect 16572 8186 16628 8188
rect 16652 8186 16708 8188
rect 16732 8186 16788 8188
rect 16492 8134 16538 8186
rect 16538 8134 16548 8186
rect 16572 8134 16602 8186
rect 16602 8134 16614 8186
rect 16614 8134 16628 8186
rect 16652 8134 16666 8186
rect 16666 8134 16678 8186
rect 16678 8134 16708 8186
rect 16732 8134 16742 8186
rect 16742 8134 16788 8186
rect 16492 8132 16548 8134
rect 16572 8132 16628 8134
rect 16652 8132 16708 8134
rect 16732 8132 16788 8134
rect 14272 6554 14328 6556
rect 14352 6554 14408 6556
rect 14432 6554 14488 6556
rect 14512 6554 14568 6556
rect 14272 6502 14318 6554
rect 14318 6502 14328 6554
rect 14352 6502 14382 6554
rect 14382 6502 14394 6554
rect 14394 6502 14408 6554
rect 14432 6502 14446 6554
rect 14446 6502 14458 6554
rect 14458 6502 14488 6554
rect 14512 6502 14522 6554
rect 14522 6502 14568 6554
rect 14272 6500 14328 6502
rect 14352 6500 14408 6502
rect 14432 6500 14488 6502
rect 14512 6500 14568 6502
rect 14272 5466 14328 5468
rect 14352 5466 14408 5468
rect 14432 5466 14488 5468
rect 14512 5466 14568 5468
rect 14272 5414 14318 5466
rect 14318 5414 14328 5466
rect 14352 5414 14382 5466
rect 14382 5414 14394 5466
rect 14394 5414 14408 5466
rect 14432 5414 14446 5466
rect 14446 5414 14458 5466
rect 14458 5414 14488 5466
rect 14512 5414 14522 5466
rect 14522 5414 14568 5466
rect 14272 5412 14328 5414
rect 14352 5412 14408 5414
rect 14432 5412 14488 5414
rect 14512 5412 14568 5414
rect 14272 4378 14328 4380
rect 14352 4378 14408 4380
rect 14432 4378 14488 4380
rect 14512 4378 14568 4380
rect 14272 4326 14318 4378
rect 14318 4326 14328 4378
rect 14352 4326 14382 4378
rect 14382 4326 14394 4378
rect 14394 4326 14408 4378
rect 14432 4326 14446 4378
rect 14446 4326 14458 4378
rect 14458 4326 14488 4378
rect 14512 4326 14522 4378
rect 14522 4326 14568 4378
rect 14272 4324 14328 4326
rect 14352 4324 14408 4326
rect 14432 4324 14488 4326
rect 14512 4324 14568 4326
rect 12053 2746 12109 2748
rect 12133 2746 12189 2748
rect 12213 2746 12269 2748
rect 12293 2746 12349 2748
rect 12053 2694 12099 2746
rect 12099 2694 12109 2746
rect 12133 2694 12163 2746
rect 12163 2694 12175 2746
rect 12175 2694 12189 2746
rect 12213 2694 12227 2746
rect 12227 2694 12239 2746
rect 12239 2694 12269 2746
rect 12293 2694 12303 2746
rect 12303 2694 12349 2746
rect 12053 2692 12109 2694
rect 12133 2692 12189 2694
rect 12213 2692 12269 2694
rect 12293 2692 12349 2694
rect 16492 7098 16548 7100
rect 16572 7098 16628 7100
rect 16652 7098 16708 7100
rect 16732 7098 16788 7100
rect 16492 7046 16538 7098
rect 16538 7046 16548 7098
rect 16572 7046 16602 7098
rect 16602 7046 16614 7098
rect 16614 7046 16628 7098
rect 16652 7046 16666 7098
rect 16666 7046 16678 7098
rect 16678 7046 16708 7098
rect 16732 7046 16742 7098
rect 16742 7046 16788 7098
rect 16492 7044 16548 7046
rect 16572 7044 16628 7046
rect 16652 7044 16708 7046
rect 16732 7044 16788 7046
rect 18711 9818 18767 9820
rect 18791 9818 18847 9820
rect 18871 9818 18927 9820
rect 18951 9818 19007 9820
rect 18711 9766 18757 9818
rect 18757 9766 18767 9818
rect 18791 9766 18821 9818
rect 18821 9766 18833 9818
rect 18833 9766 18847 9818
rect 18871 9766 18885 9818
rect 18885 9766 18897 9818
rect 18897 9766 18927 9818
rect 18951 9766 18961 9818
rect 18961 9766 19007 9818
rect 18711 9764 18767 9766
rect 18791 9764 18847 9766
rect 18871 9764 18927 9766
rect 18951 9764 19007 9766
rect 16492 6010 16548 6012
rect 16572 6010 16628 6012
rect 16652 6010 16708 6012
rect 16732 6010 16788 6012
rect 16492 5958 16538 6010
rect 16538 5958 16548 6010
rect 16572 5958 16602 6010
rect 16602 5958 16614 6010
rect 16614 5958 16628 6010
rect 16652 5958 16666 6010
rect 16666 5958 16678 6010
rect 16678 5958 16708 6010
rect 16732 5958 16742 6010
rect 16742 5958 16788 6010
rect 16492 5956 16548 5958
rect 16572 5956 16628 5958
rect 16652 5956 16708 5958
rect 16732 5956 16788 5958
rect 16492 4922 16548 4924
rect 16572 4922 16628 4924
rect 16652 4922 16708 4924
rect 16732 4922 16788 4924
rect 16492 4870 16538 4922
rect 16538 4870 16548 4922
rect 16572 4870 16602 4922
rect 16602 4870 16614 4922
rect 16614 4870 16628 4922
rect 16652 4870 16666 4922
rect 16666 4870 16678 4922
rect 16678 4870 16708 4922
rect 16732 4870 16742 4922
rect 16742 4870 16788 4922
rect 16492 4868 16548 4870
rect 16572 4868 16628 4870
rect 16652 4868 16708 4870
rect 16732 4868 16788 4870
rect 16492 3834 16548 3836
rect 16572 3834 16628 3836
rect 16652 3834 16708 3836
rect 16732 3834 16788 3836
rect 16492 3782 16538 3834
rect 16538 3782 16548 3834
rect 16572 3782 16602 3834
rect 16602 3782 16614 3834
rect 16614 3782 16628 3834
rect 16652 3782 16666 3834
rect 16666 3782 16678 3834
rect 16678 3782 16708 3834
rect 16732 3782 16742 3834
rect 16742 3782 16788 3834
rect 16492 3780 16548 3782
rect 16572 3780 16628 3782
rect 16652 3780 16708 3782
rect 16732 3780 16788 3782
rect 14272 3290 14328 3292
rect 14352 3290 14408 3292
rect 14432 3290 14488 3292
rect 14512 3290 14568 3292
rect 14272 3238 14318 3290
rect 14318 3238 14328 3290
rect 14352 3238 14382 3290
rect 14382 3238 14394 3290
rect 14394 3238 14408 3290
rect 14432 3238 14446 3290
rect 14446 3238 14458 3290
rect 14458 3238 14488 3290
rect 14512 3238 14522 3290
rect 14522 3238 14568 3290
rect 14272 3236 14328 3238
rect 14352 3236 14408 3238
rect 14432 3236 14488 3238
rect 14512 3236 14568 3238
rect 14272 2202 14328 2204
rect 14352 2202 14408 2204
rect 14432 2202 14488 2204
rect 14512 2202 14568 2204
rect 14272 2150 14318 2202
rect 14318 2150 14328 2202
rect 14352 2150 14382 2202
rect 14382 2150 14394 2202
rect 14394 2150 14408 2202
rect 14432 2150 14446 2202
rect 14446 2150 14458 2202
rect 14458 2150 14488 2202
rect 14512 2150 14522 2202
rect 14522 2150 14568 2202
rect 14272 2148 14328 2150
rect 14352 2148 14408 2150
rect 14432 2148 14488 2150
rect 14512 2148 14568 2150
rect 16492 2746 16548 2748
rect 16572 2746 16628 2748
rect 16652 2746 16708 2748
rect 16732 2746 16788 2748
rect 16492 2694 16538 2746
rect 16538 2694 16548 2746
rect 16572 2694 16602 2746
rect 16602 2694 16614 2746
rect 16614 2694 16628 2746
rect 16652 2694 16666 2746
rect 16666 2694 16678 2746
rect 16678 2694 16708 2746
rect 16732 2694 16742 2746
rect 16742 2694 16788 2746
rect 16492 2692 16548 2694
rect 16572 2692 16628 2694
rect 16652 2692 16708 2694
rect 16732 2692 16788 2694
rect 18711 8730 18767 8732
rect 18791 8730 18847 8732
rect 18871 8730 18927 8732
rect 18951 8730 19007 8732
rect 18711 8678 18757 8730
rect 18757 8678 18767 8730
rect 18791 8678 18821 8730
rect 18821 8678 18833 8730
rect 18833 8678 18847 8730
rect 18871 8678 18885 8730
rect 18885 8678 18897 8730
rect 18897 8678 18927 8730
rect 18951 8678 18961 8730
rect 18961 8678 19007 8730
rect 18711 8676 18767 8678
rect 18791 8676 18847 8678
rect 18871 8676 18927 8678
rect 18951 8676 19007 8678
rect 18711 7642 18767 7644
rect 18791 7642 18847 7644
rect 18871 7642 18927 7644
rect 18951 7642 19007 7644
rect 18711 7590 18757 7642
rect 18757 7590 18767 7642
rect 18791 7590 18821 7642
rect 18821 7590 18833 7642
rect 18833 7590 18847 7642
rect 18871 7590 18885 7642
rect 18885 7590 18897 7642
rect 18897 7590 18927 7642
rect 18951 7590 18961 7642
rect 18961 7590 19007 7642
rect 18711 7588 18767 7590
rect 18791 7588 18847 7590
rect 18871 7588 18927 7590
rect 18951 7588 19007 7590
rect 18711 6554 18767 6556
rect 18791 6554 18847 6556
rect 18871 6554 18927 6556
rect 18951 6554 19007 6556
rect 18711 6502 18757 6554
rect 18757 6502 18767 6554
rect 18791 6502 18821 6554
rect 18821 6502 18833 6554
rect 18833 6502 18847 6554
rect 18871 6502 18885 6554
rect 18885 6502 18897 6554
rect 18897 6502 18927 6554
rect 18951 6502 18961 6554
rect 18961 6502 19007 6554
rect 18711 6500 18767 6502
rect 18791 6500 18847 6502
rect 18871 6500 18927 6502
rect 18951 6500 19007 6502
rect 18711 5466 18767 5468
rect 18791 5466 18847 5468
rect 18871 5466 18927 5468
rect 18951 5466 19007 5468
rect 18711 5414 18757 5466
rect 18757 5414 18767 5466
rect 18791 5414 18821 5466
rect 18821 5414 18833 5466
rect 18833 5414 18847 5466
rect 18871 5414 18885 5466
rect 18885 5414 18897 5466
rect 18897 5414 18927 5466
rect 18951 5414 18961 5466
rect 18961 5414 19007 5466
rect 18711 5412 18767 5414
rect 18791 5412 18847 5414
rect 18871 5412 18927 5414
rect 18951 5412 19007 5414
rect 18711 4378 18767 4380
rect 18791 4378 18847 4380
rect 18871 4378 18927 4380
rect 18951 4378 19007 4380
rect 18711 4326 18757 4378
rect 18757 4326 18767 4378
rect 18791 4326 18821 4378
rect 18821 4326 18833 4378
rect 18833 4326 18847 4378
rect 18871 4326 18885 4378
rect 18885 4326 18897 4378
rect 18897 4326 18927 4378
rect 18951 4326 18961 4378
rect 18961 4326 19007 4378
rect 18711 4324 18767 4326
rect 18791 4324 18847 4326
rect 18871 4324 18927 4326
rect 18951 4324 19007 4326
rect 18711 3290 18767 3292
rect 18791 3290 18847 3292
rect 18871 3290 18927 3292
rect 18951 3290 19007 3292
rect 18711 3238 18757 3290
rect 18757 3238 18767 3290
rect 18791 3238 18821 3290
rect 18821 3238 18833 3290
rect 18833 3238 18847 3290
rect 18871 3238 18885 3290
rect 18885 3238 18897 3290
rect 18897 3238 18927 3290
rect 18951 3238 18961 3290
rect 18961 3238 19007 3290
rect 18711 3236 18767 3238
rect 18791 3236 18847 3238
rect 18871 3236 18927 3238
rect 18951 3236 19007 3238
rect 18711 2202 18767 2204
rect 18791 2202 18847 2204
rect 18871 2202 18927 2204
rect 18951 2202 19007 2204
rect 18711 2150 18757 2202
rect 18757 2150 18767 2202
rect 18791 2150 18821 2202
rect 18821 2150 18833 2202
rect 18833 2150 18847 2202
rect 18871 2150 18885 2202
rect 18885 2150 18897 2202
rect 18897 2150 18927 2202
rect 18951 2150 18961 2202
rect 18961 2150 19007 2202
rect 18711 2148 18767 2150
rect 18791 2148 18847 2150
rect 18871 2148 18927 2150
rect 18951 2148 19007 2150
<< metal3 >>
rect 5384 17440 5700 17441
rect 5384 17376 5390 17440
rect 5454 17376 5470 17440
rect 5534 17376 5550 17440
rect 5614 17376 5630 17440
rect 5694 17376 5700 17440
rect 5384 17375 5700 17376
rect 9823 17440 10139 17441
rect 9823 17376 9829 17440
rect 9893 17376 9909 17440
rect 9973 17376 9989 17440
rect 10053 17376 10069 17440
rect 10133 17376 10139 17440
rect 9823 17375 10139 17376
rect 14262 17440 14578 17441
rect 14262 17376 14268 17440
rect 14332 17376 14348 17440
rect 14412 17376 14428 17440
rect 14492 17376 14508 17440
rect 14572 17376 14578 17440
rect 14262 17375 14578 17376
rect 18701 17440 19017 17441
rect 18701 17376 18707 17440
rect 18771 17376 18787 17440
rect 18851 17376 18867 17440
rect 18931 17376 18947 17440
rect 19011 17376 19017 17440
rect 18701 17375 19017 17376
rect 3165 16896 3481 16897
rect 3165 16832 3171 16896
rect 3235 16832 3251 16896
rect 3315 16832 3331 16896
rect 3395 16832 3411 16896
rect 3475 16832 3481 16896
rect 3165 16831 3481 16832
rect 7604 16896 7920 16897
rect 7604 16832 7610 16896
rect 7674 16832 7690 16896
rect 7754 16832 7770 16896
rect 7834 16832 7850 16896
rect 7914 16832 7920 16896
rect 7604 16831 7920 16832
rect 12043 16896 12359 16897
rect 12043 16832 12049 16896
rect 12113 16832 12129 16896
rect 12193 16832 12209 16896
rect 12273 16832 12289 16896
rect 12353 16832 12359 16896
rect 12043 16831 12359 16832
rect 16482 16896 16798 16897
rect 16482 16832 16488 16896
rect 16552 16832 16568 16896
rect 16632 16832 16648 16896
rect 16712 16832 16728 16896
rect 16792 16832 16798 16896
rect 16482 16831 16798 16832
rect 5384 16352 5700 16353
rect 5384 16288 5390 16352
rect 5454 16288 5470 16352
rect 5534 16288 5550 16352
rect 5614 16288 5630 16352
rect 5694 16288 5700 16352
rect 5384 16287 5700 16288
rect 9823 16352 10139 16353
rect 9823 16288 9829 16352
rect 9893 16288 9909 16352
rect 9973 16288 9989 16352
rect 10053 16288 10069 16352
rect 10133 16288 10139 16352
rect 9823 16287 10139 16288
rect 14262 16352 14578 16353
rect 14262 16288 14268 16352
rect 14332 16288 14348 16352
rect 14412 16288 14428 16352
rect 14492 16288 14508 16352
rect 14572 16288 14578 16352
rect 14262 16287 14578 16288
rect 18701 16352 19017 16353
rect 18701 16288 18707 16352
rect 18771 16288 18787 16352
rect 18851 16288 18867 16352
rect 18931 16288 18947 16352
rect 19011 16288 19017 16352
rect 18701 16287 19017 16288
rect 3165 15808 3481 15809
rect 3165 15744 3171 15808
rect 3235 15744 3251 15808
rect 3315 15744 3331 15808
rect 3395 15744 3411 15808
rect 3475 15744 3481 15808
rect 3165 15743 3481 15744
rect 7604 15808 7920 15809
rect 7604 15744 7610 15808
rect 7674 15744 7690 15808
rect 7754 15744 7770 15808
rect 7834 15744 7850 15808
rect 7914 15744 7920 15808
rect 7604 15743 7920 15744
rect 12043 15808 12359 15809
rect 12043 15744 12049 15808
rect 12113 15744 12129 15808
rect 12193 15744 12209 15808
rect 12273 15744 12289 15808
rect 12353 15744 12359 15808
rect 12043 15743 12359 15744
rect 16482 15808 16798 15809
rect 16482 15744 16488 15808
rect 16552 15744 16568 15808
rect 16632 15744 16648 15808
rect 16712 15744 16728 15808
rect 16792 15744 16798 15808
rect 16482 15743 16798 15744
rect 5384 15264 5700 15265
rect 5384 15200 5390 15264
rect 5454 15200 5470 15264
rect 5534 15200 5550 15264
rect 5614 15200 5630 15264
rect 5694 15200 5700 15264
rect 5384 15199 5700 15200
rect 9823 15264 10139 15265
rect 9823 15200 9829 15264
rect 9893 15200 9909 15264
rect 9973 15200 9989 15264
rect 10053 15200 10069 15264
rect 10133 15200 10139 15264
rect 9823 15199 10139 15200
rect 14262 15264 14578 15265
rect 14262 15200 14268 15264
rect 14332 15200 14348 15264
rect 14412 15200 14428 15264
rect 14492 15200 14508 15264
rect 14572 15200 14578 15264
rect 14262 15199 14578 15200
rect 18701 15264 19017 15265
rect 18701 15200 18707 15264
rect 18771 15200 18787 15264
rect 18851 15200 18867 15264
rect 18931 15200 18947 15264
rect 19011 15200 19017 15264
rect 18701 15199 19017 15200
rect 3165 14720 3481 14721
rect 3165 14656 3171 14720
rect 3235 14656 3251 14720
rect 3315 14656 3331 14720
rect 3395 14656 3411 14720
rect 3475 14656 3481 14720
rect 3165 14655 3481 14656
rect 7604 14720 7920 14721
rect 7604 14656 7610 14720
rect 7674 14656 7690 14720
rect 7754 14656 7770 14720
rect 7834 14656 7850 14720
rect 7914 14656 7920 14720
rect 7604 14655 7920 14656
rect 12043 14720 12359 14721
rect 12043 14656 12049 14720
rect 12113 14656 12129 14720
rect 12193 14656 12209 14720
rect 12273 14656 12289 14720
rect 12353 14656 12359 14720
rect 12043 14655 12359 14656
rect 16482 14720 16798 14721
rect 16482 14656 16488 14720
rect 16552 14656 16568 14720
rect 16632 14656 16648 14720
rect 16712 14656 16728 14720
rect 16792 14656 16798 14720
rect 16482 14655 16798 14656
rect 5384 14176 5700 14177
rect 5384 14112 5390 14176
rect 5454 14112 5470 14176
rect 5534 14112 5550 14176
rect 5614 14112 5630 14176
rect 5694 14112 5700 14176
rect 5384 14111 5700 14112
rect 9823 14176 10139 14177
rect 9823 14112 9829 14176
rect 9893 14112 9909 14176
rect 9973 14112 9989 14176
rect 10053 14112 10069 14176
rect 10133 14112 10139 14176
rect 9823 14111 10139 14112
rect 14262 14176 14578 14177
rect 14262 14112 14268 14176
rect 14332 14112 14348 14176
rect 14412 14112 14428 14176
rect 14492 14112 14508 14176
rect 14572 14112 14578 14176
rect 14262 14111 14578 14112
rect 18701 14176 19017 14177
rect 18701 14112 18707 14176
rect 18771 14112 18787 14176
rect 18851 14112 18867 14176
rect 18931 14112 18947 14176
rect 19011 14112 19017 14176
rect 18701 14111 19017 14112
rect 3165 13632 3481 13633
rect 3165 13568 3171 13632
rect 3235 13568 3251 13632
rect 3315 13568 3331 13632
rect 3395 13568 3411 13632
rect 3475 13568 3481 13632
rect 3165 13567 3481 13568
rect 7604 13632 7920 13633
rect 7604 13568 7610 13632
rect 7674 13568 7690 13632
rect 7754 13568 7770 13632
rect 7834 13568 7850 13632
rect 7914 13568 7920 13632
rect 7604 13567 7920 13568
rect 12043 13632 12359 13633
rect 12043 13568 12049 13632
rect 12113 13568 12129 13632
rect 12193 13568 12209 13632
rect 12273 13568 12289 13632
rect 12353 13568 12359 13632
rect 12043 13567 12359 13568
rect 16482 13632 16798 13633
rect 16482 13568 16488 13632
rect 16552 13568 16568 13632
rect 16632 13568 16648 13632
rect 16712 13568 16728 13632
rect 16792 13568 16798 13632
rect 16482 13567 16798 13568
rect 5384 13088 5700 13089
rect 5384 13024 5390 13088
rect 5454 13024 5470 13088
rect 5534 13024 5550 13088
rect 5614 13024 5630 13088
rect 5694 13024 5700 13088
rect 5384 13023 5700 13024
rect 9823 13088 10139 13089
rect 9823 13024 9829 13088
rect 9893 13024 9909 13088
rect 9973 13024 9989 13088
rect 10053 13024 10069 13088
rect 10133 13024 10139 13088
rect 9823 13023 10139 13024
rect 14262 13088 14578 13089
rect 14262 13024 14268 13088
rect 14332 13024 14348 13088
rect 14412 13024 14428 13088
rect 14492 13024 14508 13088
rect 14572 13024 14578 13088
rect 14262 13023 14578 13024
rect 18701 13088 19017 13089
rect 18701 13024 18707 13088
rect 18771 13024 18787 13088
rect 18851 13024 18867 13088
rect 18931 13024 18947 13088
rect 19011 13024 19017 13088
rect 18701 13023 19017 13024
rect 3165 12544 3481 12545
rect 3165 12480 3171 12544
rect 3235 12480 3251 12544
rect 3315 12480 3331 12544
rect 3395 12480 3411 12544
rect 3475 12480 3481 12544
rect 3165 12479 3481 12480
rect 7604 12544 7920 12545
rect 7604 12480 7610 12544
rect 7674 12480 7690 12544
rect 7754 12480 7770 12544
rect 7834 12480 7850 12544
rect 7914 12480 7920 12544
rect 7604 12479 7920 12480
rect 12043 12544 12359 12545
rect 12043 12480 12049 12544
rect 12113 12480 12129 12544
rect 12193 12480 12209 12544
rect 12273 12480 12289 12544
rect 12353 12480 12359 12544
rect 12043 12479 12359 12480
rect 16482 12544 16798 12545
rect 16482 12480 16488 12544
rect 16552 12480 16568 12544
rect 16632 12480 16648 12544
rect 16712 12480 16728 12544
rect 16792 12480 16798 12544
rect 16482 12479 16798 12480
rect 7005 12338 7071 12341
rect 9213 12338 9279 12341
rect 7005 12336 9279 12338
rect 7005 12280 7010 12336
rect 7066 12280 9218 12336
rect 9274 12280 9279 12336
rect 7005 12278 9279 12280
rect 7005 12275 7071 12278
rect 9213 12275 9279 12278
rect 5384 12000 5700 12001
rect 5384 11936 5390 12000
rect 5454 11936 5470 12000
rect 5534 11936 5550 12000
rect 5614 11936 5630 12000
rect 5694 11936 5700 12000
rect 5384 11935 5700 11936
rect 9823 12000 10139 12001
rect 9823 11936 9829 12000
rect 9893 11936 9909 12000
rect 9973 11936 9989 12000
rect 10053 11936 10069 12000
rect 10133 11936 10139 12000
rect 9823 11935 10139 11936
rect 14262 12000 14578 12001
rect 14262 11936 14268 12000
rect 14332 11936 14348 12000
rect 14412 11936 14428 12000
rect 14492 11936 14508 12000
rect 14572 11936 14578 12000
rect 14262 11935 14578 11936
rect 18701 12000 19017 12001
rect 18701 11936 18707 12000
rect 18771 11936 18787 12000
rect 18851 11936 18867 12000
rect 18931 11936 18947 12000
rect 19011 11936 19017 12000
rect 18701 11935 19017 11936
rect 3165 11456 3481 11457
rect 3165 11392 3171 11456
rect 3235 11392 3251 11456
rect 3315 11392 3331 11456
rect 3395 11392 3411 11456
rect 3475 11392 3481 11456
rect 3165 11391 3481 11392
rect 7604 11456 7920 11457
rect 7604 11392 7610 11456
rect 7674 11392 7690 11456
rect 7754 11392 7770 11456
rect 7834 11392 7850 11456
rect 7914 11392 7920 11456
rect 7604 11391 7920 11392
rect 12043 11456 12359 11457
rect 12043 11392 12049 11456
rect 12113 11392 12129 11456
rect 12193 11392 12209 11456
rect 12273 11392 12289 11456
rect 12353 11392 12359 11456
rect 12043 11391 12359 11392
rect 16482 11456 16798 11457
rect 16482 11392 16488 11456
rect 16552 11392 16568 11456
rect 16632 11392 16648 11456
rect 16712 11392 16728 11456
rect 16792 11392 16798 11456
rect 16482 11391 16798 11392
rect 5384 10912 5700 10913
rect 5384 10848 5390 10912
rect 5454 10848 5470 10912
rect 5534 10848 5550 10912
rect 5614 10848 5630 10912
rect 5694 10848 5700 10912
rect 5384 10847 5700 10848
rect 9823 10912 10139 10913
rect 9823 10848 9829 10912
rect 9893 10848 9909 10912
rect 9973 10848 9989 10912
rect 10053 10848 10069 10912
rect 10133 10848 10139 10912
rect 9823 10847 10139 10848
rect 14262 10912 14578 10913
rect 14262 10848 14268 10912
rect 14332 10848 14348 10912
rect 14412 10848 14428 10912
rect 14492 10848 14508 10912
rect 14572 10848 14578 10912
rect 14262 10847 14578 10848
rect 18701 10912 19017 10913
rect 18701 10848 18707 10912
rect 18771 10848 18787 10912
rect 18851 10848 18867 10912
rect 18931 10848 18947 10912
rect 19011 10848 19017 10912
rect 18701 10847 19017 10848
rect 3165 10368 3481 10369
rect 3165 10304 3171 10368
rect 3235 10304 3251 10368
rect 3315 10304 3331 10368
rect 3395 10304 3411 10368
rect 3475 10304 3481 10368
rect 3165 10303 3481 10304
rect 7604 10368 7920 10369
rect 7604 10304 7610 10368
rect 7674 10304 7690 10368
rect 7754 10304 7770 10368
rect 7834 10304 7850 10368
rect 7914 10304 7920 10368
rect 7604 10303 7920 10304
rect 12043 10368 12359 10369
rect 12043 10304 12049 10368
rect 12113 10304 12129 10368
rect 12193 10304 12209 10368
rect 12273 10304 12289 10368
rect 12353 10304 12359 10368
rect 12043 10303 12359 10304
rect 16482 10368 16798 10369
rect 16482 10304 16488 10368
rect 16552 10304 16568 10368
rect 16632 10304 16648 10368
rect 16712 10304 16728 10368
rect 16792 10304 16798 10368
rect 16482 10303 16798 10304
rect 5384 9824 5700 9825
rect 5384 9760 5390 9824
rect 5454 9760 5470 9824
rect 5534 9760 5550 9824
rect 5614 9760 5630 9824
rect 5694 9760 5700 9824
rect 5384 9759 5700 9760
rect 9823 9824 10139 9825
rect 9823 9760 9829 9824
rect 9893 9760 9909 9824
rect 9973 9760 9989 9824
rect 10053 9760 10069 9824
rect 10133 9760 10139 9824
rect 9823 9759 10139 9760
rect 14262 9824 14578 9825
rect 14262 9760 14268 9824
rect 14332 9760 14348 9824
rect 14412 9760 14428 9824
rect 14492 9760 14508 9824
rect 14572 9760 14578 9824
rect 14262 9759 14578 9760
rect 18701 9824 19017 9825
rect 18701 9760 18707 9824
rect 18771 9760 18787 9824
rect 18851 9760 18867 9824
rect 18931 9760 18947 9824
rect 19011 9760 19017 9824
rect 18701 9759 19017 9760
rect 11973 9618 12039 9621
rect 15929 9618 15995 9621
rect 11973 9616 15995 9618
rect 11973 9560 11978 9616
rect 12034 9560 15934 9616
rect 15990 9560 15995 9616
rect 11973 9558 15995 9560
rect 11973 9555 12039 9558
rect 15929 9555 15995 9558
rect 3165 9280 3481 9281
rect 3165 9216 3171 9280
rect 3235 9216 3251 9280
rect 3315 9216 3331 9280
rect 3395 9216 3411 9280
rect 3475 9216 3481 9280
rect 3165 9215 3481 9216
rect 7604 9280 7920 9281
rect 7604 9216 7610 9280
rect 7674 9216 7690 9280
rect 7754 9216 7770 9280
rect 7834 9216 7850 9280
rect 7914 9216 7920 9280
rect 7604 9215 7920 9216
rect 12043 9280 12359 9281
rect 12043 9216 12049 9280
rect 12113 9216 12129 9280
rect 12193 9216 12209 9280
rect 12273 9216 12289 9280
rect 12353 9216 12359 9280
rect 12043 9215 12359 9216
rect 16482 9280 16798 9281
rect 16482 9216 16488 9280
rect 16552 9216 16568 9280
rect 16632 9216 16648 9280
rect 16712 9216 16728 9280
rect 16792 9216 16798 9280
rect 16482 9215 16798 9216
rect 12249 8802 12315 8805
rect 13997 8802 14063 8805
rect 12249 8800 14063 8802
rect 12249 8744 12254 8800
rect 12310 8744 14002 8800
rect 14058 8744 14063 8800
rect 12249 8742 14063 8744
rect 12249 8739 12315 8742
rect 13997 8739 14063 8742
rect 5384 8736 5700 8737
rect 5384 8672 5390 8736
rect 5454 8672 5470 8736
rect 5534 8672 5550 8736
rect 5614 8672 5630 8736
rect 5694 8672 5700 8736
rect 5384 8671 5700 8672
rect 9823 8736 10139 8737
rect 9823 8672 9829 8736
rect 9893 8672 9909 8736
rect 9973 8672 9989 8736
rect 10053 8672 10069 8736
rect 10133 8672 10139 8736
rect 9823 8671 10139 8672
rect 14262 8736 14578 8737
rect 14262 8672 14268 8736
rect 14332 8672 14348 8736
rect 14412 8672 14428 8736
rect 14492 8672 14508 8736
rect 14572 8672 14578 8736
rect 14262 8671 14578 8672
rect 18701 8736 19017 8737
rect 18701 8672 18707 8736
rect 18771 8672 18787 8736
rect 18851 8672 18867 8736
rect 18931 8672 18947 8736
rect 19011 8672 19017 8736
rect 18701 8671 19017 8672
rect 3165 8192 3481 8193
rect 3165 8128 3171 8192
rect 3235 8128 3251 8192
rect 3315 8128 3331 8192
rect 3395 8128 3411 8192
rect 3475 8128 3481 8192
rect 3165 8127 3481 8128
rect 7604 8192 7920 8193
rect 7604 8128 7610 8192
rect 7674 8128 7690 8192
rect 7754 8128 7770 8192
rect 7834 8128 7850 8192
rect 7914 8128 7920 8192
rect 7604 8127 7920 8128
rect 12043 8192 12359 8193
rect 12043 8128 12049 8192
rect 12113 8128 12129 8192
rect 12193 8128 12209 8192
rect 12273 8128 12289 8192
rect 12353 8128 12359 8192
rect 12043 8127 12359 8128
rect 16482 8192 16798 8193
rect 16482 8128 16488 8192
rect 16552 8128 16568 8192
rect 16632 8128 16648 8192
rect 16712 8128 16728 8192
rect 16792 8128 16798 8192
rect 16482 8127 16798 8128
rect 5384 7648 5700 7649
rect 5384 7584 5390 7648
rect 5454 7584 5470 7648
rect 5534 7584 5550 7648
rect 5614 7584 5630 7648
rect 5694 7584 5700 7648
rect 5384 7583 5700 7584
rect 9823 7648 10139 7649
rect 9823 7584 9829 7648
rect 9893 7584 9909 7648
rect 9973 7584 9989 7648
rect 10053 7584 10069 7648
rect 10133 7584 10139 7648
rect 9823 7583 10139 7584
rect 14262 7648 14578 7649
rect 14262 7584 14268 7648
rect 14332 7584 14348 7648
rect 14412 7584 14428 7648
rect 14492 7584 14508 7648
rect 14572 7584 14578 7648
rect 14262 7583 14578 7584
rect 18701 7648 19017 7649
rect 18701 7584 18707 7648
rect 18771 7584 18787 7648
rect 18851 7584 18867 7648
rect 18931 7584 18947 7648
rect 19011 7584 19017 7648
rect 18701 7583 19017 7584
rect 3165 7104 3481 7105
rect 3165 7040 3171 7104
rect 3235 7040 3251 7104
rect 3315 7040 3331 7104
rect 3395 7040 3411 7104
rect 3475 7040 3481 7104
rect 3165 7039 3481 7040
rect 7604 7104 7920 7105
rect 7604 7040 7610 7104
rect 7674 7040 7690 7104
rect 7754 7040 7770 7104
rect 7834 7040 7850 7104
rect 7914 7040 7920 7104
rect 7604 7039 7920 7040
rect 12043 7104 12359 7105
rect 12043 7040 12049 7104
rect 12113 7040 12129 7104
rect 12193 7040 12209 7104
rect 12273 7040 12289 7104
rect 12353 7040 12359 7104
rect 12043 7039 12359 7040
rect 16482 7104 16798 7105
rect 16482 7040 16488 7104
rect 16552 7040 16568 7104
rect 16632 7040 16648 7104
rect 16712 7040 16728 7104
rect 16792 7040 16798 7104
rect 16482 7039 16798 7040
rect 5384 6560 5700 6561
rect 5384 6496 5390 6560
rect 5454 6496 5470 6560
rect 5534 6496 5550 6560
rect 5614 6496 5630 6560
rect 5694 6496 5700 6560
rect 5384 6495 5700 6496
rect 9823 6560 10139 6561
rect 9823 6496 9829 6560
rect 9893 6496 9909 6560
rect 9973 6496 9989 6560
rect 10053 6496 10069 6560
rect 10133 6496 10139 6560
rect 9823 6495 10139 6496
rect 14262 6560 14578 6561
rect 14262 6496 14268 6560
rect 14332 6496 14348 6560
rect 14412 6496 14428 6560
rect 14492 6496 14508 6560
rect 14572 6496 14578 6560
rect 14262 6495 14578 6496
rect 18701 6560 19017 6561
rect 18701 6496 18707 6560
rect 18771 6496 18787 6560
rect 18851 6496 18867 6560
rect 18931 6496 18947 6560
rect 19011 6496 19017 6560
rect 18701 6495 19017 6496
rect 3165 6016 3481 6017
rect 3165 5952 3171 6016
rect 3235 5952 3251 6016
rect 3315 5952 3331 6016
rect 3395 5952 3411 6016
rect 3475 5952 3481 6016
rect 3165 5951 3481 5952
rect 7604 6016 7920 6017
rect 7604 5952 7610 6016
rect 7674 5952 7690 6016
rect 7754 5952 7770 6016
rect 7834 5952 7850 6016
rect 7914 5952 7920 6016
rect 7604 5951 7920 5952
rect 12043 6016 12359 6017
rect 12043 5952 12049 6016
rect 12113 5952 12129 6016
rect 12193 5952 12209 6016
rect 12273 5952 12289 6016
rect 12353 5952 12359 6016
rect 12043 5951 12359 5952
rect 16482 6016 16798 6017
rect 16482 5952 16488 6016
rect 16552 5952 16568 6016
rect 16632 5952 16648 6016
rect 16712 5952 16728 6016
rect 16792 5952 16798 6016
rect 16482 5951 16798 5952
rect 5384 5472 5700 5473
rect 5384 5408 5390 5472
rect 5454 5408 5470 5472
rect 5534 5408 5550 5472
rect 5614 5408 5630 5472
rect 5694 5408 5700 5472
rect 5384 5407 5700 5408
rect 9823 5472 10139 5473
rect 9823 5408 9829 5472
rect 9893 5408 9909 5472
rect 9973 5408 9989 5472
rect 10053 5408 10069 5472
rect 10133 5408 10139 5472
rect 9823 5407 10139 5408
rect 14262 5472 14578 5473
rect 14262 5408 14268 5472
rect 14332 5408 14348 5472
rect 14412 5408 14428 5472
rect 14492 5408 14508 5472
rect 14572 5408 14578 5472
rect 14262 5407 14578 5408
rect 18701 5472 19017 5473
rect 18701 5408 18707 5472
rect 18771 5408 18787 5472
rect 18851 5408 18867 5472
rect 18931 5408 18947 5472
rect 19011 5408 19017 5472
rect 18701 5407 19017 5408
rect 3165 4928 3481 4929
rect 3165 4864 3171 4928
rect 3235 4864 3251 4928
rect 3315 4864 3331 4928
rect 3395 4864 3411 4928
rect 3475 4864 3481 4928
rect 3165 4863 3481 4864
rect 7604 4928 7920 4929
rect 7604 4864 7610 4928
rect 7674 4864 7690 4928
rect 7754 4864 7770 4928
rect 7834 4864 7850 4928
rect 7914 4864 7920 4928
rect 7604 4863 7920 4864
rect 12043 4928 12359 4929
rect 12043 4864 12049 4928
rect 12113 4864 12129 4928
rect 12193 4864 12209 4928
rect 12273 4864 12289 4928
rect 12353 4864 12359 4928
rect 12043 4863 12359 4864
rect 16482 4928 16798 4929
rect 16482 4864 16488 4928
rect 16552 4864 16568 4928
rect 16632 4864 16648 4928
rect 16712 4864 16728 4928
rect 16792 4864 16798 4928
rect 16482 4863 16798 4864
rect 5384 4384 5700 4385
rect 5384 4320 5390 4384
rect 5454 4320 5470 4384
rect 5534 4320 5550 4384
rect 5614 4320 5630 4384
rect 5694 4320 5700 4384
rect 5384 4319 5700 4320
rect 9823 4384 10139 4385
rect 9823 4320 9829 4384
rect 9893 4320 9909 4384
rect 9973 4320 9989 4384
rect 10053 4320 10069 4384
rect 10133 4320 10139 4384
rect 9823 4319 10139 4320
rect 14262 4384 14578 4385
rect 14262 4320 14268 4384
rect 14332 4320 14348 4384
rect 14412 4320 14428 4384
rect 14492 4320 14508 4384
rect 14572 4320 14578 4384
rect 14262 4319 14578 4320
rect 18701 4384 19017 4385
rect 18701 4320 18707 4384
rect 18771 4320 18787 4384
rect 18851 4320 18867 4384
rect 18931 4320 18947 4384
rect 19011 4320 19017 4384
rect 18701 4319 19017 4320
rect 3165 3840 3481 3841
rect 3165 3776 3171 3840
rect 3235 3776 3251 3840
rect 3315 3776 3331 3840
rect 3395 3776 3411 3840
rect 3475 3776 3481 3840
rect 3165 3775 3481 3776
rect 7604 3840 7920 3841
rect 7604 3776 7610 3840
rect 7674 3776 7690 3840
rect 7754 3776 7770 3840
rect 7834 3776 7850 3840
rect 7914 3776 7920 3840
rect 7604 3775 7920 3776
rect 12043 3840 12359 3841
rect 12043 3776 12049 3840
rect 12113 3776 12129 3840
rect 12193 3776 12209 3840
rect 12273 3776 12289 3840
rect 12353 3776 12359 3840
rect 12043 3775 12359 3776
rect 16482 3840 16798 3841
rect 16482 3776 16488 3840
rect 16552 3776 16568 3840
rect 16632 3776 16648 3840
rect 16712 3776 16728 3840
rect 16792 3776 16798 3840
rect 16482 3775 16798 3776
rect 5384 3296 5700 3297
rect 5384 3232 5390 3296
rect 5454 3232 5470 3296
rect 5534 3232 5550 3296
rect 5614 3232 5630 3296
rect 5694 3232 5700 3296
rect 5384 3231 5700 3232
rect 9823 3296 10139 3297
rect 9823 3232 9829 3296
rect 9893 3232 9909 3296
rect 9973 3232 9989 3296
rect 10053 3232 10069 3296
rect 10133 3232 10139 3296
rect 9823 3231 10139 3232
rect 14262 3296 14578 3297
rect 14262 3232 14268 3296
rect 14332 3232 14348 3296
rect 14412 3232 14428 3296
rect 14492 3232 14508 3296
rect 14572 3232 14578 3296
rect 14262 3231 14578 3232
rect 18701 3296 19017 3297
rect 18701 3232 18707 3296
rect 18771 3232 18787 3296
rect 18851 3232 18867 3296
rect 18931 3232 18947 3296
rect 19011 3232 19017 3296
rect 18701 3231 19017 3232
rect 3165 2752 3481 2753
rect 3165 2688 3171 2752
rect 3235 2688 3251 2752
rect 3315 2688 3331 2752
rect 3395 2688 3411 2752
rect 3475 2688 3481 2752
rect 3165 2687 3481 2688
rect 7604 2752 7920 2753
rect 7604 2688 7610 2752
rect 7674 2688 7690 2752
rect 7754 2688 7770 2752
rect 7834 2688 7850 2752
rect 7914 2688 7920 2752
rect 7604 2687 7920 2688
rect 12043 2752 12359 2753
rect 12043 2688 12049 2752
rect 12113 2688 12129 2752
rect 12193 2688 12209 2752
rect 12273 2688 12289 2752
rect 12353 2688 12359 2752
rect 12043 2687 12359 2688
rect 16482 2752 16798 2753
rect 16482 2688 16488 2752
rect 16552 2688 16568 2752
rect 16632 2688 16648 2752
rect 16712 2688 16728 2752
rect 16792 2688 16798 2752
rect 16482 2687 16798 2688
rect 5384 2208 5700 2209
rect 5384 2144 5390 2208
rect 5454 2144 5470 2208
rect 5534 2144 5550 2208
rect 5614 2144 5630 2208
rect 5694 2144 5700 2208
rect 5384 2143 5700 2144
rect 9823 2208 10139 2209
rect 9823 2144 9829 2208
rect 9893 2144 9909 2208
rect 9973 2144 9989 2208
rect 10053 2144 10069 2208
rect 10133 2144 10139 2208
rect 9823 2143 10139 2144
rect 14262 2208 14578 2209
rect 14262 2144 14268 2208
rect 14332 2144 14348 2208
rect 14412 2144 14428 2208
rect 14492 2144 14508 2208
rect 14572 2144 14578 2208
rect 14262 2143 14578 2144
rect 18701 2208 19017 2209
rect 18701 2144 18707 2208
rect 18771 2144 18787 2208
rect 18851 2144 18867 2208
rect 18931 2144 18947 2208
rect 19011 2144 19017 2208
rect 18701 2143 19017 2144
<< via3 >>
rect 5390 17436 5454 17440
rect 5390 17380 5394 17436
rect 5394 17380 5450 17436
rect 5450 17380 5454 17436
rect 5390 17376 5454 17380
rect 5470 17436 5534 17440
rect 5470 17380 5474 17436
rect 5474 17380 5530 17436
rect 5530 17380 5534 17436
rect 5470 17376 5534 17380
rect 5550 17436 5614 17440
rect 5550 17380 5554 17436
rect 5554 17380 5610 17436
rect 5610 17380 5614 17436
rect 5550 17376 5614 17380
rect 5630 17436 5694 17440
rect 5630 17380 5634 17436
rect 5634 17380 5690 17436
rect 5690 17380 5694 17436
rect 5630 17376 5694 17380
rect 9829 17436 9893 17440
rect 9829 17380 9833 17436
rect 9833 17380 9889 17436
rect 9889 17380 9893 17436
rect 9829 17376 9893 17380
rect 9909 17436 9973 17440
rect 9909 17380 9913 17436
rect 9913 17380 9969 17436
rect 9969 17380 9973 17436
rect 9909 17376 9973 17380
rect 9989 17436 10053 17440
rect 9989 17380 9993 17436
rect 9993 17380 10049 17436
rect 10049 17380 10053 17436
rect 9989 17376 10053 17380
rect 10069 17436 10133 17440
rect 10069 17380 10073 17436
rect 10073 17380 10129 17436
rect 10129 17380 10133 17436
rect 10069 17376 10133 17380
rect 14268 17436 14332 17440
rect 14268 17380 14272 17436
rect 14272 17380 14328 17436
rect 14328 17380 14332 17436
rect 14268 17376 14332 17380
rect 14348 17436 14412 17440
rect 14348 17380 14352 17436
rect 14352 17380 14408 17436
rect 14408 17380 14412 17436
rect 14348 17376 14412 17380
rect 14428 17436 14492 17440
rect 14428 17380 14432 17436
rect 14432 17380 14488 17436
rect 14488 17380 14492 17436
rect 14428 17376 14492 17380
rect 14508 17436 14572 17440
rect 14508 17380 14512 17436
rect 14512 17380 14568 17436
rect 14568 17380 14572 17436
rect 14508 17376 14572 17380
rect 18707 17436 18771 17440
rect 18707 17380 18711 17436
rect 18711 17380 18767 17436
rect 18767 17380 18771 17436
rect 18707 17376 18771 17380
rect 18787 17436 18851 17440
rect 18787 17380 18791 17436
rect 18791 17380 18847 17436
rect 18847 17380 18851 17436
rect 18787 17376 18851 17380
rect 18867 17436 18931 17440
rect 18867 17380 18871 17436
rect 18871 17380 18927 17436
rect 18927 17380 18931 17436
rect 18867 17376 18931 17380
rect 18947 17436 19011 17440
rect 18947 17380 18951 17436
rect 18951 17380 19007 17436
rect 19007 17380 19011 17436
rect 18947 17376 19011 17380
rect 3171 16892 3235 16896
rect 3171 16836 3175 16892
rect 3175 16836 3231 16892
rect 3231 16836 3235 16892
rect 3171 16832 3235 16836
rect 3251 16892 3315 16896
rect 3251 16836 3255 16892
rect 3255 16836 3311 16892
rect 3311 16836 3315 16892
rect 3251 16832 3315 16836
rect 3331 16892 3395 16896
rect 3331 16836 3335 16892
rect 3335 16836 3391 16892
rect 3391 16836 3395 16892
rect 3331 16832 3395 16836
rect 3411 16892 3475 16896
rect 3411 16836 3415 16892
rect 3415 16836 3471 16892
rect 3471 16836 3475 16892
rect 3411 16832 3475 16836
rect 7610 16892 7674 16896
rect 7610 16836 7614 16892
rect 7614 16836 7670 16892
rect 7670 16836 7674 16892
rect 7610 16832 7674 16836
rect 7690 16892 7754 16896
rect 7690 16836 7694 16892
rect 7694 16836 7750 16892
rect 7750 16836 7754 16892
rect 7690 16832 7754 16836
rect 7770 16892 7834 16896
rect 7770 16836 7774 16892
rect 7774 16836 7830 16892
rect 7830 16836 7834 16892
rect 7770 16832 7834 16836
rect 7850 16892 7914 16896
rect 7850 16836 7854 16892
rect 7854 16836 7910 16892
rect 7910 16836 7914 16892
rect 7850 16832 7914 16836
rect 12049 16892 12113 16896
rect 12049 16836 12053 16892
rect 12053 16836 12109 16892
rect 12109 16836 12113 16892
rect 12049 16832 12113 16836
rect 12129 16892 12193 16896
rect 12129 16836 12133 16892
rect 12133 16836 12189 16892
rect 12189 16836 12193 16892
rect 12129 16832 12193 16836
rect 12209 16892 12273 16896
rect 12209 16836 12213 16892
rect 12213 16836 12269 16892
rect 12269 16836 12273 16892
rect 12209 16832 12273 16836
rect 12289 16892 12353 16896
rect 12289 16836 12293 16892
rect 12293 16836 12349 16892
rect 12349 16836 12353 16892
rect 12289 16832 12353 16836
rect 16488 16892 16552 16896
rect 16488 16836 16492 16892
rect 16492 16836 16548 16892
rect 16548 16836 16552 16892
rect 16488 16832 16552 16836
rect 16568 16892 16632 16896
rect 16568 16836 16572 16892
rect 16572 16836 16628 16892
rect 16628 16836 16632 16892
rect 16568 16832 16632 16836
rect 16648 16892 16712 16896
rect 16648 16836 16652 16892
rect 16652 16836 16708 16892
rect 16708 16836 16712 16892
rect 16648 16832 16712 16836
rect 16728 16892 16792 16896
rect 16728 16836 16732 16892
rect 16732 16836 16788 16892
rect 16788 16836 16792 16892
rect 16728 16832 16792 16836
rect 5390 16348 5454 16352
rect 5390 16292 5394 16348
rect 5394 16292 5450 16348
rect 5450 16292 5454 16348
rect 5390 16288 5454 16292
rect 5470 16348 5534 16352
rect 5470 16292 5474 16348
rect 5474 16292 5530 16348
rect 5530 16292 5534 16348
rect 5470 16288 5534 16292
rect 5550 16348 5614 16352
rect 5550 16292 5554 16348
rect 5554 16292 5610 16348
rect 5610 16292 5614 16348
rect 5550 16288 5614 16292
rect 5630 16348 5694 16352
rect 5630 16292 5634 16348
rect 5634 16292 5690 16348
rect 5690 16292 5694 16348
rect 5630 16288 5694 16292
rect 9829 16348 9893 16352
rect 9829 16292 9833 16348
rect 9833 16292 9889 16348
rect 9889 16292 9893 16348
rect 9829 16288 9893 16292
rect 9909 16348 9973 16352
rect 9909 16292 9913 16348
rect 9913 16292 9969 16348
rect 9969 16292 9973 16348
rect 9909 16288 9973 16292
rect 9989 16348 10053 16352
rect 9989 16292 9993 16348
rect 9993 16292 10049 16348
rect 10049 16292 10053 16348
rect 9989 16288 10053 16292
rect 10069 16348 10133 16352
rect 10069 16292 10073 16348
rect 10073 16292 10129 16348
rect 10129 16292 10133 16348
rect 10069 16288 10133 16292
rect 14268 16348 14332 16352
rect 14268 16292 14272 16348
rect 14272 16292 14328 16348
rect 14328 16292 14332 16348
rect 14268 16288 14332 16292
rect 14348 16348 14412 16352
rect 14348 16292 14352 16348
rect 14352 16292 14408 16348
rect 14408 16292 14412 16348
rect 14348 16288 14412 16292
rect 14428 16348 14492 16352
rect 14428 16292 14432 16348
rect 14432 16292 14488 16348
rect 14488 16292 14492 16348
rect 14428 16288 14492 16292
rect 14508 16348 14572 16352
rect 14508 16292 14512 16348
rect 14512 16292 14568 16348
rect 14568 16292 14572 16348
rect 14508 16288 14572 16292
rect 18707 16348 18771 16352
rect 18707 16292 18711 16348
rect 18711 16292 18767 16348
rect 18767 16292 18771 16348
rect 18707 16288 18771 16292
rect 18787 16348 18851 16352
rect 18787 16292 18791 16348
rect 18791 16292 18847 16348
rect 18847 16292 18851 16348
rect 18787 16288 18851 16292
rect 18867 16348 18931 16352
rect 18867 16292 18871 16348
rect 18871 16292 18927 16348
rect 18927 16292 18931 16348
rect 18867 16288 18931 16292
rect 18947 16348 19011 16352
rect 18947 16292 18951 16348
rect 18951 16292 19007 16348
rect 19007 16292 19011 16348
rect 18947 16288 19011 16292
rect 3171 15804 3235 15808
rect 3171 15748 3175 15804
rect 3175 15748 3231 15804
rect 3231 15748 3235 15804
rect 3171 15744 3235 15748
rect 3251 15804 3315 15808
rect 3251 15748 3255 15804
rect 3255 15748 3311 15804
rect 3311 15748 3315 15804
rect 3251 15744 3315 15748
rect 3331 15804 3395 15808
rect 3331 15748 3335 15804
rect 3335 15748 3391 15804
rect 3391 15748 3395 15804
rect 3331 15744 3395 15748
rect 3411 15804 3475 15808
rect 3411 15748 3415 15804
rect 3415 15748 3471 15804
rect 3471 15748 3475 15804
rect 3411 15744 3475 15748
rect 7610 15804 7674 15808
rect 7610 15748 7614 15804
rect 7614 15748 7670 15804
rect 7670 15748 7674 15804
rect 7610 15744 7674 15748
rect 7690 15804 7754 15808
rect 7690 15748 7694 15804
rect 7694 15748 7750 15804
rect 7750 15748 7754 15804
rect 7690 15744 7754 15748
rect 7770 15804 7834 15808
rect 7770 15748 7774 15804
rect 7774 15748 7830 15804
rect 7830 15748 7834 15804
rect 7770 15744 7834 15748
rect 7850 15804 7914 15808
rect 7850 15748 7854 15804
rect 7854 15748 7910 15804
rect 7910 15748 7914 15804
rect 7850 15744 7914 15748
rect 12049 15804 12113 15808
rect 12049 15748 12053 15804
rect 12053 15748 12109 15804
rect 12109 15748 12113 15804
rect 12049 15744 12113 15748
rect 12129 15804 12193 15808
rect 12129 15748 12133 15804
rect 12133 15748 12189 15804
rect 12189 15748 12193 15804
rect 12129 15744 12193 15748
rect 12209 15804 12273 15808
rect 12209 15748 12213 15804
rect 12213 15748 12269 15804
rect 12269 15748 12273 15804
rect 12209 15744 12273 15748
rect 12289 15804 12353 15808
rect 12289 15748 12293 15804
rect 12293 15748 12349 15804
rect 12349 15748 12353 15804
rect 12289 15744 12353 15748
rect 16488 15804 16552 15808
rect 16488 15748 16492 15804
rect 16492 15748 16548 15804
rect 16548 15748 16552 15804
rect 16488 15744 16552 15748
rect 16568 15804 16632 15808
rect 16568 15748 16572 15804
rect 16572 15748 16628 15804
rect 16628 15748 16632 15804
rect 16568 15744 16632 15748
rect 16648 15804 16712 15808
rect 16648 15748 16652 15804
rect 16652 15748 16708 15804
rect 16708 15748 16712 15804
rect 16648 15744 16712 15748
rect 16728 15804 16792 15808
rect 16728 15748 16732 15804
rect 16732 15748 16788 15804
rect 16788 15748 16792 15804
rect 16728 15744 16792 15748
rect 5390 15260 5454 15264
rect 5390 15204 5394 15260
rect 5394 15204 5450 15260
rect 5450 15204 5454 15260
rect 5390 15200 5454 15204
rect 5470 15260 5534 15264
rect 5470 15204 5474 15260
rect 5474 15204 5530 15260
rect 5530 15204 5534 15260
rect 5470 15200 5534 15204
rect 5550 15260 5614 15264
rect 5550 15204 5554 15260
rect 5554 15204 5610 15260
rect 5610 15204 5614 15260
rect 5550 15200 5614 15204
rect 5630 15260 5694 15264
rect 5630 15204 5634 15260
rect 5634 15204 5690 15260
rect 5690 15204 5694 15260
rect 5630 15200 5694 15204
rect 9829 15260 9893 15264
rect 9829 15204 9833 15260
rect 9833 15204 9889 15260
rect 9889 15204 9893 15260
rect 9829 15200 9893 15204
rect 9909 15260 9973 15264
rect 9909 15204 9913 15260
rect 9913 15204 9969 15260
rect 9969 15204 9973 15260
rect 9909 15200 9973 15204
rect 9989 15260 10053 15264
rect 9989 15204 9993 15260
rect 9993 15204 10049 15260
rect 10049 15204 10053 15260
rect 9989 15200 10053 15204
rect 10069 15260 10133 15264
rect 10069 15204 10073 15260
rect 10073 15204 10129 15260
rect 10129 15204 10133 15260
rect 10069 15200 10133 15204
rect 14268 15260 14332 15264
rect 14268 15204 14272 15260
rect 14272 15204 14328 15260
rect 14328 15204 14332 15260
rect 14268 15200 14332 15204
rect 14348 15260 14412 15264
rect 14348 15204 14352 15260
rect 14352 15204 14408 15260
rect 14408 15204 14412 15260
rect 14348 15200 14412 15204
rect 14428 15260 14492 15264
rect 14428 15204 14432 15260
rect 14432 15204 14488 15260
rect 14488 15204 14492 15260
rect 14428 15200 14492 15204
rect 14508 15260 14572 15264
rect 14508 15204 14512 15260
rect 14512 15204 14568 15260
rect 14568 15204 14572 15260
rect 14508 15200 14572 15204
rect 18707 15260 18771 15264
rect 18707 15204 18711 15260
rect 18711 15204 18767 15260
rect 18767 15204 18771 15260
rect 18707 15200 18771 15204
rect 18787 15260 18851 15264
rect 18787 15204 18791 15260
rect 18791 15204 18847 15260
rect 18847 15204 18851 15260
rect 18787 15200 18851 15204
rect 18867 15260 18931 15264
rect 18867 15204 18871 15260
rect 18871 15204 18927 15260
rect 18927 15204 18931 15260
rect 18867 15200 18931 15204
rect 18947 15260 19011 15264
rect 18947 15204 18951 15260
rect 18951 15204 19007 15260
rect 19007 15204 19011 15260
rect 18947 15200 19011 15204
rect 3171 14716 3235 14720
rect 3171 14660 3175 14716
rect 3175 14660 3231 14716
rect 3231 14660 3235 14716
rect 3171 14656 3235 14660
rect 3251 14716 3315 14720
rect 3251 14660 3255 14716
rect 3255 14660 3311 14716
rect 3311 14660 3315 14716
rect 3251 14656 3315 14660
rect 3331 14716 3395 14720
rect 3331 14660 3335 14716
rect 3335 14660 3391 14716
rect 3391 14660 3395 14716
rect 3331 14656 3395 14660
rect 3411 14716 3475 14720
rect 3411 14660 3415 14716
rect 3415 14660 3471 14716
rect 3471 14660 3475 14716
rect 3411 14656 3475 14660
rect 7610 14716 7674 14720
rect 7610 14660 7614 14716
rect 7614 14660 7670 14716
rect 7670 14660 7674 14716
rect 7610 14656 7674 14660
rect 7690 14716 7754 14720
rect 7690 14660 7694 14716
rect 7694 14660 7750 14716
rect 7750 14660 7754 14716
rect 7690 14656 7754 14660
rect 7770 14716 7834 14720
rect 7770 14660 7774 14716
rect 7774 14660 7830 14716
rect 7830 14660 7834 14716
rect 7770 14656 7834 14660
rect 7850 14716 7914 14720
rect 7850 14660 7854 14716
rect 7854 14660 7910 14716
rect 7910 14660 7914 14716
rect 7850 14656 7914 14660
rect 12049 14716 12113 14720
rect 12049 14660 12053 14716
rect 12053 14660 12109 14716
rect 12109 14660 12113 14716
rect 12049 14656 12113 14660
rect 12129 14716 12193 14720
rect 12129 14660 12133 14716
rect 12133 14660 12189 14716
rect 12189 14660 12193 14716
rect 12129 14656 12193 14660
rect 12209 14716 12273 14720
rect 12209 14660 12213 14716
rect 12213 14660 12269 14716
rect 12269 14660 12273 14716
rect 12209 14656 12273 14660
rect 12289 14716 12353 14720
rect 12289 14660 12293 14716
rect 12293 14660 12349 14716
rect 12349 14660 12353 14716
rect 12289 14656 12353 14660
rect 16488 14716 16552 14720
rect 16488 14660 16492 14716
rect 16492 14660 16548 14716
rect 16548 14660 16552 14716
rect 16488 14656 16552 14660
rect 16568 14716 16632 14720
rect 16568 14660 16572 14716
rect 16572 14660 16628 14716
rect 16628 14660 16632 14716
rect 16568 14656 16632 14660
rect 16648 14716 16712 14720
rect 16648 14660 16652 14716
rect 16652 14660 16708 14716
rect 16708 14660 16712 14716
rect 16648 14656 16712 14660
rect 16728 14716 16792 14720
rect 16728 14660 16732 14716
rect 16732 14660 16788 14716
rect 16788 14660 16792 14716
rect 16728 14656 16792 14660
rect 5390 14172 5454 14176
rect 5390 14116 5394 14172
rect 5394 14116 5450 14172
rect 5450 14116 5454 14172
rect 5390 14112 5454 14116
rect 5470 14172 5534 14176
rect 5470 14116 5474 14172
rect 5474 14116 5530 14172
rect 5530 14116 5534 14172
rect 5470 14112 5534 14116
rect 5550 14172 5614 14176
rect 5550 14116 5554 14172
rect 5554 14116 5610 14172
rect 5610 14116 5614 14172
rect 5550 14112 5614 14116
rect 5630 14172 5694 14176
rect 5630 14116 5634 14172
rect 5634 14116 5690 14172
rect 5690 14116 5694 14172
rect 5630 14112 5694 14116
rect 9829 14172 9893 14176
rect 9829 14116 9833 14172
rect 9833 14116 9889 14172
rect 9889 14116 9893 14172
rect 9829 14112 9893 14116
rect 9909 14172 9973 14176
rect 9909 14116 9913 14172
rect 9913 14116 9969 14172
rect 9969 14116 9973 14172
rect 9909 14112 9973 14116
rect 9989 14172 10053 14176
rect 9989 14116 9993 14172
rect 9993 14116 10049 14172
rect 10049 14116 10053 14172
rect 9989 14112 10053 14116
rect 10069 14172 10133 14176
rect 10069 14116 10073 14172
rect 10073 14116 10129 14172
rect 10129 14116 10133 14172
rect 10069 14112 10133 14116
rect 14268 14172 14332 14176
rect 14268 14116 14272 14172
rect 14272 14116 14328 14172
rect 14328 14116 14332 14172
rect 14268 14112 14332 14116
rect 14348 14172 14412 14176
rect 14348 14116 14352 14172
rect 14352 14116 14408 14172
rect 14408 14116 14412 14172
rect 14348 14112 14412 14116
rect 14428 14172 14492 14176
rect 14428 14116 14432 14172
rect 14432 14116 14488 14172
rect 14488 14116 14492 14172
rect 14428 14112 14492 14116
rect 14508 14172 14572 14176
rect 14508 14116 14512 14172
rect 14512 14116 14568 14172
rect 14568 14116 14572 14172
rect 14508 14112 14572 14116
rect 18707 14172 18771 14176
rect 18707 14116 18711 14172
rect 18711 14116 18767 14172
rect 18767 14116 18771 14172
rect 18707 14112 18771 14116
rect 18787 14172 18851 14176
rect 18787 14116 18791 14172
rect 18791 14116 18847 14172
rect 18847 14116 18851 14172
rect 18787 14112 18851 14116
rect 18867 14172 18931 14176
rect 18867 14116 18871 14172
rect 18871 14116 18927 14172
rect 18927 14116 18931 14172
rect 18867 14112 18931 14116
rect 18947 14172 19011 14176
rect 18947 14116 18951 14172
rect 18951 14116 19007 14172
rect 19007 14116 19011 14172
rect 18947 14112 19011 14116
rect 3171 13628 3235 13632
rect 3171 13572 3175 13628
rect 3175 13572 3231 13628
rect 3231 13572 3235 13628
rect 3171 13568 3235 13572
rect 3251 13628 3315 13632
rect 3251 13572 3255 13628
rect 3255 13572 3311 13628
rect 3311 13572 3315 13628
rect 3251 13568 3315 13572
rect 3331 13628 3395 13632
rect 3331 13572 3335 13628
rect 3335 13572 3391 13628
rect 3391 13572 3395 13628
rect 3331 13568 3395 13572
rect 3411 13628 3475 13632
rect 3411 13572 3415 13628
rect 3415 13572 3471 13628
rect 3471 13572 3475 13628
rect 3411 13568 3475 13572
rect 7610 13628 7674 13632
rect 7610 13572 7614 13628
rect 7614 13572 7670 13628
rect 7670 13572 7674 13628
rect 7610 13568 7674 13572
rect 7690 13628 7754 13632
rect 7690 13572 7694 13628
rect 7694 13572 7750 13628
rect 7750 13572 7754 13628
rect 7690 13568 7754 13572
rect 7770 13628 7834 13632
rect 7770 13572 7774 13628
rect 7774 13572 7830 13628
rect 7830 13572 7834 13628
rect 7770 13568 7834 13572
rect 7850 13628 7914 13632
rect 7850 13572 7854 13628
rect 7854 13572 7910 13628
rect 7910 13572 7914 13628
rect 7850 13568 7914 13572
rect 12049 13628 12113 13632
rect 12049 13572 12053 13628
rect 12053 13572 12109 13628
rect 12109 13572 12113 13628
rect 12049 13568 12113 13572
rect 12129 13628 12193 13632
rect 12129 13572 12133 13628
rect 12133 13572 12189 13628
rect 12189 13572 12193 13628
rect 12129 13568 12193 13572
rect 12209 13628 12273 13632
rect 12209 13572 12213 13628
rect 12213 13572 12269 13628
rect 12269 13572 12273 13628
rect 12209 13568 12273 13572
rect 12289 13628 12353 13632
rect 12289 13572 12293 13628
rect 12293 13572 12349 13628
rect 12349 13572 12353 13628
rect 12289 13568 12353 13572
rect 16488 13628 16552 13632
rect 16488 13572 16492 13628
rect 16492 13572 16548 13628
rect 16548 13572 16552 13628
rect 16488 13568 16552 13572
rect 16568 13628 16632 13632
rect 16568 13572 16572 13628
rect 16572 13572 16628 13628
rect 16628 13572 16632 13628
rect 16568 13568 16632 13572
rect 16648 13628 16712 13632
rect 16648 13572 16652 13628
rect 16652 13572 16708 13628
rect 16708 13572 16712 13628
rect 16648 13568 16712 13572
rect 16728 13628 16792 13632
rect 16728 13572 16732 13628
rect 16732 13572 16788 13628
rect 16788 13572 16792 13628
rect 16728 13568 16792 13572
rect 5390 13084 5454 13088
rect 5390 13028 5394 13084
rect 5394 13028 5450 13084
rect 5450 13028 5454 13084
rect 5390 13024 5454 13028
rect 5470 13084 5534 13088
rect 5470 13028 5474 13084
rect 5474 13028 5530 13084
rect 5530 13028 5534 13084
rect 5470 13024 5534 13028
rect 5550 13084 5614 13088
rect 5550 13028 5554 13084
rect 5554 13028 5610 13084
rect 5610 13028 5614 13084
rect 5550 13024 5614 13028
rect 5630 13084 5694 13088
rect 5630 13028 5634 13084
rect 5634 13028 5690 13084
rect 5690 13028 5694 13084
rect 5630 13024 5694 13028
rect 9829 13084 9893 13088
rect 9829 13028 9833 13084
rect 9833 13028 9889 13084
rect 9889 13028 9893 13084
rect 9829 13024 9893 13028
rect 9909 13084 9973 13088
rect 9909 13028 9913 13084
rect 9913 13028 9969 13084
rect 9969 13028 9973 13084
rect 9909 13024 9973 13028
rect 9989 13084 10053 13088
rect 9989 13028 9993 13084
rect 9993 13028 10049 13084
rect 10049 13028 10053 13084
rect 9989 13024 10053 13028
rect 10069 13084 10133 13088
rect 10069 13028 10073 13084
rect 10073 13028 10129 13084
rect 10129 13028 10133 13084
rect 10069 13024 10133 13028
rect 14268 13084 14332 13088
rect 14268 13028 14272 13084
rect 14272 13028 14328 13084
rect 14328 13028 14332 13084
rect 14268 13024 14332 13028
rect 14348 13084 14412 13088
rect 14348 13028 14352 13084
rect 14352 13028 14408 13084
rect 14408 13028 14412 13084
rect 14348 13024 14412 13028
rect 14428 13084 14492 13088
rect 14428 13028 14432 13084
rect 14432 13028 14488 13084
rect 14488 13028 14492 13084
rect 14428 13024 14492 13028
rect 14508 13084 14572 13088
rect 14508 13028 14512 13084
rect 14512 13028 14568 13084
rect 14568 13028 14572 13084
rect 14508 13024 14572 13028
rect 18707 13084 18771 13088
rect 18707 13028 18711 13084
rect 18711 13028 18767 13084
rect 18767 13028 18771 13084
rect 18707 13024 18771 13028
rect 18787 13084 18851 13088
rect 18787 13028 18791 13084
rect 18791 13028 18847 13084
rect 18847 13028 18851 13084
rect 18787 13024 18851 13028
rect 18867 13084 18931 13088
rect 18867 13028 18871 13084
rect 18871 13028 18927 13084
rect 18927 13028 18931 13084
rect 18867 13024 18931 13028
rect 18947 13084 19011 13088
rect 18947 13028 18951 13084
rect 18951 13028 19007 13084
rect 19007 13028 19011 13084
rect 18947 13024 19011 13028
rect 3171 12540 3235 12544
rect 3171 12484 3175 12540
rect 3175 12484 3231 12540
rect 3231 12484 3235 12540
rect 3171 12480 3235 12484
rect 3251 12540 3315 12544
rect 3251 12484 3255 12540
rect 3255 12484 3311 12540
rect 3311 12484 3315 12540
rect 3251 12480 3315 12484
rect 3331 12540 3395 12544
rect 3331 12484 3335 12540
rect 3335 12484 3391 12540
rect 3391 12484 3395 12540
rect 3331 12480 3395 12484
rect 3411 12540 3475 12544
rect 3411 12484 3415 12540
rect 3415 12484 3471 12540
rect 3471 12484 3475 12540
rect 3411 12480 3475 12484
rect 7610 12540 7674 12544
rect 7610 12484 7614 12540
rect 7614 12484 7670 12540
rect 7670 12484 7674 12540
rect 7610 12480 7674 12484
rect 7690 12540 7754 12544
rect 7690 12484 7694 12540
rect 7694 12484 7750 12540
rect 7750 12484 7754 12540
rect 7690 12480 7754 12484
rect 7770 12540 7834 12544
rect 7770 12484 7774 12540
rect 7774 12484 7830 12540
rect 7830 12484 7834 12540
rect 7770 12480 7834 12484
rect 7850 12540 7914 12544
rect 7850 12484 7854 12540
rect 7854 12484 7910 12540
rect 7910 12484 7914 12540
rect 7850 12480 7914 12484
rect 12049 12540 12113 12544
rect 12049 12484 12053 12540
rect 12053 12484 12109 12540
rect 12109 12484 12113 12540
rect 12049 12480 12113 12484
rect 12129 12540 12193 12544
rect 12129 12484 12133 12540
rect 12133 12484 12189 12540
rect 12189 12484 12193 12540
rect 12129 12480 12193 12484
rect 12209 12540 12273 12544
rect 12209 12484 12213 12540
rect 12213 12484 12269 12540
rect 12269 12484 12273 12540
rect 12209 12480 12273 12484
rect 12289 12540 12353 12544
rect 12289 12484 12293 12540
rect 12293 12484 12349 12540
rect 12349 12484 12353 12540
rect 12289 12480 12353 12484
rect 16488 12540 16552 12544
rect 16488 12484 16492 12540
rect 16492 12484 16548 12540
rect 16548 12484 16552 12540
rect 16488 12480 16552 12484
rect 16568 12540 16632 12544
rect 16568 12484 16572 12540
rect 16572 12484 16628 12540
rect 16628 12484 16632 12540
rect 16568 12480 16632 12484
rect 16648 12540 16712 12544
rect 16648 12484 16652 12540
rect 16652 12484 16708 12540
rect 16708 12484 16712 12540
rect 16648 12480 16712 12484
rect 16728 12540 16792 12544
rect 16728 12484 16732 12540
rect 16732 12484 16788 12540
rect 16788 12484 16792 12540
rect 16728 12480 16792 12484
rect 5390 11996 5454 12000
rect 5390 11940 5394 11996
rect 5394 11940 5450 11996
rect 5450 11940 5454 11996
rect 5390 11936 5454 11940
rect 5470 11996 5534 12000
rect 5470 11940 5474 11996
rect 5474 11940 5530 11996
rect 5530 11940 5534 11996
rect 5470 11936 5534 11940
rect 5550 11996 5614 12000
rect 5550 11940 5554 11996
rect 5554 11940 5610 11996
rect 5610 11940 5614 11996
rect 5550 11936 5614 11940
rect 5630 11996 5694 12000
rect 5630 11940 5634 11996
rect 5634 11940 5690 11996
rect 5690 11940 5694 11996
rect 5630 11936 5694 11940
rect 9829 11996 9893 12000
rect 9829 11940 9833 11996
rect 9833 11940 9889 11996
rect 9889 11940 9893 11996
rect 9829 11936 9893 11940
rect 9909 11996 9973 12000
rect 9909 11940 9913 11996
rect 9913 11940 9969 11996
rect 9969 11940 9973 11996
rect 9909 11936 9973 11940
rect 9989 11996 10053 12000
rect 9989 11940 9993 11996
rect 9993 11940 10049 11996
rect 10049 11940 10053 11996
rect 9989 11936 10053 11940
rect 10069 11996 10133 12000
rect 10069 11940 10073 11996
rect 10073 11940 10129 11996
rect 10129 11940 10133 11996
rect 10069 11936 10133 11940
rect 14268 11996 14332 12000
rect 14268 11940 14272 11996
rect 14272 11940 14328 11996
rect 14328 11940 14332 11996
rect 14268 11936 14332 11940
rect 14348 11996 14412 12000
rect 14348 11940 14352 11996
rect 14352 11940 14408 11996
rect 14408 11940 14412 11996
rect 14348 11936 14412 11940
rect 14428 11996 14492 12000
rect 14428 11940 14432 11996
rect 14432 11940 14488 11996
rect 14488 11940 14492 11996
rect 14428 11936 14492 11940
rect 14508 11996 14572 12000
rect 14508 11940 14512 11996
rect 14512 11940 14568 11996
rect 14568 11940 14572 11996
rect 14508 11936 14572 11940
rect 18707 11996 18771 12000
rect 18707 11940 18711 11996
rect 18711 11940 18767 11996
rect 18767 11940 18771 11996
rect 18707 11936 18771 11940
rect 18787 11996 18851 12000
rect 18787 11940 18791 11996
rect 18791 11940 18847 11996
rect 18847 11940 18851 11996
rect 18787 11936 18851 11940
rect 18867 11996 18931 12000
rect 18867 11940 18871 11996
rect 18871 11940 18927 11996
rect 18927 11940 18931 11996
rect 18867 11936 18931 11940
rect 18947 11996 19011 12000
rect 18947 11940 18951 11996
rect 18951 11940 19007 11996
rect 19007 11940 19011 11996
rect 18947 11936 19011 11940
rect 3171 11452 3235 11456
rect 3171 11396 3175 11452
rect 3175 11396 3231 11452
rect 3231 11396 3235 11452
rect 3171 11392 3235 11396
rect 3251 11452 3315 11456
rect 3251 11396 3255 11452
rect 3255 11396 3311 11452
rect 3311 11396 3315 11452
rect 3251 11392 3315 11396
rect 3331 11452 3395 11456
rect 3331 11396 3335 11452
rect 3335 11396 3391 11452
rect 3391 11396 3395 11452
rect 3331 11392 3395 11396
rect 3411 11452 3475 11456
rect 3411 11396 3415 11452
rect 3415 11396 3471 11452
rect 3471 11396 3475 11452
rect 3411 11392 3475 11396
rect 7610 11452 7674 11456
rect 7610 11396 7614 11452
rect 7614 11396 7670 11452
rect 7670 11396 7674 11452
rect 7610 11392 7674 11396
rect 7690 11452 7754 11456
rect 7690 11396 7694 11452
rect 7694 11396 7750 11452
rect 7750 11396 7754 11452
rect 7690 11392 7754 11396
rect 7770 11452 7834 11456
rect 7770 11396 7774 11452
rect 7774 11396 7830 11452
rect 7830 11396 7834 11452
rect 7770 11392 7834 11396
rect 7850 11452 7914 11456
rect 7850 11396 7854 11452
rect 7854 11396 7910 11452
rect 7910 11396 7914 11452
rect 7850 11392 7914 11396
rect 12049 11452 12113 11456
rect 12049 11396 12053 11452
rect 12053 11396 12109 11452
rect 12109 11396 12113 11452
rect 12049 11392 12113 11396
rect 12129 11452 12193 11456
rect 12129 11396 12133 11452
rect 12133 11396 12189 11452
rect 12189 11396 12193 11452
rect 12129 11392 12193 11396
rect 12209 11452 12273 11456
rect 12209 11396 12213 11452
rect 12213 11396 12269 11452
rect 12269 11396 12273 11452
rect 12209 11392 12273 11396
rect 12289 11452 12353 11456
rect 12289 11396 12293 11452
rect 12293 11396 12349 11452
rect 12349 11396 12353 11452
rect 12289 11392 12353 11396
rect 16488 11452 16552 11456
rect 16488 11396 16492 11452
rect 16492 11396 16548 11452
rect 16548 11396 16552 11452
rect 16488 11392 16552 11396
rect 16568 11452 16632 11456
rect 16568 11396 16572 11452
rect 16572 11396 16628 11452
rect 16628 11396 16632 11452
rect 16568 11392 16632 11396
rect 16648 11452 16712 11456
rect 16648 11396 16652 11452
rect 16652 11396 16708 11452
rect 16708 11396 16712 11452
rect 16648 11392 16712 11396
rect 16728 11452 16792 11456
rect 16728 11396 16732 11452
rect 16732 11396 16788 11452
rect 16788 11396 16792 11452
rect 16728 11392 16792 11396
rect 5390 10908 5454 10912
rect 5390 10852 5394 10908
rect 5394 10852 5450 10908
rect 5450 10852 5454 10908
rect 5390 10848 5454 10852
rect 5470 10908 5534 10912
rect 5470 10852 5474 10908
rect 5474 10852 5530 10908
rect 5530 10852 5534 10908
rect 5470 10848 5534 10852
rect 5550 10908 5614 10912
rect 5550 10852 5554 10908
rect 5554 10852 5610 10908
rect 5610 10852 5614 10908
rect 5550 10848 5614 10852
rect 5630 10908 5694 10912
rect 5630 10852 5634 10908
rect 5634 10852 5690 10908
rect 5690 10852 5694 10908
rect 5630 10848 5694 10852
rect 9829 10908 9893 10912
rect 9829 10852 9833 10908
rect 9833 10852 9889 10908
rect 9889 10852 9893 10908
rect 9829 10848 9893 10852
rect 9909 10908 9973 10912
rect 9909 10852 9913 10908
rect 9913 10852 9969 10908
rect 9969 10852 9973 10908
rect 9909 10848 9973 10852
rect 9989 10908 10053 10912
rect 9989 10852 9993 10908
rect 9993 10852 10049 10908
rect 10049 10852 10053 10908
rect 9989 10848 10053 10852
rect 10069 10908 10133 10912
rect 10069 10852 10073 10908
rect 10073 10852 10129 10908
rect 10129 10852 10133 10908
rect 10069 10848 10133 10852
rect 14268 10908 14332 10912
rect 14268 10852 14272 10908
rect 14272 10852 14328 10908
rect 14328 10852 14332 10908
rect 14268 10848 14332 10852
rect 14348 10908 14412 10912
rect 14348 10852 14352 10908
rect 14352 10852 14408 10908
rect 14408 10852 14412 10908
rect 14348 10848 14412 10852
rect 14428 10908 14492 10912
rect 14428 10852 14432 10908
rect 14432 10852 14488 10908
rect 14488 10852 14492 10908
rect 14428 10848 14492 10852
rect 14508 10908 14572 10912
rect 14508 10852 14512 10908
rect 14512 10852 14568 10908
rect 14568 10852 14572 10908
rect 14508 10848 14572 10852
rect 18707 10908 18771 10912
rect 18707 10852 18711 10908
rect 18711 10852 18767 10908
rect 18767 10852 18771 10908
rect 18707 10848 18771 10852
rect 18787 10908 18851 10912
rect 18787 10852 18791 10908
rect 18791 10852 18847 10908
rect 18847 10852 18851 10908
rect 18787 10848 18851 10852
rect 18867 10908 18931 10912
rect 18867 10852 18871 10908
rect 18871 10852 18927 10908
rect 18927 10852 18931 10908
rect 18867 10848 18931 10852
rect 18947 10908 19011 10912
rect 18947 10852 18951 10908
rect 18951 10852 19007 10908
rect 19007 10852 19011 10908
rect 18947 10848 19011 10852
rect 3171 10364 3235 10368
rect 3171 10308 3175 10364
rect 3175 10308 3231 10364
rect 3231 10308 3235 10364
rect 3171 10304 3235 10308
rect 3251 10364 3315 10368
rect 3251 10308 3255 10364
rect 3255 10308 3311 10364
rect 3311 10308 3315 10364
rect 3251 10304 3315 10308
rect 3331 10364 3395 10368
rect 3331 10308 3335 10364
rect 3335 10308 3391 10364
rect 3391 10308 3395 10364
rect 3331 10304 3395 10308
rect 3411 10364 3475 10368
rect 3411 10308 3415 10364
rect 3415 10308 3471 10364
rect 3471 10308 3475 10364
rect 3411 10304 3475 10308
rect 7610 10364 7674 10368
rect 7610 10308 7614 10364
rect 7614 10308 7670 10364
rect 7670 10308 7674 10364
rect 7610 10304 7674 10308
rect 7690 10364 7754 10368
rect 7690 10308 7694 10364
rect 7694 10308 7750 10364
rect 7750 10308 7754 10364
rect 7690 10304 7754 10308
rect 7770 10364 7834 10368
rect 7770 10308 7774 10364
rect 7774 10308 7830 10364
rect 7830 10308 7834 10364
rect 7770 10304 7834 10308
rect 7850 10364 7914 10368
rect 7850 10308 7854 10364
rect 7854 10308 7910 10364
rect 7910 10308 7914 10364
rect 7850 10304 7914 10308
rect 12049 10364 12113 10368
rect 12049 10308 12053 10364
rect 12053 10308 12109 10364
rect 12109 10308 12113 10364
rect 12049 10304 12113 10308
rect 12129 10364 12193 10368
rect 12129 10308 12133 10364
rect 12133 10308 12189 10364
rect 12189 10308 12193 10364
rect 12129 10304 12193 10308
rect 12209 10364 12273 10368
rect 12209 10308 12213 10364
rect 12213 10308 12269 10364
rect 12269 10308 12273 10364
rect 12209 10304 12273 10308
rect 12289 10364 12353 10368
rect 12289 10308 12293 10364
rect 12293 10308 12349 10364
rect 12349 10308 12353 10364
rect 12289 10304 12353 10308
rect 16488 10364 16552 10368
rect 16488 10308 16492 10364
rect 16492 10308 16548 10364
rect 16548 10308 16552 10364
rect 16488 10304 16552 10308
rect 16568 10364 16632 10368
rect 16568 10308 16572 10364
rect 16572 10308 16628 10364
rect 16628 10308 16632 10364
rect 16568 10304 16632 10308
rect 16648 10364 16712 10368
rect 16648 10308 16652 10364
rect 16652 10308 16708 10364
rect 16708 10308 16712 10364
rect 16648 10304 16712 10308
rect 16728 10364 16792 10368
rect 16728 10308 16732 10364
rect 16732 10308 16788 10364
rect 16788 10308 16792 10364
rect 16728 10304 16792 10308
rect 5390 9820 5454 9824
rect 5390 9764 5394 9820
rect 5394 9764 5450 9820
rect 5450 9764 5454 9820
rect 5390 9760 5454 9764
rect 5470 9820 5534 9824
rect 5470 9764 5474 9820
rect 5474 9764 5530 9820
rect 5530 9764 5534 9820
rect 5470 9760 5534 9764
rect 5550 9820 5614 9824
rect 5550 9764 5554 9820
rect 5554 9764 5610 9820
rect 5610 9764 5614 9820
rect 5550 9760 5614 9764
rect 5630 9820 5694 9824
rect 5630 9764 5634 9820
rect 5634 9764 5690 9820
rect 5690 9764 5694 9820
rect 5630 9760 5694 9764
rect 9829 9820 9893 9824
rect 9829 9764 9833 9820
rect 9833 9764 9889 9820
rect 9889 9764 9893 9820
rect 9829 9760 9893 9764
rect 9909 9820 9973 9824
rect 9909 9764 9913 9820
rect 9913 9764 9969 9820
rect 9969 9764 9973 9820
rect 9909 9760 9973 9764
rect 9989 9820 10053 9824
rect 9989 9764 9993 9820
rect 9993 9764 10049 9820
rect 10049 9764 10053 9820
rect 9989 9760 10053 9764
rect 10069 9820 10133 9824
rect 10069 9764 10073 9820
rect 10073 9764 10129 9820
rect 10129 9764 10133 9820
rect 10069 9760 10133 9764
rect 14268 9820 14332 9824
rect 14268 9764 14272 9820
rect 14272 9764 14328 9820
rect 14328 9764 14332 9820
rect 14268 9760 14332 9764
rect 14348 9820 14412 9824
rect 14348 9764 14352 9820
rect 14352 9764 14408 9820
rect 14408 9764 14412 9820
rect 14348 9760 14412 9764
rect 14428 9820 14492 9824
rect 14428 9764 14432 9820
rect 14432 9764 14488 9820
rect 14488 9764 14492 9820
rect 14428 9760 14492 9764
rect 14508 9820 14572 9824
rect 14508 9764 14512 9820
rect 14512 9764 14568 9820
rect 14568 9764 14572 9820
rect 14508 9760 14572 9764
rect 18707 9820 18771 9824
rect 18707 9764 18711 9820
rect 18711 9764 18767 9820
rect 18767 9764 18771 9820
rect 18707 9760 18771 9764
rect 18787 9820 18851 9824
rect 18787 9764 18791 9820
rect 18791 9764 18847 9820
rect 18847 9764 18851 9820
rect 18787 9760 18851 9764
rect 18867 9820 18931 9824
rect 18867 9764 18871 9820
rect 18871 9764 18927 9820
rect 18927 9764 18931 9820
rect 18867 9760 18931 9764
rect 18947 9820 19011 9824
rect 18947 9764 18951 9820
rect 18951 9764 19007 9820
rect 19007 9764 19011 9820
rect 18947 9760 19011 9764
rect 3171 9276 3235 9280
rect 3171 9220 3175 9276
rect 3175 9220 3231 9276
rect 3231 9220 3235 9276
rect 3171 9216 3235 9220
rect 3251 9276 3315 9280
rect 3251 9220 3255 9276
rect 3255 9220 3311 9276
rect 3311 9220 3315 9276
rect 3251 9216 3315 9220
rect 3331 9276 3395 9280
rect 3331 9220 3335 9276
rect 3335 9220 3391 9276
rect 3391 9220 3395 9276
rect 3331 9216 3395 9220
rect 3411 9276 3475 9280
rect 3411 9220 3415 9276
rect 3415 9220 3471 9276
rect 3471 9220 3475 9276
rect 3411 9216 3475 9220
rect 7610 9276 7674 9280
rect 7610 9220 7614 9276
rect 7614 9220 7670 9276
rect 7670 9220 7674 9276
rect 7610 9216 7674 9220
rect 7690 9276 7754 9280
rect 7690 9220 7694 9276
rect 7694 9220 7750 9276
rect 7750 9220 7754 9276
rect 7690 9216 7754 9220
rect 7770 9276 7834 9280
rect 7770 9220 7774 9276
rect 7774 9220 7830 9276
rect 7830 9220 7834 9276
rect 7770 9216 7834 9220
rect 7850 9276 7914 9280
rect 7850 9220 7854 9276
rect 7854 9220 7910 9276
rect 7910 9220 7914 9276
rect 7850 9216 7914 9220
rect 12049 9276 12113 9280
rect 12049 9220 12053 9276
rect 12053 9220 12109 9276
rect 12109 9220 12113 9276
rect 12049 9216 12113 9220
rect 12129 9276 12193 9280
rect 12129 9220 12133 9276
rect 12133 9220 12189 9276
rect 12189 9220 12193 9276
rect 12129 9216 12193 9220
rect 12209 9276 12273 9280
rect 12209 9220 12213 9276
rect 12213 9220 12269 9276
rect 12269 9220 12273 9276
rect 12209 9216 12273 9220
rect 12289 9276 12353 9280
rect 12289 9220 12293 9276
rect 12293 9220 12349 9276
rect 12349 9220 12353 9276
rect 12289 9216 12353 9220
rect 16488 9276 16552 9280
rect 16488 9220 16492 9276
rect 16492 9220 16548 9276
rect 16548 9220 16552 9276
rect 16488 9216 16552 9220
rect 16568 9276 16632 9280
rect 16568 9220 16572 9276
rect 16572 9220 16628 9276
rect 16628 9220 16632 9276
rect 16568 9216 16632 9220
rect 16648 9276 16712 9280
rect 16648 9220 16652 9276
rect 16652 9220 16708 9276
rect 16708 9220 16712 9276
rect 16648 9216 16712 9220
rect 16728 9276 16792 9280
rect 16728 9220 16732 9276
rect 16732 9220 16788 9276
rect 16788 9220 16792 9276
rect 16728 9216 16792 9220
rect 5390 8732 5454 8736
rect 5390 8676 5394 8732
rect 5394 8676 5450 8732
rect 5450 8676 5454 8732
rect 5390 8672 5454 8676
rect 5470 8732 5534 8736
rect 5470 8676 5474 8732
rect 5474 8676 5530 8732
rect 5530 8676 5534 8732
rect 5470 8672 5534 8676
rect 5550 8732 5614 8736
rect 5550 8676 5554 8732
rect 5554 8676 5610 8732
rect 5610 8676 5614 8732
rect 5550 8672 5614 8676
rect 5630 8732 5694 8736
rect 5630 8676 5634 8732
rect 5634 8676 5690 8732
rect 5690 8676 5694 8732
rect 5630 8672 5694 8676
rect 9829 8732 9893 8736
rect 9829 8676 9833 8732
rect 9833 8676 9889 8732
rect 9889 8676 9893 8732
rect 9829 8672 9893 8676
rect 9909 8732 9973 8736
rect 9909 8676 9913 8732
rect 9913 8676 9969 8732
rect 9969 8676 9973 8732
rect 9909 8672 9973 8676
rect 9989 8732 10053 8736
rect 9989 8676 9993 8732
rect 9993 8676 10049 8732
rect 10049 8676 10053 8732
rect 9989 8672 10053 8676
rect 10069 8732 10133 8736
rect 10069 8676 10073 8732
rect 10073 8676 10129 8732
rect 10129 8676 10133 8732
rect 10069 8672 10133 8676
rect 14268 8732 14332 8736
rect 14268 8676 14272 8732
rect 14272 8676 14328 8732
rect 14328 8676 14332 8732
rect 14268 8672 14332 8676
rect 14348 8732 14412 8736
rect 14348 8676 14352 8732
rect 14352 8676 14408 8732
rect 14408 8676 14412 8732
rect 14348 8672 14412 8676
rect 14428 8732 14492 8736
rect 14428 8676 14432 8732
rect 14432 8676 14488 8732
rect 14488 8676 14492 8732
rect 14428 8672 14492 8676
rect 14508 8732 14572 8736
rect 14508 8676 14512 8732
rect 14512 8676 14568 8732
rect 14568 8676 14572 8732
rect 14508 8672 14572 8676
rect 18707 8732 18771 8736
rect 18707 8676 18711 8732
rect 18711 8676 18767 8732
rect 18767 8676 18771 8732
rect 18707 8672 18771 8676
rect 18787 8732 18851 8736
rect 18787 8676 18791 8732
rect 18791 8676 18847 8732
rect 18847 8676 18851 8732
rect 18787 8672 18851 8676
rect 18867 8732 18931 8736
rect 18867 8676 18871 8732
rect 18871 8676 18927 8732
rect 18927 8676 18931 8732
rect 18867 8672 18931 8676
rect 18947 8732 19011 8736
rect 18947 8676 18951 8732
rect 18951 8676 19007 8732
rect 19007 8676 19011 8732
rect 18947 8672 19011 8676
rect 3171 8188 3235 8192
rect 3171 8132 3175 8188
rect 3175 8132 3231 8188
rect 3231 8132 3235 8188
rect 3171 8128 3235 8132
rect 3251 8188 3315 8192
rect 3251 8132 3255 8188
rect 3255 8132 3311 8188
rect 3311 8132 3315 8188
rect 3251 8128 3315 8132
rect 3331 8188 3395 8192
rect 3331 8132 3335 8188
rect 3335 8132 3391 8188
rect 3391 8132 3395 8188
rect 3331 8128 3395 8132
rect 3411 8188 3475 8192
rect 3411 8132 3415 8188
rect 3415 8132 3471 8188
rect 3471 8132 3475 8188
rect 3411 8128 3475 8132
rect 7610 8188 7674 8192
rect 7610 8132 7614 8188
rect 7614 8132 7670 8188
rect 7670 8132 7674 8188
rect 7610 8128 7674 8132
rect 7690 8188 7754 8192
rect 7690 8132 7694 8188
rect 7694 8132 7750 8188
rect 7750 8132 7754 8188
rect 7690 8128 7754 8132
rect 7770 8188 7834 8192
rect 7770 8132 7774 8188
rect 7774 8132 7830 8188
rect 7830 8132 7834 8188
rect 7770 8128 7834 8132
rect 7850 8188 7914 8192
rect 7850 8132 7854 8188
rect 7854 8132 7910 8188
rect 7910 8132 7914 8188
rect 7850 8128 7914 8132
rect 12049 8188 12113 8192
rect 12049 8132 12053 8188
rect 12053 8132 12109 8188
rect 12109 8132 12113 8188
rect 12049 8128 12113 8132
rect 12129 8188 12193 8192
rect 12129 8132 12133 8188
rect 12133 8132 12189 8188
rect 12189 8132 12193 8188
rect 12129 8128 12193 8132
rect 12209 8188 12273 8192
rect 12209 8132 12213 8188
rect 12213 8132 12269 8188
rect 12269 8132 12273 8188
rect 12209 8128 12273 8132
rect 12289 8188 12353 8192
rect 12289 8132 12293 8188
rect 12293 8132 12349 8188
rect 12349 8132 12353 8188
rect 12289 8128 12353 8132
rect 16488 8188 16552 8192
rect 16488 8132 16492 8188
rect 16492 8132 16548 8188
rect 16548 8132 16552 8188
rect 16488 8128 16552 8132
rect 16568 8188 16632 8192
rect 16568 8132 16572 8188
rect 16572 8132 16628 8188
rect 16628 8132 16632 8188
rect 16568 8128 16632 8132
rect 16648 8188 16712 8192
rect 16648 8132 16652 8188
rect 16652 8132 16708 8188
rect 16708 8132 16712 8188
rect 16648 8128 16712 8132
rect 16728 8188 16792 8192
rect 16728 8132 16732 8188
rect 16732 8132 16788 8188
rect 16788 8132 16792 8188
rect 16728 8128 16792 8132
rect 5390 7644 5454 7648
rect 5390 7588 5394 7644
rect 5394 7588 5450 7644
rect 5450 7588 5454 7644
rect 5390 7584 5454 7588
rect 5470 7644 5534 7648
rect 5470 7588 5474 7644
rect 5474 7588 5530 7644
rect 5530 7588 5534 7644
rect 5470 7584 5534 7588
rect 5550 7644 5614 7648
rect 5550 7588 5554 7644
rect 5554 7588 5610 7644
rect 5610 7588 5614 7644
rect 5550 7584 5614 7588
rect 5630 7644 5694 7648
rect 5630 7588 5634 7644
rect 5634 7588 5690 7644
rect 5690 7588 5694 7644
rect 5630 7584 5694 7588
rect 9829 7644 9893 7648
rect 9829 7588 9833 7644
rect 9833 7588 9889 7644
rect 9889 7588 9893 7644
rect 9829 7584 9893 7588
rect 9909 7644 9973 7648
rect 9909 7588 9913 7644
rect 9913 7588 9969 7644
rect 9969 7588 9973 7644
rect 9909 7584 9973 7588
rect 9989 7644 10053 7648
rect 9989 7588 9993 7644
rect 9993 7588 10049 7644
rect 10049 7588 10053 7644
rect 9989 7584 10053 7588
rect 10069 7644 10133 7648
rect 10069 7588 10073 7644
rect 10073 7588 10129 7644
rect 10129 7588 10133 7644
rect 10069 7584 10133 7588
rect 14268 7644 14332 7648
rect 14268 7588 14272 7644
rect 14272 7588 14328 7644
rect 14328 7588 14332 7644
rect 14268 7584 14332 7588
rect 14348 7644 14412 7648
rect 14348 7588 14352 7644
rect 14352 7588 14408 7644
rect 14408 7588 14412 7644
rect 14348 7584 14412 7588
rect 14428 7644 14492 7648
rect 14428 7588 14432 7644
rect 14432 7588 14488 7644
rect 14488 7588 14492 7644
rect 14428 7584 14492 7588
rect 14508 7644 14572 7648
rect 14508 7588 14512 7644
rect 14512 7588 14568 7644
rect 14568 7588 14572 7644
rect 14508 7584 14572 7588
rect 18707 7644 18771 7648
rect 18707 7588 18711 7644
rect 18711 7588 18767 7644
rect 18767 7588 18771 7644
rect 18707 7584 18771 7588
rect 18787 7644 18851 7648
rect 18787 7588 18791 7644
rect 18791 7588 18847 7644
rect 18847 7588 18851 7644
rect 18787 7584 18851 7588
rect 18867 7644 18931 7648
rect 18867 7588 18871 7644
rect 18871 7588 18927 7644
rect 18927 7588 18931 7644
rect 18867 7584 18931 7588
rect 18947 7644 19011 7648
rect 18947 7588 18951 7644
rect 18951 7588 19007 7644
rect 19007 7588 19011 7644
rect 18947 7584 19011 7588
rect 3171 7100 3235 7104
rect 3171 7044 3175 7100
rect 3175 7044 3231 7100
rect 3231 7044 3235 7100
rect 3171 7040 3235 7044
rect 3251 7100 3315 7104
rect 3251 7044 3255 7100
rect 3255 7044 3311 7100
rect 3311 7044 3315 7100
rect 3251 7040 3315 7044
rect 3331 7100 3395 7104
rect 3331 7044 3335 7100
rect 3335 7044 3391 7100
rect 3391 7044 3395 7100
rect 3331 7040 3395 7044
rect 3411 7100 3475 7104
rect 3411 7044 3415 7100
rect 3415 7044 3471 7100
rect 3471 7044 3475 7100
rect 3411 7040 3475 7044
rect 7610 7100 7674 7104
rect 7610 7044 7614 7100
rect 7614 7044 7670 7100
rect 7670 7044 7674 7100
rect 7610 7040 7674 7044
rect 7690 7100 7754 7104
rect 7690 7044 7694 7100
rect 7694 7044 7750 7100
rect 7750 7044 7754 7100
rect 7690 7040 7754 7044
rect 7770 7100 7834 7104
rect 7770 7044 7774 7100
rect 7774 7044 7830 7100
rect 7830 7044 7834 7100
rect 7770 7040 7834 7044
rect 7850 7100 7914 7104
rect 7850 7044 7854 7100
rect 7854 7044 7910 7100
rect 7910 7044 7914 7100
rect 7850 7040 7914 7044
rect 12049 7100 12113 7104
rect 12049 7044 12053 7100
rect 12053 7044 12109 7100
rect 12109 7044 12113 7100
rect 12049 7040 12113 7044
rect 12129 7100 12193 7104
rect 12129 7044 12133 7100
rect 12133 7044 12189 7100
rect 12189 7044 12193 7100
rect 12129 7040 12193 7044
rect 12209 7100 12273 7104
rect 12209 7044 12213 7100
rect 12213 7044 12269 7100
rect 12269 7044 12273 7100
rect 12209 7040 12273 7044
rect 12289 7100 12353 7104
rect 12289 7044 12293 7100
rect 12293 7044 12349 7100
rect 12349 7044 12353 7100
rect 12289 7040 12353 7044
rect 16488 7100 16552 7104
rect 16488 7044 16492 7100
rect 16492 7044 16548 7100
rect 16548 7044 16552 7100
rect 16488 7040 16552 7044
rect 16568 7100 16632 7104
rect 16568 7044 16572 7100
rect 16572 7044 16628 7100
rect 16628 7044 16632 7100
rect 16568 7040 16632 7044
rect 16648 7100 16712 7104
rect 16648 7044 16652 7100
rect 16652 7044 16708 7100
rect 16708 7044 16712 7100
rect 16648 7040 16712 7044
rect 16728 7100 16792 7104
rect 16728 7044 16732 7100
rect 16732 7044 16788 7100
rect 16788 7044 16792 7100
rect 16728 7040 16792 7044
rect 5390 6556 5454 6560
rect 5390 6500 5394 6556
rect 5394 6500 5450 6556
rect 5450 6500 5454 6556
rect 5390 6496 5454 6500
rect 5470 6556 5534 6560
rect 5470 6500 5474 6556
rect 5474 6500 5530 6556
rect 5530 6500 5534 6556
rect 5470 6496 5534 6500
rect 5550 6556 5614 6560
rect 5550 6500 5554 6556
rect 5554 6500 5610 6556
rect 5610 6500 5614 6556
rect 5550 6496 5614 6500
rect 5630 6556 5694 6560
rect 5630 6500 5634 6556
rect 5634 6500 5690 6556
rect 5690 6500 5694 6556
rect 5630 6496 5694 6500
rect 9829 6556 9893 6560
rect 9829 6500 9833 6556
rect 9833 6500 9889 6556
rect 9889 6500 9893 6556
rect 9829 6496 9893 6500
rect 9909 6556 9973 6560
rect 9909 6500 9913 6556
rect 9913 6500 9969 6556
rect 9969 6500 9973 6556
rect 9909 6496 9973 6500
rect 9989 6556 10053 6560
rect 9989 6500 9993 6556
rect 9993 6500 10049 6556
rect 10049 6500 10053 6556
rect 9989 6496 10053 6500
rect 10069 6556 10133 6560
rect 10069 6500 10073 6556
rect 10073 6500 10129 6556
rect 10129 6500 10133 6556
rect 10069 6496 10133 6500
rect 14268 6556 14332 6560
rect 14268 6500 14272 6556
rect 14272 6500 14328 6556
rect 14328 6500 14332 6556
rect 14268 6496 14332 6500
rect 14348 6556 14412 6560
rect 14348 6500 14352 6556
rect 14352 6500 14408 6556
rect 14408 6500 14412 6556
rect 14348 6496 14412 6500
rect 14428 6556 14492 6560
rect 14428 6500 14432 6556
rect 14432 6500 14488 6556
rect 14488 6500 14492 6556
rect 14428 6496 14492 6500
rect 14508 6556 14572 6560
rect 14508 6500 14512 6556
rect 14512 6500 14568 6556
rect 14568 6500 14572 6556
rect 14508 6496 14572 6500
rect 18707 6556 18771 6560
rect 18707 6500 18711 6556
rect 18711 6500 18767 6556
rect 18767 6500 18771 6556
rect 18707 6496 18771 6500
rect 18787 6556 18851 6560
rect 18787 6500 18791 6556
rect 18791 6500 18847 6556
rect 18847 6500 18851 6556
rect 18787 6496 18851 6500
rect 18867 6556 18931 6560
rect 18867 6500 18871 6556
rect 18871 6500 18927 6556
rect 18927 6500 18931 6556
rect 18867 6496 18931 6500
rect 18947 6556 19011 6560
rect 18947 6500 18951 6556
rect 18951 6500 19007 6556
rect 19007 6500 19011 6556
rect 18947 6496 19011 6500
rect 3171 6012 3235 6016
rect 3171 5956 3175 6012
rect 3175 5956 3231 6012
rect 3231 5956 3235 6012
rect 3171 5952 3235 5956
rect 3251 6012 3315 6016
rect 3251 5956 3255 6012
rect 3255 5956 3311 6012
rect 3311 5956 3315 6012
rect 3251 5952 3315 5956
rect 3331 6012 3395 6016
rect 3331 5956 3335 6012
rect 3335 5956 3391 6012
rect 3391 5956 3395 6012
rect 3331 5952 3395 5956
rect 3411 6012 3475 6016
rect 3411 5956 3415 6012
rect 3415 5956 3471 6012
rect 3471 5956 3475 6012
rect 3411 5952 3475 5956
rect 7610 6012 7674 6016
rect 7610 5956 7614 6012
rect 7614 5956 7670 6012
rect 7670 5956 7674 6012
rect 7610 5952 7674 5956
rect 7690 6012 7754 6016
rect 7690 5956 7694 6012
rect 7694 5956 7750 6012
rect 7750 5956 7754 6012
rect 7690 5952 7754 5956
rect 7770 6012 7834 6016
rect 7770 5956 7774 6012
rect 7774 5956 7830 6012
rect 7830 5956 7834 6012
rect 7770 5952 7834 5956
rect 7850 6012 7914 6016
rect 7850 5956 7854 6012
rect 7854 5956 7910 6012
rect 7910 5956 7914 6012
rect 7850 5952 7914 5956
rect 12049 6012 12113 6016
rect 12049 5956 12053 6012
rect 12053 5956 12109 6012
rect 12109 5956 12113 6012
rect 12049 5952 12113 5956
rect 12129 6012 12193 6016
rect 12129 5956 12133 6012
rect 12133 5956 12189 6012
rect 12189 5956 12193 6012
rect 12129 5952 12193 5956
rect 12209 6012 12273 6016
rect 12209 5956 12213 6012
rect 12213 5956 12269 6012
rect 12269 5956 12273 6012
rect 12209 5952 12273 5956
rect 12289 6012 12353 6016
rect 12289 5956 12293 6012
rect 12293 5956 12349 6012
rect 12349 5956 12353 6012
rect 12289 5952 12353 5956
rect 16488 6012 16552 6016
rect 16488 5956 16492 6012
rect 16492 5956 16548 6012
rect 16548 5956 16552 6012
rect 16488 5952 16552 5956
rect 16568 6012 16632 6016
rect 16568 5956 16572 6012
rect 16572 5956 16628 6012
rect 16628 5956 16632 6012
rect 16568 5952 16632 5956
rect 16648 6012 16712 6016
rect 16648 5956 16652 6012
rect 16652 5956 16708 6012
rect 16708 5956 16712 6012
rect 16648 5952 16712 5956
rect 16728 6012 16792 6016
rect 16728 5956 16732 6012
rect 16732 5956 16788 6012
rect 16788 5956 16792 6012
rect 16728 5952 16792 5956
rect 5390 5468 5454 5472
rect 5390 5412 5394 5468
rect 5394 5412 5450 5468
rect 5450 5412 5454 5468
rect 5390 5408 5454 5412
rect 5470 5468 5534 5472
rect 5470 5412 5474 5468
rect 5474 5412 5530 5468
rect 5530 5412 5534 5468
rect 5470 5408 5534 5412
rect 5550 5468 5614 5472
rect 5550 5412 5554 5468
rect 5554 5412 5610 5468
rect 5610 5412 5614 5468
rect 5550 5408 5614 5412
rect 5630 5468 5694 5472
rect 5630 5412 5634 5468
rect 5634 5412 5690 5468
rect 5690 5412 5694 5468
rect 5630 5408 5694 5412
rect 9829 5468 9893 5472
rect 9829 5412 9833 5468
rect 9833 5412 9889 5468
rect 9889 5412 9893 5468
rect 9829 5408 9893 5412
rect 9909 5468 9973 5472
rect 9909 5412 9913 5468
rect 9913 5412 9969 5468
rect 9969 5412 9973 5468
rect 9909 5408 9973 5412
rect 9989 5468 10053 5472
rect 9989 5412 9993 5468
rect 9993 5412 10049 5468
rect 10049 5412 10053 5468
rect 9989 5408 10053 5412
rect 10069 5468 10133 5472
rect 10069 5412 10073 5468
rect 10073 5412 10129 5468
rect 10129 5412 10133 5468
rect 10069 5408 10133 5412
rect 14268 5468 14332 5472
rect 14268 5412 14272 5468
rect 14272 5412 14328 5468
rect 14328 5412 14332 5468
rect 14268 5408 14332 5412
rect 14348 5468 14412 5472
rect 14348 5412 14352 5468
rect 14352 5412 14408 5468
rect 14408 5412 14412 5468
rect 14348 5408 14412 5412
rect 14428 5468 14492 5472
rect 14428 5412 14432 5468
rect 14432 5412 14488 5468
rect 14488 5412 14492 5468
rect 14428 5408 14492 5412
rect 14508 5468 14572 5472
rect 14508 5412 14512 5468
rect 14512 5412 14568 5468
rect 14568 5412 14572 5468
rect 14508 5408 14572 5412
rect 18707 5468 18771 5472
rect 18707 5412 18711 5468
rect 18711 5412 18767 5468
rect 18767 5412 18771 5468
rect 18707 5408 18771 5412
rect 18787 5468 18851 5472
rect 18787 5412 18791 5468
rect 18791 5412 18847 5468
rect 18847 5412 18851 5468
rect 18787 5408 18851 5412
rect 18867 5468 18931 5472
rect 18867 5412 18871 5468
rect 18871 5412 18927 5468
rect 18927 5412 18931 5468
rect 18867 5408 18931 5412
rect 18947 5468 19011 5472
rect 18947 5412 18951 5468
rect 18951 5412 19007 5468
rect 19007 5412 19011 5468
rect 18947 5408 19011 5412
rect 3171 4924 3235 4928
rect 3171 4868 3175 4924
rect 3175 4868 3231 4924
rect 3231 4868 3235 4924
rect 3171 4864 3235 4868
rect 3251 4924 3315 4928
rect 3251 4868 3255 4924
rect 3255 4868 3311 4924
rect 3311 4868 3315 4924
rect 3251 4864 3315 4868
rect 3331 4924 3395 4928
rect 3331 4868 3335 4924
rect 3335 4868 3391 4924
rect 3391 4868 3395 4924
rect 3331 4864 3395 4868
rect 3411 4924 3475 4928
rect 3411 4868 3415 4924
rect 3415 4868 3471 4924
rect 3471 4868 3475 4924
rect 3411 4864 3475 4868
rect 7610 4924 7674 4928
rect 7610 4868 7614 4924
rect 7614 4868 7670 4924
rect 7670 4868 7674 4924
rect 7610 4864 7674 4868
rect 7690 4924 7754 4928
rect 7690 4868 7694 4924
rect 7694 4868 7750 4924
rect 7750 4868 7754 4924
rect 7690 4864 7754 4868
rect 7770 4924 7834 4928
rect 7770 4868 7774 4924
rect 7774 4868 7830 4924
rect 7830 4868 7834 4924
rect 7770 4864 7834 4868
rect 7850 4924 7914 4928
rect 7850 4868 7854 4924
rect 7854 4868 7910 4924
rect 7910 4868 7914 4924
rect 7850 4864 7914 4868
rect 12049 4924 12113 4928
rect 12049 4868 12053 4924
rect 12053 4868 12109 4924
rect 12109 4868 12113 4924
rect 12049 4864 12113 4868
rect 12129 4924 12193 4928
rect 12129 4868 12133 4924
rect 12133 4868 12189 4924
rect 12189 4868 12193 4924
rect 12129 4864 12193 4868
rect 12209 4924 12273 4928
rect 12209 4868 12213 4924
rect 12213 4868 12269 4924
rect 12269 4868 12273 4924
rect 12209 4864 12273 4868
rect 12289 4924 12353 4928
rect 12289 4868 12293 4924
rect 12293 4868 12349 4924
rect 12349 4868 12353 4924
rect 12289 4864 12353 4868
rect 16488 4924 16552 4928
rect 16488 4868 16492 4924
rect 16492 4868 16548 4924
rect 16548 4868 16552 4924
rect 16488 4864 16552 4868
rect 16568 4924 16632 4928
rect 16568 4868 16572 4924
rect 16572 4868 16628 4924
rect 16628 4868 16632 4924
rect 16568 4864 16632 4868
rect 16648 4924 16712 4928
rect 16648 4868 16652 4924
rect 16652 4868 16708 4924
rect 16708 4868 16712 4924
rect 16648 4864 16712 4868
rect 16728 4924 16792 4928
rect 16728 4868 16732 4924
rect 16732 4868 16788 4924
rect 16788 4868 16792 4924
rect 16728 4864 16792 4868
rect 5390 4380 5454 4384
rect 5390 4324 5394 4380
rect 5394 4324 5450 4380
rect 5450 4324 5454 4380
rect 5390 4320 5454 4324
rect 5470 4380 5534 4384
rect 5470 4324 5474 4380
rect 5474 4324 5530 4380
rect 5530 4324 5534 4380
rect 5470 4320 5534 4324
rect 5550 4380 5614 4384
rect 5550 4324 5554 4380
rect 5554 4324 5610 4380
rect 5610 4324 5614 4380
rect 5550 4320 5614 4324
rect 5630 4380 5694 4384
rect 5630 4324 5634 4380
rect 5634 4324 5690 4380
rect 5690 4324 5694 4380
rect 5630 4320 5694 4324
rect 9829 4380 9893 4384
rect 9829 4324 9833 4380
rect 9833 4324 9889 4380
rect 9889 4324 9893 4380
rect 9829 4320 9893 4324
rect 9909 4380 9973 4384
rect 9909 4324 9913 4380
rect 9913 4324 9969 4380
rect 9969 4324 9973 4380
rect 9909 4320 9973 4324
rect 9989 4380 10053 4384
rect 9989 4324 9993 4380
rect 9993 4324 10049 4380
rect 10049 4324 10053 4380
rect 9989 4320 10053 4324
rect 10069 4380 10133 4384
rect 10069 4324 10073 4380
rect 10073 4324 10129 4380
rect 10129 4324 10133 4380
rect 10069 4320 10133 4324
rect 14268 4380 14332 4384
rect 14268 4324 14272 4380
rect 14272 4324 14328 4380
rect 14328 4324 14332 4380
rect 14268 4320 14332 4324
rect 14348 4380 14412 4384
rect 14348 4324 14352 4380
rect 14352 4324 14408 4380
rect 14408 4324 14412 4380
rect 14348 4320 14412 4324
rect 14428 4380 14492 4384
rect 14428 4324 14432 4380
rect 14432 4324 14488 4380
rect 14488 4324 14492 4380
rect 14428 4320 14492 4324
rect 14508 4380 14572 4384
rect 14508 4324 14512 4380
rect 14512 4324 14568 4380
rect 14568 4324 14572 4380
rect 14508 4320 14572 4324
rect 18707 4380 18771 4384
rect 18707 4324 18711 4380
rect 18711 4324 18767 4380
rect 18767 4324 18771 4380
rect 18707 4320 18771 4324
rect 18787 4380 18851 4384
rect 18787 4324 18791 4380
rect 18791 4324 18847 4380
rect 18847 4324 18851 4380
rect 18787 4320 18851 4324
rect 18867 4380 18931 4384
rect 18867 4324 18871 4380
rect 18871 4324 18927 4380
rect 18927 4324 18931 4380
rect 18867 4320 18931 4324
rect 18947 4380 19011 4384
rect 18947 4324 18951 4380
rect 18951 4324 19007 4380
rect 19007 4324 19011 4380
rect 18947 4320 19011 4324
rect 3171 3836 3235 3840
rect 3171 3780 3175 3836
rect 3175 3780 3231 3836
rect 3231 3780 3235 3836
rect 3171 3776 3235 3780
rect 3251 3836 3315 3840
rect 3251 3780 3255 3836
rect 3255 3780 3311 3836
rect 3311 3780 3315 3836
rect 3251 3776 3315 3780
rect 3331 3836 3395 3840
rect 3331 3780 3335 3836
rect 3335 3780 3391 3836
rect 3391 3780 3395 3836
rect 3331 3776 3395 3780
rect 3411 3836 3475 3840
rect 3411 3780 3415 3836
rect 3415 3780 3471 3836
rect 3471 3780 3475 3836
rect 3411 3776 3475 3780
rect 7610 3836 7674 3840
rect 7610 3780 7614 3836
rect 7614 3780 7670 3836
rect 7670 3780 7674 3836
rect 7610 3776 7674 3780
rect 7690 3836 7754 3840
rect 7690 3780 7694 3836
rect 7694 3780 7750 3836
rect 7750 3780 7754 3836
rect 7690 3776 7754 3780
rect 7770 3836 7834 3840
rect 7770 3780 7774 3836
rect 7774 3780 7830 3836
rect 7830 3780 7834 3836
rect 7770 3776 7834 3780
rect 7850 3836 7914 3840
rect 7850 3780 7854 3836
rect 7854 3780 7910 3836
rect 7910 3780 7914 3836
rect 7850 3776 7914 3780
rect 12049 3836 12113 3840
rect 12049 3780 12053 3836
rect 12053 3780 12109 3836
rect 12109 3780 12113 3836
rect 12049 3776 12113 3780
rect 12129 3836 12193 3840
rect 12129 3780 12133 3836
rect 12133 3780 12189 3836
rect 12189 3780 12193 3836
rect 12129 3776 12193 3780
rect 12209 3836 12273 3840
rect 12209 3780 12213 3836
rect 12213 3780 12269 3836
rect 12269 3780 12273 3836
rect 12209 3776 12273 3780
rect 12289 3836 12353 3840
rect 12289 3780 12293 3836
rect 12293 3780 12349 3836
rect 12349 3780 12353 3836
rect 12289 3776 12353 3780
rect 16488 3836 16552 3840
rect 16488 3780 16492 3836
rect 16492 3780 16548 3836
rect 16548 3780 16552 3836
rect 16488 3776 16552 3780
rect 16568 3836 16632 3840
rect 16568 3780 16572 3836
rect 16572 3780 16628 3836
rect 16628 3780 16632 3836
rect 16568 3776 16632 3780
rect 16648 3836 16712 3840
rect 16648 3780 16652 3836
rect 16652 3780 16708 3836
rect 16708 3780 16712 3836
rect 16648 3776 16712 3780
rect 16728 3836 16792 3840
rect 16728 3780 16732 3836
rect 16732 3780 16788 3836
rect 16788 3780 16792 3836
rect 16728 3776 16792 3780
rect 5390 3292 5454 3296
rect 5390 3236 5394 3292
rect 5394 3236 5450 3292
rect 5450 3236 5454 3292
rect 5390 3232 5454 3236
rect 5470 3292 5534 3296
rect 5470 3236 5474 3292
rect 5474 3236 5530 3292
rect 5530 3236 5534 3292
rect 5470 3232 5534 3236
rect 5550 3292 5614 3296
rect 5550 3236 5554 3292
rect 5554 3236 5610 3292
rect 5610 3236 5614 3292
rect 5550 3232 5614 3236
rect 5630 3292 5694 3296
rect 5630 3236 5634 3292
rect 5634 3236 5690 3292
rect 5690 3236 5694 3292
rect 5630 3232 5694 3236
rect 9829 3292 9893 3296
rect 9829 3236 9833 3292
rect 9833 3236 9889 3292
rect 9889 3236 9893 3292
rect 9829 3232 9893 3236
rect 9909 3292 9973 3296
rect 9909 3236 9913 3292
rect 9913 3236 9969 3292
rect 9969 3236 9973 3292
rect 9909 3232 9973 3236
rect 9989 3292 10053 3296
rect 9989 3236 9993 3292
rect 9993 3236 10049 3292
rect 10049 3236 10053 3292
rect 9989 3232 10053 3236
rect 10069 3292 10133 3296
rect 10069 3236 10073 3292
rect 10073 3236 10129 3292
rect 10129 3236 10133 3292
rect 10069 3232 10133 3236
rect 14268 3292 14332 3296
rect 14268 3236 14272 3292
rect 14272 3236 14328 3292
rect 14328 3236 14332 3292
rect 14268 3232 14332 3236
rect 14348 3292 14412 3296
rect 14348 3236 14352 3292
rect 14352 3236 14408 3292
rect 14408 3236 14412 3292
rect 14348 3232 14412 3236
rect 14428 3292 14492 3296
rect 14428 3236 14432 3292
rect 14432 3236 14488 3292
rect 14488 3236 14492 3292
rect 14428 3232 14492 3236
rect 14508 3292 14572 3296
rect 14508 3236 14512 3292
rect 14512 3236 14568 3292
rect 14568 3236 14572 3292
rect 14508 3232 14572 3236
rect 18707 3292 18771 3296
rect 18707 3236 18711 3292
rect 18711 3236 18767 3292
rect 18767 3236 18771 3292
rect 18707 3232 18771 3236
rect 18787 3292 18851 3296
rect 18787 3236 18791 3292
rect 18791 3236 18847 3292
rect 18847 3236 18851 3292
rect 18787 3232 18851 3236
rect 18867 3292 18931 3296
rect 18867 3236 18871 3292
rect 18871 3236 18927 3292
rect 18927 3236 18931 3292
rect 18867 3232 18931 3236
rect 18947 3292 19011 3296
rect 18947 3236 18951 3292
rect 18951 3236 19007 3292
rect 19007 3236 19011 3292
rect 18947 3232 19011 3236
rect 3171 2748 3235 2752
rect 3171 2692 3175 2748
rect 3175 2692 3231 2748
rect 3231 2692 3235 2748
rect 3171 2688 3235 2692
rect 3251 2748 3315 2752
rect 3251 2692 3255 2748
rect 3255 2692 3311 2748
rect 3311 2692 3315 2748
rect 3251 2688 3315 2692
rect 3331 2748 3395 2752
rect 3331 2692 3335 2748
rect 3335 2692 3391 2748
rect 3391 2692 3395 2748
rect 3331 2688 3395 2692
rect 3411 2748 3475 2752
rect 3411 2692 3415 2748
rect 3415 2692 3471 2748
rect 3471 2692 3475 2748
rect 3411 2688 3475 2692
rect 7610 2748 7674 2752
rect 7610 2692 7614 2748
rect 7614 2692 7670 2748
rect 7670 2692 7674 2748
rect 7610 2688 7674 2692
rect 7690 2748 7754 2752
rect 7690 2692 7694 2748
rect 7694 2692 7750 2748
rect 7750 2692 7754 2748
rect 7690 2688 7754 2692
rect 7770 2748 7834 2752
rect 7770 2692 7774 2748
rect 7774 2692 7830 2748
rect 7830 2692 7834 2748
rect 7770 2688 7834 2692
rect 7850 2748 7914 2752
rect 7850 2692 7854 2748
rect 7854 2692 7910 2748
rect 7910 2692 7914 2748
rect 7850 2688 7914 2692
rect 12049 2748 12113 2752
rect 12049 2692 12053 2748
rect 12053 2692 12109 2748
rect 12109 2692 12113 2748
rect 12049 2688 12113 2692
rect 12129 2748 12193 2752
rect 12129 2692 12133 2748
rect 12133 2692 12189 2748
rect 12189 2692 12193 2748
rect 12129 2688 12193 2692
rect 12209 2748 12273 2752
rect 12209 2692 12213 2748
rect 12213 2692 12269 2748
rect 12269 2692 12273 2748
rect 12209 2688 12273 2692
rect 12289 2748 12353 2752
rect 12289 2692 12293 2748
rect 12293 2692 12349 2748
rect 12349 2692 12353 2748
rect 12289 2688 12353 2692
rect 16488 2748 16552 2752
rect 16488 2692 16492 2748
rect 16492 2692 16548 2748
rect 16548 2692 16552 2748
rect 16488 2688 16552 2692
rect 16568 2748 16632 2752
rect 16568 2692 16572 2748
rect 16572 2692 16628 2748
rect 16628 2692 16632 2748
rect 16568 2688 16632 2692
rect 16648 2748 16712 2752
rect 16648 2692 16652 2748
rect 16652 2692 16708 2748
rect 16708 2692 16712 2748
rect 16648 2688 16712 2692
rect 16728 2748 16792 2752
rect 16728 2692 16732 2748
rect 16732 2692 16788 2748
rect 16788 2692 16792 2748
rect 16728 2688 16792 2692
rect 5390 2204 5454 2208
rect 5390 2148 5394 2204
rect 5394 2148 5450 2204
rect 5450 2148 5454 2204
rect 5390 2144 5454 2148
rect 5470 2204 5534 2208
rect 5470 2148 5474 2204
rect 5474 2148 5530 2204
rect 5530 2148 5534 2204
rect 5470 2144 5534 2148
rect 5550 2204 5614 2208
rect 5550 2148 5554 2204
rect 5554 2148 5610 2204
rect 5610 2148 5614 2204
rect 5550 2144 5614 2148
rect 5630 2204 5694 2208
rect 5630 2148 5634 2204
rect 5634 2148 5690 2204
rect 5690 2148 5694 2204
rect 5630 2144 5694 2148
rect 9829 2204 9893 2208
rect 9829 2148 9833 2204
rect 9833 2148 9889 2204
rect 9889 2148 9893 2204
rect 9829 2144 9893 2148
rect 9909 2204 9973 2208
rect 9909 2148 9913 2204
rect 9913 2148 9969 2204
rect 9969 2148 9973 2204
rect 9909 2144 9973 2148
rect 9989 2204 10053 2208
rect 9989 2148 9993 2204
rect 9993 2148 10049 2204
rect 10049 2148 10053 2204
rect 9989 2144 10053 2148
rect 10069 2204 10133 2208
rect 10069 2148 10073 2204
rect 10073 2148 10129 2204
rect 10129 2148 10133 2204
rect 10069 2144 10133 2148
rect 14268 2204 14332 2208
rect 14268 2148 14272 2204
rect 14272 2148 14328 2204
rect 14328 2148 14332 2204
rect 14268 2144 14332 2148
rect 14348 2204 14412 2208
rect 14348 2148 14352 2204
rect 14352 2148 14408 2204
rect 14408 2148 14412 2204
rect 14348 2144 14412 2148
rect 14428 2204 14492 2208
rect 14428 2148 14432 2204
rect 14432 2148 14488 2204
rect 14488 2148 14492 2204
rect 14428 2144 14492 2148
rect 14508 2204 14572 2208
rect 14508 2148 14512 2204
rect 14512 2148 14568 2204
rect 14568 2148 14572 2204
rect 14508 2144 14572 2148
rect 18707 2204 18771 2208
rect 18707 2148 18711 2204
rect 18711 2148 18767 2204
rect 18767 2148 18771 2204
rect 18707 2144 18771 2148
rect 18787 2204 18851 2208
rect 18787 2148 18791 2204
rect 18791 2148 18847 2204
rect 18847 2148 18851 2204
rect 18787 2144 18851 2148
rect 18867 2204 18931 2208
rect 18867 2148 18871 2204
rect 18871 2148 18927 2204
rect 18927 2148 18931 2204
rect 18867 2144 18931 2148
rect 18947 2204 19011 2208
rect 18947 2148 18951 2204
rect 18951 2148 19007 2204
rect 19007 2148 19011 2204
rect 18947 2144 19011 2148
<< metal4 >>
rect 3163 16896 3483 17456
rect 3163 16832 3171 16896
rect 3235 16832 3251 16896
rect 3315 16832 3331 16896
rect 3395 16832 3411 16896
rect 3475 16832 3483 16896
rect 3163 15808 3483 16832
rect 3163 15744 3171 15808
rect 3235 15744 3251 15808
rect 3315 15744 3331 15808
rect 3395 15744 3411 15808
rect 3475 15744 3483 15808
rect 3163 14720 3483 15744
rect 3163 14656 3171 14720
rect 3235 14656 3251 14720
rect 3315 14656 3331 14720
rect 3395 14656 3411 14720
rect 3475 14656 3483 14720
rect 3163 13632 3483 14656
rect 3163 13568 3171 13632
rect 3235 13568 3251 13632
rect 3315 13568 3331 13632
rect 3395 13568 3411 13632
rect 3475 13568 3483 13632
rect 3163 12544 3483 13568
rect 3163 12480 3171 12544
rect 3235 12480 3251 12544
rect 3315 12480 3331 12544
rect 3395 12480 3411 12544
rect 3475 12480 3483 12544
rect 3163 11456 3483 12480
rect 3163 11392 3171 11456
rect 3235 11392 3251 11456
rect 3315 11392 3331 11456
rect 3395 11392 3411 11456
rect 3475 11392 3483 11456
rect 3163 10368 3483 11392
rect 3163 10304 3171 10368
rect 3235 10304 3251 10368
rect 3315 10304 3331 10368
rect 3395 10304 3411 10368
rect 3475 10304 3483 10368
rect 3163 9280 3483 10304
rect 3163 9216 3171 9280
rect 3235 9216 3251 9280
rect 3315 9216 3331 9280
rect 3395 9216 3411 9280
rect 3475 9216 3483 9280
rect 3163 8192 3483 9216
rect 3163 8128 3171 8192
rect 3235 8128 3251 8192
rect 3315 8128 3331 8192
rect 3395 8128 3411 8192
rect 3475 8128 3483 8192
rect 3163 7104 3483 8128
rect 3163 7040 3171 7104
rect 3235 7040 3251 7104
rect 3315 7040 3331 7104
rect 3395 7040 3411 7104
rect 3475 7040 3483 7104
rect 3163 6016 3483 7040
rect 3163 5952 3171 6016
rect 3235 5952 3251 6016
rect 3315 5952 3331 6016
rect 3395 5952 3411 6016
rect 3475 5952 3483 6016
rect 3163 4928 3483 5952
rect 3163 4864 3171 4928
rect 3235 4864 3251 4928
rect 3315 4864 3331 4928
rect 3395 4864 3411 4928
rect 3475 4864 3483 4928
rect 3163 3840 3483 4864
rect 3163 3776 3171 3840
rect 3235 3776 3251 3840
rect 3315 3776 3331 3840
rect 3395 3776 3411 3840
rect 3475 3776 3483 3840
rect 3163 2752 3483 3776
rect 3163 2688 3171 2752
rect 3235 2688 3251 2752
rect 3315 2688 3331 2752
rect 3395 2688 3411 2752
rect 3475 2688 3483 2752
rect 3163 2128 3483 2688
rect 5382 17440 5702 17456
rect 5382 17376 5390 17440
rect 5454 17376 5470 17440
rect 5534 17376 5550 17440
rect 5614 17376 5630 17440
rect 5694 17376 5702 17440
rect 5382 16352 5702 17376
rect 5382 16288 5390 16352
rect 5454 16288 5470 16352
rect 5534 16288 5550 16352
rect 5614 16288 5630 16352
rect 5694 16288 5702 16352
rect 5382 15264 5702 16288
rect 5382 15200 5390 15264
rect 5454 15200 5470 15264
rect 5534 15200 5550 15264
rect 5614 15200 5630 15264
rect 5694 15200 5702 15264
rect 5382 14176 5702 15200
rect 5382 14112 5390 14176
rect 5454 14112 5470 14176
rect 5534 14112 5550 14176
rect 5614 14112 5630 14176
rect 5694 14112 5702 14176
rect 5382 13088 5702 14112
rect 5382 13024 5390 13088
rect 5454 13024 5470 13088
rect 5534 13024 5550 13088
rect 5614 13024 5630 13088
rect 5694 13024 5702 13088
rect 5382 12000 5702 13024
rect 5382 11936 5390 12000
rect 5454 11936 5470 12000
rect 5534 11936 5550 12000
rect 5614 11936 5630 12000
rect 5694 11936 5702 12000
rect 5382 10912 5702 11936
rect 5382 10848 5390 10912
rect 5454 10848 5470 10912
rect 5534 10848 5550 10912
rect 5614 10848 5630 10912
rect 5694 10848 5702 10912
rect 5382 9824 5702 10848
rect 5382 9760 5390 9824
rect 5454 9760 5470 9824
rect 5534 9760 5550 9824
rect 5614 9760 5630 9824
rect 5694 9760 5702 9824
rect 5382 8736 5702 9760
rect 5382 8672 5390 8736
rect 5454 8672 5470 8736
rect 5534 8672 5550 8736
rect 5614 8672 5630 8736
rect 5694 8672 5702 8736
rect 5382 7648 5702 8672
rect 5382 7584 5390 7648
rect 5454 7584 5470 7648
rect 5534 7584 5550 7648
rect 5614 7584 5630 7648
rect 5694 7584 5702 7648
rect 5382 6560 5702 7584
rect 5382 6496 5390 6560
rect 5454 6496 5470 6560
rect 5534 6496 5550 6560
rect 5614 6496 5630 6560
rect 5694 6496 5702 6560
rect 5382 5472 5702 6496
rect 5382 5408 5390 5472
rect 5454 5408 5470 5472
rect 5534 5408 5550 5472
rect 5614 5408 5630 5472
rect 5694 5408 5702 5472
rect 5382 4384 5702 5408
rect 5382 4320 5390 4384
rect 5454 4320 5470 4384
rect 5534 4320 5550 4384
rect 5614 4320 5630 4384
rect 5694 4320 5702 4384
rect 5382 3296 5702 4320
rect 5382 3232 5390 3296
rect 5454 3232 5470 3296
rect 5534 3232 5550 3296
rect 5614 3232 5630 3296
rect 5694 3232 5702 3296
rect 5382 2208 5702 3232
rect 5382 2144 5390 2208
rect 5454 2144 5470 2208
rect 5534 2144 5550 2208
rect 5614 2144 5630 2208
rect 5694 2144 5702 2208
rect 5382 2128 5702 2144
rect 7602 16896 7922 17456
rect 7602 16832 7610 16896
rect 7674 16832 7690 16896
rect 7754 16832 7770 16896
rect 7834 16832 7850 16896
rect 7914 16832 7922 16896
rect 7602 15808 7922 16832
rect 7602 15744 7610 15808
rect 7674 15744 7690 15808
rect 7754 15744 7770 15808
rect 7834 15744 7850 15808
rect 7914 15744 7922 15808
rect 7602 14720 7922 15744
rect 7602 14656 7610 14720
rect 7674 14656 7690 14720
rect 7754 14656 7770 14720
rect 7834 14656 7850 14720
rect 7914 14656 7922 14720
rect 7602 13632 7922 14656
rect 7602 13568 7610 13632
rect 7674 13568 7690 13632
rect 7754 13568 7770 13632
rect 7834 13568 7850 13632
rect 7914 13568 7922 13632
rect 7602 12544 7922 13568
rect 7602 12480 7610 12544
rect 7674 12480 7690 12544
rect 7754 12480 7770 12544
rect 7834 12480 7850 12544
rect 7914 12480 7922 12544
rect 7602 11456 7922 12480
rect 7602 11392 7610 11456
rect 7674 11392 7690 11456
rect 7754 11392 7770 11456
rect 7834 11392 7850 11456
rect 7914 11392 7922 11456
rect 7602 10368 7922 11392
rect 7602 10304 7610 10368
rect 7674 10304 7690 10368
rect 7754 10304 7770 10368
rect 7834 10304 7850 10368
rect 7914 10304 7922 10368
rect 7602 9280 7922 10304
rect 7602 9216 7610 9280
rect 7674 9216 7690 9280
rect 7754 9216 7770 9280
rect 7834 9216 7850 9280
rect 7914 9216 7922 9280
rect 7602 8192 7922 9216
rect 7602 8128 7610 8192
rect 7674 8128 7690 8192
rect 7754 8128 7770 8192
rect 7834 8128 7850 8192
rect 7914 8128 7922 8192
rect 7602 7104 7922 8128
rect 7602 7040 7610 7104
rect 7674 7040 7690 7104
rect 7754 7040 7770 7104
rect 7834 7040 7850 7104
rect 7914 7040 7922 7104
rect 7602 6016 7922 7040
rect 7602 5952 7610 6016
rect 7674 5952 7690 6016
rect 7754 5952 7770 6016
rect 7834 5952 7850 6016
rect 7914 5952 7922 6016
rect 7602 4928 7922 5952
rect 7602 4864 7610 4928
rect 7674 4864 7690 4928
rect 7754 4864 7770 4928
rect 7834 4864 7850 4928
rect 7914 4864 7922 4928
rect 7602 3840 7922 4864
rect 7602 3776 7610 3840
rect 7674 3776 7690 3840
rect 7754 3776 7770 3840
rect 7834 3776 7850 3840
rect 7914 3776 7922 3840
rect 7602 2752 7922 3776
rect 7602 2688 7610 2752
rect 7674 2688 7690 2752
rect 7754 2688 7770 2752
rect 7834 2688 7850 2752
rect 7914 2688 7922 2752
rect 7602 2128 7922 2688
rect 9821 17440 10141 17456
rect 9821 17376 9829 17440
rect 9893 17376 9909 17440
rect 9973 17376 9989 17440
rect 10053 17376 10069 17440
rect 10133 17376 10141 17440
rect 9821 16352 10141 17376
rect 9821 16288 9829 16352
rect 9893 16288 9909 16352
rect 9973 16288 9989 16352
rect 10053 16288 10069 16352
rect 10133 16288 10141 16352
rect 9821 15264 10141 16288
rect 9821 15200 9829 15264
rect 9893 15200 9909 15264
rect 9973 15200 9989 15264
rect 10053 15200 10069 15264
rect 10133 15200 10141 15264
rect 9821 14176 10141 15200
rect 9821 14112 9829 14176
rect 9893 14112 9909 14176
rect 9973 14112 9989 14176
rect 10053 14112 10069 14176
rect 10133 14112 10141 14176
rect 9821 13088 10141 14112
rect 9821 13024 9829 13088
rect 9893 13024 9909 13088
rect 9973 13024 9989 13088
rect 10053 13024 10069 13088
rect 10133 13024 10141 13088
rect 9821 12000 10141 13024
rect 9821 11936 9829 12000
rect 9893 11936 9909 12000
rect 9973 11936 9989 12000
rect 10053 11936 10069 12000
rect 10133 11936 10141 12000
rect 9821 10912 10141 11936
rect 9821 10848 9829 10912
rect 9893 10848 9909 10912
rect 9973 10848 9989 10912
rect 10053 10848 10069 10912
rect 10133 10848 10141 10912
rect 9821 9824 10141 10848
rect 9821 9760 9829 9824
rect 9893 9760 9909 9824
rect 9973 9760 9989 9824
rect 10053 9760 10069 9824
rect 10133 9760 10141 9824
rect 9821 8736 10141 9760
rect 9821 8672 9829 8736
rect 9893 8672 9909 8736
rect 9973 8672 9989 8736
rect 10053 8672 10069 8736
rect 10133 8672 10141 8736
rect 9821 7648 10141 8672
rect 9821 7584 9829 7648
rect 9893 7584 9909 7648
rect 9973 7584 9989 7648
rect 10053 7584 10069 7648
rect 10133 7584 10141 7648
rect 9821 6560 10141 7584
rect 9821 6496 9829 6560
rect 9893 6496 9909 6560
rect 9973 6496 9989 6560
rect 10053 6496 10069 6560
rect 10133 6496 10141 6560
rect 9821 5472 10141 6496
rect 9821 5408 9829 5472
rect 9893 5408 9909 5472
rect 9973 5408 9989 5472
rect 10053 5408 10069 5472
rect 10133 5408 10141 5472
rect 9821 4384 10141 5408
rect 9821 4320 9829 4384
rect 9893 4320 9909 4384
rect 9973 4320 9989 4384
rect 10053 4320 10069 4384
rect 10133 4320 10141 4384
rect 9821 3296 10141 4320
rect 9821 3232 9829 3296
rect 9893 3232 9909 3296
rect 9973 3232 9989 3296
rect 10053 3232 10069 3296
rect 10133 3232 10141 3296
rect 9821 2208 10141 3232
rect 9821 2144 9829 2208
rect 9893 2144 9909 2208
rect 9973 2144 9989 2208
rect 10053 2144 10069 2208
rect 10133 2144 10141 2208
rect 9821 2128 10141 2144
rect 12041 16896 12361 17456
rect 12041 16832 12049 16896
rect 12113 16832 12129 16896
rect 12193 16832 12209 16896
rect 12273 16832 12289 16896
rect 12353 16832 12361 16896
rect 12041 15808 12361 16832
rect 12041 15744 12049 15808
rect 12113 15744 12129 15808
rect 12193 15744 12209 15808
rect 12273 15744 12289 15808
rect 12353 15744 12361 15808
rect 12041 14720 12361 15744
rect 12041 14656 12049 14720
rect 12113 14656 12129 14720
rect 12193 14656 12209 14720
rect 12273 14656 12289 14720
rect 12353 14656 12361 14720
rect 12041 13632 12361 14656
rect 12041 13568 12049 13632
rect 12113 13568 12129 13632
rect 12193 13568 12209 13632
rect 12273 13568 12289 13632
rect 12353 13568 12361 13632
rect 12041 12544 12361 13568
rect 12041 12480 12049 12544
rect 12113 12480 12129 12544
rect 12193 12480 12209 12544
rect 12273 12480 12289 12544
rect 12353 12480 12361 12544
rect 12041 11456 12361 12480
rect 12041 11392 12049 11456
rect 12113 11392 12129 11456
rect 12193 11392 12209 11456
rect 12273 11392 12289 11456
rect 12353 11392 12361 11456
rect 12041 10368 12361 11392
rect 12041 10304 12049 10368
rect 12113 10304 12129 10368
rect 12193 10304 12209 10368
rect 12273 10304 12289 10368
rect 12353 10304 12361 10368
rect 12041 9280 12361 10304
rect 12041 9216 12049 9280
rect 12113 9216 12129 9280
rect 12193 9216 12209 9280
rect 12273 9216 12289 9280
rect 12353 9216 12361 9280
rect 12041 8192 12361 9216
rect 12041 8128 12049 8192
rect 12113 8128 12129 8192
rect 12193 8128 12209 8192
rect 12273 8128 12289 8192
rect 12353 8128 12361 8192
rect 12041 7104 12361 8128
rect 12041 7040 12049 7104
rect 12113 7040 12129 7104
rect 12193 7040 12209 7104
rect 12273 7040 12289 7104
rect 12353 7040 12361 7104
rect 12041 6016 12361 7040
rect 12041 5952 12049 6016
rect 12113 5952 12129 6016
rect 12193 5952 12209 6016
rect 12273 5952 12289 6016
rect 12353 5952 12361 6016
rect 12041 4928 12361 5952
rect 12041 4864 12049 4928
rect 12113 4864 12129 4928
rect 12193 4864 12209 4928
rect 12273 4864 12289 4928
rect 12353 4864 12361 4928
rect 12041 3840 12361 4864
rect 12041 3776 12049 3840
rect 12113 3776 12129 3840
rect 12193 3776 12209 3840
rect 12273 3776 12289 3840
rect 12353 3776 12361 3840
rect 12041 2752 12361 3776
rect 12041 2688 12049 2752
rect 12113 2688 12129 2752
rect 12193 2688 12209 2752
rect 12273 2688 12289 2752
rect 12353 2688 12361 2752
rect 12041 2128 12361 2688
rect 14260 17440 14580 17456
rect 14260 17376 14268 17440
rect 14332 17376 14348 17440
rect 14412 17376 14428 17440
rect 14492 17376 14508 17440
rect 14572 17376 14580 17440
rect 14260 16352 14580 17376
rect 14260 16288 14268 16352
rect 14332 16288 14348 16352
rect 14412 16288 14428 16352
rect 14492 16288 14508 16352
rect 14572 16288 14580 16352
rect 14260 15264 14580 16288
rect 14260 15200 14268 15264
rect 14332 15200 14348 15264
rect 14412 15200 14428 15264
rect 14492 15200 14508 15264
rect 14572 15200 14580 15264
rect 14260 14176 14580 15200
rect 14260 14112 14268 14176
rect 14332 14112 14348 14176
rect 14412 14112 14428 14176
rect 14492 14112 14508 14176
rect 14572 14112 14580 14176
rect 14260 13088 14580 14112
rect 14260 13024 14268 13088
rect 14332 13024 14348 13088
rect 14412 13024 14428 13088
rect 14492 13024 14508 13088
rect 14572 13024 14580 13088
rect 14260 12000 14580 13024
rect 14260 11936 14268 12000
rect 14332 11936 14348 12000
rect 14412 11936 14428 12000
rect 14492 11936 14508 12000
rect 14572 11936 14580 12000
rect 14260 10912 14580 11936
rect 14260 10848 14268 10912
rect 14332 10848 14348 10912
rect 14412 10848 14428 10912
rect 14492 10848 14508 10912
rect 14572 10848 14580 10912
rect 14260 9824 14580 10848
rect 14260 9760 14268 9824
rect 14332 9760 14348 9824
rect 14412 9760 14428 9824
rect 14492 9760 14508 9824
rect 14572 9760 14580 9824
rect 14260 8736 14580 9760
rect 14260 8672 14268 8736
rect 14332 8672 14348 8736
rect 14412 8672 14428 8736
rect 14492 8672 14508 8736
rect 14572 8672 14580 8736
rect 14260 7648 14580 8672
rect 14260 7584 14268 7648
rect 14332 7584 14348 7648
rect 14412 7584 14428 7648
rect 14492 7584 14508 7648
rect 14572 7584 14580 7648
rect 14260 6560 14580 7584
rect 14260 6496 14268 6560
rect 14332 6496 14348 6560
rect 14412 6496 14428 6560
rect 14492 6496 14508 6560
rect 14572 6496 14580 6560
rect 14260 5472 14580 6496
rect 14260 5408 14268 5472
rect 14332 5408 14348 5472
rect 14412 5408 14428 5472
rect 14492 5408 14508 5472
rect 14572 5408 14580 5472
rect 14260 4384 14580 5408
rect 14260 4320 14268 4384
rect 14332 4320 14348 4384
rect 14412 4320 14428 4384
rect 14492 4320 14508 4384
rect 14572 4320 14580 4384
rect 14260 3296 14580 4320
rect 14260 3232 14268 3296
rect 14332 3232 14348 3296
rect 14412 3232 14428 3296
rect 14492 3232 14508 3296
rect 14572 3232 14580 3296
rect 14260 2208 14580 3232
rect 14260 2144 14268 2208
rect 14332 2144 14348 2208
rect 14412 2144 14428 2208
rect 14492 2144 14508 2208
rect 14572 2144 14580 2208
rect 14260 2128 14580 2144
rect 16480 16896 16800 17456
rect 16480 16832 16488 16896
rect 16552 16832 16568 16896
rect 16632 16832 16648 16896
rect 16712 16832 16728 16896
rect 16792 16832 16800 16896
rect 16480 15808 16800 16832
rect 16480 15744 16488 15808
rect 16552 15744 16568 15808
rect 16632 15744 16648 15808
rect 16712 15744 16728 15808
rect 16792 15744 16800 15808
rect 16480 14720 16800 15744
rect 16480 14656 16488 14720
rect 16552 14656 16568 14720
rect 16632 14656 16648 14720
rect 16712 14656 16728 14720
rect 16792 14656 16800 14720
rect 16480 13632 16800 14656
rect 16480 13568 16488 13632
rect 16552 13568 16568 13632
rect 16632 13568 16648 13632
rect 16712 13568 16728 13632
rect 16792 13568 16800 13632
rect 16480 12544 16800 13568
rect 16480 12480 16488 12544
rect 16552 12480 16568 12544
rect 16632 12480 16648 12544
rect 16712 12480 16728 12544
rect 16792 12480 16800 12544
rect 16480 11456 16800 12480
rect 16480 11392 16488 11456
rect 16552 11392 16568 11456
rect 16632 11392 16648 11456
rect 16712 11392 16728 11456
rect 16792 11392 16800 11456
rect 16480 10368 16800 11392
rect 16480 10304 16488 10368
rect 16552 10304 16568 10368
rect 16632 10304 16648 10368
rect 16712 10304 16728 10368
rect 16792 10304 16800 10368
rect 16480 9280 16800 10304
rect 16480 9216 16488 9280
rect 16552 9216 16568 9280
rect 16632 9216 16648 9280
rect 16712 9216 16728 9280
rect 16792 9216 16800 9280
rect 16480 8192 16800 9216
rect 16480 8128 16488 8192
rect 16552 8128 16568 8192
rect 16632 8128 16648 8192
rect 16712 8128 16728 8192
rect 16792 8128 16800 8192
rect 16480 7104 16800 8128
rect 16480 7040 16488 7104
rect 16552 7040 16568 7104
rect 16632 7040 16648 7104
rect 16712 7040 16728 7104
rect 16792 7040 16800 7104
rect 16480 6016 16800 7040
rect 16480 5952 16488 6016
rect 16552 5952 16568 6016
rect 16632 5952 16648 6016
rect 16712 5952 16728 6016
rect 16792 5952 16800 6016
rect 16480 4928 16800 5952
rect 16480 4864 16488 4928
rect 16552 4864 16568 4928
rect 16632 4864 16648 4928
rect 16712 4864 16728 4928
rect 16792 4864 16800 4928
rect 16480 3840 16800 4864
rect 16480 3776 16488 3840
rect 16552 3776 16568 3840
rect 16632 3776 16648 3840
rect 16712 3776 16728 3840
rect 16792 3776 16800 3840
rect 16480 2752 16800 3776
rect 16480 2688 16488 2752
rect 16552 2688 16568 2752
rect 16632 2688 16648 2752
rect 16712 2688 16728 2752
rect 16792 2688 16800 2752
rect 16480 2128 16800 2688
rect 18699 17440 19019 17456
rect 18699 17376 18707 17440
rect 18771 17376 18787 17440
rect 18851 17376 18867 17440
rect 18931 17376 18947 17440
rect 19011 17376 19019 17440
rect 18699 16352 19019 17376
rect 18699 16288 18707 16352
rect 18771 16288 18787 16352
rect 18851 16288 18867 16352
rect 18931 16288 18947 16352
rect 19011 16288 19019 16352
rect 18699 15264 19019 16288
rect 18699 15200 18707 15264
rect 18771 15200 18787 15264
rect 18851 15200 18867 15264
rect 18931 15200 18947 15264
rect 19011 15200 19019 15264
rect 18699 14176 19019 15200
rect 18699 14112 18707 14176
rect 18771 14112 18787 14176
rect 18851 14112 18867 14176
rect 18931 14112 18947 14176
rect 19011 14112 19019 14176
rect 18699 13088 19019 14112
rect 18699 13024 18707 13088
rect 18771 13024 18787 13088
rect 18851 13024 18867 13088
rect 18931 13024 18947 13088
rect 19011 13024 19019 13088
rect 18699 12000 19019 13024
rect 18699 11936 18707 12000
rect 18771 11936 18787 12000
rect 18851 11936 18867 12000
rect 18931 11936 18947 12000
rect 19011 11936 19019 12000
rect 18699 10912 19019 11936
rect 18699 10848 18707 10912
rect 18771 10848 18787 10912
rect 18851 10848 18867 10912
rect 18931 10848 18947 10912
rect 19011 10848 19019 10912
rect 18699 9824 19019 10848
rect 18699 9760 18707 9824
rect 18771 9760 18787 9824
rect 18851 9760 18867 9824
rect 18931 9760 18947 9824
rect 19011 9760 19019 9824
rect 18699 8736 19019 9760
rect 18699 8672 18707 8736
rect 18771 8672 18787 8736
rect 18851 8672 18867 8736
rect 18931 8672 18947 8736
rect 19011 8672 19019 8736
rect 18699 7648 19019 8672
rect 18699 7584 18707 7648
rect 18771 7584 18787 7648
rect 18851 7584 18867 7648
rect 18931 7584 18947 7648
rect 19011 7584 19019 7648
rect 18699 6560 19019 7584
rect 18699 6496 18707 6560
rect 18771 6496 18787 6560
rect 18851 6496 18867 6560
rect 18931 6496 18947 6560
rect 19011 6496 19019 6560
rect 18699 5472 19019 6496
rect 18699 5408 18707 5472
rect 18771 5408 18787 5472
rect 18851 5408 18867 5472
rect 18931 5408 18947 5472
rect 19011 5408 19019 5472
rect 18699 4384 19019 5408
rect 18699 4320 18707 4384
rect 18771 4320 18787 4384
rect 18851 4320 18867 4384
rect 18931 4320 18947 4384
rect 19011 4320 19019 4384
rect 18699 3296 19019 4320
rect 18699 3232 18707 3296
rect 18771 3232 18787 3296
rect 18851 3232 18867 3296
rect 18931 3232 18947 3296
rect 19011 3232 19019 3296
rect 18699 2208 19019 3232
rect 18699 2144 18707 2208
rect 18771 2144 18787 2208
rect 18851 2144 18867 2208
rect 18931 2144 18947 2208
rect 19011 2144 19019 2208
rect 18699 2128 19019 2144
use sky130_fd_sc_hd__diode_2  ANTENNA__277__A $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 9108 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__279__A
timestamp 1666464484
transform -1 0 15916 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__300__A
timestamp 1666464484
transform -1 0 18308 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__307__A_N
timestamp 1666464484
transform 1 0 13616 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__311__A_N
timestamp 1666464484
transform 1 0 16836 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__322__A
timestamp 1666464484
transform 1 0 8648 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__356__A
timestamp 1666464484
transform -1 0 18400 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__357__A_N
timestamp 1666464484
transform -1 0 18400 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__370__A
timestamp 1666464484
transform 1 0 3956 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__384__A
timestamp 1666464484
transform 1 0 5888 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__385__B
timestamp 1666464484
transform 1 0 4232 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__387__B1
timestamp 1666464484
transform 1 0 2208 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__390__B1
timestamp 1666464484
transform -1 0 1840 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__392__B1
timestamp 1666464484
transform 1 0 12144 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__394__B1
timestamp 1666464484
transform 1 0 10764 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__398__A
timestamp 1666464484
transform 1 0 7360 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__401__A
timestamp 1666464484
transform 1 0 5520 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__415__B1
timestamp 1666464484
transform 1 0 11040 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__417__C1
timestamp 1666464484
transform 1 0 10856 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__431__A
timestamp 1666464484
transform 1 0 14168 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__433__A
timestamp 1666464484
transform 1 0 13616 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__436__A
timestamp 1666464484
transform 1 0 13892 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__439__A
timestamp 1666464484
transform 1 0 14352 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__442__A
timestamp 1666464484
transform 1 0 13616 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__444__A
timestamp 1666464484
transform 1 0 10396 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__448__A
timestamp 1666464484
transform 1 0 13340 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__454__B
timestamp 1666464484
transform 1 0 11408 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__458__B1
timestamp 1666464484
transform 1 0 11868 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__462__A
timestamp 1666464484
transform 1 0 14720 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__464__C1
timestamp 1666464484
transform 1 0 17756 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__467__A
timestamp 1666464484
transform 1 0 16192 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__469__A
timestamp 1666464484
transform 1 0 11684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__472__B
timestamp 1666464484
transform 1 0 3956 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__476__A
timestamp 1666464484
transform 1 0 3956 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__478__A
timestamp 1666464484
transform 1 0 7360 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__482__A
timestamp 1666464484
transform -1 0 13248 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__484__A
timestamp 1666464484
transform 1 0 12880 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__490__B1
timestamp 1666464484
transform -1 0 5796 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__494__B1
timestamp 1666464484
transform 1 0 3128 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__496__B1
timestamp 1666464484
transform -1 0 1840 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A
timestamp 1666464484
transform 1 0 8464 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1666464484
transform -1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1666464484
transform -1 0 12512 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1932 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3036 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1666464484
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 4324 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 5336 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1666464484
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1666464484
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65
timestamp 1666464484
transform 1 0 7084 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72
timestamp 1666464484
transform 1 0 7728 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1666464484
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1666464484
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_103
timestamp 1666464484
transform 1 0 10580 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1666464484
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1666464484
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_117
timestamp 1666464484
transform 1 0 11868 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1666464484
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_159
timestamp 1666464484
transform 1 0 15732 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1666464484
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_169
timestamp 1666464484
transform 1 0 16652 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_181
timestamp 1666464484
transform 1 0 17756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_187
timestamp 1666464484
transform 1 0 18308 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1666464484
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_15
timestamp 1666464484
transform 1 0 2484 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_34
timestamp 1666464484
transform 1 0 4232 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1666464484
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1666464484
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_66
timestamp 1666464484
transform 1 0 7176 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_88
timestamp 1666464484
transform 1 0 9200 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1666464484
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_113
timestamp 1666464484
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_131
timestamp 1666464484
transform 1 0 13156 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_139
timestamp 1666464484
transform 1 0 13892 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_156
timestamp 1666464484
transform 1 0 15456 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_160
timestamp 1666464484
transform 1 0 15824 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1666464484
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1666464484
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_180
timestamp 1666464484
transform 1 0 17664 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_188
timestamp 1666464484
transform 1 0 18400 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1666464484
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1666464484
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1666464484
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_29
timestamp 1666464484
transform 1 0 3772 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_47
timestamp 1666464484
transform 1 0 5428 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_62
timestamp 1666464484
transform 1 0 6808 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_74
timestamp 1666464484
transform 1 0 7912 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_78
timestamp 1666464484
transform 1 0 8280 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp 1666464484
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_85
timestamp 1666464484
transform 1 0 8924 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_92
timestamp 1666464484
transform 1 0 9568 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_99
timestamp 1666464484
transform 1 0 10212 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_107
timestamp 1666464484
transform 1 0 10948 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_114
timestamp 1666464484
transform 1 0 11592 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_122
timestamp 1666464484
transform 1 0 12328 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1666464484
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1666464484
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 1666464484
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_147
timestamp 1666464484
transform 1 0 14628 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_155
timestamp 1666464484
transform 1 0 15364 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_160
timestamp 1666464484
transform 1 0 15824 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_168
timestamp 1666464484
transform 1 0 16560 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_177
timestamp 1666464484
transform 1 0 17388 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_183
timestamp 1666464484
transform 1 0 17940 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_188
timestamp 1666464484
transform 1 0 18400 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1666464484
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1666464484
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_27
timestamp 1666464484
transform 1 0 3588 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_35
timestamp 1666464484
transform 1 0 4324 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_40
timestamp 1666464484
transform 1 0 4784 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_49
timestamp 1666464484
transform 1 0 5612 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1666464484
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp 1666464484
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_65
timestamp 1666464484
transform 1 0 7084 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_75
timestamp 1666464484
transform 1 0 8004 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_84
timestamp 1666464484
transform 1 0 8832 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_88
timestamp 1666464484
transform 1 0 9200 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1666464484
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1666464484
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_113
timestamp 1666464484
transform 1 0 11500 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_131
timestamp 1666464484
transform 1 0 13156 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_155
timestamp 1666464484
transform 1 0 15364 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1666464484
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_169
timestamp 1666464484
transform 1 0 16652 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_177
timestamp 1666464484
transform 1 0 17388 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_183
timestamp 1666464484
transform 1 0 17940 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_189
timestamp 1666464484
transform 1 0 18492 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1666464484
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_15
timestamp 1666464484
transform 1 0 2484 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_25
timestamp 1666464484
transform 1 0 3404 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_29
timestamp 1666464484
transform 1 0 3772 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_33
timestamp 1666464484
transform 1 0 4140 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_36
timestamp 1666464484
transform 1 0 4416 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_4_50
timestamp 1666464484
transform 1 0 5704 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_56
timestamp 1666464484
transform 1 0 6256 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_62
timestamp 1666464484
transform 1 0 6808 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_82
timestamp 1666464484
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_85
timestamp 1666464484
transform 1 0 8924 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_90
timestamp 1666464484
transform 1 0 9384 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_99
timestamp 1666464484
transform 1 0 10212 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_108
timestamp 1666464484
transform 1 0 11040 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_115
timestamp 1666464484
transform 1 0 11684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_127
timestamp 1666464484
transform 1 0 12788 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_135
timestamp 1666464484
transform 1 0 13524 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp 1666464484
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_141
timestamp 1666464484
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_151
timestamp 1666464484
transform 1 0 14996 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_163
timestamp 1666464484
transform 1 0 16100 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_172
timestamp 1666464484
transform 1 0 16928 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_186
timestamp 1666464484
transform 1 0 18216 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_3
timestamp 1666464484
transform 1 0 1380 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_11
timestamp 1666464484
transform 1 0 2116 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_28
timestamp 1666464484
transform 1 0 3680 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_48
timestamp 1666464484
transform 1 0 5520 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp 1666464484
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_57
timestamp 1666464484
transform 1 0 6348 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_68
timestamp 1666464484
transform 1 0 7360 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_72
timestamp 1666464484
transform 1 0 7728 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_93
timestamp 1666464484
transform 1 0 9660 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_101
timestamp 1666464484
transform 1 0 10396 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_110
timestamp 1666464484
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_113
timestamp 1666464484
transform 1 0 11500 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_133
timestamp 1666464484
transform 1 0 13340 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_5_155
timestamp 1666464484
transform 1 0 15364 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_161
timestamp 1666464484
transform 1 0 15916 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp 1666464484
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_169
timestamp 1666464484
transform 1 0 16652 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_182
timestamp 1666464484
transform 1 0 17848 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_188
timestamp 1666464484
transform 1 0 18400 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_3
timestamp 1666464484
transform 1 0 1380 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_11
timestamp 1666464484
transform 1 0 2116 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_14
timestamp 1666464484
transform 1 0 2392 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_22
timestamp 1666464484
transform 1 0 3128 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1666464484
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_33
timestamp 1666464484
transform 1 0 4140 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_41
timestamp 1666464484
transform 1 0 4876 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_65
timestamp 1666464484
transform 1 0 7084 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_74
timestamp 1666464484
transform 1 0 7912 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82
timestamp 1666464484
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_85
timestamp 1666464484
transform 1 0 8924 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_97
timestamp 1666464484
transform 1 0 10028 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_108
timestamp 1666464484
transform 1 0 11040 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_114
timestamp 1666464484
transform 1 0 11592 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_118
timestamp 1666464484
transform 1 0 11960 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_125
timestamp 1666464484
transform 1 0 12604 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_129
timestamp 1666464484
transform 1 0 12972 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 1666464484
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_141
timestamp 1666464484
transform 1 0 14076 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_147
timestamp 1666464484
transform 1 0 14628 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_150
timestamp 1666464484
transform 1 0 14904 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_162
timestamp 1666464484
transform 1 0 16008 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_166
timestamp 1666464484
transform 1 0 16376 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_173
timestamp 1666464484
transform 1 0 17020 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_182
timestamp 1666464484
transform 1 0 17848 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_188
timestamp 1666464484
transform 1 0 18400 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1666464484
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_15
timestamp 1666464484
transform 1 0 2484 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_22
timestamp 1666464484
transform 1 0 3128 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_30
timestamp 1666464484
transform 1 0 3864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_34
timestamp 1666464484
transform 1 0 4232 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1666464484
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_57
timestamp 1666464484
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_62
timestamp 1666464484
transform 1 0 6808 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_70
timestamp 1666464484
transform 1 0 7544 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_81
timestamp 1666464484
transform 1 0 8556 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_92
timestamp 1666464484
transform 1 0 9568 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_102
timestamp 1666464484
transform 1 0 10488 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_109
timestamp 1666464484
transform 1 0 11132 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_113
timestamp 1666464484
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_119
timestamp 1666464484
transform 1 0 12052 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_125
timestamp 1666464484
transform 1 0 12604 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_129
timestamp 1666464484
transform 1 0 12972 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_135
timestamp 1666464484
transform 1 0 13524 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_147
timestamp 1666464484
transform 1 0 14628 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_157
timestamp 1666464484
transform 1 0 15548 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_163
timestamp 1666464484
transform 1 0 16100 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1666464484
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_169
timestamp 1666464484
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_174
timestamp 1666464484
transform 1 0 17112 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_185
timestamp 1666464484
transform 1 0 18124 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_189
timestamp 1666464484
transform 1 0 18492 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_3
timestamp 1666464484
transform 1 0 1380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_8
timestamp 1666464484
transform 1 0 1840 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_15
timestamp 1666464484
transform 1 0 2484 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_26
timestamp 1666464484
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1666464484
transform 1 0 3772 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_47
timestamp 1666464484
transform 1 0 5428 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_55
timestamp 1666464484
transform 1 0 6164 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_72
timestamp 1666464484
transform 1 0 7728 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_76
timestamp 1666464484
transform 1 0 8096 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_82
timestamp 1666464484
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_85
timestamp 1666464484
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_90
timestamp 1666464484
transform 1 0 9384 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_110
timestamp 1666464484
transform 1 0 11224 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_116
timestamp 1666464484
transform 1 0 11776 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_119
timestamp 1666464484
transform 1 0 12052 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_130
timestamp 1666464484
transform 1 0 13064 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1666464484
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_141
timestamp 1666464484
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_159
timestamp 1666464484
transform 1 0 15732 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_169
timestamp 1666464484
transform 1 0 16652 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_178
timestamp 1666464484
transform 1 0 17480 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_186
timestamp 1666464484
transform 1 0 18216 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_3
timestamp 1666464484
transform 1 0 1380 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_11
timestamp 1666464484
transform 1 0 2116 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_21
timestamp 1666464484
transform 1 0 3036 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_30
timestamp 1666464484
transform 1 0 3864 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_36
timestamp 1666464484
transform 1 0 4416 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_42
timestamp 1666464484
transform 1 0 4968 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_50
timestamp 1666464484
transform 1 0 5704 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1666464484
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_57
timestamp 1666464484
transform 1 0 6348 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_65
timestamp 1666464484
transform 1 0 7084 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_85
timestamp 1666464484
transform 1 0 8924 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_89
timestamp 1666464484
transform 1 0 9292 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_96
timestamp 1666464484
transform 1 0 9936 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_100
timestamp 1666464484
transform 1 0 10304 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_103
timestamp 1666464484
transform 1 0 10580 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_110
timestamp 1666464484
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_113
timestamp 1666464484
transform 1 0 11500 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_131
timestamp 1666464484
transform 1 0 13156 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_139
timestamp 1666464484
transform 1 0 13892 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_151
timestamp 1666464484
transform 1 0 14996 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_163
timestamp 1666464484
transform 1 0 16100 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1666464484
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_169
timestamp 1666464484
transform 1 0 16652 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_9_184
timestamp 1666464484
transform 1 0 18032 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1666464484
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_12
timestamp 1666464484
transform 1 0 2208 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_23
timestamp 1666464484
transform 1 0 3220 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1666464484
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_29
timestamp 1666464484
transform 1 0 3772 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_36
timestamp 1666464484
transform 1 0 4416 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_45
timestamp 1666464484
transform 1 0 5244 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_55
timestamp 1666464484
transform 1 0 6164 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_64
timestamp 1666464484
transform 1 0 6992 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_70
timestamp 1666464484
transform 1 0 7544 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_81
timestamp 1666464484
transform 1 0 8556 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_85
timestamp 1666464484
transform 1 0 8924 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_93
timestamp 1666464484
transform 1 0 9660 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_101
timestamp 1666464484
transform 1 0 10396 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_107
timestamp 1666464484
transform 1 0 10948 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_115
timestamp 1666464484
transform 1 0 11684 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1666464484
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_136
timestamp 1666464484
transform 1 0 13616 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1666464484
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_153
timestamp 1666464484
transform 1 0 15180 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_157
timestamp 1666464484
transform 1 0 15548 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_162
timestamp 1666464484
transform 1 0 16008 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_171
timestamp 1666464484
transform 1 0 16836 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_177
timestamp 1666464484
transform 1 0 17388 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_186
timestamp 1666464484
transform 1 0 18216 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_3
timestamp 1666464484
transform 1 0 1380 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_16
timestamp 1666464484
transform 1 0 2576 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_20
timestamp 1666464484
transform 1 0 2944 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_37
timestamp 1666464484
transform 1 0 4508 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_48
timestamp 1666464484
transform 1 0 5520 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1666464484
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_68
timestamp 1666464484
transform 1 0 7360 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_74
timestamp 1666464484
transform 1 0 7912 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_83
timestamp 1666464484
transform 1 0 8740 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_89
timestamp 1666464484
transform 1 0 9292 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_96
timestamp 1666464484
transform 1 0 9936 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1666464484
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_113
timestamp 1666464484
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_122
timestamp 1666464484
transform 1 0 12328 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_136
timestamp 1666464484
transform 1 0 13616 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_156
timestamp 1666464484
transform 1 0 15456 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1666464484
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp 1666464484
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_173
timestamp 1666464484
transform 1 0 17020 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_183
timestamp 1666464484
transform 1 0 17940 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_189
timestamp 1666464484
transform 1 0 18492 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1666464484
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1666464484
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1666464484
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_29
timestamp 1666464484
transform 1 0 3772 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_37
timestamp 1666464484
transform 1 0 4508 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_44
timestamp 1666464484
transform 1 0 5152 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_51
timestamp 1666464484
transform 1 0 5796 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_60
timestamp 1666464484
transform 1 0 6624 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_68
timestamp 1666464484
transform 1 0 7360 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_74
timestamp 1666464484
transform 1 0 7912 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1666464484
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_85
timestamp 1666464484
transform 1 0 8924 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_89
timestamp 1666464484
transform 1 0 9292 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_100
timestamp 1666464484
transform 1 0 10304 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_113
timestamp 1666464484
transform 1 0 11500 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_127
timestamp 1666464484
transform 1 0 12788 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1666464484
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_141
timestamp 1666464484
transform 1 0 14076 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_147
timestamp 1666464484
transform 1 0 14628 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_156
timestamp 1666464484
transform 1 0 15456 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_169
timestamp 1666464484
transform 1 0 16652 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_181
timestamp 1666464484
transform 1 0 17756 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_188
timestamp 1666464484
transform 1 0 18400 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1666464484
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_15
timestamp 1666464484
transform 1 0 2484 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_33
timestamp 1666464484
transform 1 0 4140 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1666464484
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_57
timestamp 1666464484
transform 1 0 6348 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_64
timestamp 1666464484
transform 1 0 6992 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_84
timestamp 1666464484
transform 1 0 8832 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_13_95
timestamp 1666464484
transform 1 0 9844 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_101
timestamp 1666464484
transform 1 0 10396 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_109
timestamp 1666464484
transform 1 0 11132 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_113
timestamp 1666464484
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_119
timestamp 1666464484
transform 1 0 12052 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_131
timestamp 1666464484
transform 1 0 13156 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_140
timestamp 1666464484
transform 1 0 13984 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_146
timestamp 1666464484
transform 1 0 14536 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_150
timestamp 1666464484
transform 1 0 14904 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_158
timestamp 1666464484
transform 1 0 15640 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_162
timestamp 1666464484
transform 1 0 16008 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1666464484
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_174
timestamp 1666464484
transform 1 0 17112 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_182
timestamp 1666464484
transform 1 0 17848 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_3
timestamp 1666464484
transform 1 0 1380 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_11
timestamp 1666464484
transform 1 0 2116 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_18
timestamp 1666464484
transform 1 0 2760 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_25
timestamp 1666464484
transform 1 0 3404 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1666464484
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_33
timestamp 1666464484
transform 1 0 4140 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_65
timestamp 1666464484
transform 1 0 7084 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_75
timestamp 1666464484
transform 1 0 8004 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_79
timestamp 1666464484
transform 1 0 8372 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1666464484
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_85
timestamp 1666464484
transform 1 0 8924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_107
timestamp 1666464484
transform 1 0 10948 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_117
timestamp 1666464484
transform 1 0 11868 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_132
timestamp 1666464484
transform 1 0 13248 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_138
timestamp 1666464484
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_141
timestamp 1666464484
transform 1 0 14076 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_14_146
timestamp 1666464484
transform 1 0 14536 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_14_160
timestamp 1666464484
transform 1 0 15824 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_174
timestamp 1666464484
transform 1 0 17112 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_185
timestamp 1666464484
transform 1 0 18124 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_189
timestamp 1666464484
transform 1 0 18492 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1666464484
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_15
timestamp 1666464484
transform 1 0 2484 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_19
timestamp 1666464484
transform 1 0 2852 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_27
timestamp 1666464484
transform 1 0 3588 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_36
timestamp 1666464484
transform 1 0 4416 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_43
timestamp 1666464484
transform 1 0 5060 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_54
timestamp 1666464484
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp 1666464484
transform 1 0 6348 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_75
timestamp 1666464484
transform 1 0 8004 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_83
timestamp 1666464484
transform 1 0 8740 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_94
timestamp 1666464484
transform 1 0 9752 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_98
timestamp 1666464484
transform 1 0 10120 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_106
timestamp 1666464484
transform 1 0 10856 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_113
timestamp 1666464484
transform 1 0 11500 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_118
timestamp 1666464484
transform 1 0 11960 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_15_131
timestamp 1666464484
transform 1 0 13156 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_139
timestamp 1666464484
transform 1 0 13892 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_156
timestamp 1666464484
transform 1 0 15456 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_163
timestamp 1666464484
transform 1 0 16100 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1666464484
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1666464484
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_179
timestamp 1666464484
transform 1 0 17572 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_188
timestamp 1666464484
transform 1 0 18400 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1666464484
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_20
timestamp 1666464484
transform 1 0 2944 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1666464484
transform 1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_36
timestamp 1666464484
transform 1 0 4416 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_50
timestamp 1666464484
transform 1 0 5704 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_58
timestamp 1666464484
transform 1 0 6440 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_67
timestamp 1666464484
transform 1 0 7268 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_78
timestamp 1666464484
transform 1 0 8280 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_85
timestamp 1666464484
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_92
timestamp 1666464484
transform 1 0 9568 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_100
timestamp 1666464484
transform 1 0 10304 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_106
timestamp 1666464484
transform 1 0 10856 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_118
timestamp 1666464484
transform 1 0 11960 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_128
timestamp 1666464484
transform 1 0 12880 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1666464484
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_141
timestamp 1666464484
transform 1 0 14076 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_145
timestamp 1666464484
transform 1 0 14444 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_149
timestamp 1666464484
transform 1 0 14812 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_158
timestamp 1666464484
transform 1 0 15640 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_170
timestamp 1666464484
transform 1 0 16744 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_16_183
timestamp 1666464484
transform 1 0 17940 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_189
timestamp 1666464484
transform 1 0 18492 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1666464484
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_15
timestamp 1666464484
transform 1 0 2484 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_34
timestamp 1666464484
transform 1 0 4232 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1666464484
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_57
timestamp 1666464484
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_66
timestamp 1666464484
transform 1 0 7176 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_74
timestamp 1666464484
transform 1 0 7912 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_82
timestamp 1666464484
transform 1 0 8648 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_91
timestamp 1666464484
transform 1 0 9476 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_99
timestamp 1666464484
transform 1 0 10212 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_103
timestamp 1666464484
transform 1 0 10580 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1666464484
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_113
timestamp 1666464484
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_120
timestamp 1666464484
transform 1 0 12144 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_128
timestamp 1666464484
transform 1 0 12880 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_135
timestamp 1666464484
transform 1 0 13524 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_141
timestamp 1666464484
transform 1 0 14076 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_148
timestamp 1666464484
transform 1 0 14720 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_152
timestamp 1666464484
transform 1 0 15088 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1666464484
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1666464484
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1666464484
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_174
timestamp 1666464484
transform 1 0 17112 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_183
timestamp 1666464484
transform 1 0 17940 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_189
timestamp 1666464484
transform 1 0 18492 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_3
timestamp 1666464484
transform 1 0 1380 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_8
timestamp 1666464484
transform 1 0 1840 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_16
timestamp 1666464484
transform 1 0 2576 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_23
timestamp 1666464484
transform 1 0 3220 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1666464484
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_29
timestamp 1666464484
transform 1 0 3772 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_35
timestamp 1666464484
transform 1 0 4324 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_47
timestamp 1666464484
transform 1 0 5428 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_60
timestamp 1666464484
transform 1 0 6624 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_68
timestamp 1666464484
transform 1 0 7360 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1666464484
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_85
timestamp 1666464484
transform 1 0 8924 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_93
timestamp 1666464484
transform 1 0 9660 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_107
timestamp 1666464484
transform 1 0 10948 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_118
timestamp 1666464484
transform 1 0 11960 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_18_130
timestamp 1666464484
transform 1 0 13064 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1666464484
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1666464484
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_159
timestamp 1666464484
transform 1 0 15732 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_174
timestamp 1666464484
transform 1 0 17112 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_184
timestamp 1666464484
transform 1 0 18032 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_19_3
timestamp 1666464484
transform 1 0 1380 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_11
timestamp 1666464484
transform 1 0 2116 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_18
timestamp 1666464484
transform 1 0 2760 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_26
timestamp 1666464484
transform 1 0 3496 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_43
timestamp 1666464484
transform 1 0 5060 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_54
timestamp 1666464484
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_57
timestamp 1666464484
transform 1 0 6348 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_63
timestamp 1666464484
transform 1 0 6900 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_69
timestamp 1666464484
transform 1 0 7452 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_93
timestamp 1666464484
transform 1 0 9660 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_97
timestamp 1666464484
transform 1 0 10028 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_104
timestamp 1666464484
transform 1 0 10672 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1666464484
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_113
timestamp 1666464484
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_118
timestamp 1666464484
transform 1 0 11960 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_130
timestamp 1666464484
transform 1 0 13064 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_144
timestamp 1666464484
transform 1 0 14352 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_156
timestamp 1666464484
transform 1 0 15456 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_160
timestamp 1666464484
transform 1 0 15824 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_164
timestamp 1666464484
transform 1 0 16192 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_169
timestamp 1666464484
transform 1 0 16652 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_180
timestamp 1666464484
transform 1 0 17664 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_188
timestamp 1666464484
transform 1 0 18400 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_3
timestamp 1666464484
transform 1 0 1380 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_11
timestamp 1666464484
transform 1 0 2116 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_18
timestamp 1666464484
transform 1 0 2760 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_24
timestamp 1666464484
transform 1 0 3312 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1666464484
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_41
timestamp 1666464484
transform 1 0 4876 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_65
timestamp 1666464484
transform 1 0 7084 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_72
timestamp 1666464484
transform 1 0 7728 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_78
timestamp 1666464484
transform 1 0 8280 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1666464484
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_85
timestamp 1666464484
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_92
timestamp 1666464484
transform 1 0 9568 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_102
timestamp 1666464484
transform 1 0 10488 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_110
timestamp 1666464484
transform 1 0 11224 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_125
timestamp 1666464484
transform 1 0 12604 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_137
timestamp 1666464484
transform 1 0 13708 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1666464484
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_159
timestamp 1666464484
transform 1 0 15732 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_167
timestamp 1666464484
transform 1 0 16468 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_173
timestamp 1666464484
transform 1 0 17020 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_180
timestamp 1666464484
transform 1 0 17664 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_187
timestamp 1666464484
transform 1 0 18308 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_3
timestamp 1666464484
transform 1 0 1380 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_17
timestamp 1666464484
transform 1 0 2668 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_37
timestamp 1666464484
transform 1 0 4508 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_21_49
timestamp 1666464484
transform 1 0 5612 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1666464484
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_57
timestamp 1666464484
transform 1 0 6348 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_63
timestamp 1666464484
transform 1 0 6900 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_72
timestamp 1666464484
transform 1 0 7728 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_80
timestamp 1666464484
transform 1 0 8464 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_89
timestamp 1666464484
transform 1 0 9292 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_102
timestamp 1666464484
transform 1 0 10488 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_108
timestamp 1666464484
transform 1 0 11040 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_113
timestamp 1666464484
transform 1 0 11500 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_21_130
timestamp 1666464484
transform 1 0 13064 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_138
timestamp 1666464484
transform 1 0 13800 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_145
timestamp 1666464484
transform 1 0 14444 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_152
timestamp 1666464484
transform 1 0 15088 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_160
timestamp 1666464484
transform 1 0 15824 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1666464484
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1666464484
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_178
timestamp 1666464484
transform 1 0 17480 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_186
timestamp 1666464484
transform 1 0 18216 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1666464484
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_15
timestamp 1666464484
transform 1 0 2484 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1666464484
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_29
timestamp 1666464484
transform 1 0 3772 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_49
timestamp 1666464484
transform 1 0 5612 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_59
timestamp 1666464484
transform 1 0 6532 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_79
timestamp 1666464484
transform 1 0 8372 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1666464484
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_85
timestamp 1666464484
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_103
timestamp 1666464484
transform 1 0 10580 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_107
timestamp 1666464484
transform 1 0 10948 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_111
timestamp 1666464484
transform 1 0 11316 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_123
timestamp 1666464484
transform 1 0 12420 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1666464484
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1666464484
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_141
timestamp 1666464484
transform 1 0 14076 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_150
timestamp 1666464484
transform 1 0 14904 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_158
timestamp 1666464484
transform 1 0 15640 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_168
timestamp 1666464484
transform 1 0 16560 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_180
timestamp 1666464484
transform 1 0 17664 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_188
timestamp 1666464484
transform 1 0 18400 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1666464484
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_15
timestamp 1666464484
transform 1 0 2484 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_19
timestamp 1666464484
transform 1 0 2852 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_36
timestamp 1666464484
transform 1 0 4416 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_48
timestamp 1666464484
transform 1 0 5520 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1666464484
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1666464484
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_57
timestamp 1666464484
transform 1 0 6348 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_65
timestamp 1666464484
transform 1 0 7084 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_72
timestamp 1666464484
transform 1 0 7728 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_80
timestamp 1666464484
transform 1 0 8464 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_84
timestamp 1666464484
transform 1 0 8832 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_91
timestamp 1666464484
transform 1 0 9476 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_100
timestamp 1666464484
transform 1 0 10304 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_107
timestamp 1666464484
transform 1 0 10948 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1666464484
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_113
timestamp 1666464484
transform 1 0 11500 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_117
timestamp 1666464484
transform 1 0 11868 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_134
timestamp 1666464484
transform 1 0 13432 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_154
timestamp 1666464484
transform 1 0 15272 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1666464484
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1666464484
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_178
timestamp 1666464484
transform 1 0 17480 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1666464484
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_15
timestamp 1666464484
transform 1 0 2484 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_26
timestamp 1666464484
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1666464484
transform 1 0 3772 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_36
timestamp 1666464484
transform 1 0 4416 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_44
timestamp 1666464484
transform 1 0 5152 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_61
timestamp 1666464484
transform 1 0 6716 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_81
timestamp 1666464484
transform 1 0 8556 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_24_85
timestamp 1666464484
transform 1 0 8924 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_107
timestamp 1666464484
transform 1 0 10948 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_122
timestamp 1666464484
transform 1 0 12328 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_129
timestamp 1666464484
transform 1 0 12972 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_137
timestamp 1666464484
transform 1 0 13708 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_141
timestamp 1666464484
transform 1 0 14076 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_145
timestamp 1666464484
transform 1 0 14444 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_151
timestamp 1666464484
transform 1 0 14996 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_161
timestamp 1666464484
transform 1 0 15916 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_173
timestamp 1666464484
transform 1 0 17020 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_185
timestamp 1666464484
transform 1 0 18124 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_189
timestamp 1666464484
transform 1 0 18492 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1666464484
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_15
timestamp 1666464484
transform 1 0 2484 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_21
timestamp 1666464484
transform 1 0 3036 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_38
timestamp 1666464484
transform 1 0 4600 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_50
timestamp 1666464484
transform 1 0 5704 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 1666464484
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_57
timestamp 1666464484
transform 1 0 6348 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_64
timestamp 1666464484
transform 1 0 6992 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_72
timestamp 1666464484
transform 1 0 7728 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_78
timestamp 1666464484
transform 1 0 8280 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_98
timestamp 1666464484
transform 1 0 10120 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1666464484
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1666464484
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_113
timestamp 1666464484
transform 1 0 11500 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_125
timestamp 1666464484
transform 1 0 12604 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_132
timestamp 1666464484
transform 1 0 13248 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_136
timestamp 1666464484
transform 1 0 13616 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_153
timestamp 1666464484
transform 1 0 15180 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_165
timestamp 1666464484
transform 1 0 16284 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1666464484
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_181
timestamp 1666464484
transform 1 0 17756 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_189
timestamp 1666464484
transform 1 0 18492 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1666464484
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_15
timestamp 1666464484
transform 1 0 2484 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_23
timestamp 1666464484
transform 1 0 3220 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1666464484
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1666464484
transform 1 0 3772 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_33
timestamp 1666464484
transform 1 0 4140 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_45
timestamp 1666464484
transform 1 0 5244 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_62
timestamp 1666464484
transform 1 0 6808 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1666464484
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_85
timestamp 1666464484
transform 1 0 8924 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_97
timestamp 1666464484
transform 1 0 10028 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_117
timestamp 1666464484
transform 1 0 11868 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_126
timestamp 1666464484
transform 1 0 12696 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_132
timestamp 1666464484
transform 1 0 13248 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1666464484
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1666464484
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1666464484
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1666464484
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_189
timestamp 1666464484
transform 1 0 18492 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1666464484
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_15
timestamp 1666464484
transform 1 0 2484 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_24
timestamp 1666464484
transform 1 0 3312 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_29
timestamp 1666464484
transform 1 0 3772 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_47
timestamp 1666464484
transform 1 0 5428 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1666464484
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_57
timestamp 1666464484
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_64
timestamp 1666464484
transform 1 0 6992 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_70
timestamp 1666464484
transform 1 0 7544 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_82
timestamp 1666464484
transform 1 0 8648 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_85
timestamp 1666464484
transform 1 0 8924 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_90
timestamp 1666464484
transform 1 0 9384 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_96
timestamp 1666464484
transform 1 0 9936 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_102
timestamp 1666464484
transform 1 0 10488 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_109
timestamp 1666464484
transform 1 0 11132 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1666464484
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_118
timestamp 1666464484
transform 1 0 11960 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_124
timestamp 1666464484
transform 1 0 12512 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_130
timestamp 1666464484
transform 1 0 13064 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_138
timestamp 1666464484
transform 1 0 13800 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_141
timestamp 1666464484
transform 1 0 14076 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_153
timestamp 1666464484
transform 1 0 15180 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_161
timestamp 1666464484
transform 1 0 15916 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1666464484
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1666464484
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_181
timestamp 1666464484
transform 1 0 17756 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_189
timestamp 1666464484
transform 1 0 18492 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1666464484
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1666464484
transform -1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1666464484
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1666464484
transform -1 0 18860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1666464484
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1666464484
transform -1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1666464484
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1666464484
transform -1 0 18860 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1666464484
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1666464484
transform -1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1666464484
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1666464484
transform -1 0 18860 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1666464484
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1666464484
transform -1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1666464484
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1666464484
transform -1 0 18860 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1666464484
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1666464484
transform -1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1666464484
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1666464484
transform -1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1666464484
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1666464484
transform -1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1666464484
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1666464484
transform -1 0 18860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1666464484
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1666464484
transform -1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1666464484
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1666464484
transform -1 0 18860 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1666464484
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1666464484
transform -1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1666464484
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1666464484
transform -1 0 18860 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1666464484
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1666464484
transform -1 0 18860 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1666464484
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1666464484
transform -1 0 18860 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1666464484
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1666464484
transform -1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1666464484
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1666464484
transform -1 0 18860 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1666464484
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1666464484
transform -1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1666464484
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1666464484
transform -1 0 18860 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1666464484
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1666464484
transform -1 0 18860 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1666464484
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1666464484
transform -1 0 18860 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1666464484
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1666464484
transform -1 0 18860 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1666464484
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1666464484
transform -1 0 18860 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1666464484
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1666464484
transform -1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1666464484
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1666464484
transform -1 0 18860 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1666464484
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1666464484
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1666464484
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1666464484
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1666464484
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1666464484
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1666464484
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1666464484
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1666464484
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1666464484
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1666464484
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1666464484
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1666464484
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1666464484
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1666464484
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1666464484
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1666464484
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1666464484
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1666464484
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1666464484
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1666464484
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1666464484
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1666464484
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1666464484
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1666464484
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1666464484
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1666464484
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1666464484
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1666464484
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1666464484
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1666464484
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1666464484
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1666464484
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1666464484
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1666464484
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1666464484
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1666464484
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1666464484
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1666464484
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1666464484
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1666464484
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1666464484
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1666464484
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1666464484
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1666464484
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1666464484
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1666464484
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1666464484
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1666464484
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1666464484
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1666464484
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1666464484
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1666464484
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1666464484
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1666464484
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1666464484
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1666464484
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1666464484
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1666464484
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1666464484
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1666464484
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1666464484
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1666464484
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1666464484
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1666464484
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1666464484
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1666464484
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1666464484
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1666464484
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1666464484
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1666464484
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1666464484
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1666464484
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1666464484
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1666464484
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1666464484
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1666464484
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1666464484
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1666464484
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1666464484
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1666464484
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1666464484
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1666464484
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1666464484
transform 1 0 3680 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1666464484
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1666464484
transform 1 0 8832 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1666464484
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1666464484
transform 1 0 13984 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1666464484
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _252_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 4140 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _253_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2392 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _254_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 4876 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _255_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 3864 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _256_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2576 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _257_
timestamp 1666464484
transform 1 0 1564 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _258_
timestamp 1666464484
transform 1 0 1932 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _259_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 6532 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _260_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 17664 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _261_
timestamp 1666464484
transform -1 0 9568 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _262_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 17664 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _263_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 17848 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nor2b_1  _264_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 17020 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _265_
timestamp 1666464484
transform -1 0 17664 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _266_
timestamp 1666464484
transform 1 0 11960 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _267_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 16376 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _268_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 17480 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _269_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 15732 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _270_
timestamp 1666464484
transform -1 0 9568 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _271_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 7544 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _272_
timestamp 1666464484
transform 1 0 12604 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _273_
timestamp 1666464484
transform -1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nor2b_2  _274_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 13064 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _275_
timestamp 1666464484
transform -1 0 13064 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _276_
timestamp 1666464484
transform 1 0 13524 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _277_
timestamp 1666464484
transform 1 0 9384 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _278_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 18032 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _279_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 16376 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _280_
timestamp 1666464484
transform 1 0 10212 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _281_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 13248 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _282_
timestamp 1666464484
transform 1 0 16836 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _283_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 17480 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nand4b_1  _284_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 16836 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _285_
timestamp 1666464484
transform 1 0 17480 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _286_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 18124 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _287_
timestamp 1666464484
transform 1 0 16008 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _288_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 16008 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _289_
timestamp 1666464484
transform 1 0 10948 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _290_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 12788 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _291_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 13984 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _292_
timestamp 1666464484
transform -1 0 13616 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _293_
timestamp 1666464484
transform -1 0 17940 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _294_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 17112 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _295_
timestamp 1666464484
transform -1 0 12144 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _296_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 12512 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _297_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 12880 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _298_
timestamp 1666464484
transform -1 0 13524 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _299_
timestamp 1666464484
transform -1 0 16836 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2b_1  _300_
timestamp 1666464484
transform 1 0 15916 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _301_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 17020 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _302_
timestamp 1666464484
transform 1 0 14996 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _303_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 16008 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _304_
timestamp 1666464484
transform -1 0 13800 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _305_
timestamp 1666464484
transform 1 0 16100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _306_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 17848 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__and4b_1  _307_
timestamp 1666464484
transform -1 0 14996 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _308_
timestamp 1666464484
transform 1 0 17388 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _309_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 17480 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _310_
timestamp 1666464484
transform 1 0 18124 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _311_
timestamp 1666464484
transform -1 0 17756 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nor3b_1  _312_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 17388 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _313_
timestamp 1666464484
transform 1 0 17204 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and4b_1  _314_
timestamp 1666464484
transform -1 0 13616 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nand3b_1  _315_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 16560 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _316_
timestamp 1666464484
transform -1 0 17940 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _317_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 16836 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_1  _318_
timestamp 1666464484
transform -1 0 12052 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _319_
timestamp 1666464484
transform 1 0 10396 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _320_
timestamp 1666464484
transform -1 0 11868 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _321_
timestamp 1666464484
transform -1 0 10948 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _322_
timestamp 1666464484
transform -1 0 8648 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _323_
timestamp 1666464484
transform -1 0 12236 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _324_
timestamp 1666464484
transform 1 0 10672 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _325_
timestamp 1666464484
transform 1 0 10488 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _326_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 12328 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _327_
timestamp 1666464484
transform 1 0 9016 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _328_
timestamp 1666464484
transform 1 0 9200 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _329_
timestamp 1666464484
transform 1 0 10120 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _330_
timestamp 1666464484
transform 1 0 10856 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _331_
timestamp 1666464484
transform 1 0 4508 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _332_
timestamp 1666464484
transform 1 0 4692 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _333_
timestamp 1666464484
transform 1 0 5796 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _334_
timestamp 1666464484
transform 1 0 7912 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a31oi_2  _335_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 8556 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  _336_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 10028 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_4  _337_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 8924 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__and2_1  _338_
timestamp 1666464484
transform 1 0 4784 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _339_
timestamp 1666464484
transform -1 0 5796 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _340_
timestamp 1666464484
transform 1 0 5796 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _341_
timestamp 1666464484
transform 1 0 6532 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _342_
timestamp 1666464484
transform -1 0 6624 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _343_
timestamp 1666464484
transform 1 0 8188 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _344_
timestamp 1666464484
transform -1 0 7360 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _345_
timestamp 1666464484
transform 1 0 9108 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _346_
timestamp 1666464484
transform 1 0 8924 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_2  _347_
timestamp 1666464484
transform 1 0 6624 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_1  _348_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 11960 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _349_
timestamp 1666464484
transform -1 0 10580 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _350_
timestamp 1666464484
transform 1 0 11684 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and4bb_2  _351_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 10028 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__or3_1  _352_
timestamp 1666464484
transform -1 0 17480 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_1  _353_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 18400 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _354_
timestamp 1666464484
transform -1 0 17112 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _355_
timestamp 1666464484
transform 1 0 16836 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _356_
timestamp 1666464484
transform 1 0 17204 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _357_
timestamp 1666464484
transform 1 0 17204 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_1  _358_
timestamp 1666464484
transform 1 0 17664 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _359_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 17480 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _360_
timestamp 1666464484
transform -1 0 16100 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a2111o_1  _361_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 15824 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _362_
timestamp 1666464484
transform 1 0 12512 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _363_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 12236 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _364_
timestamp 1666464484
transform 1 0 13156 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nor4_2  _365_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 11868 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__or4b_1  _366_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 8740 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _367_
timestamp 1666464484
transform 1 0 8280 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _368_
timestamp 1666464484
transform 1 0 6532 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _369_
timestamp 1666464484
transform 1 0 9936 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _370_
timestamp 1666464484
transform -1 0 4876 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _371_
timestamp 1666464484
transform 1 0 6532 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_1  _372_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 6532 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _373_
timestamp 1666464484
transform 1 0 8372 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _374_
timestamp 1666464484
transform -1 0 7912 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _375_
timestamp 1666464484
transform -1 0 6808 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _376_
timestamp 1666464484
transform 1 0 6348 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _377_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 6532 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a31oi_1  _378_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 8832 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _379_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 7176 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _380_
timestamp 1666464484
transform 1 0 7452 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _381_
timestamp 1666464484
transform 1 0 7452 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _382_
timestamp 1666464484
transform -1 0 10212 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _383_
timestamp 1666464484
transform -1 0 5336 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _384_
timestamp 1666464484
transform -1 0 5704 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _385_
timestamp 1666464484
transform -1 0 4232 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _386_
timestamp 1666464484
transform 1 0 9384 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _387_
timestamp 1666464484
transform -1 0 3128 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _388_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 3404 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _389_
timestamp 1666464484
transform 1 0 2760 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _390_
timestamp 1666464484
transform 1 0 2852 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _391_
timestamp 1666464484
transform -1 0 2484 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _392_
timestamp 1666464484
transform 1 0 12696 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _393_
timestamp 1666464484
transform 1 0 9200 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _394_
timestamp 1666464484
transform -1 0 10396 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _395_
timestamp 1666464484
transform -1 0 9936 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _396_
timestamp 1666464484
transform 1 0 8372 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _397_
timestamp 1666464484
transform -1 0 7268 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _398_
timestamp 1666464484
transform -1 0 7084 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _399_
timestamp 1666464484
transform -1 0 9752 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _400_
timestamp 1666464484
transform -1 0 8648 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _401_
timestamp 1666464484
transform -1 0 6072 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _402_
timestamp 1666464484
transform 1 0 7452 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _403_
timestamp 1666464484
transform 1 0 7452 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _404_
timestamp 1666464484
transform 1 0 10856 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _405_
timestamp 1666464484
transform 1 0 3220 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _406_
timestamp 1666464484
transform 1 0 6992 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _407_
timestamp 1666464484
transform 1 0 7636 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _408_
timestamp 1666464484
transform 1 0 6992 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _409_
timestamp 1666464484
transform 1 0 6992 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _410_
timestamp 1666464484
transform -1 0 6624 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _411_
timestamp 1666464484
transform 1 0 5796 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _412_
timestamp 1666464484
transform -1 0 7176 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _413_
timestamp 1666464484
transform 1 0 6072 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _414_
timestamp 1666464484
transform 1 0 8004 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _415_
timestamp 1666464484
transform -1 0 8648 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _416_
timestamp 1666464484
transform -1 0 9292 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a211oi_1  _417_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 10488 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _418_
timestamp 1666464484
transform 1 0 9844 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _419_
timestamp 1666464484
transform 1 0 9844 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _420_
timestamp 1666464484
transform -1 0 9476 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_2  _421_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 9660 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _422_
timestamp 1666464484
transform 1 0 11040 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _423_
timestamp 1666464484
transform -1 0 12420 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _424_
timestamp 1666464484
transform -1 0 11960 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _425_
timestamp 1666464484
transform -1 0 12972 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _426_
timestamp 1666464484
transform 1 0 12052 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _427_
timestamp 1666464484
transform -1 0 13248 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _428_
timestamp 1666464484
transform -1 0 12604 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _429_
timestamp 1666464484
transform 1 0 14536 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _430_
timestamp 1666464484
transform -1 0 14904 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _431_
timestamp 1666464484
transform 1 0 14812 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _432_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 14720 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _433_
timestamp 1666464484
transform -1 0 14444 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _434_
timestamp 1666464484
transform -1 0 16192 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _435_
timestamp 1666464484
transform 1 0 15180 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _436_
timestamp 1666464484
transform -1 0 14720 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _437_
timestamp 1666464484
transform 1 0 15364 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _438_
timestamp 1666464484
transform 1 0 15088 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _439_
timestamp 1666464484
transform -1 0 14812 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _440_
timestamp 1666464484
transform -1 0 16008 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _441_
timestamp 1666464484
transform 1 0 14720 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _442_
timestamp 1666464484
transform 1 0 14628 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _443_
timestamp 1666464484
transform -1 0 11224 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _444_
timestamp 1666464484
transform -1 0 11224 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _445_
timestamp 1666464484
transform -1 0 14996 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and4b_1  _446_
timestamp 1666464484
transform 1 0 15364 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _447_
timestamp 1666464484
transform -1 0 16008 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _448_
timestamp 1666464484
transform -1 0 13800 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _449_
timestamp 1666464484
transform -1 0 10028 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _450_
timestamp 1666464484
transform 1 0 9108 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _451_
timestamp 1666464484
transform -1 0 10212 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _452_
timestamp 1666464484
transform -1 0 9568 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _453_
timestamp 1666464484
transform 1 0 10396 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _454_
timestamp 1666464484
transform -1 0 11224 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _455_
timestamp 1666464484
transform 1 0 10580 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _456_
timestamp 1666464484
transform -1 0 11684 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _457_
timestamp 1666464484
transform -1 0 12972 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _458_
timestamp 1666464484
transform 1 0 12052 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _459_
timestamp 1666464484
transform -1 0 12052 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _460_
timestamp 1666464484
transform -1 0 16376 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _461_
timestamp 1666464484
transform -1 0 16928 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _462_
timestamp 1666464484
transform -1 0 16100 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _463_
timestamp 1666464484
transform 1 0 16100 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _464_
timestamp 1666464484
transform -1 0 17388 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _465_
timestamp 1666464484
transform -1 0 16560 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _466_
timestamp 1666464484
transform 1 0 16928 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _467_
timestamp 1666464484
transform 1 0 18032 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _468_
timestamp 1666464484
transform 1 0 16836 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _469_
timestamp 1666464484
transform -1 0 16376 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _470_
timestamp 1666464484
transform 1 0 3956 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _471_
timestamp 1666464484
transform 1 0 4784 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _472_
timestamp 1666464484
transform 1 0 2300 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _473_
timestamp 1666464484
transform -1 0 3404 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _474_
timestamp 1666464484
transform -1 0 3496 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _475_
timestamp 1666464484
transform -1 0 2852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _476_
timestamp 1666464484
transform -1 0 3220 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _477_
timestamp 1666464484
transform -1 0 3312 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _478_
timestamp 1666464484
transform -1 0 6992 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _479_
timestamp 1666464484
transform 1 0 5796 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _480_
timestamp 1666464484
transform -1 0 6992 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _481_
timestamp 1666464484
transform 1 0 5796 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _482_
timestamp 1666464484
transform 1 0 12236 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _483_
timestamp 1666464484
transform 1 0 11684 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _484_
timestamp 1666464484
transform 1 0 10028 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _485_
timestamp 1666464484
transform -1 0 10764 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _486_
timestamp 1666464484
transform 1 0 7820 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _487_
timestamp 1666464484
transform 1 0 9108 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _488_
timestamp 1666464484
transform 1 0 6624 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _489_
timestamp 1666464484
transform 1 0 7452 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _490_
timestamp 1666464484
transform 1 0 5244 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _491_
timestamp 1666464484
transform -1 0 6532 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _492_
timestamp 1666464484
transform -1 0 4416 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _493_
timestamp 1666464484
transform -1 0 3496 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _494_
timestamp 1666464484
transform 1 0 2392 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _495_
timestamp 1666464484
transform 1 0 2116 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _496_
timestamp 1666464484
transform 1 0 2208 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _497_
timestamp 1666464484
transform -1 0 2760 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _498_
timestamp 1666464484
transform -1 0 4416 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _499_
timestamp 1666464484
transform -1 0 4324 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _500_
timestamp 1666464484
transform 1 0 2484 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _501_
timestamp 1666464484
transform -1 0 3220 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _502_
timestamp 1666464484
transform -1 0 5612 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _503_
timestamp 1666464484
transform -1 0 4784 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _504_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2760 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _505_
timestamp 1666464484
transform -1 0 5428 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _506_
timestamp 1666464484
transform 1 0 7728 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _507_
timestamp 1666464484
transform 1 0 9108 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _508_
timestamp 1666464484
transform 1 0 11684 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _509_
timestamp 1666464484
transform 1 0 9752 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _510_
timestamp 1666464484
transform 1 0 4048 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _511_
timestamp 1666464484
transform -1 0 3680 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _512_
timestamp 1666464484
transform -1 0 5428 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _513_
timestamp 1666464484
transform 1 0 12236 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _514_
timestamp 1666464484
transform 1 0 9752 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _515_
timestamp 1666464484
transform 1 0 7360 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _516_
timestamp 1666464484
transform 1 0 6532 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _517_
timestamp 1666464484
transform 1 0 6900 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _518_
timestamp 1666464484
transform 1 0 5612 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _519_
timestamp 1666464484
transform 1 0 4600 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _520_
timestamp 1666464484
transform 1 0 9108 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _521_
timestamp 1666464484
transform 1 0 9476 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _522_
timestamp 1666464484
transform 1 0 11960 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _523_
timestamp 1666464484
transform 1 0 13708 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _524_
timestamp 1666464484
transform 1 0 13800 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _525_
timestamp 1666464484
transform 1 0 14260 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _526_
timestamp 1666464484
transform 1 0 14260 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _527_
timestamp 1666464484
transform 1 0 13984 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _528_
timestamp 1666464484
transform 1 0 13984 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _529_
timestamp 1666464484
transform 1 0 11684 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _530_
timestamp 1666464484
transform 1 0 14260 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _531_
timestamp 1666464484
transform 1 0 9292 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _532_
timestamp 1666464484
transform 1 0 11684 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _533_
timestamp 1666464484
transform 1 0 11868 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _534_
timestamp 1666464484
transform 1 0 13892 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _535_
timestamp 1666464484
transform 1 0 13892 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _536_
timestamp 1666464484
transform 1 0 14260 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _537_
timestamp 1666464484
transform 1 0 13984 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _538_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 4508 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _539_
timestamp 1666464484
transform 1 0 3036 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _540_
timestamp 1666464484
transform -1 0 4140 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _541_
timestamp 1666464484
transform -1 0 4600 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _542_
timestamp 1666464484
transform -1 0 5428 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _543_
timestamp 1666464484
transform 1 0 5336 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _544_
timestamp 1666464484
transform -1 0 8648 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _545_
timestamp 1666464484
transform 1 0 10396 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _546_
timestamp 1666464484
transform 1 0 8648 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _547_
timestamp 1666464484
transform 1 0 7084 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _548_
timestamp 1666464484
transform 1 0 5244 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _549_
timestamp 1666464484
transform 1 0 4140 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _550_
timestamp 1666464484
transform 1 0 2944 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _551_
timestamp 1666464484
transform -1 0 4508 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _552_
timestamp 1666464484
transform -1 0 5060 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _553_
timestamp 1666464484
transform 1 0 2760 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _554_
timestamp 1666464484
transform 1 0 4600 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _555_
timestamp 1666464484
transform 1 0 7176 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _556_
timestamp 1666464484
transform 1 0 6256 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _557_
timestamp 1666464484
transform 1 0 4600 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 9108 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1666464484
transform -1 0 7084 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1666464484
transform 1 0 7820 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1666464484
transform -1 0 7084 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1666464484
transform -1 0 9660 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 16836 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1666464484
transform 1 0 10856 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output3
timestamp 1666464484
transform -1 0 1932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output4
timestamp 1666464484
transform -1 0 4324 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output5
timestamp 1666464484
transform -1 0 6072 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp 1666464484
transform -1 0 8648 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp 1666464484
transform 1 0 11224 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp 1666464484
transform 1 0 14260 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 1666464484
transform 1 0 15456 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 1666464484
transform 1 0 18032 0 1 3264
box -38 -48 406 592
<< labels >>
flabel metal2 s 3330 19200 3386 20000 0 FreeSans 224 90 0 0 clk
port 0 nsew signal input
flabel metal2 s 16578 19200 16634 20000 0 FreeSans 224 90 0 0 io_in
port 1 nsew signal input
flabel metal2 s 1214 0 1270 800 0 FreeSans 224 90 0 0 io_out[0]
port 2 nsew signal tristate
flabel metal2 s 3698 0 3754 800 0 FreeSans 224 90 0 0 io_out[1]
port 3 nsew signal tristate
flabel metal2 s 6182 0 6238 800 0 FreeSans 224 90 0 0 io_out[2]
port 4 nsew signal tristate
flabel metal2 s 8666 0 8722 800 0 FreeSans 224 90 0 0 io_out[3]
port 5 nsew signal tristate
flabel metal2 s 11150 0 11206 800 0 FreeSans 224 90 0 0 io_out[4]
port 6 nsew signal tristate
flabel metal2 s 13634 0 13690 800 0 FreeSans 224 90 0 0 io_out[5]
port 7 nsew signal tristate
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 io_out[6]
port 8 nsew signal tristate
flabel metal2 s 18602 0 18658 800 0 FreeSans 224 90 0 0 io_out[7]
port 9 nsew signal tristate
flabel metal2 s 9954 19200 10010 20000 0 FreeSans 224 90 0 0 rst
port 10 nsew signal input
flabel metal4 s 3163 2128 3483 17456 0 FreeSans 1920 90 0 0 vccd1
port 11 nsew power bidirectional
flabel metal4 s 7602 2128 7922 17456 0 FreeSans 1920 90 0 0 vccd1
port 11 nsew power bidirectional
flabel metal4 s 12041 2128 12361 17456 0 FreeSans 1920 90 0 0 vccd1
port 11 nsew power bidirectional
flabel metal4 s 16480 2128 16800 17456 0 FreeSans 1920 90 0 0 vccd1
port 11 nsew power bidirectional
flabel metal4 s 5382 2128 5702 17456 0 FreeSans 1920 90 0 0 vssd1
port 12 nsew ground bidirectional
flabel metal4 s 9821 2128 10141 17456 0 FreeSans 1920 90 0 0 vssd1
port 12 nsew ground bidirectional
flabel metal4 s 14260 2128 14580 17456 0 FreeSans 1920 90 0 0 vssd1
port 12 nsew ground bidirectional
flabel metal4 s 18699 2128 19019 17456 0 FreeSans 1920 90 0 0 vssd1
port 12 nsew ground bidirectional
rlabel metal1 9982 16864 9982 16864 0 vccd1
rlabel via1 10061 17408 10061 17408 0 vssd1
rlabel metal1 6486 3162 6486 3162 0 _000_
rlabel metal1 7482 3094 7482 3094 0 _001_
rlabel metal1 9230 2346 9230 2346 0 _002_
rlabel metal1 8832 2618 8832 2618 0 _003_
rlabel metal1 10207 3026 10207 3026 0 _004_
rlabel metal1 4876 2618 4876 2618 0 _005_
rlabel metal1 4268 5202 4268 5202 0 _006_
rlabel metal1 3450 4794 3450 4794 0 _007_
rlabel metal1 3730 6698 3730 6698 0 _008_
rlabel metal1 12645 2346 12645 2346 0 _009_
rlabel metal1 9972 6766 9972 6766 0 _010_
rlabel metal1 7268 7514 7268 7514 0 _011_
rlabel metal1 7452 10234 7452 10234 0 _012_
rlabel metal2 7038 14178 7038 14178 0 _013_
rlabel metal1 5888 12954 5888 12954 0 _014_
rlabel metal1 5515 11730 5515 11730 0 _015_
rlabel metal2 9246 14178 9246 14178 0 _016_
rlabel metal1 9568 15130 9568 15130 0 _017_
rlabel metal2 12558 14790 12558 14790 0 _018_
rlabel metal1 13646 16150 13646 16150 0 _019_
rlabel metal2 14950 14518 14950 14518 0 _020_
rlabel metal1 14480 13294 14480 13294 0 _021_
rlabel metal1 14628 11866 14628 11866 0 _022_
rlabel metal1 14485 10710 14485 10710 0 _023_
rlabel metal1 14485 8534 14485 8534 0 _024_
rlabel metal1 11530 7446 11530 7446 0 _025_
rlabel metal1 14152 6698 14152 6698 0 _026_
rlabel metal1 9568 3706 9568 3706 0 _027_
rlabel metal1 11806 4182 11806 4182 0 _028_
rlabel metal1 12088 5202 12088 5202 0 _029_
rlabel metal2 15870 4998 15870 4998 0 _030_
rlabel metal1 14853 4114 14853 4114 0 _031_
rlabel metal1 16325 2346 16325 2346 0 _032_
rlabel metal1 16008 2482 16008 2482 0 _033_
rlabel via1 4825 9554 4825 9554 0 _034_
rlabel metal1 3491 8466 3491 8466 0 _035_
rlabel metal1 3316 9622 3316 9622 0 _036_
rlabel via1 4282 16150 4282 16150 0 _037_
rlabel metal1 5489 17238 5489 17238 0 _038_
rlabel metal2 5842 16354 5842 16354 0 _039_
rlabel metal1 9031 16490 9031 16490 0 _040_
rlabel metal2 10718 16354 10718 16354 0 _041_
rlabel via1 8965 16082 8965 16082 0 _042_
rlabel metal2 7498 15266 7498 15266 0 _043_
rlabel metal2 6486 14994 6486 14994 0 _044_
rlabel metal1 3940 14314 3940 14314 0 _045_
rlabel metal2 3082 14382 3082 14382 0 _046_
rlabel metal2 4186 13430 4186 13430 0 _047_
rlabel metal1 4512 12818 4512 12818 0 _048_
rlabel via1 3077 11730 3077 11730 0 _049_
rlabel metal1 5382 4148 5382 4148 0 _050_
rlabel metal1 7723 4590 7723 4590 0 _051_
rlabel via1 6573 6766 6573 6766 0 _052_
rlabel metal1 4820 3026 4820 3026 0 _053_
rlabel metal1 4554 7922 4554 7922 0 _054_
rlabel metal2 5014 8772 5014 8772 0 _055_
rlabel metal1 6118 8330 6118 8330 0 _056_
rlabel metal2 3450 7684 3450 7684 0 _057_
rlabel metal2 2622 8262 2622 8262 0 _058_
rlabel metal1 2116 8058 2116 8058 0 _059_
rlabel metal2 6026 7888 6026 7888 0 _060_
rlabel metal1 8326 7412 8326 7412 0 _061_
rlabel metal1 16422 11526 16422 11526 0 _062_
rlabel metal2 7222 13362 7222 13362 0 _063_
rlabel metal1 17204 12818 17204 12818 0 _064_
rlabel metal1 16836 13294 16836 13294 0 _065_
rlabel metal1 16974 12750 16974 12750 0 _066_
rlabel metal1 16192 12682 16192 12682 0 _067_
rlabel metal1 12650 13158 12650 13158 0 _068_
rlabel metal2 15870 15266 15870 15266 0 _069_
rlabel metal1 16606 13702 16606 13702 0 _070_
rlabel metal1 15824 14246 15824 14246 0 _071_
rlabel metal1 8004 8942 8004 8942 0 _072_
rlabel metal1 14444 10098 14444 10098 0 _073_
rlabel metal2 13202 10744 13202 10744 0 _074_
rlabel metal2 12650 14246 12650 14246 0 _075_
rlabel metal2 12466 13328 12466 13328 0 _076_
rlabel metal1 13202 11186 13202 11186 0 _077_
rlabel metal1 17158 2618 17158 2618 0 _078_
rlabel metal1 10396 10642 10396 10642 0 _079_
rlabel metal2 18078 13668 18078 13668 0 _080_
rlabel metal1 15732 14042 15732 14042 0 _081_
rlabel metal1 14720 11050 14720 11050 0 _082_
rlabel metal1 13662 8466 13662 8466 0 _083_
rlabel metal1 17342 11730 17342 11730 0 _084_
rlabel metal2 17802 9928 17802 9928 0 _085_
rlabel metal1 17572 14926 17572 14926 0 _086_
rlabel metal1 17940 11730 17940 11730 0 _087_
rlabel metal2 17618 9180 17618 9180 0 _088_
rlabel metal1 16882 11118 16882 11118 0 _089_
rlabel metal1 15410 11152 15410 11152 0 _090_
rlabel metal1 12742 9384 12742 9384 0 _091_
rlabel metal2 13662 9197 13662 9197 0 _092_
rlabel metal1 13754 8976 13754 8976 0 _093_
rlabel metal1 13432 8058 13432 8058 0 _094_
rlabel metal1 16744 11866 16744 11866 0 _095_
rlabel metal1 16330 12410 16330 12410 0 _096_
rlabel metal1 12581 12206 12581 12206 0 _097_
rlabel metal1 13294 11764 13294 11764 0 _098_
rlabel metal1 13110 11594 13110 11594 0 _099_
rlabel metal1 13294 8602 13294 8602 0 _100_
rlabel metal1 17204 6766 17204 6766 0 _101_
rlabel metal1 16560 3434 16560 3434 0 _102_
rlabel metal1 16422 5542 16422 5542 0 _103_
rlabel metal1 15364 7378 15364 7378 0 _104_
rlabel metal2 15962 6324 15962 6324 0 _105_
rlabel metal1 14214 5882 14214 5882 0 _106_
rlabel metal1 17434 6732 17434 6732 0 _107_
rlabel metal1 17940 6970 17940 6970 0 _108_
rlabel metal1 14260 4794 14260 4794 0 _109_
rlabel metal1 17848 5882 17848 5882 0 _110_
rlabel metal2 18078 6936 18078 6936 0 _111_
rlabel metal1 17986 8466 17986 8466 0 _112_
rlabel metal1 17158 9146 17158 9146 0 _113_
rlabel metal1 17250 7310 17250 7310 0 _114_
rlabel metal2 17250 8058 17250 8058 0 _115_
rlabel metal1 12673 8602 12673 8602 0 _116_
rlabel metal1 17710 11050 17710 11050 0 _117_
rlabel metal1 15778 9588 15778 9588 0 _118_
rlabel metal1 16376 9554 16376 9554 0 _119_
rlabel metal1 13478 8908 13478 8908 0 _120_
rlabel metal1 10166 13804 10166 13804 0 _121_
rlabel via1 12466 9027 12466 9027 0 _122_
rlabel metal1 10534 13906 10534 13906 0 _123_
rlabel metal1 10994 9622 10994 9622 0 _124_
rlabel metal1 12006 8058 12006 8058 0 _125_
rlabel metal1 10672 9146 10672 9146 0 _126_
rlabel metal1 11454 8942 11454 8942 0 _127_
rlabel metal2 9430 8092 9430 8092 0 _128_
rlabel metal1 9338 11866 9338 11866 0 _129_
rlabel metal1 9844 12886 9844 12886 0 _130_
rlabel metal2 10626 13124 10626 13124 0 _131_
rlabel metal2 13846 7854 13846 7854 0 _132_
rlabel metal1 4968 7854 4968 7854 0 _133_
rlabel metal1 6900 8602 6900 8602 0 _134_
rlabel metal1 7590 7854 7590 7854 0 _135_
rlabel metal2 8510 7582 8510 7582 0 _136_
rlabel metal1 7958 6358 7958 6358 0 _137_
rlabel metal2 10350 15300 10350 15300 0 _138_
rlabel metal1 5796 7854 5796 7854 0 _139_
rlabel metal2 6394 8704 6394 8704 0 _140_
rlabel metal1 6486 8058 6486 8058 0 _141_
rlabel metal2 6578 8738 6578 8738 0 _142_
rlabel metal1 6992 5202 6992 5202 0 _143_
rlabel metal1 8648 6630 8648 6630 0 _144_
rlabel metal1 7176 2346 7176 2346 0 _145_
rlabel metal2 9430 6460 9430 6460 0 _146_
rlabel metal2 8510 5882 8510 5882 0 _147_
rlabel metal1 8188 8466 8188 8466 0 _148_
rlabel metal1 11086 12138 11086 12138 0 _149_
rlabel metal2 10442 11968 10442 11968 0 _150_
rlabel metal1 11454 12614 11454 12614 0 _151_
rlabel metal1 15318 7310 15318 7310 0 _152_
rlabel metal2 17066 7718 17066 7718 0 _153_
rlabel metal1 18216 7854 18216 7854 0 _154_
rlabel metal1 16790 8942 16790 8942 0 _155_
rlabel metal1 17434 6426 17434 6426 0 _156_
rlabel metal1 17480 2550 17480 2550 0 _157_
rlabel viali 17884 4590 17884 4590 0 _158_
rlabel metal2 18170 6256 18170 6256 0 _159_
rlabel metal2 17526 8534 17526 8534 0 _160_
rlabel metal1 16146 9146 16146 9146 0 _161_
rlabel metal1 12190 9010 12190 9010 0 _162_
rlabel metal1 12604 10778 12604 10778 0 _163_
rlabel metal1 12374 8976 12374 8976 0 _164_
rlabel metal1 12926 8942 12926 8942 0 _165_
rlabel metal2 12558 9724 12558 9724 0 _166_
rlabel metal2 8602 7004 8602 7004 0 _167_
rlabel metal2 7038 3468 7038 3468 0 _168_
rlabel metal1 2484 10030 2484 10030 0 _169_
rlabel metal2 6210 4522 6210 4522 0 _170_
rlabel metal1 5934 2550 5934 2550 0 _171_
rlabel metal1 8050 5678 8050 5678 0 _172_
rlabel metal1 5290 2448 5290 2448 0 _173_
rlabel metal2 6762 5542 6762 5542 0 _174_
rlabel metal1 7820 2414 7820 2414 0 _175_
rlabel metal1 7958 4114 7958 4114 0 _176_
rlabel metal1 15732 2414 15732 2414 0 _177_
rlabel metal1 2438 13328 2438 13328 0 _178_
rlabel metal1 3128 4590 3128 4590 0 _179_
rlabel metal2 2254 6460 2254 6460 0 _180_
rlabel metal1 2438 6800 2438 6800 0 _181_
rlabel metal1 9568 8942 9568 8942 0 _182_
rlabel metal2 9706 7684 9706 7684 0 _183_
rlabel metal1 6946 7208 6946 7208 0 _184_
rlabel metal1 7590 10166 7590 10166 0 _185_
rlabel metal1 8832 8942 8832 8942 0 _186_
rlabel metal1 7406 13294 7406 13294 0 _187_
rlabel metal1 7590 10030 7590 10030 0 _188_
rlabel metal2 7498 13702 7498 13702 0 _189_
rlabel metal2 3266 10880 3266 10880 0 _190_
rlabel metal2 4278 14433 4278 14433 0 _191_
rlabel metal1 7452 11322 7452 11322 0 _192_
rlabel metal2 7958 12036 7958 12036 0 _193_
rlabel metal2 6394 11662 6394 11662 0 _194_
rlabel metal1 6118 12410 6118 12410 0 _195_
rlabel metal1 6164 11118 6164 11118 0 _196_
rlabel metal1 9430 13838 9430 13838 0 _197_
rlabel metal1 8832 12410 8832 12410 0 _198_
rlabel metal1 10166 13498 10166 13498 0 _199_
rlabel metal1 9798 14042 9798 14042 0 _200_
rlabel metal1 9246 15028 9246 15028 0 _201_
rlabel metal2 15410 13634 15410 13634 0 _202_
rlabel metal1 11914 14348 11914 14348 0 _203_
rlabel metal2 12282 16014 12282 16014 0 _204_
rlabel metal1 12558 15470 12558 15470 0 _205_
rlabel metal1 13202 16150 13202 16150 0 _206_
rlabel metal1 12098 16048 12098 16048 0 _207_
rlabel metal2 14674 14858 14674 14858 0 _208_
rlabel metal2 14858 14076 14858 14076 0 _209_
rlabel metal1 14720 12954 14720 12954 0 _210_
rlabel metal1 15916 12614 15916 12614 0 _211_
rlabel metal1 14950 11730 14950 11730 0 _212_
rlabel metal1 15640 10234 15640 10234 0 _213_
rlabel metal1 14950 10234 14950 10234 0 _214_
rlabel metal2 15318 9248 15318 9248 0 _215_
rlabel metal2 14766 9350 14766 9350 0 _216_
rlabel metal2 11178 7820 11178 7820 0 _217_
rlabel metal1 13754 6834 13754 6834 0 _218_
rlabel metal2 16054 7650 16054 7650 0 _219_
rlabel metal2 16054 4964 16054 4964 0 _220_
rlabel metal1 10120 4794 10120 4794 0 _221_
rlabel via1 9974 4522 9974 4522 0 _222_
rlabel metal1 9522 3502 9522 3502 0 _223_
rlabel metal2 10810 5168 10810 5168 0 _224_
rlabel metal1 11178 5338 11178 5338 0 _225_
rlabel metal1 11224 4590 11224 4590 0 _226_
rlabel metal1 12282 6426 12282 6426 0 _227_
rlabel metal1 12006 5882 12006 5882 0 _228_
rlabel metal2 15962 4862 15962 4862 0 _229_
rlabel metal1 17250 4182 17250 4182 0 _230_
rlabel metal1 16606 3978 16606 3978 0 _231_
rlabel metal2 18170 3332 18170 3332 0 _232_
rlabel metal2 17434 3162 17434 3162 0 _233_
rlabel metal1 16606 2414 16606 2414 0 _234_
rlabel metal1 4692 10642 4692 10642 0 _235_
rlabel metal1 2944 10030 2944 10030 0 _236_
rlabel metal1 2944 15334 2944 15334 0 _237_
rlabel metal2 2806 16966 2806 16966 0 _238_
rlabel metal2 6578 16694 6578 16694 0 _239_
rlabel metal2 6026 16524 6026 16524 0 _240_
rlabel metal2 12650 16966 12650 16966 0 _241_
rlabel metal2 10534 16524 10534 16524 0 _242_
rlabel metal1 8786 16218 8786 16218 0 _243_
rlabel metal1 7360 14994 7360 14994 0 _244_
rlabel metal1 5845 14042 5845 14042 0 _245_
rlabel metal1 3634 14382 3634 14382 0 _246_
rlabel metal2 2346 13702 2346 13702 0 _247_
rlabel metal2 2530 12614 2530 12614 0 _248_
rlabel metal2 4002 11764 4002 11764 0 _249_
rlabel metal2 2898 11764 2898 11764 0 _250_
rlabel metal1 4876 4114 4876 4114 0 _251_
rlabel metal1 6118 15878 6118 15878 0 clk
rlabel metal1 9660 12818 9660 12818 0 clknet_0_clk
rlabel metal2 4646 7412 4646 7412 0 clknet_2_0__leaf_clk
rlabel metal1 14168 2482 14168 2482 0 clknet_2_1__leaf_clk
rlabel metal1 5014 12682 5014 12682 0 clknet_2_2__leaf_clk
rlabel metal1 14076 13294 14076 13294 0 clknet_2_3__leaf_clk
rlabel metal2 6946 5746 6946 5746 0 dice.bcd\[0\]
rlabel metal1 8878 4794 8878 4794 0 dice.bcd\[1\]
rlabel metal2 7682 6460 7682 6460 0 dice.bcd\[2\]
rlabel metal1 12466 6732 12466 6732 0 dice.clkdiv\[0\]
rlabel metal1 9476 10710 9476 10710 0 dice.clkdiv\[1\]
rlabel metal2 12834 10812 12834 10812 0 dice.clkdiv\[2\]
rlabel metal1 7820 13294 7820 13294 0 dice.clkdiv\[3\]
rlabel metal1 11040 12818 11040 12818 0 dice.clkdiv\[4\]
rlabel metal1 9522 11662 9522 11662 0 dice.clkdiv\[5\]
rlabel metal1 10442 13294 10442 13294 0 dice.clkdiv\[6\]
rlabel metal2 10902 15164 10902 15164 0 dice.clkdiv\[7\]
rlabel metal2 17066 13532 17066 13532 0 dice.counter\[0\]
rlabel metal1 14628 4658 14628 4658 0 dice.counter\[10\]
rlabel metal2 13294 4828 13294 4828 0 dice.counter\[11\]
rlabel metal2 17066 5814 17066 5814 0 dice.counter\[12\]
rlabel metal1 17434 4250 17434 4250 0 dice.counter\[13\]
rlabel metal1 15824 2618 15824 2618 0 dice.counter\[14\]
rlabel metal1 17296 2414 17296 2414 0 dice.counter\[15\]
rlabel metal2 17158 15470 17158 15470 0 dice.counter\[1\]
rlabel metal1 15778 14994 15778 14994 0 dice.counter\[2\]
rlabel metal1 17066 13226 17066 13226 0 dice.counter\[3\]
rlabel via1 16422 11101 16422 11101 0 dice.counter\[4\]
rlabel metal1 17204 10030 17204 10030 0 dice.counter\[5\]
rlabel metal2 17342 9520 17342 9520 0 dice.counter\[6\]
rlabel via1 15882 7310 15882 7310 0 dice.counter\[7\]
rlabel metal2 17434 5304 17434 5304 0 dice.counter\[8\]
rlabel metal2 13110 5100 13110 5100 0 dice.counter\[9\]
rlabel metal2 2622 13532 2622 13532 0 dice.lfsr\[0\]
rlabel metal2 6854 15164 6854 15164 0 dice.lfsr\[10\]
rlabel metal1 5842 14518 5842 14518 0 dice.lfsr\[11\]
rlabel metal1 4278 15130 4278 15130 0 dice.lfsr\[12\]
rlabel metal2 2714 13600 2714 13600 0 dice.lfsr\[13\]
rlabel metal1 2576 12206 2576 12206 0 dice.lfsr\[14\]
rlabel metal2 4186 11322 4186 11322 0 dice.lfsr\[15\]
rlabel metal1 2622 7412 2622 7412 0 dice.lfsr\[1\]
rlabel metal1 2300 9350 2300 9350 0 dice.lfsr\[2\]
rlabel metal1 3174 15470 3174 15470 0 dice.lfsr\[3\]
rlabel metal1 3588 16558 3588 16558 0 dice.lfsr\[4\]
rlabel metal2 6946 16286 6946 16286 0 dice.lfsr\[5\]
rlabel metal2 7222 16966 7222 16966 0 dice.lfsr\[6\]
rlabel metal1 12282 16456 12282 16456 0 dice.lfsr\[7\]
rlabel metal1 10166 16218 10166 16218 0 dice.lfsr\[8\]
rlabel metal1 8280 15334 8280 15334 0 dice.lfsr\[9\]
rlabel metal2 4002 5814 4002 5814 0 dice.r_counter\[0\]
rlabel metal1 2806 7344 2806 7344 0 dice.r_counter\[1\]
rlabel metal1 1794 7786 1794 7786 0 dice.r_counter\[2\]
rlabel metal1 16468 17306 16468 17306 0 io_in
rlabel metal2 1242 1520 1242 1520 0 io_out[0]
rlabel metal2 3726 1520 3726 1520 0 io_out[1]
rlabel metal2 6210 1520 6210 1520 0 io_out[2]
rlabel metal2 8694 1520 8694 1520 0 io_out[3]
rlabel metal1 11316 3366 11316 3366 0 io_out[4]
rlabel metal1 14076 3366 14076 3366 0 io_out[5]
rlabel metal1 15916 3366 15916 3366 0 io_out[6]
rlabel metal1 18446 3366 18446 3366 0 io_out[7]
rlabel metal2 16974 16048 16974 16048 0 net1
rlabel metal1 13708 2618 13708 2618 0 net10
rlabel metal2 9890 16762 9890 16762 0 net2
rlabel metal1 2944 2414 2944 2414 0 net3
rlabel metal1 4232 2822 4232 2822 0 net4
rlabel metal2 6026 2618 6026 2618 0 net5
rlabel metal1 8648 2414 8648 2414 0 net6
rlabel metal1 10902 2618 10902 2618 0 net7
rlabel metal1 13294 3162 13294 3162 0 net8
rlabel metal1 15502 3468 15502 3468 0 net9
rlabel metal1 10718 17170 10718 17170 0 rst
<< properties >>
string FIXED_BBOX 0 0 20000 20000
<< end >>
