VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tholin_avalonsemi_tbb1143
  CLASS BLOCK ;
  FOREIGN tholin_avalonsemi_tbb1143 ;
  ORIGIN 0.000 0.000 ;
  SIZE 160.000 BY 160.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.670 156.000 10.950 160.000 ;
    END
  END clk
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.230 156.000 50.510 160.000 ;
    END
  END io_in[0]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.010 156.000 70.290 160.000 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 156.000 90.070 160.000 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 156.000 109.850 160.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.350 156.000 129.630 160.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.130 156.000 149.410 160.000 ;
    END
  END io_in[5]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 10.240 160.000 10.840 ;
    END
  END io_out[0]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 29.960 160.000 30.560 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 49.680 160.000 50.280 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 69.400 160.000 70.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 89.120 160.000 89.720 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 108.840 160.000 109.440 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 128.560 160.000 129.160 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 148.280 160.000 148.880 ;
    END
  END io_out[7]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 156.000 30.730 160.000 ;
    END
  END rst
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 23.290 10.640 24.890 147.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 60.430 10.640 62.030 147.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 97.570 10.640 99.170 147.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 134.710 10.640 136.310 147.120 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 41.860 10.640 43.460 147.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 79.000 10.640 80.600 147.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 116.140 10.640 117.740 147.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 153.280 10.640 154.880 147.120 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 142.745 154.290 145.575 ;
        RECT 5.330 137.305 154.290 140.135 ;
        RECT 5.330 131.865 154.290 134.695 ;
        RECT 5.330 126.425 154.290 129.255 ;
        RECT 5.330 120.985 154.290 123.815 ;
        RECT 5.330 115.545 154.290 118.375 ;
        RECT 5.330 110.105 154.290 112.935 ;
        RECT 5.330 104.665 154.290 107.495 ;
        RECT 5.330 99.225 154.290 102.055 ;
        RECT 5.330 93.785 154.290 96.615 ;
        RECT 5.330 88.345 154.290 91.175 ;
        RECT 5.330 82.905 154.290 85.735 ;
        RECT 5.330 77.465 154.290 80.295 ;
        RECT 5.330 72.025 154.290 74.855 ;
        RECT 5.330 66.585 154.290 69.415 ;
        RECT 5.330 61.145 154.290 63.975 ;
        RECT 5.330 55.705 154.290 58.535 ;
        RECT 5.330 50.265 154.290 53.095 ;
        RECT 5.330 44.825 154.290 47.655 ;
        RECT 5.330 39.385 154.290 42.215 ;
        RECT 5.330 33.945 154.290 36.775 ;
        RECT 5.330 28.505 154.290 31.335 ;
        RECT 5.330 23.065 154.290 25.895 ;
        RECT 5.330 17.625 154.290 20.455 ;
        RECT 5.330 12.185 154.290 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 154.100 146.965 ;
      LAYER met1 ;
        RECT 5.520 10.640 155.410 147.120 ;
      LAYER met2 ;
        RECT 9.300 155.720 10.390 156.810 ;
        RECT 11.230 155.720 30.170 156.810 ;
        RECT 31.010 155.720 49.950 156.810 ;
        RECT 50.790 155.720 69.730 156.810 ;
        RECT 70.570 155.720 89.510 156.810 ;
        RECT 90.350 155.720 109.290 156.810 ;
        RECT 110.130 155.720 129.070 156.810 ;
        RECT 129.910 155.720 148.850 156.810 ;
        RECT 149.690 155.720 155.390 156.810 ;
        RECT 9.300 9.675 155.390 155.720 ;
      LAYER met3 ;
        RECT 23.300 147.880 155.600 148.745 ;
        RECT 23.300 129.560 156.090 147.880 ;
        RECT 23.300 128.160 155.600 129.560 ;
        RECT 23.300 109.840 156.090 128.160 ;
        RECT 23.300 108.440 155.600 109.840 ;
        RECT 23.300 90.120 156.090 108.440 ;
        RECT 23.300 88.720 155.600 90.120 ;
        RECT 23.300 70.400 156.090 88.720 ;
        RECT 23.300 69.000 155.600 70.400 ;
        RECT 23.300 50.680 156.090 69.000 ;
        RECT 23.300 49.280 155.600 50.680 ;
        RECT 23.300 30.960 156.090 49.280 ;
        RECT 23.300 29.560 155.600 30.960 ;
        RECT 23.300 11.240 156.090 29.560 ;
        RECT 23.300 9.840 155.600 11.240 ;
        RECT 23.300 9.695 156.090 9.840 ;
  END
END tholin_avalonsemi_tbb1143
END LIBRARY

