* NGSPICE file created from wrapped_as2650.ext - technology: sky130B

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_4 abstract view
.subckt sky130_fd_sc_hd__nor4b_4 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_4 abstract view
.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_4 abstract view
.subckt sky130_fd_sc_hd__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_4 abstract view
.subckt sky130_fd_sc_hd__o21ba_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

.subckt wrapped_as2650 clk io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_oeb io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[2] io_out[3] io_out[4]
+ io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] rst vccd1 vssd1
X_3155_ _3869_/B _5165_/B vssd1 vssd1 vccd1 vccd1 _3744_/B sky130_fd_sc_hd__nand2_1
XFILLER_39_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5417__B1 _5507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3086_ _5179_/A _3092_/B _5162_/B _4046_/A vssd1 vssd1 vccd1 vccd1 _3107_/B sky130_fd_sc_hd__or4_4
XANTENNA__4654__B _5203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5766__A _5767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4670__A _4672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3988_ _3021_/Y _3197_/B _5428_/A vssd1 vssd1 vccd1 vccd1 _3988_/X sky130_fd_sc_hd__mux2_1
X_5727_ _3974_/C _3998_/C _5726_/Y _3615_/B _3958_/Y vssd1 vssd1 vccd1 vccd1 _5728_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_136_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5658_ _5710_/S _3713_/X _3950_/C vssd1 vssd1 vccd1 vccd1 _5658_/X sky130_fd_sc_hd__o21a_1
XFILLER_136_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4609_ _5241_/A _3966_/B _4608_/X vssd1 vssd1 vccd1 vccd1 _5876_/B sky130_fd_sc_hd__a21oi_2
X_5589_ _5512_/A _5598_/B _5579_/B _3122_/A vssd1 vssd1 vccd1 vccd1 _5589_/X sky130_fd_sc_hd__a31o_1
XFILLER_117_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4459__A1 _4891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5006__A _5547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout75_A _5943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4616__D1 _5048_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3895__S _4819_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4919__C1 _3116_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4580__A _5239_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5187__A2 _5244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3196__A _3941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5615__S _5703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3370__A1 _3960_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3135__S _3135_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4870__A1 _4872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4870__B2 _5463_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4960_ _6193_/Q _4647_/B _4648_/Y _6004_/Q _4826_/Y vssd1 vssd1 vccd1 vccd1 _4960_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_64_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3911_ _3913_/A _5766_/C vssd1 vssd1 vccd1 vccd1 _4438_/S sky130_fd_sc_hd__or2_4
XFILLER_44_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4891_ _4891_/A _4979_/B vssd1 vssd1 vccd1 vccd1 _4892_/B sky130_fd_sc_hd__nor2_2
XFILLER_32_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3842_ _3855_/S _3842_/B vssd1 vssd1 vccd1 vccd1 _3842_/Y sky130_fd_sc_hd__nor2_1
X_3773_ _6034_/Q _3771_/X _3770_/X _3764_/Y vssd1 vssd1 vccd1 vccd1 _6034_/D sky130_fd_sc_hd__a211o_1
XFILLER_9_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5512_ _5512_/A _5512_/B vssd1 vssd1 vccd1 vccd1 _5512_/Y sky130_fd_sc_hd__nor2_1
XFILLER_118_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5443_ _5943_/C _5421_/Y _5442_/X _5513_/A vssd1 vssd1 vccd1 vccd1 _5443_/X sky130_fd_sc_hd__o211a_1
XANTENNA__5335__C1 _5058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5350__A2 _3243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5374_ _5387_/B _5385_/C vssd1 vssd1 vccd1 vccd1 _5374_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__4649__B _5509_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4325_ _4325_/A _4325_/B vssd1 vssd1 vccd1 vccd1 _4328_/A sky130_fd_sc_hd__xnor2_2
XFILLER_113_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout105 _4022_/D vssd1 vssd1 vccd1 vccd1 _3975_/C sky130_fd_sc_hd__clkbuf_8
Xfanout116 _5848_/A0 vssd1 vssd1 vccd1 vccd1 _3410_/B sky130_fd_sc_hd__buf_4
XFILLER_99_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout127 _5903_/A vssd1 vssd1 vccd1 vccd1 _5707_/A sky130_fd_sc_hd__buf_4
XFILLER_101_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout138 _5503_/A vssd1 vssd1 vccd1 vccd1 _5934_/A sky130_fd_sc_hd__buf_6
Xfanout149 _5476_/A vssd1 vssd1 vccd1 vccd1 _5330_/B sky130_fd_sc_hd__buf_12
X_4256_ _6097_/Q _3721_/X _4259_/S vssd1 vssd1 vccd1 vccd1 _6097_/D sky130_fd_sc_hd__mux2_1
XANTENNA__5102__A2 _3869_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3207_ _5054_/A _5840_/B vssd1 vssd1 vccd1 vccd1 _4886_/B sky130_fd_sc_hd__or2_4
XFILLER_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4665__A _5264_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4187_ _4183_/Y _4184_/X _4149_/Y _4151_/Y vssd1 vssd1 vccd1 vccd1 _4187_/X sky130_fd_sc_hd__o211a_2
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3138_ _3766_/A _3257_/B vssd1 vssd1 vccd1 vccd1 _3227_/A sky130_fd_sc_hd__nor2_1
XFILLER_103_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3069_ _3107_/A _3126_/A vssd1 vssd1 vccd1 vccd1 _3069_/Y sky130_fd_sc_hd__nor2_8
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4613__A1 _4577_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5943__B _5943_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3744__A _5124_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5877__B1 _3164_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3888__C1 _5138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3352__A1 _4010_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_31_clk_A clkbuf_3_5__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3104__A1 _5731_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3104__B2 _5075_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4294__B _4294_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_46_clk_A _6230_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3407__A2 _4697_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4907__A2 _4883_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3591__A1 _4410_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3591__B2 _3590_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5868__A0 _5136_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4110_ _4110_/A _4110_/B vssd1 vssd1 vccd1 vccd1 _4117_/A sky130_fd_sc_hd__xor2_2
XFILLER_110_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5090_ _5090_/A _5090_/B vssd1 vssd1 vccd1 vccd1 _5090_/Y sky130_fd_sc_hd__nand2_1
XFILLER_68_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4041_ _6062_/Q _3721_/X _4044_/S vssd1 vssd1 vccd1 vccd1 _6062_/D sky130_fd_sc_hd__mux2_1
XFILLER_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4843__A1 _4842_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5992_ _6106_/Q vssd1 vssd1 vccd1 vccd1 _6106_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_24_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4943_ _4943_/A _4943_/B vssd1 vssd1 vccd1 vccd1 _5509_/B sky130_fd_sc_hd__nor2_1
XANTENNA__3829__A _5888_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4874_ _6190_/Q _5046_/B _4873_/Y _5047_/C1 vssd1 vssd1 vccd1 vccd1 _6190_/D sky130_fd_sc_hd__o211a_1
XANTENNA__5556__C1 _5556_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3825_ _3513_/B _3746_/A _3824_/X _3849_/B vssd1 vssd1 vccd1 vccd1 _3825_/X sky130_fd_sc_hd__a211o_1
XANTENNA__5020__B2 _5069_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3756_ _5226_/A _3845_/B _3737_/Y _3755_/Y vssd1 vssd1 vccd1 vccd1 _3756_/X sky130_fd_sc_hd__a211o_1
XFILLER_119_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3687_ _5503_/A _5943_/B vssd1 vssd1 vccd1 vccd1 _4462_/B sky130_fd_sc_hd__nand2_4
XFILLER_106_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5426_ _5428_/A _5428_/B vssd1 vssd1 vccd1 vccd1 _5452_/A sky130_fd_sc_hd__and2_1
XANTENNA__3334__A1 _3599_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5357_ _5333_/A _5556_/A2 _5354_/Y _5356_/Y _5556_/C1 vssd1 vssd1 vccd1 vccd1 _6222_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_102_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4308_ _4308_/A _4308_/B vssd1 vssd1 vccd1 vccd1 _4315_/A sky130_fd_sc_hd__xnor2_4
XFILLER_99_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5288_ _5595_/A _5257_/Y _5250_/X vssd1 vssd1 vccd1 vccd1 _5288_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_101_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5087__A1 _5227_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4239_ _4239_/A _4239_/B vssd1 vssd1 vccd1 vccd1 _4246_/S sky130_fd_sc_hd__nand2_8
XFILLER_101_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_556 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4842__B _4842_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3458__B _3458_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5562__A2 _5360_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4770__A0 _4767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3325__A1 _6011_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5078__A1 _5258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4825__A1 _6189_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4825__B2 _4819_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output19_A _6193_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4244__S _4246_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3610_ _3563_/S _4846_/B _3605_/X _3227_/X vssd1 vssd1 vccd1 vccd1 _3610_/X sky130_fd_sc_hd__a211o_2
XANTENNA__5553__A2 _5442_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4590_ _4604_/A _5635_/A _5634_/C _3978_/B vssd1 vssd1 vccd1 vccd1 _5104_/B sky130_fd_sc_hd__or4b_4
X_3541_ _3541_/A _3561_/B vssd1 vssd1 vccd1 vccd1 _3541_/X sky130_fd_sc_hd__or2_1
XFILLER_116_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6260_ _6260_/CLK _6260_/D vssd1 vssd1 vccd1 vccd1 _6260_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3472_ _3960_/B _3456_/X _3471_/X _3511_/A vssd1 vssd1 vccd1 vccd1 _3472_/X sky130_fd_sc_hd__o211a_1
X_5211_ _5960_/C1 _5209_/X _5210_/X _5956_/A vssd1 vssd1 vccd1 vccd1 _6218_/D sky130_fd_sc_hd__o211a_1
XFILLER_103_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6191_ _6217_/CLK _6191_/D vssd1 vssd1 vccd1 vccd1 _6191_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_124_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5142_ _5095_/A _5136_/X _5141_/Y _5075_/C _5131_/A vssd1 vssd1 vccd1 vccd1 _5142_/Y
+ sky130_fd_sc_hd__o32ai_4
XFILLER_123_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5608__A3 _5108_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5073_ _5244_/A _4638_/Y _4644_/B _5072_/X vssd1 vssd1 vccd1 vccd1 _5074_/A sky130_fd_sc_hd__a31o_1
XFILLER_84_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4024_ _3020_/Y _5207_/S _3883_/X _4023_/X vssd1 vssd1 vccd1 vccd1 _4025_/B sky130_fd_sc_hd__o31a_1
XFILLER_49_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4662__B _4663_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5975_ _5959_/A _5692_/B _3960_/C vssd1 vssd1 vccd1 vccd1 _5976_/D sky130_fd_sc_hd__o21ai_1
XFILLER_52_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4926_ _4926_/A vssd1 vssd1 vccd1 vccd1 _4926_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5529__C1 _5403_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4857_ _4872_/A _4979_/B vssd1 vssd1 vccd1 vccd1 _4925_/B sky130_fd_sc_hd__and2_4
XFILLER_138_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3808_ _4301_/A _3832_/A2 _3432_/Y _3765_/X _3772_/X vssd1 vssd1 vccd1 vccd1 _3808_/X
+ sky130_fd_sc_hd__o221a_1
X_4788_ _5367_/A _5172_/B _4787_/X _4646_/Y vssd1 vssd1 vccd1 vccd1 _4788_/X sky130_fd_sc_hd__o211a_1
XFILLER_119_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3739_ _5707_/A _4614_/A _3744_/C vssd1 vssd1 vccd1 vccd1 _3801_/B sky130_fd_sc_hd__or3_4
XFILLER_119_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4504__A0 _4672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3307__A1 _3575_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5409_ _5929_/B2 _5408_/X _5407_/X vssd1 vssd1 vccd1 vccd1 _5409_/X sky130_fd_sc_hd__a21o_2
XFILLER_106_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4837__B _4837_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3741__B _3741_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4853__A _6190_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4064__S _4066_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3188__B _5617_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5535__A2 _5251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4747__B _5344_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5859__A _5859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5471__B2 _5943_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5223__A1 _3156_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4026__A2 _5148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5760_ _3942_/B _5742_/Y _5758_/X _5759_/X vssd1 vssd1 vccd1 vccd1 _6247_/D sky130_fd_sc_hd__a22o_1
XFILLER_50_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4711_ _5034_/A _4750_/B _4710_/Y _4701_/X _3116_/B vssd1 vssd1 vccd1 vccd1 _4711_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__4982__B1 _4979_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5691_ _5730_/A _3937_/D _5690_/X _5732_/C1 vssd1 vssd1 vccd1 vccd1 _5691_/X sky130_fd_sc_hd__o211a_1
X_4642_ _4642_/A _4646_/A vssd1 vssd1 vccd1 vccd1 _4642_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__3537__A1 _4362_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3537__B2 _3536_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4573_ _5238_/B _5617_/C _5839_/A _4572_/X vssd1 vssd1 vccd1 vccd1 _4575_/S sky130_fd_sc_hd__o211a_2
XFILLER_116_612 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4003__A _5840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3524_ _3516_/Y _3517_/X _3521_/X _3523_/X vssd1 vssd1 vccd1 vccd1 _3524_/X sky130_fd_sc_hd__a211o_1
XFILLER_116_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6243_ _6256_/CLK _6243_/D vssd1 vssd1 vccd1 vccd1 _6243_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_131_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3455_ _3646_/B _3450_/D _3448_/Y _3541_/A _3454_/X vssd1 vssd1 vccd1 vccd1 _4734_/B
+ sky130_fd_sc_hd__o221a_4
X_6174_ _6179_/CLK _6174_/D vssd1 vssd1 vccd1 vccd1 _6174_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4657__B _4658_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3386_ _3801_/A _3500_/B vssd1 vssd1 vccd1 vccd1 _3448_/A sky130_fd_sc_hd__nand2_1
XFILLER_69_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5125_ _5124_/X _6206_/Q _5129_/S vssd1 vssd1 vccd1 vccd1 _6206_/D sky130_fd_sc_hd__mux2_1
XFILLER_85_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout192_A _3241_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5056_ _5090_/A _4745_/A _5638_/C _5055_/X _4581_/X vssd1 vssd1 vccd1 vccd1 _5059_/B
+ sky130_fd_sc_hd__o2111a_1
XANTENNA__3988__S _5428_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4007_ _6058_/Q _5561_/S _3032_/Y _6296_/Q _4004_/X vssd1 vssd1 vccd1 vccd1 _4009_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_25_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4017__A2 _3033_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5958_ _3112_/B _3975_/C _5131_/B _5960_/C1 vssd1 vssd1 vccd1 vccd1 _5976_/B sky130_fd_sc_hd__a211o_1
XFILLER_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4909_ _4945_/A _4945_/B vssd1 vssd1 vccd1 vccd1 _4910_/B sky130_fd_sc_hd__or2_1
X_5889_ _5889_/A _5889_/B vssd1 vssd1 vccd1 vccd1 _5889_/X sky130_fd_sc_hd__or2_1
XFILLER_138_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5060__A1_N _5065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4567__B _5075_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_724 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_74 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3199__A _5734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5205__A1 _5097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3767__A1 _5210_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3240_ _3240_/A _3241_/B vssd1 vssd1 vccd1 vccd1 _3240_/Y sky130_fd_sc_hd__nand2_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5141__B1 _5136_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3171_ _6200_/Q _6199_/Q vssd1 vssd1 vccd1 vccd1 _4842_/B sky130_fd_sc_hd__nor2_8
XFILLER_39_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5444__A1 _5058_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4652__C1 _5090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5812_ _3583_/X _5801_/B _5801_/Y _6270_/Q vssd1 vssd1 vccd1 vccd1 _5812_/X sky130_fd_sc_hd__a22o_1
XFILLER_90_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3758__A1 _3287_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5743_ _5767_/A _5743_/B _5743_/C vssd1 vssd1 vccd1 vccd1 _5791_/A sky130_fd_sc_hd__or3_4
XFILLER_31_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5674_ _5075_/A _3390_/Y _5203_/A _3410_/B _5728_/A vssd1 vssd1 vccd1 vccd1 _5675_/C
+ sky130_fd_sc_hd__a221o_1
X_4625_ _4625_/A _5093_/A vssd1 vssd1 vccd1 vccd1 _4625_/Y sky130_fd_sc_hd__nor2_1
XFILLER_135_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4556_ _6178_/Q _4562_/B vssd1 vssd1 vccd1 vccd1 _4556_/X sky130_fd_sc_hd__or2_1
XFILLER_116_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3507_ _3507_/A _3507_/B vssd1 vssd1 vccd1 vccd1 _3507_/Y sky130_fd_sc_hd__nand2_1
XFILLER_116_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4487_ _6136_/Q _4499_/B vssd1 vssd1 vccd1 vccd1 _4487_/X sky130_fd_sc_hd__or2_1
XFILLER_104_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6226_ _6254_/CLK _6226_/D vssd1 vssd1 vccd1 vccd1 _6226_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3438_ _6277_/Q _6113_/Q _3551_/S vssd1 vssd1 vccd1 vccd1 _5367_/B sky130_fd_sc_hd__mux2_8
XFILLER_103_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4387__B _4410_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3291__B _6009_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6157_ _6263_/CLK _6157_/D vssd1 vssd1 vccd1 vccd1 _6157_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3694__A0 _3942_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3369_ _3362_/X _3365_/Y _3367_/X _3368_/Y vssd1 vssd1 vccd1 vccd1 _3369_/X sky130_fd_sc_hd__a31o_1
XFILLER_85_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5108_ _5108_/A _5108_/B vssd1 vssd1 vccd1 vccd1 _5110_/A sky130_fd_sc_hd__nand2_2
XFILLER_111_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6088_ _6248_/CLK _6088_/D vssd1 vssd1 vccd1 vccd1 _6088_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5499__A _5504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5039_ _4981_/A _4988_/B _5015_/A _5031_/Y vssd1 vssd1 vccd1 vccd1 _5040_/B sky130_fd_sc_hd__o31a_1
XFILLER_73_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4850__B _4886_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3921__A1 _3730_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput20 _6194_/Q vssd1 vssd1 vccd1 vccd1 io_out[18] sky130_fd_sc_hd__buf_4
Xoutput31 _6284_/Q vssd1 vssd1 vccd1 vccd1 io_out[3] sky130_fd_sc_hd__buf_4
XFILLER_1_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5674__A1 _5075_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5674__B2 _3410_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5729__A2 _5649_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4937__B1 _5172_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4410_ _4426_/A _4410_/B _4426_/B _4410_/D vssd1 vssd1 vccd1 vccd1 _4411_/B sky130_fd_sc_hd__and4_1
X_5390_ _5392_/A _5392_/B vssd1 vssd1 vccd1 vccd1 _5391_/A sky130_fd_sc_hd__nand2_2
XFILLER_132_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4341_ _4426_/A _4309_/B _4342_/B _4410_/B vssd1 vssd1 vccd1 vccd1 _4341_/X sky130_fd_sc_hd__a22o_1
XFILLER_99_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4272_ _4272_/A _4272_/B vssd1 vssd1 vccd1 vccd1 _4274_/A sky130_fd_sc_hd__nor2_4
Xfanout309 _6010_/Q vssd1 vssd1 vccd1 vccd1 _5054_/A sky130_fd_sc_hd__buf_12
X_6011_ _6258_/CLK _6011_/D vssd1 vssd1 vccd1 vccd1 _6011_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__5665__A1 _4690_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3223_ _3706_/A _3747_/A vssd1 vssd1 vccd1 vccd1 _3476_/A sky130_fd_sc_hd__or2_4
XFILLER_39_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3154_ _3922_/S _5104_/A vssd1 vssd1 vccd1 vccd1 _3980_/B sky130_fd_sc_hd__nor2_4
XFILLER_55_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3428__B1 _5743_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3085_ _3085_/A _3123_/A _5058_/A vssd1 vssd1 vccd1 vccd1 _4612_/B sky130_fd_sc_hd__or3_2
XANTENNA__5968__A2 _5970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4951__A _6193_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout155_A _3069_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5766__B _5767_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4670__B _5263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3987_ _5712_/S _3987_/B _3986_/X vssd1 vssd1 vccd1 vccd1 _3987_/X sky130_fd_sc_hd__or3b_1
XFILLER_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout322_A input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5726_ _5726_/A _5726_/B vssd1 vssd1 vccd1 vccd1 _5726_/Y sky130_fd_sc_hd__nand2_1
XFILLER_109_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5657_ _5940_/A0 _4615_/A _3772_/B vssd1 vssd1 vccd1 vccd1 _5657_/X sky130_fd_sc_hd__a21o_1
X_4608_ _5976_/A _5241_/A _4608_/C vssd1 vssd1 vccd1 vccd1 _4608_/X sky130_fd_sc_hd__and3_1
X_5588_ _6232_/Q _5454_/A _5072_/B _5587_/X vssd1 vssd1 vccd1 vccd1 _5588_/X sky130_fd_sc_hd__a31o_1
XANTENNA__3903__A1 _3711_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4539_ _4539_/A _6172_/Q vssd1 vssd1 vccd1 vccd1 _6171_/D sky130_fd_sc_hd__and2_1
XFILLER_116_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4459__A2 _4438_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5006__B _5029_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6209_ _6209_/CLK _6209_/D vssd1 vssd1 vccd1 vccd1 _6209_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout68_A _5494_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6230__CLK _6230_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_6__f_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _6233_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5957__A _5976_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4580__B _5238_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5187__A3 _4648_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3196__B _4003_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_5_clk_A clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5692__A _6301_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3940__A _3940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3910_ _3913_/A _5766_/C vssd1 vssd1 vccd1 vccd1 _4458_/B sky130_fd_sc_hd__nor2_8
XANTENNA__4771__A _5119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4890_ _4891_/A _4979_/B vssd1 vssd1 vccd1 vccd1 _4924_/A sky130_fd_sc_hd__and2_2
X_3841_ _5898_/B _3840_/Y _3841_/S vssd1 vssd1 vccd1 vccd1 _3842_/B sky130_fd_sc_hd__mux2_4
XFILLER_60_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3387__A _3387_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4386__A1 _3807_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3772_ _3766_/Y _3772_/B _4539_/A _5191_/A vssd1 vssd1 vccd1 vccd1 _3772_/X sky130_fd_sc_hd__and4b_4
XFILLER_118_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5511_ _5312_/B _5513_/B _5507_/X _5510_/X vssd1 vssd1 vccd1 vccd1 _5511_/X sky130_fd_sc_hd__o211a_1
XFILLER_8_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5442_ _5442_/A _5442_/B vssd1 vssd1 vccd1 vccd1 _5442_/X sky130_fd_sc_hd__or2_1
XFILLER_133_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5373_ _3081_/Y _5371_/X _5372_/X vssd1 vssd1 vccd1 vccd1 _5373_/X sky130_fd_sc_hd__a21o_1
XFILLER_126_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4324_ _4325_/A _4325_/B vssd1 vssd1 vccd1 vccd1 _4355_/B sky130_fd_sc_hd__and2_1
XFILLER_113_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout106 _3557_/X vssd1 vssd1 vccd1 vccd1 _3615_/B sky130_fd_sc_hd__buf_6
Xfanout117 _3340_/X vssd1 vssd1 vccd1 vccd1 _5848_/A0 sky130_fd_sc_hd__buf_4
XANTENNA__5099__C1 _5192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout128 _5882_/S vssd1 vssd1 vccd1 vccd1 _5712_/S sky130_fd_sc_hd__buf_6
XFILLER_99_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4255_ _6096_/Q _3718_/X _4259_/S vssd1 vssd1 vccd1 vccd1 _6096_/D sky130_fd_sc_hd__mux2_1
Xfanout139 _5957_/B vssd1 vssd1 vccd1 vccd1 _5503_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_113_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4946__A _4946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5102__A3 _5634_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3206_ _5054_/A _5840_/B vssd1 vssd1 vccd1 vccd1 _4812_/S sky130_fd_sc_hd__nor2_8
XFILLER_101_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4186_ _4149_/Y _4151_/Y _4183_/Y _4184_/X vssd1 vssd1 vccd1 vccd1 _4193_/A sky130_fd_sc_hd__a211oi_4
XANTENNA__4665__B _4665_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3137_ _5800_/A _3869_/A vssd1 vssd1 vccd1 vccd1 _3137_/X sky130_fd_sc_hd__or2_1
XFILLER_27_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3068_ _3111_/B _6213_/Q _3092_/B vssd1 vssd1 vccd1 vccd1 _3126_/A sky130_fd_sc_hd__or3b_4
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5271__C1 _5507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5810__A1 _3529_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3297__A _6200_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5709_ _5409_/X _5708_/X _5734_/A vssd1 vssd1 vccd1 vccd1 _5709_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4129__A1 _4437_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5943__C _5943_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5877__A1 _6298_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5629__A1 _5710_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5629__B2 _5734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5687__A _5728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3812__A0 _3450_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3935__A _5241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5317__B1 _5349_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5868__A1 _5114_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3343__A2 _3410_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4766__A _5367_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3670__A _5054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4040_ _6061_/Q _3718_/X _4044_/S vssd1 vssd1 vccd1 vccd1 _6061_/D sky130_fd_sc_hd__mux2_1
XFILLER_80_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5991_ _6105_/Q vssd1 vssd1 vccd1 vccd1 _6105_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_80_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4942_ _6192_/Q _5046_/B _4941_/X _5047_/C1 vssd1 vssd1 vccd1 vccd1 _6192_/D sky130_fd_sc_hd__o211a_1
XFILLER_91_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4873_ _4871_/Y _4872_/Y _5046_/B vssd1 vssd1 vccd1 vccd1 _4873_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_20_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3824_ _3594_/B _3738_/X _3801_/B _3823_/X vssd1 vssd1 vccd1 vccd1 _3824_/X sky130_fd_sc_hd__o211a_1
X_3755_ _4620_/A _3845_/B vssd1 vssd1 vccd1 vccd1 _3755_/Y sky130_fd_sc_hd__nor2_1
XFILLER_134_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3686_ _5768_/A0 _6019_/Q _3902_/A vssd1 vssd1 vccd1 vccd1 _3686_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout118_A _3643_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3319__C1 _3145_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5425_ _5428_/A _5653_/A vssd1 vssd1 vccd1 vccd1 _5425_/Y sky130_fd_sc_hd__nand2_1
XFILLER_133_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5356_ _5058_/C _5355_/X _5556_/A2 vssd1 vssd1 vccd1 vccd1 _5356_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4307_ _4308_/A _4308_/B vssd1 vssd1 vccd1 vccd1 _4347_/A sky130_fd_sc_hd__and2_1
XFILLER_101_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4676__A _5034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5287_ _5276_/X _5286_/X _5058_/C vssd1 vssd1 vccd1 vccd1 _5287_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_59_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4238_ _5742_/C _4238_/B vssd1 vssd1 vccd1 vccd1 _4239_/B sky130_fd_sc_hd__or2_4
XFILLER_74_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5492__C1 _3122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_844 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4169_ _4169_/A _4169_/B _4169_/C vssd1 vssd1 vccd1 vccd1 _4210_/A sky130_fd_sc_hd__nand3_4
XFILLER_67_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4598__A1 _5148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3739__B _4614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3270__A1 _6012_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5970__A _5970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4586__A _4643_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3490__A _5818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5078__A2 _3059_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4825__A2 _4647_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3649__B _3649_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5538__B1 _3059_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3540_ _3594_/A _3540_/B vssd1 vssd1 vccd1 vccd1 _3561_/B sky130_fd_sc_hd__nor2_1
XFILLER_116_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4761__B2 _4638_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3471_ _3462_/X _3463_/Y _3470_/X vssd1 vssd1 vccd1 vccd1 _3471_/X sky130_fd_sc_hd__a21o_1
XFILLER_115_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5210_ _6218_/Q _5210_/B vssd1 vssd1 vccd1 vccd1 _5210_/X sky130_fd_sc_hd__or2_1
XANTENNA__4513__A1 _3010_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5710__A0 _3488_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6190_ _6288_/CLK _6190_/D vssd1 vssd1 vccd1 vccd1 _6190_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_130_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5141_ _5139_/X _5140_/Y _5136_/C vssd1 vssd1 vccd1 vccd1 _5141_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_124_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5072_ _5072_/A _5072_/B _5072_/C vssd1 vssd1 vccd1 vccd1 _5072_/X sky130_fd_sc_hd__and3_1
XANTENNA__5474__C1 _5948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4023_ _4023_/A _4023_/B _4022_/X vssd1 vssd1 vccd1 vccd1 _4023_/X sky130_fd_sc_hd__or3b_1
XFILLER_37_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4029__A0 _5128_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5974_ _5970_/A _5973_/X _5972_/X _5956_/A vssd1 vssd1 vccd1 vccd1 _6299_/D sky130_fd_sc_hd__o211a_1
XANTENNA__5120__A _6238_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4925_ _4925_/A _4925_/B _4925_/C _4900_/A vssd1 vssd1 vccd1 vccd1 _4926_/A sky130_fd_sc_hd__or4b_2
XFILLER_21_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4856_ _4705_/A _4864_/B _4753_/A vssd1 vssd1 vccd1 vccd1 _4856_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout235_A _4577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_30_clk_A clkbuf_3_5__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3807_ _3855_/S _3807_/B vssd1 vssd1 vccd1 vccd1 _3807_/Y sky130_fd_sc_hd__nor2_1
X_4787_ _5360_/S _4777_/Y _3671_/Y _6188_/Q vssd1 vssd1 vccd1 vccd1 _4787_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_119_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3738_ _3738_/A _3744_/C vssd1 vssd1 vccd1 vccd1 _3738_/X sky130_fd_sc_hd__or2_4
XFILLER_118_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3669_ _4046_/A _3669_/B vssd1 vssd1 vccd1 vccd1 _5158_/B sky130_fd_sc_hd__nor2_4
XFILLER_118_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_45_clk_A _6233_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5408_ _6255_/Q _6122_/Q _6024_/Q _6247_/Q _3241_/A _3241_/B vssd1 vssd1 vccd1 vccd1
+ _5408_/X sky130_fd_sc_hd__mux4_2
XFILLER_133_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5339_ _4644_/A _5329_/Y _5354_/B _5464_/A _5607_/B1 vssd1 vssd1 vccd1 vccd1 _5347_/B
+ sky130_fd_sc_hd__o221a_1
XANTENNA__3741__C _4886_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5768__A0 _5768_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_644 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5232__A2 _3243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4991__A1 _6194_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3188__C _3940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5940__A0 _5940_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3482__B2 _3236_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4710_ _4710_/A _4710_/B _4713_/A vssd1 vssd1 vccd1 vccd1 _4710_/Y sky130_fd_sc_hd__nand3_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4982__A1 _5504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5690_ _5718_/A _5690_/B vssd1 vssd1 vccd1 vccd1 _5690_/X sky130_fd_sc_hd__or2_1
X_4641_ _5218_/B _4646_/A vssd1 vssd1 vccd1 vccd1 _4644_/B sky130_fd_sc_hd__and2_4
XANTENNA__5931__A0 _5767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4572_ _4569_/X _4572_/B _4572_/C vssd1 vssd1 vccd1 vccd1 _4572_/X sky130_fd_sc_hd__and3b_1
XFILLER_116_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3523_ _3365_/B _3510_/Y _3522_/X _3312_/B _3145_/C vssd1 vssd1 vccd1 vccd1 _3523_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4003__B _4003_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6242_ _6293_/CLK _6242_/D vssd1 vssd1 vccd1 vccd1 _6242_/Q sky130_fd_sc_hd__dfxtp_1
X_3454_ _3611_/A _3599_/B _3454_/C vssd1 vssd1 vccd1 vccd1 _3454_/X sky130_fd_sc_hd__or3_1
XFILLER_115_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3842__B _3842_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6173_ _6177_/CLK _6173_/D vssd1 vssd1 vccd1 vccd1 _6173_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3385_ _3387_/A _3500_/B _3347_/Y _3599_/A vssd1 vssd1 vccd1 vccd1 _3389_/B sky130_fd_sc_hd__a22o_2
XANTENNA__3334__S _4010_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5115__A _6237_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5124_ _5859_/A _4819_/B _5124_/S vssd1 vssd1 vccd1 vccd1 _5124_/X sky130_fd_sc_hd__mux2_2
XFILLER_57_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5055_ _5072_/A _5870_/A _5075_/C _4596_/B vssd1 vssd1 vccd1 vccd1 _5055_/X sky130_fd_sc_hd__o31a_1
XFILLER_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_49_clk _6230_/CLK vssd1 vssd1 vccd1 vccd1 _6155_/CLK sky130_fd_sc_hd__clkbuf_16
X_4006_ _3766_/A _4767_/A _5714_/A _6291_/Q _4005_/X vssd1 vssd1 vccd1 vccd1 _4009_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_65_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3473__A1 _3422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5957_ _5976_/A _5957_/B vssd1 vssd1 vccd1 vccd1 _5961_/C sky130_fd_sc_hd__nor2_1
XFILLER_111_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4973__A1 _5731_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4908_ _5454_/A _4883_/B _4812_/S vssd1 vssd1 vccd1 vccd1 _4945_/B sky130_fd_sc_hd__o21ai_4
XFILLER_33_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5888_ _5888_/A _5888_/B vssd1 vssd1 vccd1 vccd1 _5888_/Y sky130_fd_sc_hd__nor2_1
XFILLER_138_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4839_ _5392_/A _5703_/B _4769_/A _4769_/B _4766_/X vssd1 vssd1 vccd1 vccd1 _4840_/B
+ sky130_fd_sc_hd__a221o_2
XANTENNA__3509__S _3922_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5922__B1 _5921_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5150__A1 _5191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4864__A _5330_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4661__A0 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3199__B _5710_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5610__C1 _5513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3767__A2 _3772_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3943__A _3943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3170_ _3170_/A _3170_/B vssd1 vssd1 vccd1 vccd1 _5617_/A sky130_fd_sc_hd__nand2_8
XFILLER_121_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3455__B2 _3541_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5811_ _5817_/A1 _4127_/Y _5810_/X vssd1 vssd1 vccd1 vccd1 _6269_/D sky130_fd_sc_hd__a21o_1
XFILLER_23_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5742_ _5742_/A _5742_/B _5742_/C vssd1 vssd1 vccd1 vccd1 _5742_/Y sky130_fd_sc_hd__nor3_4
XFILLER_50_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5673_ input3/X _3179_/X _5671_/X _5672_/X _3974_/C vssd1 vssd1 vccd1 vccd1 _5675_/B
+ sky130_fd_sc_hd__o221a_1
X_4624_ _5640_/B _5063_/A vssd1 vssd1 vccd1 vccd1 _5093_/A sky130_fd_sc_hd__nand2_8
XANTENNA__5380__A1 _5929_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4555_ _5856_/A _4564_/A2 _4553_/X _4554_/Y vssd1 vssd1 vccd1 vccd1 _6177_/D sky130_fd_sc_hd__a22o_1
XFILLER_116_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout100_A _5238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3506_ _3499_/X _4772_/B _3563_/S vssd1 vssd1 vccd1 vccd1 _3506_/X sky130_fd_sc_hd__mux2_1
XFILLER_116_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4486_ _5926_/A0 _4501_/A2 _4484_/X _4485_/Y vssd1 vssd1 vccd1 vccd1 _6135_/D sky130_fd_sc_hd__a22o_1
X_6225_ _6295_/CLK _6225_/D vssd1 vssd1 vccd1 vccd1 _6225_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3437_ _5114_/A _3549_/B _3398_/A _3436_/X vssd1 vssd1 vccd1 vccd1 _3437_/X sky130_fd_sc_hd__o211a_1
XFILLER_98_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5683__A2 _5848_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6156_ _6179_/CLK _6156_/D vssd1 vssd1 vccd1 vccd1 _6156_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3368_ _4003_/B _3358_/B _3881_/A vssd1 vssd1 vccd1 vccd1 _3368_/Y sky130_fd_sc_hd__a21oi_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5107_ _5903_/B _6201_/Q _5129_/S vssd1 vssd1 vccd1 vccd1 _6201_/D sky130_fd_sc_hd__mux2_1
X_6087_ _6260_/CLK _6087_/D vssd1 vssd1 vccd1 vccd1 _6087_/Q sky130_fd_sc_hd__dfxtp_1
X_3299_ _4010_/B _3646_/B vssd1 vssd1 vccd1 vccd1 _4665_/B sky130_fd_sc_hd__xnor2_4
XFILLER_111_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5038_ _5567_/A _4645_/B _5036_/Y _5037_/X vssd1 vssd1 vccd1 vccd1 _5038_/X sky130_fd_sc_hd__o22a_1
XFILLER_85_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5719__S _5731_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5371__A1 _3059_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput10 _3019_/Y vssd1 vssd1 vccd1 vccd1 io_oeb sky130_fd_sc_hd__buf_4
XFILLER_134_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput21 _6195_/Q vssd1 vssd1 vccd1 vccd1 io_out[19] sky130_fd_sc_hd__buf_4
Xoutput32 _6285_/Q vssd1 vssd1 vccd1 vccd1 io_out[4] sky130_fd_sc_hd__buf_4
XFILLER_107_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3134__A0 _4846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3702__S _3705_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3437__A1 _5114_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3938__A _5888_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4937__A1 _6192_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4937__B2 _4974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5362__A1 _4642_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5362__B2 _4646_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3673__A _5158_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4340_ _4340_/A _4340_/B vssd1 vssd1 vccd1 vccd1 _4345_/A sky130_fd_sc_hd__xnor2_1
XFILLER_125_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4271_ _5109_/A _3280_/X _4410_/D _4270_/A vssd1 vssd1 vccd1 vccd1 _4272_/B sky130_fd_sc_hd__a22oi_4
XFILLER_98_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3125__B1 _5239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3222_ _3706_/A _3747_/A vssd1 vssd1 vccd1 vccd1 _3583_/S sky130_fd_sc_hd__nor2_4
X_6010_ _6217_/CLK _6010_/D vssd1 vssd1 vccd1 vccd1 _6010_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_98_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3153_ _5634_/A _5143_/B vssd1 vssd1 vccd1 vccd1 _5104_/A sky130_fd_sc_hd__or2_4
XFILLER_95_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_419 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3084_ _5075_/B _3084_/B vssd1 vssd1 vccd1 vccd1 _3084_/X sky130_fd_sc_hd__or2_4
XFILLER_48_780 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4009__A _5976_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5539__S _5539_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5766__C _5766_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout148_A _5456_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3986_ _3986_/A _3986_/B _3986_/C _3599_/C vssd1 vssd1 vccd1 vccd1 _3986_/X sky130_fd_sc_hd__or4b_1
XFILLER_22_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3567__B _3567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5725_ _5882_/S _3649_/B _3597_/B _5903_/A _3179_/X vssd1 vssd1 vccd1 vccd1 _5726_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_31_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout315_A _3028_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5656_ _5656_/A _5735_/S vssd1 vssd1 vccd1 vccd1 _5656_/Y sky130_fd_sc_hd__nor2_1
XFILLER_108_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4607_ _4615_/B _5634_/C _5148_/A vssd1 vssd1 vccd1 vccd1 _5080_/A sky130_fd_sc_hd__o21a_1
XFILLER_117_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5587_ _5512_/A _5585_/X _5586_/X vssd1 vssd1 vccd1 vccd1 _5587_/X sky130_fd_sc_hd__a21o_1
XFILLER_116_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4538_ _3042_/Y _6171_/Q _4537_/Y vssd1 vssd1 vccd1 vccd1 _6170_/D sky130_fd_sc_hd__o21ai_1
XFILLER_117_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4469_ _3942_/D _4468_/X _4477_/S vssd1 vssd1 vccd1 vccd1 _6128_/D sky130_fd_sc_hd__mux2_1
XFILLER_89_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6208_ _6302_/CLK _6208_/D vssd1 vssd1 vccd1 vccd1 _6208_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_58_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6139_ _6179_/CLK _6139_/D vssd1 vssd1 vccd1 vccd1 _6139_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3522__S _3658_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3419__A1 _3621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5957__B _5957_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4919__B2 _4705_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5041__A0 _6196_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5592__A1 _6008_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3196__C _3312_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3658__A1 _3649_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4607__B1 _5148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5280__B1 _5742_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4771__B _4772_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5359__S _5539_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3840_ _4837_/B _3816_/B _3839_/X vssd1 vssd1 vccd1 vccd1 _3840_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_32_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3387__B _3500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3771_ _3855_/S _3771_/B vssd1 vssd1 vccd1 vccd1 _3771_/X sky130_fd_sc_hd__and2_4
XANTENNA__5883__A _5883_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5510_ _5510_/A _5537_/B _5227_/Y vssd1 vssd1 vccd1 vccd1 _5510_/X sky130_fd_sc_hd__or3b_2
XFILLER_12_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5441_ _5929_/B2 _5439_/X _5440_/X _5438_/X vssd1 vssd1 vccd1 vccd1 _5442_/B sky130_fd_sc_hd__a31o_4
XANTENNA__5335__A1 _4644_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5372_ _5464_/A _5358_/Y _5359_/X _4644_/A _5607_/B1 vssd1 vssd1 vccd1 vccd1 _5372_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__3441__S0 _4067_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4323_ _4323_/A _4323_/B vssd1 vssd1 vccd1 vccd1 _4325_/B sky130_fd_sc_hd__xnor2_2
XFILLER_114_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout107 _3557_/X vssd1 vssd1 vccd1 vccd1 _3594_/B sky130_fd_sc_hd__buf_4
XFILLER_87_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout118 _3643_/A vssd1 vssd1 vccd1 vccd1 _3986_/B sky130_fd_sc_hd__buf_8
XFILLER_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout129 _3111_/X vssd1 vssd1 vccd1 vccd1 _5069_/A sky130_fd_sc_hd__buf_6
X_4254_ _6095_/Q _3715_/X _4259_/S vssd1 vssd1 vccd1 vccd1 _6095_/D sky130_fd_sc_hd__mux2_1
XFILLER_87_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4438__S _4438_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3205_ _3205_/A _3257_/B _3744_/B _3706_/A vssd1 vssd1 vccd1 vccd1 _3210_/B sky130_fd_sc_hd__or4_4
XFILLER_101_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4185_ _4185_/A _4185_/B _4185_/C vssd1 vssd1 vccd1 vccd1 _4185_/Y sky130_fd_sc_hd__nand3_4
XFILLER_67_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3136_ _4067_/A _3869_/A vssd1 vssd1 vccd1 vccd1 _3136_/Y sky130_fd_sc_hd__nor2_4
XFILLER_83_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3067_ _3111_/B _3067_/B vssd1 vssd1 vccd1 vccd1 _5244_/B sky130_fd_sc_hd__nor2_2
XFILLER_103_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout265_A _4085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5269__S _5360_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3297__B _3297_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5574__A1 _3484_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3969_ _4596_/B _4605_/A _5617_/C vssd1 vssd1 vccd1 vccd1 _3969_/X sky130_fd_sc_hd__and3_1
XFILLER_50_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5708_ _6291_/Q _6042_/Q _5735_/S vssd1 vssd1 vccd1 vccd1 _5708_/X sky130_fd_sc_hd__mux2_1
XFILLER_109_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5639_ _5647_/B _5639_/B _5647_/D vssd1 vssd1 vccd1 vccd1 _5640_/D sky130_fd_sc_hd__and3_1
XFILLER_136_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3337__A0 _6013_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4202__A _4202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3888__A1 _5241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5629__A2 _3709_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout80_A _3103_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3104__A3 _4753_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4872__A _4872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4065__A1 _3727_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5565__A1 _3059_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4112__A _4197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3951__A _4022_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4766__B _4767_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3670__B _5330_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5990_ _6104_/Q vssd1 vssd1 vccd1 vccd1 _6104_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_18_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5253__B1 _4576_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4941_ _4931_/X _4940_/X _5046_/B vssd1 vssd1 vccd1 vccd1 _4941_/X sky130_fd_sc_hd__a21bo_1
XFILLER_64_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3803__A1 _4162_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4872_ _4872_/A _4872_/B vssd1 vssd1 vccd1 vccd1 _4872_/Y sky130_fd_sc_hd__nor2_1
XFILLER_33_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5556__A1 _5547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3823_ _5392_/A _3845_/B _3737_/Y _3822_/Y vssd1 vssd1 vccd1 vccd1 _3823_/X sky130_fd_sc_hd__a211o_1
XFILLER_32_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3754_ _6067_/Q _4294_/B vssd1 vssd1 vccd1 vccd1 _3855_/S sky130_fd_sc_hd__or2_4
XFILLER_118_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3685_ _5767_/A _3704_/B _5743_/C vssd1 vssd1 vccd1 vccd1 _3705_/A sky130_fd_sc_hd__or3_4
XANTENNA__3337__S _3551_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5424_ _5072_/B _5418_/X _5423_/X vssd1 vssd1 vccd1 vccd1 _5424_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_133_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5355_ _5943_/C _5354_/B _5353_/Y _5442_/A _5347_/X vssd1 vssd1 vccd1 vccd1 _5355_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_99_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4306_ _4301_/A _4389_/B _4274_/A _4272_/A vssd1 vssd1 vccd1 vccd1 _4308_/B sky130_fd_sc_hd__a31o_2
XFILLER_87_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4128__A1_N _3819_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5286_ _3949_/Y _5257_/Y _5283_/Y _5442_/A _5285_/X vssd1 vssd1 vccd1 vccd1 _5286_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_101_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4237_ _5742_/C _4238_/B vssd1 vssd1 vccd1 vccd1 _4237_/Y sky130_fd_sc_hd__nor2_1
XFILLER_102_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4168_ _4168_/A _4200_/A vssd1 vssd1 vccd1 vccd1 _4169_/C sky130_fd_sc_hd__nor2_2
XFILLER_56_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_4_clk_A clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3119_ _5050_/B _5050_/C vssd1 vssd1 vccd1 vccd1 _5647_/B sky130_fd_sc_hd__nand2_2
XFILLER_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4099_ _4099_/A _4099_/B vssd1 vssd1 vccd1 vccd1 _4099_/X sky130_fd_sc_hd__xor2_4
XANTENNA__5795__A1 _3721_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4598__A2 _5096_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3101__A _3101_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4586__B _4586_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3490__B _3555_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_555 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5483__A0 _4633_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5698__A _5714_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4806__S _4806_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4038__A1 _3711_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5786__A1 _5446_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5210__B _5210_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4107__A _4162_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3011__A _5333_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4746__C1 _5034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3470_ _3312_/Y _3466_/Y _3469_/X vssd1 vssd1 vccd1 vccd1 _3470_/X sky130_fd_sc_hd__a21o_1
XFILLER_131_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3681__A _5767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5140_ _5131_/B _4594_/B _3856_/X _5131_/A vssd1 vssd1 vccd1 vccd1 _5140_/Y sky130_fd_sc_hd__o211ai_2
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5071_ _5071_/A _5071_/B vssd1 vssd1 vccd1 vccd1 _6197_/D sky130_fd_sc_hd__and2_1
X_4022_ _6058_/Q _5207_/S _4022_/C _4022_/D vssd1 vssd1 vccd1 vccd1 _4022_/X sky130_fd_sc_hd__or4_1
XFILLER_96_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4029__A1 _3986_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5777__A1 _3011_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5973_ _5108_/A _5503_/A _3883_/X _5110_/B vssd1 vssd1 vccd1 vccd1 _5973_/X sky130_fd_sc_hd__o31a_1
XFILLER_92_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5120__B _5934_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4924_ _4924_/A _4924_/B vssd1 vssd1 vccd1 vccd1 _4924_/X sky130_fd_sc_hd__or2_1
XFILLER_33_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4855_ _4916_/C _4855_/B vssd1 vssd1 vccd1 vccd1 _4864_/B sky130_fd_sc_hd__or2_1
XFILLER_21_745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3856__A _4642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3806_ _5677_/B _3805_/Y _3841_/S vssd1 vssd1 vccd1 vccd1 _3807_/B sky130_fd_sc_hd__mux2_4
XANTENNA_fanout130_A _4654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout228_A _6293_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4786_ _3116_/B _4776_/X _4785_/Y vssd1 vssd1 vccd1 vccd1 _4786_/X sky130_fd_sc_hd__a21o_1
XFILLER_20_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3575__B _3575_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3737_ _3738_/A _3744_/C vssd1 vssd1 vccd1 vccd1 _3737_/Y sky130_fd_sc_hd__nor2_2
XFILLER_106_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3668_ _6018_/Q _3231_/Y _3667_/X vssd1 vssd1 vccd1 vccd1 _6018_/D sky130_fd_sc_hd__o21a_1
XFILLER_106_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5407_ _6130_/Q _5767_/B _5405_/X _3236_/Y _5406_/X vssd1 vssd1 vccd1 vccd1 _5407_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_134_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5701__A1 _3513_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3307__A3 _3267_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3599_ _3599_/A _3599_/B _3599_/C vssd1 vssd1 vccd1 vccd1 _3599_/X sky130_fd_sc_hd__and3_1
XFILLER_88_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5338_ _5338_/A _5338_/B vssd1 vssd1 vccd1 vccd1 _5338_/Y sky130_fd_sc_hd__nand2_1
XFILLER_87_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5269_ _4657_/A _6004_/Q _5360_/S vssd1 vssd1 vccd1 vccd1 _5269_/X sky130_fd_sc_hd__mux2_1
XFILLER_75_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5311__A _5605_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout43_A _5867_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4991__A2 _4990_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3766__A _3766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4259__A1 _3730_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5456__A0 _6010_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3006__A _4216_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout290 _6212_/Q vssd1 vssd1 vccd1 vccd1 _3092_/B sky130_fd_sc_hd__buf_4
XFILLER_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3440__S _3551_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3482__A2 _5743_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5221__A _5221_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5759__A1 _5387_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output24_A _6197_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4982__A2 _5488_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3676__A _3948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4640_ _4640_/A _4644_/A vssd1 vssd1 vccd1 vccd1 _4640_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__4719__C1 _4963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4571_ _3974_/C _3865_/Y _5203_/A vssd1 vssd1 vccd1 vccd1 _4572_/C sky130_fd_sc_hd__a21oi_1
X_3522_ _6205_/Q _3513_/B _3658_/S vssd1 vssd1 vccd1 vccd1 _3522_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4003__C _4003_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6241_ _6241_/CLK _6241_/D vssd1 vssd1 vccd1 vccd1 _6241_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3453_ _3644_/B _3450_/D _3448_/Y _3561_/A _3452_/X vssd1 vssd1 vccd1 vccd1 _4726_/B
+ sky130_fd_sc_hd__o221a_4
XFILLER_131_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4498__A1 _3942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4300__A _4301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6172_ _6264_/CLK _6172_/D vssd1 vssd1 vccd1 vccd1 _6172_/Q sky130_fd_sc_hd__dfxtp_1
X_3384_ _3592_/A _3384_/B vssd1 vssd1 vccd1 vccd1 _3384_/X sky130_fd_sc_hd__or2_1
XFILLER_97_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5115__B _5158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5123_ _5122_/Y _6205_/Q _5129_/S vssd1 vssd1 vccd1 vccd1 _6205_/D sky130_fd_sc_hd__mux2_1
XANTENNA__5447__B1 _5480_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5054_ _5054_/A _5203_/C vssd1 vssd1 vccd1 vccd1 _5638_/C sky130_fd_sc_hd__nand2_2
XFILLER_38_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4005_ _6299_/Q _5108_/A _4850_/A _6057_/Q vssd1 vssd1 vccd1 vccd1 _4005_/X sky130_fd_sc_hd__o22a_1
XFILLER_84_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout178_A _4167_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4970__A _6193_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5956_ _5956_/A _5956_/B _5956_/C vssd1 vssd1 vccd1 vccd1 _6296_/D sky130_fd_sc_hd__and3_1
XANTENNA_fanout345_A _4657_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4907_ _5454_/A _4883_/B _4847_/B _4849_/B _4845_/Y vssd1 vssd1 vccd1 vccd1 _4945_/A
+ sky130_fd_sc_hd__a221oi_4
XANTENNA__4973__A2 _4945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5887_ _5888_/A _5888_/B vssd1 vssd1 vccd1 vccd1 _5887_/Y sky130_fd_sc_hd__nand2_1
XFILLER_21_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4838_ _4836_/X _4838_/B vssd1 vssd1 vccd1 vccd1 _4841_/A sky130_fd_sc_hd__nand2b_2
XFILLER_138_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5922__A1 _5296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4769_ _4769_/A _4769_/B vssd1 vssd1 vccd1 vccd1 _4769_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_119_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5135__C1 _5227_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4489__A1 _3942_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5686__B1 _5203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3260__S _3551_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5976__A _5976_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5913__A1 _3880_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3943__B _5109_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4652__A1 _5255_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3455__A2 _3450_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4652__B2 _4644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5886__A _5900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5810_ _3529_/X _5801_/B _5801_/Y _6269_/Q vssd1 vssd1 vccd1 vccd1 _5810_/X sky130_fd_sc_hd__a22o_1
XFILLER_50_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_44_clk_A clkbuf_3_4__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5741_ _4216_/A _5649_/X _5740_/X _5956_/A vssd1 vssd1 vccd1 vccd1 _6241_/D sky130_fd_sc_hd__o211a_1
X_5672_ _3867_/B _3388_/B _3458_/B _3867_/A _3996_/B vssd1 vssd1 vccd1 vccd1 _5672_/X
+ sky130_fd_sc_hd__a221o_1
X_4623_ _4623_/A _5132_/B vssd1 vssd1 vccd1 vccd1 _5063_/A sky130_fd_sc_hd__nand2_4
XFILLER_129_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4554_ _3010_/Y _4562_/B _4564_/A2 vssd1 vssd1 vccd1 vccd1 _4554_/Y sky130_fd_sc_hd__a21oi_1
X_3505_ _3644_/B _3513_/B _3504_/Y _3608_/A _3503_/Y vssd1 vssd1 vccd1 vccd1 _4772_/B
+ sky130_fd_sc_hd__o221a_4
X_4485_ _5305_/A _4499_/B _4501_/A2 vssd1 vssd1 vccd1 vccd1 _4485_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_89_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6224_ _6227_/CLK _6224_/D vssd1 vssd1 vccd1 vccd1 _6224_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3436_ _3636_/A _4619_/B vssd1 vssd1 vccd1 vccd1 _3436_/X sky130_fd_sc_hd__or2_1
XFILLER_131_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6155_ _6155_/CLK _6155_/D vssd1 vssd1 vccd1 vccd1 _6155_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3367_ _3313_/Y _3364_/X _3366_/X _4003_/C vssd1 vssd1 vccd1 vccd1 _3367_/X sky130_fd_sc_hd__o22a_1
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout295_A _5960_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5106_ _4085_/A _5264_/A _5124_/S vssd1 vssd1 vccd1 vccd1 _5903_/B sky130_fd_sc_hd__mux2_1
XFILLER_111_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6086_ _6272_/CLK _6086_/D vssd1 vssd1 vccd1 vccd1 _6086_/Q sky130_fd_sc_hd__dfxtp_1
X_3298_ _3541_/A _3611_/A vssd1 vssd1 vccd1 vccd1 _3646_/B sky130_fd_sc_hd__nand2_8
XFILLER_100_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5037_ _6196_/Q _4647_/B _4648_/Y _6007_/Q _5227_/B vssd1 vssd1 vccd1 vccd1 _5037_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_85_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5939_ _3948_/A _3242_/X _5938_/X vssd1 vssd1 vccd1 vccd1 _5939_/X sky130_fd_sc_hd__a21o_1
XFILLER_40_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3382__A1 _5929_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput11 _6281_/Q vssd1 vssd1 vccd1 vccd1 io_out[0] sky130_fd_sc_hd__buf_4
XFILLER_103_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput22 _6282_/Q vssd1 vssd1 vccd1 vccd1 io_out[1] sky130_fd_sc_hd__buf_4
XANTENNA__5036__A _5509_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput33 _6286_/Q vssd1 vssd1 vccd1 vccd1 io_out[5] sky130_fd_sc_hd__buf_4
XFILLER_107_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3134__A1 _6009_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5470__S _5470_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4594__B _4594_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_1__f_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3673__B _4647_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4570__B1 _3971_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4270_ _4270_/A _5109_/A _4426_/B _4410_/D vssd1 vssd1 vccd1 vccd1 _4272_/A sky130_fd_sc_hd__and4_2
XFILLER_99_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3125__A1 _5075_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3221_ _5840_/A _5360_/S _5617_/B _3221_/D vssd1 vssd1 vccd1 vccd1 _3747_/A sky130_fd_sc_hd__or4_4
XFILLER_86_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3152_ _3958_/A _5143_/B vssd1 vssd1 vccd1 vccd1 _5165_/B sky130_fd_sc_hd__nor2_4
XFILLER_67_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3083_ _5075_/B _3084_/B vssd1 vssd1 vccd1 vccd1 _3083_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__3428__A2 _3589_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5586__C1 _3058_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3985_ _5626_/B _3607_/A _3594_/B _5707_/A vssd1 vssd1 vccd1 vccd1 _3993_/A sky130_fd_sc_hd__a211o_1
XFILLER_22_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5724_ _3772_/B _5722_/X _5723_/X vssd1 vssd1 vccd1 vccd1 _5726_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__4025__A _5148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5655_ _5454_/B _5654_/X _5653_/X _5732_/C1 vssd1 vssd1 vccd1 vccd1 _5655_/X sky130_fd_sc_hd__o211a_1
XFILLER_108_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4606_ _5976_/A _5959_/A _3877_/B _5048_/C vssd1 vssd1 vccd1 vccd1 _5878_/A sky130_fd_sc_hd__o31a_2
XANTENNA_fanout210_A _5733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5586_ _6008_/Q _5454_/B _4644_/B _5580_/Y _3058_/B vssd1 vssd1 vccd1 vccd1 _5586_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout308_A _6066_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4537_ _3042_/Y _6171_/Q _4540_/A vssd1 vssd1 vccd1 vccd1 _4537_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_132_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4468_ _5333_/A _6128_/Q _4476_/S vssd1 vssd1 vccd1 vccd1 _4468_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6207_ _6302_/CLK _6207_/D vssd1 vssd1 vccd1 vccd1 _6207_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3419_ _3621_/A _3414_/Y _3418_/X vssd1 vssd1 vccd1 vccd1 _3419_/Y sky130_fd_sc_hd__o21ai_1
X_4399_ _4399_/A _4399_/B vssd1 vssd1 vccd1 vccd1 _4401_/B sky130_fd_sc_hd__xor2_1
XANTENNA__3667__A2 _3666_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6138_ _6180_/CLK _6138_/D vssd1 vssd1 vccd1 vccd1 _6138_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6069_ _6209_/CLK _6069_/D vssd1 vssd1 vccd1 vccd1 _6069_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__4616__A1 _4604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5592__A2 _5360_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4833__A2_N _4872_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3949__A _4638_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3387__C _3500_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3770_ _4197_/B _5943_/A _3250_/X _3765_/X _3769_/X vssd1 vssd1 vccd1 vccd1 _3770_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_9_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3684__A _3734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5440_ _6123_/Q _3901_/B _3704_/B _6025_/Q vssd1 vssd1 vccd1 vccd1 _5440_/X sky130_fd_sc_hd__o22a_1
XFILLER_118_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3346__A1 _3266_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5371_ _3059_/Y _5364_/Y _5370_/X _5363_/X vssd1 vssd1 vccd1 vccd1 _5371_/X sky130_fd_sc_hd__a31o_1
XFILLER_114_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3441__S1 _3551_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4322_ _4323_/B _4323_/A vssd1 vssd1 vccd1 vccd1 _4355_/A sky130_fd_sc_hd__and2b_1
XFILLER_99_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5099__A1 _3297_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout108 _3593_/A vssd1 vssd1 vccd1 vccd1 _3567_/B sky130_fd_sc_hd__buf_8
XFILLER_113_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4253_ _6094_/Q _3711_/X _4259_/S vssd1 vssd1 vccd1 vccd1 _6094_/D sky130_fd_sc_hd__mux2_1
Xfanout119 _3388_/B vssd1 vssd1 vccd1 vccd1 _3986_/A sky130_fd_sc_hd__buf_12
XFILLER_68_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3204_ _3498_/S vssd1 vssd1 vccd1 vccd1 _3204_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4184_ _4185_/A _4185_/B _4185_/C vssd1 vssd1 vccd1 vccd1 _4184_/X sky130_fd_sc_hd__and3_2
XFILLER_79_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3135_ _5072_/A _5054_/A _3135_/S vssd1 vssd1 vccd1 vccd1 _6010_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_857 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3066_ _5162_/B _3067_/B vssd1 vssd1 vccd1 vccd1 _3669_/B sky130_fd_sc_hd__or2_2
XFILLER_36_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5271__A1 _5072_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4074__A2 _4072_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout258_A _4270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5574__A2 _5909_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3968_ _5634_/A _5509_/C _5227_/B vssd1 vssd1 vccd1 vccd1 _5617_/C sky130_fd_sc_hd__or3_2
XFILLER_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5707_ _5707_/A _5707_/B vssd1 vssd1 vccd1 vccd1 _5707_/Y sky130_fd_sc_hd__nor2_1
X_3899_ _6042_/Q _3889_/X _3898_/Y vssd1 vssd1 vccd1 vccd1 _6042_/D sky130_fd_sc_hd__o21a_1
XFILLER_12_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5638_ _5638_/A _5638_/B _5638_/C vssd1 vssd1 vccd1 vccd1 _5647_/D sky130_fd_sc_hd__and3_1
XFILLER_12_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5569_ _4638_/B _5565_/Y _5568_/Y _5072_/C vssd1 vssd1 vccd1 vccd1 _5569_/X sky130_fd_sc_hd__o211a_1
XANTENNA__4202__B _4311_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4872__B _4872_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3769__A _5210_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3273__B1 _5263_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3576__A1 _3658_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5317__A2 _4234_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3328__B2 _3236_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4112__B _4197_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3009__A _5488_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3951__B _5635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3679__A _3974_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4940_ _4936_/X _4939_/X _5488_/A _4872_/B vssd1 vssd1 vccd1 vccd1 _4940_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_73_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3803__A2 _3777_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3398__B _3500_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4871_ _4863_/X _4870_/X _4931_/B vssd1 vssd1 vccd1 vccd1 _4871_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__5005__A1 _4745_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5005__B2 _4744_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3822_ _5706_/B _3845_/B vssd1 vssd1 vccd1 vccd1 _3822_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__5556__A2 _5556_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3753_ _3811_/S _3777_/S _3753_/C vssd1 vssd1 vccd1 vccd1 _4294_/B sky130_fd_sc_hd__and3_2
XFILLER_9_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4303__A _4334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5308__A2 _5300_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3684_ _3734_/A _5048_/C vssd1 vssd1 vccd1 vccd1 _3684_/X sky130_fd_sc_hd__or2_2
XANTENNA__3319__A1 _3312_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5423_ _4644_/B _5421_/Y _5422_/X _3121_/B _5507_/A vssd1 vssd1 vccd1 vccd1 _5423_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_133_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4022__B _5207_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5354_ _5595_/A _5354_/B vssd1 vssd1 vccd1 vccd1 _5354_/Y sky130_fd_sc_hd__nor2_1
XFILLER_114_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4305_ _4305_/A _4305_/B vssd1 vssd1 vccd1 vccd1 _4308_/A sky130_fd_sc_hd__nor2_4
X_5285_ _5512_/A _5257_/Y _5284_/Y _3122_/A vssd1 vssd1 vccd1 vccd1 _5285_/X sky130_fd_sc_hd__a211o_1
XFILLER_99_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4236_ _5767_/C _4238_/B vssd1 vssd1 vccd1 vccd1 _4239_/A sky130_fd_sc_hd__or2_4
XANTENNA__5492__A1 _5551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4167_ _4197_/A _4197_/B _4167_/C _4167_/D vssd1 vssd1 vccd1 vccd1 _4200_/A sky130_fd_sc_hd__and4_2
XFILLER_68_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3118_ _4963_/A _5069_/A vssd1 vssd1 vccd1 vccd1 _3118_/Y sky130_fd_sc_hd__nand2_2
XFILLER_55_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4098_ _4107_/C _4098_/B vssd1 vssd1 vccd1 vccd1 _4099_/B sky130_fd_sc_hd__or2_4
XFILLER_15_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3049_ _3107_/A _3050_/B vssd1 vssd1 vccd1 vccd1 _3049_/Y sky130_fd_sc_hd__nor2_4
XFILLER_130_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4213__A _4214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5483__A1 _6003_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4883__A _5454_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5235__B2 _5929_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4107__B _4176_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4746__B1 _4745_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout90 _3205_/A vssd1 vssd1 vccd1 vccd1 _5936_/A sky130_fd_sc_hd__buf_6
XANTENNA__3438__S _3551_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5171__B1 _5498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3681__B _3901_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5070_ _6197_/Q _5069_/X _5070_/S vssd1 vssd1 vccd1 vccd1 _5071_/B sky130_fd_sc_hd__mux2_1
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5474__A1 _4891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4021_ _4022_/C _3975_/C _4015_/X _4020_/X vssd1 vssd1 vccd1 vccd1 _4023_/B sky130_fd_sc_hd__o211a_1
XANTENNA__4793__A _4990_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5972_ _5110_/A _5963_/Y _6299_/Q vssd1 vssd1 vccd1 vccd1 _5972_/X sky130_fd_sc_hd__a21o_1
XFILLER_80_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3202__A _3880_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3788__A1 _3450_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4985__B1 _3116_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4923_ _4820_/B _4867_/A _4860_/Y _4900_/A _4925_/B vssd1 vssd1 vccd1 vccd1 _4924_/B
+ sky130_fd_sc_hd__a41o_1
XFILLER_80_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5529__A2 _5522_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4854_ _6190_/Q _4854_/B vssd1 vssd1 vccd1 vccd1 _4855_/B sky130_fd_sc_hd__nor2_1
XFILLER_21_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3856__B _5883_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3805_ _4734_/B _3816_/B _3804_/X vssd1 vssd1 vccd1 vccd1 _3805_/Y sky130_fd_sc_hd__o21ai_1
X_4785_ _4783_/Y _4784_/X _4778_/X vssd1 vssd1 vccd1 vccd1 _4785_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__4033__A _5436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3736_ _3736_/A _3744_/C vssd1 vssd1 vccd1 vccd1 _3810_/S sky130_fd_sc_hd__or2_2
XANTENNA_fanout123_A _3245_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3667_ _3631_/A _3666_/X _3633_/X vssd1 vssd1 vccd1 vccd1 _3667_/X sky130_fd_sc_hd__a21o_1
XFILLER_118_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3872__A _5943_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5406_ _6178_/Q _4234_/B _4058_/B _6138_/Q vssd1 vssd1 vccd1 vccd1 _5406_/X sky130_fd_sc_hd__o22a_1
XANTENNA__5701__A2 _3958_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3598_ _3599_/B _3599_/C vssd1 vssd1 vccd1 vccd1 _3643_/B sky130_fd_sc_hd__nand2_2
XFILLER_133_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3712__A1 _3711_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5337_ _5133_/X _5354_/B _5336_/X _5244_/A vssd1 vssd1 vccd1 vccd1 _5338_/B sky130_fd_sc_hd__o211a_1
XFILLER_114_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5268_ _4672_/A _4678_/Y _5561_/S vssd1 vssd1 vccd1 vccd1 _5284_/B sky130_fd_sc_hd__mux2_2
XFILLER_87_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5465__A1 _5607_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5799__A _5799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4219_ _4221_/A _4221_/B _4221_/C vssd1 vssd1 vccd1 vccd1 _4219_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_87_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5199_ _5202_/B _5199_/B _5199_/C vssd1 vssd1 vccd1 vccd1 _5199_/X sky130_fd_sc_hd__and3b_1
XFILLER_68_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3112__A _5065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3766__B _5503_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_466 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5456__A1 _5454_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout280 _6224_/Q vssd1 vssd1 vccd1 vccd1 _5387_/A sky130_fd_sc_hd__buf_4
XFILLER_15_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout291 _3105_/A vssd1 vssd1 vccd1 vccd1 _5162_/B sky130_fd_sc_hd__buf_6
XFILLER_46_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5208__A1 _5790_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5208__B2 _6162_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3022__A _3873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4967__B1 _5239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3676__B _5075_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4570_ _5543_/S _5625_/B _4580_/C _3971_/B _4604_/A vssd1 vssd1 vccd1 vccd1 _4572_/B
+ sky130_fd_sc_hd__o32a_1
XFILLER_128_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3521_ _3520_/X _3572_/A vssd1 vssd1 vccd1 vccd1 _3521_/X sky130_fd_sc_hd__and2b_1
XFILLER_6_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4003__D _5241_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6240_ _6241_/CLK _6240_/D vssd1 vssd1 vccd1 vccd1 _6240_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3452_ _3608_/A _3599_/B _3454_/C vssd1 vssd1 vccd1 vccd1 _3452_/X sky130_fd_sc_hd__or3_1
XANTENNA__5695__A1 _5710_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6171_ _6264_/CLK _6171_/D vssd1 vssd1 vccd1 vccd1 _6171_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4300__B _4426_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3383_ _4270_/A _3832_/A2 _3251_/B _3382_/X _3255_/Y vssd1 vssd1 vccd1 vccd1 _3384_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_124_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5122_ _5982_/A vssd1 vssd1 vccd1 vccd1 _5122_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5447__A1 _4872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5053_ _5090_/A _5731_/S vssd1 vssd1 vccd1 vccd1 _5203_/C sky130_fd_sc_hd__nor2_1
XFILLER_84_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5412__A _5412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4004_ _6292_/Q _3030_/Y _3033_/Y _6298_/Q vssd1 vssd1 vccd1 vccd1 _4004_/X sky130_fd_sc_hd__o22a_1
XFILLER_65_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5131__B _5131_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5955_ _5955_/A _5955_/B vssd1 vssd1 vccd1 vccd1 _5956_/C sky130_fd_sc_hd__nand2_1
XFILLER_34_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout240_A _4216_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4906_ _4625_/A _5093_/A _4904_/X _4905_/X _5071_/A vssd1 vssd1 vccd1 vccd1 _6191_/D
+ sky130_fd_sc_hd__o311a_1
XANTENNA_fanout338_A input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5886_ _5900_/A _5900_/B vssd1 vssd1 vccd1 vccd1 _5949_/A sky130_fd_sc_hd__nor2_1
XFILLER_21_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4837_ _5428_/A _4837_/B vssd1 vssd1 vccd1 vccd1 _4838_/B sky130_fd_sc_hd__or2_2
XFILLER_119_420 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5383__B1 _5251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5922__A2 _4586_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4768_ _4691_/A _4733_/X _4736_/X _4735_/B vssd1 vssd1 vccd1 vccd1 _4769_/B sky130_fd_sc_hd__a31o_2
XFILLER_107_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3719_ _6029_/Q _3718_/X _3731_/S vssd1 vssd1 vccd1 vccd1 _6029_/D sky130_fd_sc_hd__mux2_1
X_4699_ _4699_/A _4699_/B vssd1 vssd1 vccd1 vccd1 _4699_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_134_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5135__B1 _4648_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5686__A1 _5075_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5686__B2 _3458_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3697__A0 _5387_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5438__B2 _3236_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6233__CLK _6233_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4637__S _5041_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5610__A1 _3590_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5610__B2 _5943_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5913__A2 _4604_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3716__S _3731_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5126__A0 _5862_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3943__C _3943_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3688__A0 _3943_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3017__A _6200_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4652__A2 _4644_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5601__A1 _4645_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3687__A _5503_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5740_ _5740_/A _5740_/B _5740_/C vssd1 vssd1 vccd1 vccd1 _5740_/X sky130_fd_sc_hd__or3_2
XFILLER_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5671_ _3765_/B _5321_/X _5668_/Y _5669_/X _5670_/X vssd1 vssd1 vccd1 vccd1 _5671_/X
+ sky130_fd_sc_hd__o221a_1
X_4622_ _5625_/A _4622_/B _5220_/S vssd1 vssd1 vccd1 vccd1 _5132_/B sky130_fd_sc_hd__and3_2
XANTENNA__5904__A2 _3986_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3915__A1 _3711_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4553_ _6177_/Q _4553_/B vssd1 vssd1 vccd1 vccd1 _4553_/X sky130_fd_sc_hd__or2_1
XANTENNA__4311__A _4426_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3504_ _5707_/B _3599_/B vssd1 vssd1 vccd1 vccd1 _3504_/Y sky130_fd_sc_hd__xnor2_2
X_4484_ _6135_/Q _4499_/B vssd1 vssd1 vccd1 vccd1 _4484_/X sky130_fd_sc_hd__or2_1
X_6223_ _6254_/CLK _6223_/D vssd1 vssd1 vccd1 vccd1 _6223_/Q sky130_fd_sc_hd__dfxtp_1
X_3435_ _3450_/D _3435_/B vssd1 vssd1 vccd1 vccd1 _4619_/B sky130_fd_sc_hd__xnor2_4
XFILLER_116_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6154_ _6154_/CLK _6154_/D vssd1 vssd1 vccd1 vccd1 _6154_/Q sky130_fd_sc_hd__dfxtp_1
X_3366_ _6202_/Q _3388_/B _3658_/S vssd1 vssd1 vccd1 vccd1 _3366_/X sky130_fd_sc_hd__mux2_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5105_ _5105_/A _5105_/B _5105_/C vssd1 vssd1 vccd1 vccd1 _5129_/S sky130_fd_sc_hd__or3_4
XANTENNA_fanout190_A _3241_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6085_ _6265_/CLK _6085_/D vssd1 vssd1 vccd1 vccd1 _6085_/Q sky130_fd_sc_hd__dfxtp_1
X_3297_ _6200_/Q _3297_/B vssd1 vssd1 vccd1 vccd1 _3611_/A sky130_fd_sc_hd__nand2_8
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5036_ _5509_/C _5036_/B vssd1 vssd1 vccd1 vccd1 _5036_/Y sky130_fd_sc_hd__nor2_1
XFILLER_122_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_24 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3597__A _5707_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5938_ _3243_/Y _5928_/Y _5937_/X _5928_/B _4638_/A vssd1 vssd1 vccd1 vccd1 _5938_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__4800__C1 _5071_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5869_ _3958_/A _5119_/A _5869_/S vssd1 vssd1 vccd1 vccd1 _6290_/D sky130_fd_sc_hd__mux2_1
XANTENNA__5356__B1 _5556_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3906__A1 _3721_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput12 _6186_/Q vssd1 vssd1 vccd1 vccd1 io_out[10] sky130_fd_sc_hd__buf_4
XANTENNA__5659__A1 _5734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput23 _6196_/Q vssd1 vssd1 vccd1 vccd1 io_out[20] sky130_fd_sc_hd__buf_4
Xoutput34 _6287_/Q vssd1 vssd1 vccd1 vccd1 io_out[6] sky130_fd_sc_hd__buf_4
XFILLER_89_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5831__A1 _3583_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4891__A _4891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5926__S _5943_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5227__A _5227_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4131__A _4301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4570__A1 _5543_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4570__B2 _4604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3970__A _3970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3220_ _3231_/C vssd1 vssd1 vccd1 vccd1 _3631_/A sky130_fd_sc_hd__inv_2
XANTENNA__3125__A2 _4643_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3151_ _3312_/A _3677_/B vssd1 vssd1 vccd1 vccd1 _5143_/B sky130_fd_sc_hd__or2_4
XFILLER_39_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3082_ _5162_/B _4046_/A vssd1 vssd1 vccd1 vccd1 _3084_/B sky130_fd_sc_hd__nand2_2
XFILLER_82_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5822__A1 _5835_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5586__B1 _4644_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3984_ _5645_/A _5961_/B _3984_/C _3983_/X vssd1 vssd1 vccd1 vccd1 _3984_/X sky130_fd_sc_hd__or4b_4
X_5723_ _5710_/S _4167_/D _5442_/B _5734_/A _3950_/C vssd1 vssd1 vccd1 vccd1 _5723_/X
+ sky130_fd_sc_hd__o221a_1
X_5654_ _4658_/B _4663_/B _5703_/A vssd1 vssd1 vccd1 vccd1 _5654_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4605_ _4605_/A _4605_/B _5871_/A _4605_/D vssd1 vssd1 vccd1 vccd1 _5062_/B sky130_fd_sc_hd__and4_1
XFILLER_117_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5585_ _5603_/S _5582_/X _5602_/B _5584_/Y vssd1 vssd1 vccd1 vccd1 _5585_/X sky130_fd_sc_hd__a31o_1
XANTENNA__5137__A _5258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4561__A1 _3942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4536_ _6157_/Q _6170_/Q _4535_/Y vssd1 vssd1 vccd1 vccd1 _6169_/D sky130_fd_sc_hd__o21a_1
XANTENNA_fanout203_A _5622_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4976__A _6194_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4467_ _5926_/A0 _4466_/X _4477_/S vssd1 vssd1 vccd1 vccd1 _6127_/D sky130_fd_sc_hd__mux2_1
XFILLER_131_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3880__A _3880_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6206_ _6206_/CLK _6206_/D vssd1 vssd1 vccd1 vccd1 _6206_/Q sky130_fd_sc_hd__dfxtp_2
X_3418_ _3313_/Y _3416_/Y _3926_/B _4003_/C _3365_/Y vssd1 vssd1 vccd1 vccd1 _3418_/X
+ sky130_fd_sc_hd__o221a_1
X_4398_ _4399_/B _4399_/A vssd1 vssd1 vccd1 vccd1 _4417_/A sky130_fd_sc_hd__nand2b_1
XFILLER_86_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input8_A io_in[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6137_ _6177_/CLK _6137_/D vssd1 vssd1 vccd1 vccd1 _6137_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3349_ _3388_/A _3561_/A _3608_/A vssd1 vssd1 vccd1 vccd1 _3350_/B sky130_fd_sc_hd__a21bo_2
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_760 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6068_ _6290_/CLK _6068_/D vssd1 vssd1 vccd1 vccd1 _6068_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5019_ _4963_/A _5018_/X _5010_/X _4753_/A vssd1 vssd1 vccd1 vccd1 _5019_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_45_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4216__A _4216_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3120__A _4642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4552__A1 _3942_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4886__A _5454_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_43_clk_A clkbuf_3_4__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4304__A1 _4334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_866 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5804__A1 _3375_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5280__A2 _3243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3949__B _3964_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3030__A _4633_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3579__C1 _3145_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3965__A _4638_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3684__B _5048_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4543__A1 _3943_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3346__A2 _3266_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5370_ _5370_/A _5653_/A _5368_/X vssd1 vssd1 vccd1 vccd1 _5370_/X sky130_fd_sc_hd__or3b_2
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4321_ _4321_/A _4321_/B vssd1 vssd1 vccd1 vccd1 _4323_/B sky130_fd_sc_hd__nor2_2
XFILLER_99_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5099__A2 _5097_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4252_ _4252_/A _5769_/S vssd1 vssd1 vccd1 vccd1 _4259_/S sky130_fd_sc_hd__nand2_8
Xfanout109 _3492_/X vssd1 vssd1 vccd1 vccd1 _3593_/A sky130_fd_sc_hd__buf_6
XFILLER_113_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3203_ _3212_/A _5707_/A _4614_/A vssd1 vssd1 vccd1 vccd1 _3203_/X sky130_fd_sc_hd__or3_2
XFILLER_86_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4183_ _4185_/B _4185_/C _4185_/A vssd1 vssd1 vccd1 vccd1 _4183_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__3205__A _3205_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3134_ _4846_/A _6009_/Q _3135_/S vssd1 vssd1 vccd1 vccd1 _6009_/D sky130_fd_sc_hd__mux2_1
XFILLER_28_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3806__A0 _5677_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3065_ _5162_/B _3067_/B vssd1 vssd1 vccd1 vccd1 _5238_/B sky130_fd_sc_hd__nor2_2
XFILLER_94_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3859__B _5976_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4036__A _5767_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout153_A _3069_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3967_ _5138_/A _5943_/B _5206_/A vssd1 vssd1 vccd1 vccd1 _5961_/B sky130_fd_sc_hd__or3b_2
X_5706_ _5733_/A _5706_/B vssd1 vssd1 vccd1 vccd1 _5706_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_fanout320_A _5799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_30_clk clkbuf_3_5__f_clk/X vssd1 vssd1 vccd1 vccd1 _6263_/CLK sky130_fd_sc_hd__clkbuf_16
X_3898_ _3889_/X _3897_/Y _5192_/A vssd1 vssd1 vccd1 vccd1 _3898_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_109_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3594__B _3594_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5637_ _5645_/B _5637_/B _5632_/X vssd1 vssd1 vccd1 vccd1 _5642_/B sky130_fd_sc_hd__or3b_1
XANTENNA__5731__A0 _4883_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5568_ _5583_/B _5567_/Y _5291_/Y vssd1 vssd1 vccd1 vccd1 _5568_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_88_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_584 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4519_ _3942_/A _4518_/X _4521_/S vssd1 vssd1 vccd1 vccd1 _6155_/D sky130_fd_sc_hd__mux2_1
XFILLER_2_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5499_ _5504_/A _5500_/B vssd1 vssd1 vccd1 vccd1 _5540_/C sky130_fd_sc_hd__and2_4
XFILLER_78_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5495__C1 _5251_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout66_A _4601_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3769__B _4539_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4470__A0 _5358_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3273__A1 _4096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3273__B2 _3885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3576__A2 _3567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_21_clk _6084_/CLK vssd1 vssd1 vccd1 vccd1 _6265_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_6_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3328__A2 _5743_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4112__C _4112_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3025__A _3958_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5253__A2 _5556_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3679__B _5172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4461__A0 _5255_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3264__A1 _5818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4870_ _4872_/A _4645_/Y _4869_/X _5463_/A _4963_/A vssd1 vssd1 vccd1 vccd1 _4870_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_33_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3821_ _6038_/Q _3771_/X _3819_/Y _3820_/X vssd1 vssd1 vccd1 vccd1 _6038_/D sky130_fd_sc_hd__a211o_1
XFILLER_60_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3752_ _3156_/Y _5464_/A _3744_/C _3810_/S _3751_/X vssd1 vssd1 vccd1 vccd1 _3753_/C
+ sky130_fd_sc_hd__o311a_1
Xclkbuf_leaf_12_clk _6219_/CLK vssd1 vssd1 vccd1 vccd1 _6218_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_9_472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4303__B _4389_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3683_ _5512_/A _5943_/B vssd1 vssd1 vccd1 vccd1 _5048_/C sky130_fd_sc_hd__nand2_8
XANTENNA__4516__A1 _5385_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5422_ _6009_/Q _5428_/A _5456_/S vssd1 vssd1 vccd1 vccd1 _5422_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4022__C _4022_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5353_ _5353_/A vssd1 vssd1 vccd1 vccd1 _5353_/Y sky130_fd_sc_hd__inv_2
XFILLER_114_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5415__A _5446_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4304_ _4334_/A _4389_/B _4303_/C vssd1 vssd1 vccd1 vccd1 _4305_/B sky130_fd_sc_hd__a21oi_2
XFILLER_102_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5284_ _5512_/A _5284_/B vssd1 vssd1 vccd1 vccd1 _5284_/Y sky130_fd_sc_hd__nor2_1
XFILLER_99_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4235_ _5767_/C _4238_/B vssd1 vssd1 vccd1 vccd1 _4490_/B sky130_fd_sc_hd__nor2_2
XFILLER_87_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5492__A2 _5482_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4166_ _4197_/A _4167_/C _4167_/D _4197_/B vssd1 vssd1 vccd1 vccd1 _4168_/A sky130_fd_sc_hd__a22oi_2
XANTENNA__5229__C1 _5227_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3117_ _3958_/A _4654_/A vssd1 vssd1 vccd1 vccd1 _5050_/C sky130_fd_sc_hd__nor2_2
XFILLER_95_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout270_A _6230_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4097_ _4096_/A _4111_/B _4112_/C _4197_/B vssd1 vssd1 vccd1 vccd1 _4098_/B sky130_fd_sc_hd__a22oi_1
XFILLER_83_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3048_ _5179_/A _3092_/B _3107_/A vssd1 vssd1 vccd1 vccd1 _5075_/B sky130_fd_sc_hd__or3_4
XFILLER_24_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4999_ _6005_/Q _4999_/B vssd1 vssd1 vccd1 vccd1 _4999_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__3558__A2 _3607_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5952__B1 _3883_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4213__B _4214_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4507__A1 _5305_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5325__A _5333_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4883__B _4883_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4994__A1 _5547_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3719__S _3731_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4746__A1 _4744_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4746__B2 _4740_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout80 _3103_/Y vssd1 vssd1 vccd1 vccd1 _5051_/D sky130_fd_sc_hd__buf_6
XFILLER_128_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout91 _3080_/Y vssd1 vssd1 vccd1 vccd1 _3205_/A sky130_fd_sc_hd__buf_4
XFILLER_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5171__A1 _5172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3681__C _5766_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5474__A2 _5251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4020_ _5976_/A _4020_/B _4009_/B vssd1 vssd1 vccd1 vccd1 _4020_/X sky130_fd_sc_hd__or3b_1
XFILLER_111_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5889__B _5889_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_1_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _6196_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_84_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3485__A1 _4334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3485__B2 _3484_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5971_ _5968_/Y _5970_/X _5986_/B1 vssd1 vssd1 vccd1 vccd1 _6298_/D sky130_fd_sc_hd__a21oi_1
XFILLER_64_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5631__C1 _3974_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3202__B _5148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4922_ _4964_/A _4922_/B vssd1 vssd1 vccd1 vccd1 _4934_/A sky130_fd_sc_hd__and2_2
XFILLER_80_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4853_ _6190_/Q _4854_/B vssd1 vssd1 vccd1 vccd1 _4916_/C sky130_fd_sc_hd__and2_2
XFILLER_100_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3804_ _4726_/B _3740_/X _3749_/X _3803_/X vssd1 vssd1 vccd1 vccd1 _3804_/X sky130_fd_sc_hd__a211o_1
XANTENNA__3856__C _3952_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4784_ _4791_/A _4791_/B _4782_/Y _3116_/X vssd1 vssd1 vccd1 vccd1 _4784_/X sky130_fd_sc_hd__a31o_1
XFILLER_21_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3735_ _3736_/A _3744_/C vssd1 vssd1 vccd1 vccd1 _3834_/B sky130_fd_sc_hd__nor2_1
XANTENNA__4033__B _5742_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3666_ _3476_/A _5900_/A _3665_/X vssd1 vssd1 vccd1 vccd1 _3666_/X sky130_fd_sc_hd__o21a_4
XANTENNA_fanout116_A _5848_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5405_ _5436_/A _6154_/Q _5436_/C vssd1 vssd1 vccd1 vccd1 _5405_/X sky130_fd_sc_hd__and3_1
XFILLER_133_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3597_ _5707_/B _3597_/B _3607_/B vssd1 vssd1 vccd1 vccd1 _3599_/C sky130_fd_sc_hd__and3_1
X_5336_ _5072_/B _5329_/Y _5335_/X vssd1 vssd1 vccd1 vccd1 _5336_/X sky130_fd_sc_hd__a21o_1
XFILLER_130_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5267_ _5265_/Y _5266_/X _3059_/Y _5261_/Y vssd1 vssd1 vccd1 vccd1 _5267_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_88_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4218_ _4218_/A _4218_/B vssd1 vssd1 vccd1 vccd1 _4221_/C sky130_fd_sc_hd__nor2_2
XFILLER_56_611 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5198_ _3116_/X _3168_/Y _5617_/A _3118_/Y vssd1 vssd1 vccd1 vccd1 _5199_/C sky130_fd_sc_hd__a31o_1
XFILLER_28_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4149_ _4150_/A _4150_/B vssd1 vssd1 vccd1 vccd1 _4149_/Y sky130_fd_sc_hd__nand2b_2
XFILLER_83_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3112__B _3112_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4728__A1 _4697_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5153__A1 _5131_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout270 _6230_/Q vssd1 vssd1 vccd1 vccd1 _5547_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_59_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3467__A1 _3458_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout281 _6223_/Q vssd1 vssd1 vccd1 vccd1 _5358_/A sky130_fd_sc_hd__clkbuf_16
XANTENNA__5861__C1 _5866_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout292 _6211_/Q vssd1 vssd1 vccd1 vccd1 _3105_/A sky130_fd_sc_hd__buf_6
XFILLER_115_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5613__C1 _5948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4967__A1 _6193_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3957__B _3960_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4719__A1 _6221_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4719__B2 _5463_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3520_ _3462_/X _3935_/C _3518_/Y _3621_/A vssd1 vssd1 vccd1 vccd1 _3520_/X sky130_fd_sc_hd__a31o_1
XFILLER_6_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5144__A1 _5054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3451_ _3450_/A _3986_/A _3801_/A _3450_/D vssd1 vssd1 vccd1 vccd1 _3454_/C sky130_fd_sc_hd__o31a_1
XFILLER_115_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5695__A2 _4112_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3382_ _5929_/B2 _3381_/X _3380_/X vssd1 vssd1 vccd1 vccd1 _3382_/X sky130_fd_sc_hd__a21o_2
X_6170_ _6170_/CLK _6170_/D vssd1 vssd1 vccd1 vccd1 _6170_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5121_ _4767_/A _5241_/A _5120_/Y vssd1 vssd1 vccd1 vccd1 _5982_/A sky130_fd_sc_hd__o21a_1
XFILLER_124_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5052_ _5052_/A _5052_/B vssd1 vssd1 vccd1 vccd1 _5838_/A sky130_fd_sc_hd__or2_1
XFILLER_111_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4003_ _5840_/A _4003_/B _4003_/C _5241_/B vssd1 vssd1 vccd1 vccd1 _4009_/B sky130_fd_sc_hd__and4_2
XANTENNA__4309__A _4410_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3213__A _4638_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5604__C1 _3060_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5954_ _3941_/A _3923_/B _5949_/X _5953_/X vssd1 vssd1 vccd1 vccd1 _5956_/B sky130_fd_sc_hd__a31o_1
XFILLER_111_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4905_ _6191_/Q _4970_/B vssd1 vssd1 vccd1 vccd1 _4905_/X sky130_fd_sc_hd__or2_1
XFILLER_80_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5885_ _6291_/Q _5879_/X _5883_/X _5884_/X _5956_/A vssd1 vssd1 vccd1 vccd1 _6291_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4836_ _5428_/A _4837_/B vssd1 vssd1 vccd1 vccd1 _4836_/X sky130_fd_sc_hd__and2_1
XANTENNA_fanout233_A _6290_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5907__B1 _4576_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5383__A1 _5943_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4979__A _5547_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4767_ _4767_/A _4767_/B vssd1 vssd1 vccd1 vccd1 _4769_/A sky130_fd_sc_hd__xnor2_2
XFILLER_119_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3718_ _6013_/Q _3706_/Y _3717_/X vssd1 vssd1 vccd1 vccd1 _3718_/X sky130_fd_sc_hd__a21o_4
XFILLER_134_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4698_ _4698_/A _4698_/B vssd1 vssd1 vccd1 vccd1 _4699_/B sky130_fd_sc_hd__nand2_1
X_3649_ _3649_/A _3649_/B vssd1 vssd1 vccd1 vccd1 _3651_/B sky130_fd_sc_hd__nand2_2
XFILLER_134_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_58 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5319_ _6021_/Q _5349_/B1 _5742_/B _6244_/Q vssd1 vssd1 vccd1 vccd1 _5319_/X sky130_fd_sc_hd__o22a_1
XFILLER_29_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6299_ _6299_/CLK _6299_/D vssd1 vssd1 vccd1 vccd1 _6299_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5438__A2 _5767_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5610__A2 _5442_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3793__A _3937_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5126__A1 _4846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5513__A _5513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4637__A0 _6184_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3033__A _5344_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3687__B _5943_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3612__B2 _3541_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5670_ _5710_/S _4111_/B _3950_/C vssd1 vssd1 vccd1 vccd1 _5670_/X sky130_fd_sc_hd__o21a_1
XANTENNA_clkbuf_0_clk_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4621_ _3495_/B _5706_/B _5733_/B _4621_/D vssd1 vssd1 vccd1 vccd1 _5220_/S sky130_fd_sc_hd__and4b_4
XFILLER_129_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4552_ _3942_/D _4237_/Y _4550_/X _4551_/Y vssd1 vssd1 vccd1 vccd1 _6176_/D sky130_fd_sc_hd__a22o_1
XFILLER_7_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3503_ _3561_/A _3507_/B vssd1 vssd1 vccd1 vccd1 _3503_/Y sky130_fd_sc_hd__nand2b_1
X_4483_ _5935_/A0 _4501_/A2 _4481_/X _4482_/X vssd1 vssd1 vccd1 vccd1 _6134_/D sky130_fd_sc_hd__a22o_1
XANTENNA__4311__B _4311_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3128__A0 _4633_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3208__A _5703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6222_ _6227_/CLK _6222_/D vssd1 vssd1 vccd1 vccd1 _6222_/Q sky130_fd_sc_hd__dfxtp_4
X_3434_ _3599_/A _3405_/B _3387_/X vssd1 vssd1 vccd1 vccd1 _3435_/B sky130_fd_sc_hd__a21oi_4
XFILLER_131_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6153_ _6154_/CLK _6153_/D vssd1 vssd1 vccd1 vccd1 _6153_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3365_ _4003_/B _3365_/B vssd1 vssd1 vccd1 vccd1 _3365_/Y sky130_fd_sc_hd__nand2_2
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5532__A1_N _4586_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5104_ _5104_/A _5104_/B vssd1 vssd1 vccd1 vccd1 _5105_/C sky130_fd_sc_hd__nor2_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6084_ _6084_/CLK _6084_/D vssd1 vssd1 vccd1 vccd1 _6084_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3296_ _3296_/A _6199_/Q vssd1 vssd1 vccd1 vccd1 _3541_/A sky130_fd_sc_hd__nand2_8
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5035_ _5034_/A _5028_/X _5034_/Y vssd1 vssd1 vccd1 vccd1 _5035_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_100_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3851__A1 _4883_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3597__B _3597_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5937_ _5503_/A _5934_/B _5110_/A _5936_/X vssd1 vssd1 vccd1 vccd1 _5937_/X sky130_fd_sc_hd__o211a_1
XFILLER_80_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5868_ _5136_/C _5114_/A _5869_/S vssd1 vssd1 vccd1 vccd1 _6289_/D sky130_fd_sc_hd__mux2_1
XANTENNA__5356__A1 _5058_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4819_ _5385_/A _4819_/B vssd1 vssd1 vccd1 vccd1 _4820_/B sky130_fd_sc_hd__or2_4
X_5799_ _5799_/A _5799_/B vssd1 vssd1 vccd1 vccd1 _5819_/A sky130_fd_sc_hd__nand2_4
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3118__A _4963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput13 _6187_/Q vssd1 vssd1 vccd1 vccd1 io_out[11] sky130_fd_sc_hd__buf_4
XANTENNA__5659__A2 _5283_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput24 _6197_/Q vssd1 vssd1 vccd1 vccd1 io_out[21] sky130_fd_sc_hd__buf_4
Xoutput35 _6288_/Q vssd1 vssd1 vccd1 vccd1 io_out[7] sky130_fd_sc_hd__buf_4
XFILLER_1_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5333__A _5333_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4891__B _4979_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5479__S _5539_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_3_1__f_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _6230_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__5227__B _5227_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4131__B _4311_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3028__A _4540_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3970__B _4604_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3125__A3 _5498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3150_ _4622_/B _3970_/A vssd1 vssd1 vccd1 vccd1 _3677_/B sky130_fd_sc_hd__nand2_8
X_3081_ _5403_/A _5512_/A vssd1 vssd1 vccd1 vccd1 _3081_/Y sky130_fd_sc_hd__nor2_2
XFILLER_67_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4086__A1 _4136_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5897__B _5898_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5586__A1 _6008_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3983_ _5874_/A _5644_/A _3983_/C vssd1 vssd1 vccd1 vccd1 _3983_/X sky130_fd_sc_hd__and3_1
XFILLER_22_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5722_ _6057_/Q _6300_/Q _5735_/S vssd1 vssd1 vccd1 vccd1 _5722_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5653_ _5653_/A _5653_/B vssd1 vssd1 vccd1 vccd1 _5653_/X sky130_fd_sc_hd__or2_1
X_4604_ _4604_/A _4604_/B _4604_/C _5928_/B vssd1 vssd1 vccd1 vccd1 _5248_/A sky130_fd_sc_hd__or4_1
X_5584_ _5603_/S _5595_/B vssd1 vssd1 vccd1 vccd1 _5584_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__5137__B _5928_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4535_ _6157_/Q _6170_/Q _4540_/A vssd1 vssd1 vccd1 vccd1 _4535_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_116_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4466_ _6221_/Q _6127_/Q _4476_/S vssd1 vssd1 vccd1 vccd1 _4466_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5471__A1_N _5909_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3880__B _3880_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6205_ _6302_/CLK _6205_/D vssd1 vssd1 vccd1 vccd1 _6205_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_132_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3417_ _6203_/Q _3410_/B _3658_/S vssd1 vssd1 vccd1 vccd1 _3926_/B sky130_fd_sc_hd__mux2_1
X_4397_ _4373_/A _4373_/B _4376_/A vssd1 vssd1 vccd1 vccd1 _4399_/B sky130_fd_sc_hd__o21a_1
XFILLER_131_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6136_ _6176_/CLK _6136_/D vssd1 vssd1 vccd1 vccd1 _6136_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3348_ _3388_/A _3986_/A vssd1 vssd1 vccd1 vccd1 _3353_/A sky130_fd_sc_hd__xnor2_4
XFILLER_133_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3277__A_N _6292_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4992__A _5330_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6067_ _6209_/CLK _6067_/D vssd1 vssd1 vccd1 vccd1 _6067_/Q sky130_fd_sc_hd__dfxtp_4
X_3279_ _4216_/A _3257_/B _5450_/B _3885_/A vssd1 vssd1 vccd1 vccd1 _3284_/A sky130_fd_sc_hd__a22o_4
XFILLER_39_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5018_ _5547_/A _5463_/A _5017_/X _4638_/A vssd1 vssd1 vccd1 vccd1 _5018_/X sky130_fd_sc_hd__o22a_1
XFILLER_73_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3824__A1 _3594_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_775 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_499 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4216__B _4216_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3120__B _3121_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3588__B1 _5743_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4886__B _4886_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4304__A2 _4389_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_878 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3815__A1 _4772_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4240__A1 _3711_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3965__B _5928_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5238__A _5238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4320_ _4320_/A _4320_/B vssd1 vssd1 vccd1 vccd1 _4323_/A sky130_fd_sc_hd__xnor2_4
XFILLER_99_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4251_ _5743_/C _4251_/B vssd1 vssd1 vccd1 vccd1 _5769_/S sky130_fd_sc_hd__or2_4
XFILLER_114_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3202_ _3880_/B _5148_/A vssd1 vssd1 vccd1 vccd1 _4614_/A sky130_fd_sc_hd__nand2_4
XFILLER_113_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4182_ _4181_/B _4181_/C _4181_/A vssd1 vssd1 vccd1 vccd1 _4185_/C sky130_fd_sc_hd__a21o_2
XFILLER_67_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3205__B _3257_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3133_ _4819_/B _6008_/Q _3135_/S vssd1 vssd1 vccd1 vccd1 _6008_/D sky130_fd_sc_hd__mux2_1
XFILLER_94_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3920__S _3921_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3064_ _3092_/B _3107_/A _5179_/A vssd1 vssd1 vccd1 vccd1 _3067_/B sky130_fd_sc_hd__or3b_4
XFILLER_48_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3221__A _5840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4036__B _5925_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3966_ _5934_/A _3966_/B vssd1 vssd1 vccd1 vccd1 _5206_/A sky130_fd_sc_hd__nand2_1
XFILLER_10_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5705_ _5730_/A _5888_/B _5704_/X _5732_/C1 vssd1 vssd1 vccd1 vccd1 _5705_/X sky130_fd_sc_hd__o211a_1
X_3897_ _3964_/B _3897_/B vssd1 vssd1 vccd1 vccd1 _3897_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5148__A _5148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5636_ _5838_/B _5636_/B _5870_/B vssd1 vssd1 vccd1 vccd1 _5645_/B sky130_fd_sc_hd__or3b_1
XANTENNA_fanout313_A _5556_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5567_ _5567_/A _5567_/B vssd1 vssd1 vccd1 vccd1 _5567_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__5731__A1 _4877_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3891__A _4604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4518_ _5446_/B _6155_/Q _4520_/S vssd1 vssd1 vccd1 vccd1 _4518_/X sky130_fd_sc_hd__mux2_1
X_5498_ _5498_/A _5512_/B vssd1 vssd1 vccd1 vccd1 _5503_/B sky130_fd_sc_hd__nor2_1
XFILLER_117_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4449_ _6121_/Q _4458_/B vssd1 vssd1 vccd1 vccd1 _4449_/X sky130_fd_sc_hd__or2_1
XFILLER_77_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3115__B _3116_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6119_ _6155_/CLK _6119_/D vssd1 vssd1 vccd1 vccd1 _6119_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5798__A1 _3730_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout59_A _3958_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5330__B _5330_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3769__C _3772_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3273__A2 _3257_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4661__S _4812_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5058__A _5058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5722__A1 _6300_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4112__D _4112_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5486__B1 _5551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5789__A1 _5480_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3679__C _5330_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3264__A2 _5622_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3976__A _5097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3820_ _4334_/A _3832_/A2 _3484_/X _3765_/X _3772_/X vssd1 vssd1 vccd1 vccd1 _3820_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_60_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5410__B1 _5409_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3751_ _3751_/A _3812_/S _3841_/S _3816_/B vssd1 vssd1 vccd1 vccd1 _3751_/X sky130_fd_sc_hd__and4_1
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3682_ _5635_/A _3893_/B _3883_/A vssd1 vssd1 vccd1 vccd1 _5943_/B sky130_fd_sc_hd__nor3_4
XFILLER_9_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5421_ _5480_/C _5421_/B vssd1 vssd1 vccd1 vccd1 _5421_/Y sky130_fd_sc_hd__nor2_2
XANTENNA__3915__S _3921_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5352_ _5348_/X _5349_/X _5351_/X _5470_/S vssd1 vssd1 vccd1 vccd1 _5353_/A sky130_fd_sc_hd__a22o_4
XANTENNA__4600__A _4963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4303_ _4334_/A _4389_/B _4303_/C vssd1 vssd1 vccd1 vccd1 _4305_/A sky130_fd_sc_hd__and3_2
X_5283_ _5283_/A vssd1 vssd1 vccd1 vccd1 _5283_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3216__A _5840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4234_ _5436_/A _4234_/B vssd1 vssd1 vccd1 vccd1 _4238_/B sky130_fd_sc_hd__or2_2
XFILLER_101_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4165_ _4165_/A _4165_/B _4165_/C vssd1 vssd1 vccd1 vccd1 _4169_/B sky130_fd_sc_hd__nand3_2
XFILLER_83_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3116_ _6216_/Q _3116_/B vssd1 vssd1 vccd1 vccd1 _3116_/X sky130_fd_sc_hd__or2_4
X_4096_ _4096_/A _4136_/A _4311_/B _4309_/B vssd1 vssd1 vccd1 vccd1 _4107_/C sky130_fd_sc_hd__and4_1
XFILLER_83_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3047_ _5179_/A _3092_/B _3107_/A vssd1 vssd1 vccd1 vccd1 _5239_/B sky130_fd_sc_hd__nor3_4
XANTENNA__4047__A _4596_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout263_A _5109_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3886__A _5870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_42_clk_A clkbuf_3_4__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4998_ _6194_/Q _5046_/B _4997_/Y _5047_/C1 vssd1 vssd1 vccd1 vccd1 _6194_/D sky130_fd_sc_hd__o211a_1
XFILLER_23_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3949_ _4638_/A _3964_/B vssd1 vssd1 vccd1 vccd1 _3949_/Y sky130_fd_sc_hd__nand2_2
XANTENNA__5952__A1 _3943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5619_ _5622_/A _5840_/B _4648_/A _4946_/A vssd1 vssd1 vccd1 vccd1 _5619_/X sky130_fd_sc_hd__o211a_1
XFILLER_125_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5704__A1 _3740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5468__B1 _4058_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5341__A _5344_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4994__A2 _4644_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout70 _3868_/Y vssd1 vssd1 vccd1 vccd1 _5911_/C sky130_fd_sc_hd__clkbuf_4
Xfanout81 _3102_/Y vssd1 vssd1 vccd1 vccd1 _4753_/A sky130_fd_sc_hd__buf_8
Xfanout92 _5058_/A vssd1 vssd1 vccd1 vccd1 _5551_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_128_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3036__A _5392_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5251__A _5251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5970_ _5970_/A _5970_/B vssd1 vssd1 vccd1 vccd1 _5970_/X sky130_fd_sc_hd__or2_1
XFILLER_52_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4434__A1 _3853_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4921_ _5488_/A _4979_/B vssd1 vssd1 vccd1 vccd1 _4922_/B sky130_fd_sc_hd__or2_1
XFILLER_46_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5397__S _5539_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4852_ _4843_/X _4851_/X _3116_/B vssd1 vssd1 vccd1 vccd1 _4852_/X sky130_fd_sc_hd__o21a_2
XFILLER_60_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3803_ _4162_/A _3777_/S _3802_/Y _3751_/A vssd1 vssd1 vccd1 vccd1 _3803_/X sky130_fd_sc_hd__o211a_1
XFILLER_20_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4783_ _4791_/A _4782_/Y _4791_/B vssd1 vssd1 vccd1 vccd1 _4783_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_20_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3734_ _3734_/A _3750_/C vssd1 vssd1 vccd1 vccd1 _3744_/C sky130_fd_sc_hd__or2_4
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_17 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3665_ _3227_/X _4877_/B _3664_/X _3583_/S vssd1 vssd1 vccd1 vccd1 _3665_/X sky130_fd_sc_hd__a211o_1
XANTENNA__5426__A _5428_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5404_ _4596_/D _5389_/Y _5397_/X _5463_/A _5072_/C vssd1 vssd1 vccd1 vccd1 _5404_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_106_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3596_ _3599_/A _3607_/A _3642_/B _3387_/A vssd1 vssd1 vccd1 vccd1 _3596_/X sky130_fd_sc_hd__a22o_1
XFILLER_133_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5335_ _4644_/B _5354_/B _5331_/X _5058_/A vssd1 vssd1 vccd1 vccd1 _5335_/X sky130_fd_sc_hd__a211o_1
XFILLER_114_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5266_ _5265_/A _5265_/B _5653_/A vssd1 vssd1 vccd1 vccd1 _5266_/X sky130_fd_sc_hd__a21o_1
XFILLER_87_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4217_ _4216_/A _4216_/B _4216_/C vssd1 vssd1 vccd1 vccd1 _4218_/B sky130_fd_sc_hd__a21oi_1
XFILLER_75_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_815 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5197_ _6216_/Q _5197_/B vssd1 vssd1 vccd1 vccd1 _5199_/B sky130_fd_sc_hd__or2_1
XANTENNA__5161__A _5192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4148_ _4148_/A _4148_/B vssd1 vssd1 vccd1 vccd1 _4150_/B sky130_fd_sc_hd__xnor2_4
XFILLER_83_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4079_ _3783_/B _4069_/B _4072_/C _6080_/Q vssd1 vssd1 vccd1 vccd1 _4079_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_83_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4728__A2 _4697_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5689__A0 _4772_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4113__B1 _4112_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout260 _6236_/Q vssd1 vssd1 vccd1 vccd1 _3943_/A sky130_fd_sc_hd__buf_6
XFILLER_121_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout271 _5540_/B vssd1 vssd1 vccd1 vccd1 _5547_/B sky130_fd_sc_hd__buf_4
XFILLER_59_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5071__A _5071_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout282 _6223_/Q vssd1 vssd1 vccd1 vccd1 _5387_/B sky130_fd_sc_hd__buf_2
XFILLER_87_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5861__B1 _5860_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout293 _6210_/Q vssd1 vssd1 vccd1 vccd1 _5258_/A sky130_fd_sc_hd__buf_8
XFILLER_120_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3303__B _3388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4967__A2 _5561_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5010__S _5034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5916__A1 _4577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3450_ _3450_/A _3986_/A _3500_/A _3450_/D vssd1 vssd1 vccd1 vccd1 _3599_/B sky130_fd_sc_hd__nor4_4
XANTENNA__5144__A2 _4946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3381_ _6260_/Q _6052_/Q _6045_/Q _6029_/Q _3241_/A _3241_/B vssd1 vssd1 vccd1 vccd1
+ _3381_/X sky130_fd_sc_hd__mux4_1
XFILLER_97_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5120_ _6238_/Q _5934_/A vssd1 vssd1 vccd1 vccd1 _5120_/Y sky130_fd_sc_hd__nand2_1
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4104__B1 _4072_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5051_ _6217_/Q _5051_/B _5051_/C _5051_/D vssd1 vssd1 vccd1 vccd1 _5639_/B sky130_fd_sc_hd__or4_1
XFILLER_85_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5852__A0 _3500_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4655__A1 _5221_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4002_ _5707_/A _3615_/B _3987_/B _5712_/S _3179_/X vssd1 vssd1 vccd1 vccd1 _4002_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_84_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4309__B _4309_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3213__B _5570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4407__A1 _3819_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5953_ _5883_/A _5112_/X _5952_/X _5955_/B vssd1 vssd1 vccd1 vccd1 _5953_/X sky130_fd_sc_hd__a31o_1
XFILLER_34_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4904_ _5480_/B _5871_/C _4903_/X _4931_/B vssd1 vssd1 vccd1 vccd1 _4904_/X sky130_fd_sc_hd__o22a_1
X_5884_ _3941_/A _3937_/D _5879_/X vssd1 vssd1 vccd1 vccd1 _5884_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__3630__A2 _5898_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4835_ _6189_/Q _5046_/B _4834_/Y _5047_/C1 vssd1 vssd1 vccd1 vccd1 _6189_/D sky130_fd_sc_hd__o211a_1
XANTENNA__5907__A1 _6292_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4766_ _5367_/A _4767_/B vssd1 vssd1 vccd1 vccd1 _4766_/X sky130_fd_sc_hd__and2_1
XANTENNA__4979__B _4979_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3883__B _3975_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3717_ _4111_/B _5743_/C _3708_/Y _5540_/B vssd1 vssd1 vccd1 vccd1 _3717_/X sky130_fd_sc_hd__o22a_1
X_4697_ _4697_/A _4697_/B vssd1 vssd1 vccd1 vccd1 _4698_/B sky130_fd_sc_hd__nand2_1
XFILLER_107_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3648_ _6208_/Q _3986_/B vssd1 vssd1 vccd1 vccd1 _3651_/A sky130_fd_sc_hd__nand2_1
XFILLER_136_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3579_ _3365_/B _3618_/B _3578_/X _3312_/B _3145_/C vssd1 vssd1 vccd1 vccd1 _3579_/Y
+ sky130_fd_sc_hd__a221oi_2
X_5318_ _6127_/Q _5767_/B _5316_/X _3236_/Y _5317_/X vssd1 vssd1 vccd1 vccd1 _5318_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_102_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6298_ _6302_/CLK _6298_/D vssd1 vssd1 vccd1 vccd1 _6298_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5249_ _5172_/Y _5249_/B _5249_/C _5249_/D vssd1 vssd1 vccd1 vccd1 _5250_/D sky130_fd_sc_hd__and4b_1
XFILLER_103_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3123__B _5072_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4235__A _5767_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3385__A1 _3387_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4582__B1 _4587_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3385__B2 _3599_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4637__A1 _4634_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3968__B _5509_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3612__A2 _3594_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4620_ _4620_/A _4620_/B _5721_/B _4620_/D vssd1 vssd1 vccd1 vccd1 _4621_/D sky130_fd_sc_hd__and4_1
XFILLER_129_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4551_ _3011_/Y _4562_/B _4237_/Y vssd1 vssd1 vccd1 vccd1 _4551_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_129_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3502_ _3593_/B _3502_/B vssd1 vssd1 vccd1 vccd1 _3507_/B sky130_fd_sc_hd__nand2b_1
X_4482_ _4672_/A _4239_/A _4059_/B vssd1 vssd1 vccd1 vccd1 _4482_/X sky130_fd_sc_hd__o21a_1
XFILLER_116_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3128__A1 _4974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6221_ _6227_/CLK _6221_/D vssd1 vssd1 vccd1 vccd1 _6221_/Q sky130_fd_sc_hd__dfxtp_4
X_3433_ _4301_/A _3832_/A2 _3251_/B _3432_/Y _3255_/Y vssd1 vssd1 vccd1 vccd1 _3433_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_131_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6152_ _6176_/CLK _6152_/D vssd1 vssd1 vccd1 vccd1 _6152_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3364_ _3935_/B _3364_/B vssd1 vssd1 vccd1 vccd1 _3364_/X sky130_fd_sc_hd__xor2_1
XFILLER_106_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5103_ _5870_/A _5634_/D _5102_/X vssd1 vssd1 vccd1 vccd1 _5105_/B sky130_fd_sc_hd__a21o_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6083_ _6272_/CLK _6083_/D vssd1 vssd1 vccd1 vccd1 _6083_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3295_ _6200_/Q _3297_/B vssd1 vssd1 vccd1 vccd1 _3507_/A sky130_fd_sc_hd__nor2_1
XANTENNA__3224__A _5124_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5034_ _5034_/A _5034_/B vssd1 vssd1 vccd1 vccd1 _5034_/Y sky130_fd_sc_hd__nand2_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout176_A _4216_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3597__C _3607_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout343_A input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5936_ _5936_/A _5943_/A _5936_/C vssd1 vssd1 vccd1 vccd1 _5936_/X sky130_fd_sc_hd__or3_1
XANTENNA__4800__A1 _4625_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3603__A2 _3643_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5867_ _5867_/A1 _5865_/X _5866_/Y vssd1 vssd1 vccd1 vccd1 _6288_/D sky130_fd_sc_hd__a21oi_1
XANTENNA__3894__A _5622_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4818_ _5385_/A _4819_/B vssd1 vssd1 vccd1 vccd1 _4860_/B sky130_fd_sc_hd__nand2_2
X_5798_ _6264_/Q _3730_/X _5798_/S vssd1 vssd1 vccd1 vccd1 _6264_/D sky130_fd_sc_hd__mux2_1
XFILLER_21_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3367__B2 _4003_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4749_ _4782_/A _4791_/A vssd1 vssd1 vccd1 vccd1 _4755_/A sky130_fd_sc_hd__nand2_4
XFILLER_134_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput14 _6188_/Q vssd1 vssd1 vccd1 vccd1 io_out[12] sky130_fd_sc_hd__buf_4
XANTENNA__3118__B _5069_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput25 _6198_/Q vssd1 vssd1 vccd1 vccd1 io_out[22] sky130_fd_sc_hd__buf_4
XFILLER_122_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput36 _6184_/Q vssd1 vssd1 vccd1 vccd1 io_out[8] sky130_fd_sc_hd__buf_4
XFILLER_89_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5614__A _5653_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout89_A _3205_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5044__A1 _5051_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5044__B2 _4963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_331 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3044__A _5136_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3080_ _4046_/A _5227_/B vssd1 vssd1 vccd1 vccd1 _3080_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__4086__A2 _4311_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3979__A _5638_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5035__A1 _5034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5586__A2 _5454_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3982_ _5239_/A _3982_/B _3982_/C vssd1 vssd1 vccd1 vccd1 _3983_/C sky130_fd_sc_hd__and3_1
X_5721_ _5733_/A _5721_/B vssd1 vssd1 vccd1 vccd1 _5728_/C sky130_fd_sc_hd__nor2_1
XANTENNA__3918__S _3921_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5652_ _3251_/A _5728_/A _5651_/X _5932_/A vssd1 vssd1 vccd1 vccd1 _6234_/D sky130_fd_sc_hd__a211oi_1
XANTENNA__3349__A1 _3388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4603_ _4605_/D vssd1 vssd1 vccd1 vccd1 _4603_/Y sky130_fd_sc_hd__inv_2
XFILLER_129_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5583_ _6232_/Q _5583_/B vssd1 vssd1 vccd1 vccd1 _5602_/B sky130_fd_sc_hd__nand2_1
XANTENNA__3219__A _3869_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4534_ _4540_/A _6169_/Q vssd1 vssd1 vccd1 vccd1 _6168_/D sky130_fd_sc_hd__or2_1
XFILLER_7_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4465_ _5935_/A0 _4464_/X _4475_/S vssd1 vssd1 vccd1 vccd1 _6126_/D sky130_fd_sc_hd__mux2_1
XFILLER_116_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6204_ _6206_/CLK _6204_/D vssd1 vssd1 vccd1 vccd1 _6204_/Q sky130_fd_sc_hd__dfxtp_2
X_3416_ _3925_/A _3464_/B vssd1 vssd1 vccd1 vccd1 _3416_/Y sky130_fd_sc_hd__xnor2_1
X_4396_ _4424_/A _4424_/B vssd1 vssd1 vccd1 vccd1 _4399_/A sky130_fd_sc_hd__xor2_2
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6135_ _6284_/CLK _6135_/D vssd1 vssd1 vccd1 vccd1 _6135_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3347_ _3450_/A _3986_/A vssd1 vssd1 vccd1 vccd1 _3347_/Y sky130_fd_sc_hd__nor2_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6066_ _6290_/CLK _6066_/D vssd1 vssd1 vccd1 vccd1 _6066_/Q sky130_fd_sc_hd__dfxtp_4
X_3278_ _6280_/Q _6116_/Q _3551_/S vssd1 vssd1 vccd1 vccd1 _5450_/B sky130_fd_sc_hd__mux2_4
XFILLER_85_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5017_ _4638_/B _4640_/A _5016_/X _5013_/X _5403_/A vssd1 vssd1 vccd1 vccd1 _5017_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_73_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5919_ _5919_/A _5919_/B _5919_/C vssd1 vssd1 vccd1 vccd1 _5920_/D sky130_fd_sc_hd__and3_1
XFILLER_22_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4537__B1 _4540_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3760__A1 _4659_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5344__A _5344_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3815__A2 _3740_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5017__A1 _4638_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5017__B2 _5403_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3579__B2 _3312_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5238__B _5238_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5725__C1 _3179_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3039__A _4974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4250_ _5743_/C _4251_/B vssd1 vssd1 vccd1 vccd1 _4250_/Y sky130_fd_sc_hd__nor2_8
XFILLER_113_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3201_ _5936_/A _3706_/A _3324_/A vssd1 vssd1 vccd1 vccd1 _3255_/A sky130_fd_sc_hd__or3_4
XANTENNA__4700__A0 _4697_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4181_ _4181_/A _4181_/B _4181_/C vssd1 vssd1 vccd1 vccd1 _4185_/B sky130_fd_sc_hd__nand3_4
XFILLER_68_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3132_ _5119_/A _6007_/Q _3135_/S vssd1 vssd1 vccd1 vccd1 _6007_/D sky130_fd_sc_hd__mux2_1
X_3063_ _5162_/B _5258_/A vssd1 vssd1 vccd1 vccd1 _3111_/B sky130_fd_sc_hd__or2_4
XFILLER_94_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5008__A1 _5547_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3221__B _5360_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4740__A1_N _5703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3965_ _4638_/A _5928_/B vssd1 vssd1 vccd1 vccd1 _3965_/Y sky130_fd_sc_hd__nand2_2
XFILLER_50_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5704_ _3740_/A _4808_/B _5703_/X _5718_/A vssd1 vssd1 vccd1 vccd1 _5704_/X sky130_fd_sc_hd__a211o_1
XFILLER_31_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3896_ _5859_/A _3895_/X _4643_/A vssd1 vssd1 vccd1 vccd1 _3897_/B sky130_fd_sc_hd__mux2_1
XANTENNA_fanout139_A _5957_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4519__A0 _3942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3990__A1 _3942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5148__B _5241_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5635_ _5635_/A _5635_/B vssd1 vssd1 vccd1 vccd1 _5636_/B sky130_fd_sc_hd__nor2_1
XFILLER_128_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5566_ _5567_/A _5567_/B vssd1 vssd1 vccd1 vccd1 _5583_/B sky130_fd_sc_hd__and2_1
XANTENNA_fanout306_A _6066_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3891__B _4604_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4517_ _3942_/B _3912_/Y _4515_/X _4516_/X vssd1 vssd1 vccd1 vccd1 _6154_/D sky130_fd_sc_hd__a22o_1
X_5497_ _5504_/A _4965_/Y _5539_/S vssd1 vssd1 vccd1 vccd1 _5512_/B sky130_fd_sc_hd__mux2_2
XANTENNA_clkbuf_leaf_1_clk_A clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5164__A _5238_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4448_ _3942_/D _3900_/Y _4446_/X _4447_/Y vssd1 vssd1 vccd1 vccd1 _6120_/D sky130_fd_sc_hd__a22o_1
XANTENNA__5495__A1 _5058_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4379_ _4379_/A _4379_/B vssd1 vssd1 vccd1 vccd1 _4380_/B sky130_fd_sc_hd__nand2_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6118_ _6256_/CLK _6118_/D vssd1 vssd1 vccd1 vccd1 _6118_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5247__A1 _5158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6049_ _6260_/CLK _6049_/D vssd1 vssd1 vccd1 vccd1 _6049_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4758__B1 _4648_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3430__B1 _5924_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5058__B _5096_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5183__B1 _4946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3306__B _3575_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3249__B1 _3589_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3976__B _5096_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3468__S _3658_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5410__A1 _4586_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5410__B2 _5909_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3750_ _5617_/A _3750_/B _3750_/C vssd1 vssd1 vccd1 vccd1 _3816_/B sky130_fd_sc_hd__or3_4
XFILLER_9_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3681_ _5767_/A _3901_/B _5766_/C vssd1 vssd1 vccd1 vccd1 _3902_/A sky130_fd_sc_hd__or3_4
X_5420_ _6225_/Q _5420_/B vssd1 vssd1 vccd1 vccd1 _5421_/B sky130_fd_sc_hd__nor2_1
XFILLER_9_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5174__B1 _5494_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3724__A1 _6015_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5351_ _6176_/Q _4234_/B _4058_/B _6136_/Q _5350_/X vssd1 vssd1 vccd1 vccd1 _5351_/X
+ sky130_fd_sc_hd__o221a_2
XANTENNA__4600__B _4654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4302_ _4302_/A _4302_/B vssd1 vssd1 vccd1 vccd1 _4303_/C sky130_fd_sc_hd__xor2_2
X_5282_ _5929_/B2 _5280_/X _5281_/X _5279_/X vssd1 vssd1 vccd1 vccd1 _5283_/A sky130_fd_sc_hd__a31o_4
XANTENNA__5477__A1 _4974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4233_ _4233_/A1 _4231_/X _4232_/X vssd1 vssd1 vccd1 vccd1 _6086_/D sky130_fd_sc_hd__a21o_1
XANTENNA__3216__B _5653_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4164_ _4165_/A _4165_/B _4165_/C vssd1 vssd1 vccd1 vccd1 _4169_/A sky130_fd_sc_hd__a21o_1
XFILLER_114_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5229__A1 _5768_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3115_ _6216_/Q _3116_/B vssd1 vssd1 vccd1 vccd1 _3115_/Y sky130_fd_sc_hd__nor2_2
XFILLER_83_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4095_ _4084_/B _4093_/Y _4094_/X vssd1 vssd1 vccd1 vccd1 _4099_/A sky130_fd_sc_hd__a21o_2
XFILLER_95_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3232__A _5570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3046_ _5179_/A _4046_/A _3092_/B _5162_/B vssd1 vssd1 vccd1 vccd1 _3050_/B sky130_fd_sc_hd__or4b_4
XANTENNA__4047__B _4462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout256_A _6237_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3660__B1 _3881_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4997_ _4986_/X _4996_/Y _4721_/B vssd1 vssd1 vccd1 vccd1 _4997_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_11_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3948_ _3948_/A _5928_/B vssd1 vssd1 vccd1 vccd1 _4586_/B sky130_fd_sc_hd__nor2_8
XANTENNA__5952__A2 _5934_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3879_ _5095_/A _4587_/B vssd1 vssd1 vccd1 vccd1 _3879_/X sky130_fd_sc_hd__or2_4
XFILLER_109_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5618_ _5622_/A _4592_/B _3940_/A _5456_/S vssd1 vssd1 vccd1 vccd1 _5618_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5704__A2 _4808_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4079__A1_N _3783_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3715__A1 _6012_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5549_ _5567_/B _5548_/Y _5291_/Y vssd1 vssd1 vccd1 vccd1 _5549_/X sky130_fd_sc_hd__o21a_1
XFILLER_117_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5622__A _5622_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout71_A _3867_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5341__B _5341_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4238__A _5742_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5069__A _5069_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout60 _3793_/B vssd1 vssd1 vccd1 vccd1 _3841_/S sky130_fd_sc_hd__buf_6
XFILLER_80_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout71 _3867_/Y vssd1 vssd1 vccd1 vccd1 _3950_/C sky130_fd_sc_hd__buf_6
Xfanout82 _3102_/Y vssd1 vssd1 vccd1 vccd1 _5732_/C1 sky130_fd_sc_hd__clkbuf_4
Xfanout93 _5058_/A vssd1 vssd1 vccd1 vccd1 _5512_/A sky130_fd_sc_hd__buf_12
XFILLER_80_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3317__A _4003_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_551 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5678__S _5703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5631__A1 _5264_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3987__A _5712_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4920_ _5488_/A _4979_/B vssd1 vssd1 vccd1 vccd1 _4964_/A sky130_fd_sc_hd__nand2_1
XFILLER_61_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4851_ _4886_/B _4849_/Y _4850_/Y _3740_/A vssd1 vssd1 vccd1 vccd1 _4851_/X sky130_fd_sc_hd__o211a_1
X_3802_ _3800_/X _3801_/Y _3777_/S vssd1 vssd1 vccd1 vccd1 _3802_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__5395__B1 _5454_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4782_ _4782_/A _4782_/B vssd1 vssd1 vccd1 vccd1 _4782_/Y sky130_fd_sc_hd__nand2_2
XFILLER_14_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3733_ _3734_/A _3750_/C vssd1 vssd1 vccd1 vccd1 _3745_/C sky130_fd_sc_hd__nor2_1
X_3664_ _3563_/S _3641_/X _4883_/B _3210_/C _3210_/D vssd1 vssd1 vccd1 vccd1 _3664_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_109_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5403_ _5403_/A _5403_/B _5403_/C vssd1 vssd1 vccd1 vccd1 _5403_/X sky130_fd_sc_hd__or3_1
XANTENNA__5426__B _5428_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3595_ _3387_/A _3594_/A _3594_/B vssd1 vssd1 vccd1 vccd1 _3595_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_115_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5334_ _5387_/C _5334_/B vssd1 vssd1 vccd1 vccd1 _5354_/B sky130_fd_sc_hd__or2_4
XFILLER_88_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_17 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5265_ _5265_/A _5265_/B vssd1 vssd1 vccd1 vccd1 _5265_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__5442__A _5442_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4216_ _4216_/A _4216_/B _4216_/C vssd1 vssd1 vccd1 vccd1 _4218_/A sky130_fd_sc_hd__and3_2
XFILLER_102_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5196_ _6216_/Q _5197_/B vssd1 vssd1 vccd1 vccd1 _5202_/B sky130_fd_sc_hd__and2_1
XFILLER_29_827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4147_ _4148_/A _4148_/B vssd1 vssd1 vccd1 vccd1 _4181_/A sky130_fd_sc_hd__and2b_2
XANTENNA__4058__A _5436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4078_ _4084_/A _4076_/Y _4089_/A vssd1 vssd1 vccd1 vccd1 _4078_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_83_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3897__A _3964_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3029_ _4990_/A vssd1 vssd1 vccd1 vccd1 _3029_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_71_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_554 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5386__B1 _5387_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5617__A _5617_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5689__A1 _4767_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4897__C1 _4826_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3137__A _5800_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4361__A1 _3795_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4667__S _4806_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4113__A1 _4197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4113__B2 _4197_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout250 _6239_/Q vssd1 vssd1 vccd1 vccd1 _5859_/A sky130_fd_sc_hd__buf_6
Xfanout261 _5109_/A vssd1 vssd1 vccd1 vccd1 _5935_/A0 sky130_fd_sc_hd__buf_6
Xfanout272 _6229_/Q vssd1 vssd1 vccd1 vccd1 _5540_/B sky130_fd_sc_hd__buf_6
XFILLER_75_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout283 _6222_/Q vssd1 vssd1 vccd1 vccd1 _5333_/A sky130_fd_sc_hd__buf_8
Xfanout294 _5960_/C1 vssd1 vssd1 vccd1 vccd1 _5097_/A sky130_fd_sc_hd__buf_8
XFILLER_46_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_808 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5613__A1 _6233_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_4__f_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5916__A2 _5172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5527__A _5547_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3380_ _6074_/Q _5743_/B _3378_/X _3236_/Y _3379_/X vssd1 vssd1 vccd1 vccd1 _3380_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_108_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5262__A _5263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_41_clk_A clkbuf_3_4__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5301__A0 _5305_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5050_ _5072_/A _5050_/B _5050_/C vssd1 vssd1 vccd1 vccd1 _5052_/B sky130_fd_sc_hd__and3_1
XFILLER_111_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5852__A1 _3942_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4655__A2 _4872_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4001_ _3947_/X _3984_/X _3999_/X _4000_/Y vssd1 vssd1 vccd1 vccd1 _6057_/D sky130_fd_sc_hd__o31a_1
XFILLER_84_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_56_clk_A _6133_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5604__A1 _4638_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5952_ _3943_/A _5934_/A _3883_/X vssd1 vssd1 vccd1 vccd1 _5952_/X sky130_fd_sc_hd__a21o_1
XFILLER_52_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4903_ _4963_/A _4898_/X _4902_/X _4895_/Y vssd1 vssd1 vccd1 vccd1 _4903_/X sky130_fd_sc_hd__o211a_1
X_5883_ _5883_/A _5883_/B vssd1 vssd1 vccd1 vccd1 _5883_/X sky130_fd_sc_hd__and2_1
XFILLER_34_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4834_ _4832_/Y _4833_/X _4721_/B vssd1 vssd1 vccd1 vccd1 _4834_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_60_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3918__A1 _3721_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4765_ _4625_/A _5093_/A _4763_/X _4764_/X _5866_/B1 vssd1 vssd1 vccd1 vccd1 _6187_/D
+ sky130_fd_sc_hd__o311a_1
X_3716_ _6028_/Q _3715_/X _3731_/S vssd1 vssd1 vccd1 vccd1 _6028_/D sky130_fd_sc_hd__mux2_1
XANTENNA_fanout121_A _3450_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4696_ _4697_/A _4697_/B vssd1 vssd1 vccd1 vccd1 _4698_/A sky130_fd_sc_hd__or2_4
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3647_ _3541_/A _3642_/Y _3643_/Y _3611_/A _3646_/X vssd1 vssd1 vccd1 vccd1 _4877_/B
+ sky130_fd_sc_hd__o221a_4
XFILLER_20_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3578_ _6206_/Q _3567_/B _3658_/S vssd1 vssd1 vccd1 vccd1 _3578_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5317_ _6175_/Q _4234_/B _5349_/B1 _6135_/Q vssd1 vssd1 vccd1 vccd1 _5317_/X sky130_fd_sc_hd__o22a_1
XFILLER_102_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6297_ _6301_/CLK _6297_/D vssd1 vssd1 vccd1 vccd1 _6297_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5172__A _5172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5248_ _5248_/A _5248_/B _5248_/C _5248_/D vssd1 vssd1 vccd1 vccd1 _5249_/C sky130_fd_sc_hd__and4_1
XFILLER_102_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5179_ _5179_/A _5179_/B vssd1 vssd1 vccd1 vccd1 _5195_/C sky130_fd_sc_hd__and2_1
XFILLER_29_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5900__A _5900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5111__S _5129_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5359__A0 _3010_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3909__A1 _3730_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4251__A _5743_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4582__A1 _5605_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3385__A2 _3500_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5834__A1 _3666_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4426__A _4426_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3968__C _5227_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output15_A _6189_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3376__A2 _3375_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4573__A1 _5238_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4550_ _6176_/Q _4553_/B vssd1 vssd1 vccd1 vccd1 _4550_/X sky130_fd_sc_hd__or2_1
XFILLER_128_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3501_ _3801_/A _3500_/B _3458_/B _3513_/B vssd1 vssd1 vccd1 vccd1 _3502_/B sky130_fd_sc_hd__a31o_1
XFILLER_116_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4481_ _6134_/Q _4499_/B vssd1 vssd1 vccd1 vccd1 _4481_/X sky130_fd_sc_hd__or2_1
XFILLER_7_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6220_ _6232_/CLK _6220_/D vssd1 vssd1 vccd1 vccd1 _6220_/Q sky130_fd_sc_hd__dfxtp_2
X_3432_ _3432_/A vssd1 vssd1 vccd1 vccd1 _3432_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3208__C _3741_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3533__C1 _5470_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6151_ _6154_/CLK _6151_/D vssd1 vssd1 vccd1 vccd1 _6151_/Q sky130_fd_sc_hd__dfxtp_1
X_3363_ _3285_/Y _3316_/B _3303_/X vssd1 vssd1 vccd1 vccd1 _3364_/B sky130_fd_sc_hd__o21bai_4
XFILLER_124_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5102_ _5957_/B _3869_/B _5634_/B _3741_/B vssd1 vssd1 vccd1 vccd1 _5102_/X sky130_fd_sc_hd__a31o_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6082_ _6274_/CLK _6082_/D vssd1 vssd1 vccd1 vccd1 _6082_/Q sky130_fd_sc_hd__dfxtp_1
X_3294_ _3563_/S _4659_/B _3289_/X _3227_/X vssd1 vssd1 vccd1 vccd1 _3294_/X sky130_fd_sc_hd__a211o_1
XFILLER_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5825__A1 _3425_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3224__B _3706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5033_ _5040_/A _5033_/B vssd1 vssd1 vccd1 vccd1 _5034_/B sky130_fd_sc_hd__xnor2_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3300__A2 _4665_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4336__A _4362_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5589__B1 _3122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout169_A _3901_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5935_ _5935_/A0 _3242_/X _5943_/B vssd1 vssd1 vccd1 vccd1 _5936_/C sky130_fd_sc_hd__mux2_1
XFILLER_22_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4800__A2 _5093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4770__S _4806_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5866_ _6288_/Q _5867_/A1 _5866_/B1 vssd1 vssd1 vccd1 vccd1 _5866_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout336_A _4819_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3894__B _3975_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4817_ _4745_/A _4813_/X _4824_/B _4744_/B _5034_/A vssd1 vssd1 vccd1 vccd1 _4817_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4013__B1 _3615_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5797_ _6263_/Q _3727_/X _5798_/S vssd1 vssd1 vccd1 vccd1 _6263_/D sky130_fd_sc_hd__mux2_1
XFILLER_31_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5761__A0 _5446_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4564__A1 _5790_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4748_ _5333_/A _5344_/A vssd1 vssd1 vccd1 vccd1 _4791_/A sky130_fd_sc_hd__nand2_4
X_4679_ _6185_/Q _4678_/Y _5041_/S vssd1 vssd1 vccd1 vccd1 _4679_/X sky130_fd_sc_hd__mux2_1
XFILLER_134_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput15 _6189_/Q vssd1 vssd1 vccd1 vccd1 io_out[13] sky130_fd_sc_hd__buf_4
Xoutput26 _6181_/Q vssd1 vssd1 vccd1 vccd1 io_out[23] sky130_fd_sc_hd__buf_4
Xoutput37 _6185_/Q vssd1 vssd1 vccd1 vccd1 io_out[9] sky130_fd_sc_hd__buf_4
XFILLER_122_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5614__B _5889_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5106__S _5124_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5816__A1 _3666_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3150__A _4622_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4680__S _5054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_51_clk _6133_/CLK vssd1 vssd1 vccd1 vccd1 _6177_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_24_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_663 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4004__B1 _3033_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5201__C1 _5071_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4555__A1 _5856_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5016__S _5041_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3530__A2 _3529_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5807__A1 _5835_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3044__B _3958_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5540__A _6230_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3060__A _3060_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3981_ _3114_/C _5617_/C _5206_/B _3981_/D vssd1 vssd1 vccd1 vccd1 _3982_/C sky130_fd_sc_hd__and4b_1
XANTENNA__3995__A _5883_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5720_ _5718_/A _5719_/X _5718_/Y _5732_/C1 vssd1 vssd1 vccd1 vccd1 _5728_/B sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_42_clk clkbuf_3_4__f_clk/X vssd1 vssd1 vccd1 vccd1 _6259_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5651_ _5733_/A _4620_/A _5650_/X vssd1 vssd1 vccd1 vccd1 _5651_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__4546__A1 _5935_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4602_ _5075_/B _3123_/A _5097_/A vssd1 vssd1 vccd1 vccd1 _4605_/D sky130_fd_sc_hd__a21oi_2
X_5582_ _6232_/Q _5583_/B vssd1 vssd1 vccd1 vccd1 _5582_/X sky130_fd_sc_hd__or2_1
XFILLER_129_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3219__B _5818_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4533_ _6157_/Q _6168_/Q _4532_/Y vssd1 vssd1 vccd1 vccd1 _6167_/D sky130_fd_sc_hd__o21a_1
XFILLER_8_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4464_ _4672_/A _6126_/Q _4476_/S vssd1 vssd1 vccd1 vccd1 _4464_/X sky130_fd_sc_hd__mux2_1
XFILLER_104_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6203_ _6206_/CLK _6203_/D vssd1 vssd1 vccd1 vccd1 _6203_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_132_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3415_ _3935_/B _3364_/B _3358_/A vssd1 vssd1 vccd1 vccd1 _3464_/B sky130_fd_sc_hd__a21oi_2
XFILLER_131_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4395_ _4393_/B _4368_/B _4370_/B _4371_/B _4371_/A vssd1 vssd1 vccd1 vccd1 _4424_/B
+ sky130_fd_sc_hd__o32a_4
XANTENNA__3235__A _3241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6134_ _6179_/CLK _6134_/D vssd1 vssd1 vccd1 vccd1 _6134_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3346_ _3266_/A _3266_/B _3274_/A _3274_/B vssd1 vssd1 vccd1 vccd1 _3500_/B sky130_fd_sc_hd__o22a_4
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6065_ _6093_/CLK _6065_/D vssd1 vssd1 vccd1 vccd1 _6065_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3277_ _6292_/Q _6298_/Q vssd1 vssd1 vccd1 vccd1 _3316_/A sky130_fd_sc_hd__nand2b_2
XANTENNA__5450__A _5599_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout286_A _5768_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5016_ _6195_/Q _5015_/Y _5041_/S vssd1 vssd1 vccd1 vccd1 _5016_/X sky130_fd_sc_hd__mux2_1
XFILLER_85_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5431__C1 _3059_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3588__A2 _5439_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5918_ _5870_/A _3883_/X _5914_/X _5917_/X vssd1 vssd1 vccd1 vccd1 _5919_/C sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_33_clk clkbuf_3_5__f_clk/X vssd1 vssd1 vccd1 vccd1 _6144_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_42_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_140 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5849_ _5849_/A vssd1 vssd1 vccd1 vccd1 _5850_/B sky130_fd_sc_hd__inv_2
XFILLER_10_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5625__A _5625_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3760__A2 _3740_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5344__B _5653_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4473__A0 _3942_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5017__A2 _4640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4776__B2 _4946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_24_clk _6233_/CLK vssd1 vssd1 vccd1 vccd1 _6041_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_60_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5238__C _5238_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5725__B1 _3597_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3981__C _5206_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3055__A _5075_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3200_ _3765_/B _4604_/C vssd1 vssd1 vccd1 vccd1 _3772_/B sky130_fd_sc_hd__nand2_8
XFILLER_79_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4180_ _4180_/A _4180_/B _4180_/C vssd1 vssd1 vccd1 vccd1 _4181_/C sky130_fd_sc_hd__nand3_4
XFILLER_79_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3131_ _5344_/A _6006_/Q _3135_/S vssd1 vssd1 vccd1 vccd1 _6006_/D sky130_fd_sc_hd__mux2_1
XANTENNA__3205__D _3706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3062_ _5162_/B _3072_/A vssd1 vssd1 vccd1 vccd1 _3062_/Y sky130_fd_sc_hd__nor2_2
XANTENNA__4464__A0 _4672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5661__C1 _3974_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5008__A2 _5029_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3221__C _5617_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5413__C1 _5251_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4614__A _4614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3964_ _5911_/A _3964_/B vssd1 vssd1 vccd1 vccd1 _5909_/B sky130_fd_sc_hd__nor2_8
XANTENNA__5964__B1 _3766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_15_clk _6233_/CLK vssd1 vssd1 vccd1 vccd1 _6206_/CLK sky130_fd_sc_hd__clkbuf_16
X_5703_ _5703_/A _5703_/B vssd1 vssd1 vccd1 vccd1 _5703_/X sky130_fd_sc_hd__and2_1
XFILLER_50_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3895_ _6042_/Q _5934_/B _4819_/B vssd1 vssd1 vccd1 vccd1 _3895_/X sky130_fd_sc_hd__mux2_1
X_5634_ _5634_/A _5634_/B _5634_/C _5634_/D vssd1 vssd1 vccd1 vccd1 _5635_/B sky130_fd_sc_hd__or4_1
XFILLER_136_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5565_ _3059_/Y _5560_/Y _5564_/Y vssd1 vssd1 vccd1 vccd1 _5565_/Y sky130_fd_sc_hd__a21oi_1
X_4516_ _5385_/A _4520_/S _4521_/S vssd1 vssd1 vccd1 vccd1 _4516_/X sky130_fd_sc_hd__o21a_1
XANTENNA__3891__C _5928_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout201_A _3869_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5496_ _5488_/A _5556_/A2 _5495_/X _5556_/C1 vssd1 vssd1 vccd1 vccd1 _6227_/D sky130_fd_sc_hd__o211a_1
XFILLER_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4447_ _3011_/Y _4458_/B _3900_/Y vssd1 vssd1 vccd1 vccd1 _4447_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_132_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5495__A2 _5482_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4378_ _4379_/A _4379_/B vssd1 vssd1 vccd1 vccd1 _4401_/A sky130_fd_sc_hd__or2_1
XFILLER_98_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6117_ _6250_/CLK _6117_/D vssd1 vssd1 vccd1 vccd1 _6117_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input6_A io_in[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3329_ _6259_/Q _6051_/Q _6044_/Q _6028_/Q _3241_/A _3241_/B vssd1 vssd1 vccd1 vccd1
+ _3329_/X sky130_fd_sc_hd__mux4_2
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5247__A2 _4577_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6048_ _6262_/CLK _6048_/D vssd1 vssd1 vccd1 vccd1 _6048_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5652__C1 _5932_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4524__A _4539_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4758__B2 _5344_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5058__C _5058_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5183__A1 _5054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5090__A _5090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3680_ _3678_/X _3679_/X _4462_/A vssd1 vssd1 vccd1 vccd1 _5766_/C sky130_fd_sc_hd__a21o_4
XFILLER_127_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5350_ _6152_/Q _3243_/A _5767_/B _6128_/Q vssd1 vssd1 vccd1 vccd1 _5350_/X sky130_fd_sc_hd__o22a_1
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4301_ _4301_/A _4410_/D vssd1 vssd1 vccd1 vccd1 _4302_/B sky130_fd_sc_hd__nand2_2
X_5281_ _6118_/Q _3901_/B _3704_/B _6020_/Q vssd1 vssd1 vccd1 vccd1 _5281_/X sky130_fd_sc_hd__o22a_1
XFILLER_114_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4232_ _3853_/X _4071_/A _4072_/C _6086_/Q vssd1 vssd1 vccd1 vccd1 _4232_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3216__C _4806_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_4_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _6007_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_101_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4163_ _4163_/A _4311_/B vssd1 vssd1 vccd1 vccd1 _4165_/C sky130_fd_sc_hd__and2_1
XFILLER_68_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5229__A2 _5227_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3114_ _5096_/C _3114_/B _3114_/C vssd1 vssd1 vccd1 vccd1 _3127_/A sky130_fd_sc_hd__or3_2
X_4094_ _4162_/A _4162_/B _4216_/B _4214_/B vssd1 vssd1 vccd1 vccd1 _4094_/X sky130_fd_sc_hd__and4_1
XANTENNA__3232__B _5734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3045_ _6217_/Q _6216_/Q _6215_/Q _6214_/Q vssd1 vssd1 vccd1 vccd1 _3107_/A sky130_fd_sc_hd__or4_4
XFILLER_71_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3660__A1 _4003_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5937__B1 _5110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout151_A _5476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4996_ _5547_/B _4872_/B _4991_/X _4995_/X vssd1 vssd1 vccd1 vccd1 _4996_/Y sky130_fd_sc_hd__o22ai_1
XANTENNA_fanout249_A _5859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3947_ _3936_/X _3940_/Y _3946_/X _3941_/A vssd1 vssd1 vccd1 vccd1 _3947_/X sky130_fd_sc_hd__o211a_1
X_3878_ _3878_/A _4608_/C vssd1 vssd1 vccd1 vccd1 _5692_/B sky130_fd_sc_hd__nand2_2
X_5617_ _5617_/A _5617_/B _5617_/C vssd1 vssd1 vccd1 vccd1 _5617_/X sky130_fd_sc_hd__or3_1
XANTENNA__3394__S _3709_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5548_ _5540_/B _5547_/C _5547_/A vssd1 vssd1 vccd1 vccd1 _5548_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_3_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5479_ _3009_/Y _4934_/X _5539_/S vssd1 vssd1 vccd1 vccd1 _5491_/B sky130_fd_sc_hd__mux2_2
XFILLER_133_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5468__A2 _4234_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3884__D1 _4604_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout64_A _4638_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3142__B _6070_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout50 _4237_/Y vssd1 vssd1 vccd1 vccd1 _4564_/A2 sky130_fd_sc_hd__buf_4
Xfanout61 _3253_/Y vssd1 vssd1 vccd1 vccd1 _5835_/A1 sky130_fd_sc_hd__buf_4
XANTENNA__3403__B2 _3986_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout72 _3678_/B vssd1 vssd1 vccd1 vccd1 _5607_/B1 sky130_fd_sc_hd__clkbuf_8
Xfanout83 _5731_/S vssd1 vssd1 vccd1 vccd1 _5703_/A sky130_fd_sc_hd__buf_6
Xfanout94 _3079_/Y vssd1 vssd1 vccd1 vccd1 _5058_/A sky130_fd_sc_hd__buf_4
XFILLER_10_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_82 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5085__A _5093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4903__A1 _4963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3317__B _4003_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4667__A0 _5263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5864__C1 _5866_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5616__C1 _4753_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3052__B _3970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5092__B1 _4931_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_7__f_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _6084_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_563 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5631__A2 _3179_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3987__B _3987_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_0_clk_A _6133_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4850_ _4850_/A _4886_/B vssd1 vssd1 vccd1 vccd1 _4850_/Y sky130_fd_sc_hd__nand2_1
XFILLER_60_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3801_ _3801_/A _3801_/B vssd1 vssd1 vccd1 vccd1 _3801_/Y sky130_fd_sc_hd__nor2_1
X_4781_ _4860_/A _4781_/B vssd1 vssd1 vccd1 vccd1 _4791_/B sky130_fd_sc_hd__nand2_2
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3732_ _3732_/A _5936_/A vssd1 vssd1 vccd1 vccd1 _3769_/D sky130_fd_sc_hd__nor2_1
XANTENNA__5707__B _5707_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3663_ _3511_/A _3931_/B _3661_/Y _3662_/X vssd1 vssd1 vccd1 vccd1 _5900_/A sky130_fd_sc_hd__o22a_4
X_5402_ _5507_/A _5401_/X _5389_/Y _5310_/Y vssd1 vssd1 vccd1 vccd1 _5403_/C sky130_fd_sc_hd__a2bb2o_1
X_3594_ _3594_/A _3594_/B vssd1 vssd1 vccd1 vccd1 _3606_/B sky130_fd_sc_hd__nor2_1
XFILLER_127_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3227__B _4592_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5333_ _5333_/A _5333_/B vssd1 vssd1 vccd1 vccd1 _5334_/B sky130_fd_sc_hd__nor2_1
XFILLER_88_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5264_ _5264_/A _5264_/B vssd1 vssd1 vccd1 vccd1 _5265_/B sky130_fd_sc_hd__nand2_2
XFILLER_125_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5442__B _5442_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5855__C1 _5866_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4215_ _4215_/A _4215_/B vssd1 vssd1 vccd1 vccd1 _4216_/C sky130_fd_sc_hd__xnor2_1
XFILLER_130_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5195_ _6215_/Q _6214_/Q _5195_/C vssd1 vssd1 vccd1 vccd1 _5197_/B sky130_fd_sc_hd__and3_1
XANTENNA__3243__A _3243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout199_A _3922_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4146_ _4146_/A _4146_/B vssd1 vssd1 vccd1 vccd1 _4148_/B sky130_fd_sc_hd__xnor2_4
XFILLER_29_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4058__B _4058_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4077_ _4197_/A _4136_/A _4173_/B _4176_/B vssd1 vssd1 vccd1 vccd1 _4089_/A sky130_fd_sc_hd__and4_1
XFILLER_37_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3028_ _4540_/A vssd1 vssd1 vccd1 vccd1 _3028_/Y sky130_fd_sc_hd__inv_4
XFILLER_55_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3633__A1 _4216_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4979_ _5547_/B _4979_/B vssd1 vssd1 vccd1 vccd1 _4980_/B sky130_fd_sc_hd__or2_1
XANTENNA__3397__B1 _5341_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4802__A _5392_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5617__B _5617_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4897__B1 _4648_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3137__B _3869_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4113__A2 _4112_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4249__A _5767_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout240 _4216_/A vssd1 vssd1 vccd1 vccd1 _4426_/A sky130_fd_sc_hd__buf_6
Xfanout251 _6238_/Q vssd1 vssd1 vccd1 vccd1 _5856_/A sky130_fd_sc_hd__buf_6
Xfanout262 _4096_/A vssd1 vssd1 vccd1 vccd1 _4197_/A sky130_fd_sc_hd__buf_6
XFILLER_115_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout273 _6228_/Q vssd1 vssd1 vccd1 vccd1 _5504_/A sky130_fd_sc_hd__clkbuf_16
XANTENNA__5861__A2 _5867_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout284 _6220_/Q vssd1 vssd1 vccd1 vccd1 _4672_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_75_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout295 _5960_/C1 vssd1 vssd1 vccd1 vccd1 _3014_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_86_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5613__A2 _5250_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3624__A1 _3615_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5916__A3 _3678_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4585__C1 _5192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3483__S0 _3241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5262__B _5263_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4000_ _3021_/Y _3984_/X _5932_/A vssd1 vssd1 vccd1 vccd1 _4000_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_77_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5689__S _5703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3998__A _5226_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5951_ _5951_/A _5951_/B _5951_/C vssd1 vssd1 vccd1 vccd1 _5955_/B sky130_fd_sc_hd__nand3_2
XFILLER_46_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4812__A0 _5714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4902_ _6191_/Q _5561_/S _5239_/A _4901_/X vssd1 vssd1 vccd1 vccd1 _4902_/X sky130_fd_sc_hd__a211o_1
XFILLER_34_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5882_ _3615_/B _5881_/X _5882_/S vssd1 vssd1 vccd1 vccd1 _5883_/B sky130_fd_sc_hd__mux2_1
X_4833_ _5385_/A _4872_/B _4823_/X _5069_/A vssd1 vssd1 vccd1 vccd1 _4833_/X sky130_fd_sc_hd__a2bb2o_1
XANTENNA__3379__B1 _3589_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4622__A _5625_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4764_ _6187_/Q _4970_/B vssd1 vssd1 vccd1 vccd1 _4764_/X sky130_fd_sc_hd__or2_1
XANTENNA__4040__A1 _3718_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3715_ _6012_/Q _3706_/Y _3714_/X vssd1 vssd1 vccd1 vccd1 _3715_/X sky130_fd_sc_hd__a21o_4
XFILLER_119_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4695_ _4660_/A _4660_/B _4657_/X vssd1 vssd1 vccd1 vccd1 _4699_/A sky130_fd_sc_hd__a21o_1
XANTENNA__3238__A _5924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3646_ _3986_/B _3646_/B vssd1 vssd1 vccd1 vccd1 _3646_/X sky130_fd_sc_hd__or2_1
X_3577_ _3658_/S _3567_/B _3575_/X vssd1 vssd1 vccd1 vccd1 _5888_/A sky130_fd_sc_hd__o21ai_1
X_5316_ _5436_/A _6151_/Q _5436_/C vssd1 vssd1 vccd1 vccd1 _5316_/X sky130_fd_sc_hd__and3_1
XFILLER_0_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6296_ _6301_/CLK _6296_/D vssd1 vssd1 vccd1 vccd1 _6296_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5172__B _5172_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5247_ _5158_/A _4577_/C _3865_/Y _3879_/X vssd1 vssd1 vccd1 vccd1 _5248_/D sky130_fd_sc_hd__a211o_1
XFILLER_29_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5843__A2 _5841_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5178_ _5179_/A _5179_/B vssd1 vssd1 vccd1 vccd1 _5180_/A sky130_fd_sc_hd__nor2_1
XANTENNA__3854__A1 _5128_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4129_ _4437_/A1 _4127_/Y _4128_/X vssd1 vssd1 vccd1 vccd1 _6083_/D sky130_fd_sc_hd__a21o_1
XFILLER_84_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4251__B _4251_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4582__A2 _3996_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3148__A _3880_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4707__A _6221_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4426__B _4426_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3058__A _5218_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3500_ _3500_/A _3500_/B _3500_/C _3513_/B vssd1 vssd1 vccd1 vccd1 _3593_/B sky130_fd_sc_hd__and4_2
XFILLER_128_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4480_ _3943_/C _4057_/Y _4478_/X _4479_/Y vssd1 vssd1 vccd1 vccd1 _6133_/D sky130_fd_sc_hd__a22o_1
XFILLER_7_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3431_ _5470_/S _3428_/X _3430_/X vssd1 vssd1 vccd1 vccd1 _3432_/A sky130_fd_sc_hd__a21oi_4
XANTENNA__3208__D _4886_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3533__B1 _3704_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6150_ _6155_/CLK _6150_/D vssd1 vssd1 vccd1 vccd1 _6150_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3362_ _3360_/X _3361_/Y _3621_/A vssd1 vssd1 vccd1 vccd1 _3362_/X sky130_fd_sc_hd__a21o_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5101_ _3296_/A _5097_/X _5100_/Y _5192_/A vssd1 vssd1 vccd1 vccd1 _6200_/D sky130_fd_sc_hd__a211oi_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6081_ _6272_/CLK _6081_/D vssd1 vssd1 vccd1 vccd1 _6081_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3293_ _4010_/B _3644_/B vssd1 vssd1 vccd1 vccd1 _4659_/B sky130_fd_sc_hd__xnor2_4
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5032_ _4981_/A _4983_/X _5015_/A _5031_/Y vssd1 vssd1 vccd1 vccd1 _5033_/B sky130_fd_sc_hd__o31a_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3836__A1 _3643_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5589__A1 _5512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4336__B _4389_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3240__B _3241_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5934_ _5934_/A _5934_/B vssd1 vssd1 vccd1 vccd1 _5985_/B sky130_fd_sc_hd__nor2_1
XANTENNA__4261__A1 _4216_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5865_ _3649_/B _3944_/A _5865_/S vssd1 vssd1 vccd1 vccd1 _5865_/X sky130_fd_sc_hd__mux2_8
XFILLER_33_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5448__A _5480_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4816_ _4854_/B _4816_/B vssd1 vssd1 vccd1 vccd1 _4824_/B sky130_fd_sc_hd__or2_1
XANTENNA_fanout231_A _5625_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5796_ _6262_/Q _3724_/X _5798_/S vssd1 vssd1 vccd1 vccd1 _6262_/D sky130_fd_sc_hd__mux2_1
XANTENNA_fanout329_A _5599_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4013__B2 _4850_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4747_ _5333_/A _5344_/A vssd1 vssd1 vccd1 vccd1 _4782_/A sky130_fd_sc_hd__or2_4
XANTENNA__4071__B _4296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4678_ _4678_/A _4678_/B vssd1 vssd1 vccd1 vccd1 _4678_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_107_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3629_ _3511_/A _3923_/A _3628_/X vssd1 vssd1 vccd1 vccd1 _5898_/B sky130_fd_sc_hd__o21a_4
Xoutput16 _6190_/Q vssd1 vssd1 vccd1 vccd1 io_out[14] sky130_fd_sc_hd__buf_4
Xoutput27 _6183_/Q vssd1 vssd1 vccd1 vccd1 io_out[24] sky130_fd_sc_hd__buf_4
XFILLER_88_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6279_ _6279_/CLK _6279_/D vssd1 vssd1 vccd1 vccd1 _6279_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5911__A _5911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3827__A1 _4808_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4527__A _4540_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3150__B _3970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5160__A2_N _3105_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5358__A _5358_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_40_clk_A clkbuf_3_4__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4004__A1 _6292_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4004__B2 _6298_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5792__S _5798_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4960__C1 _4826_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_55_clk_A _6133_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5093__A _5093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5268__A0 _4672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3818__A1 _3937_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5540__B _5540_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4491__A1 _3010_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3294__A2 _4659_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3060__B _3060_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3980_ _5634_/A _3980_/B _5634_/B _5634_/D vssd1 vssd1 vccd1 vccd1 _3981_/D sky130_fd_sc_hd__or4_1
XFILLER_16_661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4243__A1 _3721_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5440__B1 _3704_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clkbuf_0_clk/X sky130_fd_sc_hd__clkbuf_16
X_5650_ _3388_/A _5203_/A _5616_/X _5631_/X _5728_/A vssd1 vssd1 vccd1 vccd1 _5650_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4601_ _5090_/A _5069_/A vssd1 vssd1 vccd1 vccd1 _4601_/Y sky130_fd_sc_hd__nand2_4
XFILLER_129_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5581_ _3536_/X _5909_/B _5580_/Y _4586_/B vssd1 vssd1 vccd1 vccd1 _5581_/X sky130_fd_sc_hd__a22o_1
X_4532_ _6157_/Q _6168_/Q _4540_/A vssd1 vssd1 vccd1 vccd1 _4532_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4463_ _3943_/C _4461_/X _4475_/S vssd1 vssd1 vccd1 vccd1 _6125_/D sky130_fd_sc_hd__mux2_1
XANTENNA__5207__S _5207_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6202_ _6234_/CLK _6202_/D vssd1 vssd1 vccd1 vccd1 _6202_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_131_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3414_ _3925_/A _3414_/B vssd1 vssd1 vccd1 vccd1 _3414_/Y sky130_fd_sc_hd__xnor2_1
X_4394_ _4394_/A _4394_/B vssd1 vssd1 vccd1 vccd1 _4424_/A sky130_fd_sc_hd__nand2_2
XFILLER_131_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3235__B _3241_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6133_ _6133_/CLK _6133_/D vssd1 vssd1 vccd1 vccd1 _6133_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3345_ _4096_/A _3560_/S _3344_/X vssd1 vssd1 vccd1 vccd1 _3345_/X sky130_fd_sc_hd__a21o_1
XFILLER_97_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6064_ _6264_/CLK _6064_/D vssd1 vssd1 vccd1 vccd1 _6064_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3276_ _3398_/A _3986_/A _3275_/X _3498_/S vssd1 vssd1 vccd1 vccd1 _3276_/X sky130_fd_sc_hd__o211a_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5015_ _5015_/A _5015_/B vssd1 vssd1 vccd1 vccd1 _5015_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__5450__B _5450_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout181_A _3488_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4482__A1 _4672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3251__A _3251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5917_ _4577_/A _3950_/C _5172_/B _5058_/D _5916_/Y vssd1 vssd1 vccd1 vccd1 _5917_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__4082__A _4162_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5848_ _5848_/A0 _5926_/A0 _5862_/B vssd1 vssd1 vccd1 vccd1 _5849_/A sky130_fd_sc_hd__mux2_8
XFILLER_21_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5779_ _6254_/Q _5788_/B vssd1 vssd1 vccd1 vccd1 _5779_/X sky130_fd_sc_hd__or2_1
XFILLER_5_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3145__B _5883_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3276__A2 _3986_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3161__A _4642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5670__B1 _3950_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5422__A0 _6009_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5489__B1 _5607_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3055__B _4003_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4161__B1 _4342_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5551__A _5551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3130_ _4707_/B _6005_/Q _3135_/S vssd1 vssd1 vccd1 vccd1 _6005_/D sky130_fd_sc_hd__mux2_1
XFILLER_94_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4167__A _4197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3061_ _3107_/A _5179_/A _3092_/B vssd1 vssd1 vccd1 vccd1 _3072_/A sky130_fd_sc_hd__or3b_4
XFILLER_48_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5697__S _5712_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3963_ _4604_/A _3978_/B vssd1 vssd1 vccd1 vccd1 _5640_/B sky130_fd_sc_hd__or2_4
XFILLER_50_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4614__B _4614_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5702_ _4163_/A _5649_/X _5701_/X _5956_/A vssd1 vssd1 vccd1 vccd1 _6238_/D sky130_fd_sc_hd__o211a_1
X_3894_ _5622_/A _3975_/C vssd1 vssd1 vccd1 vccd1 _5934_/B sky130_fd_sc_hd__or2_4
XFILLER_137_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5633_ _6217_/Q _5065_/A _4744_/B _5097_/A vssd1 vssd1 vccd1 vccd1 _5838_/B sky130_fd_sc_hd__a31o_2
XANTENNA__5716__A1 _3593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5564_ _5072_/B _5561_/X _5563_/X vssd1 vssd1 vccd1 vccd1 _5564_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_117_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4515_ _6154_/Q _4515_/B vssd1 vssd1 vccd1 vccd1 _4515_/X sky130_fd_sc_hd__or2_1
X_5495_ _5058_/C _5482_/Y _5490_/X _5494_/X _5251_/Y vssd1 vssd1 vccd1 vccd1 _5495_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_132_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4446_ _6120_/Q _4458_/B vssd1 vssd1 vccd1 vccd1 _4446_/X sky130_fd_sc_hd__or2_1
XFILLER_104_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4377_ _4348_/B _4350_/B _4348_/A vssd1 vssd1 vccd1 vccd1 _4379_/B sky130_fd_sc_hd__o21ba_1
XFILLER_98_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6116_ _6280_/CLK _6116_/D vssd1 vssd1 vccd1 vccd1 _6116_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3328_ _6073_/Q _5743_/B _3326_/X _3236_/Y _3327_/X vssd1 vssd1 vccd1 vccd1 _3328_/X
+ sky130_fd_sc_hd__o221a_2
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6047_ _6295_/CLK _6047_/D vssd1 vssd1 vccd1 vccd1 _6047_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5101__C1 _5192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3259_ _6265_/Q _6011_/Q _6079_/Q _6034_/Q _4067_/A _3709_/S vssd1 vssd1 vccd1 vccd1
+ _3259_/X sky130_fd_sc_hd__mux4_2
XANTENNA__4077__A _4197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3290__A_N _6009_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4758__A2 _4647_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3430__A2 _5439_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4540__A _4540_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5183__A2 _5143_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3156__A _5840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4694__A1 _4707_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3497__A2 _3593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3249__A2 _3589_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_778 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5946__B2 _4586_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3709__A0 _6011_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4906__C1 _5071_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4300_ _4301_/A _4426_/B vssd1 vssd1 vccd1 vccd1 _4335_/A sky130_fd_sc_hd__nand2_1
XFILLER_5_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5280_ _6251_/Q _3243_/A _5742_/B _6243_/Q vssd1 vssd1 vccd1 vccd1 _5280_/X sky130_fd_sc_hd__o22a_1
XFILLER_99_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4231_ _4231_/A _4231_/B vssd1 vssd1 vccd1 vccd1 _4231_/X sky130_fd_sc_hd__xor2_2
XANTENNA__5331__C1 _3121_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5882__A0 _3615_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4685__B2 _5069_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4162_ _4162_/A _4162_/B _4309_/B _4342_/B vssd1 vssd1 vccd1 vccd1 _4165_/B sky130_fd_sc_hd__nand4_4
XFILLER_68_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3113_ _5069_/A _4605_/A vssd1 vssd1 vccd1 vccd1 _3114_/C sky130_fd_sc_hd__nand2_1
XANTENNA__3513__B _3513_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4093_ _4162_/A _4216_/B vssd1 vssd1 vccd1 vccd1 _4093_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__4437__A1 _4437_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3044_ _5136_/C _3958_/A vssd1 vssd1 vccd1 vccd1 _3044_/Y sky130_fd_sc_hd__nand2_1
XFILLER_36_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4625__A _4625_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5220__S _5220_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5937__A1 _5503_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5398__C1 _4646_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4995_ _5547_/B _4644_/A _4994_/X _5072_/C _5058_/C vssd1 vssd1 vccd1 vccd1 _4995_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_23_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout144_A _5075_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3946_ _3649_/B _3643_/B _5634_/B _3945_/Y _5124_/S vssd1 vssd1 vccd1 vccd1 _3946_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_32_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3877_ _5976_/A _3877_/B vssd1 vssd1 vccd1 vccd1 _4615_/A sky130_fd_sc_hd__nor2_4
XFILLER_137_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout311_A _5561_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5616_ _5454_/B _5615_/X _5614_/X _4753_/A vssd1 vssd1 vccd1 vccd1 _5616_/X sky130_fd_sc_hd__o211a_1
X_5547_ _5547_/A _5547_/B _5547_/C vssd1 vssd1 vccd1 vccd1 _5567_/B sky130_fd_sc_hd__and3_1
X_5478_ _4974_/A _5476_/Y _5477_/Y vssd1 vssd1 vccd1 vccd1 _5478_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_132_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5322__C1 _5595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4429_ _4429_/A _4429_/B vssd1 vssd1 vccd1 vccd1 _4431_/C sky130_fd_sc_hd__xnor2_1
XFILLER_133_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3704__A _5767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5191__A _5191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3939__B1 _5900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout40 _4625_/Y vssd1 vssd1 vccd1 vccd1 _4970_/B sky130_fd_sc_hd__buf_2
Xfanout51 _4057_/Y vssd1 vssd1 vccd1 vccd1 _4501_/A2 sky130_fd_sc_hd__buf_4
XFILLER_120_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout62 _3253_/Y vssd1 vssd1 vccd1 vccd1 _5817_/A1 sky130_fd_sc_hd__buf_2
Xfanout73 _3195_/X vssd1 vssd1 vccd1 vccd1 _5734_/A sky130_fd_sc_hd__buf_6
Xfanout84 _3091_/Y vssd1 vssd1 vccd1 vccd1 _5731_/S sky130_fd_sc_hd__clkbuf_16
Xfanout95 _5148_/A vssd1 vssd1 vccd1 vccd1 _5241_/A sky130_fd_sc_hd__buf_6
XANTENNA__5366__A _5367_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4270__A _4270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5156__A2 _5133_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5085__B _5093_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4364__B1 _4410_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5864__B1 _5863_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5092__A1 _4596_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3800_ _3443_/Y _3738_/X _3801_/B _3799_/X vssd1 vssd1 vccd1 vccd1 _3800_/X sky130_fd_sc_hd__o211a_1
X_4780_ _5358_/A _5367_/A vssd1 vssd1 vccd1 vccd1 _4781_/B sky130_fd_sc_hd__or2_1
XFILLER_21_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3731_ _6033_/Q _3730_/X _3731_/S vssd1 vssd1 vccd1 vccd1 _6033_/D sky130_fd_sc_hd__mux2_1
XFILLER_13_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3662_ _6208_/Q _3145_/C _3986_/B _3422_/A vssd1 vssd1 vccd1 vccd1 _3662_/X sky130_fd_sc_hd__a31o_1
X_5401_ _5327_/A _5446_/C _5386_/Y _5400_/Y vssd1 vssd1 vccd1 vccd1 _5401_/X sky130_fd_sc_hd__o31a_1
XANTENNA__5552__C1 _3122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3593_ _3593_/A _3593_/B _3594_/B vssd1 vssd1 vccd1 vccd1 _3642_/B sky130_fd_sc_hd__and3_2
X_5332_ _5333_/A _5333_/B vssd1 vssd1 vccd1 vccd1 _5387_/C sky130_fd_sc_hd__and2_4
XFILLER_114_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5263_ _5263_/A _5263_/B vssd1 vssd1 vccd1 vccd1 _5265_/A sky130_fd_sc_hd__xnor2_4
XFILLER_88_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4214_ _4214_/A _4214_/B _4215_/A vssd1 vssd1 vccd1 vccd1 _4214_/X sky130_fd_sc_hd__and3_2
X_5194_ _6215_/Q _5192_/C _5193_/Y vssd1 vssd1 vccd1 vccd1 _6215_/D sky130_fd_sc_hd__o21a_1
XANTENNA__3243__B _5924_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3330__A1 _3590_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4145_ _4145_/A _4145_/B vssd1 vssd1 vccd1 vccd1 _4146_/B sky130_fd_sc_hd__xnor2_4
XFILLER_110_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4058__C _5742_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5607__B1 _5607_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4076_ _4136_/A _4176_/B vssd1 vssd1 vccd1 vccd1 _4076_/Y sky130_fd_sc_hd__nand2_1
XFILLER_95_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3027_ _5054_/A vssd1 vssd1 vccd1 vccd1 _4648_/A sky130_fd_sc_hd__inv_4
XANTENNA_fanout261_A _5109_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3633__A2 _3765_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4978_ _5547_/B _4979_/B vssd1 vssd1 vccd1 vccd1 _4980_/A sky130_fd_sc_hd__nand2_1
XANTENNA__3397__A1 _4162_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3397__B2 _3885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4802__B _5703_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3929_ _3935_/D _3928_/X _3619_/C vssd1 vssd1 vccd1 vccd1 _3929_/X sky130_fd_sc_hd__o21a_1
XFILLER_137_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4897__B2 _5072_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5125__S _5129_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout230 _5625_/A vssd1 vssd1 vccd1 vccd1 _3958_/A sky130_fd_sc_hd__clkbuf_16
XANTENNA__4249__B _4251_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout241 _5128_/A0 vssd1 vssd1 vccd1 vccd1 _4216_/A sky130_fd_sc_hd__clkbuf_16
Xfanout252 _6238_/Q vssd1 vssd1 vccd1 vccd1 _4334_/A sky130_fd_sc_hd__buf_8
XANTENNA__3153__B _5143_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout263 _5109_/A vssd1 vssd1 vccd1 vccd1 _4096_/A sky130_fd_sc_hd__buf_6
Xfanout274 _6227_/Q vssd1 vssd1 vccd1 vccd1 _5488_/A sky130_fd_sc_hd__buf_6
XFILLER_86_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout285 _6220_/Q vssd1 vssd1 vccd1 vccd1 _5292_/B sky130_fd_sc_hd__buf_6
XFILLER_101_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout296 _6209_/Q vssd1 vssd1 vccd1 vccd1 _5960_/C1 sky130_fd_sc_hd__buf_6
XFILLER_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4265__A _4362_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4821__A1 _5358_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5795__S _5798_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5096__A _5148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3483__S1 _5940_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3560__A1 _4202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3063__B _5258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3998__B _4657_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4175__A _4202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5950_ _5911_/A _3867_/Y _3972_/Y _4697_/A _5876_/A vssd1 vssd1 vccd1 vccd1 _5951_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_19_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4901_ _5041_/S _4900_/Y _4640_/A _4638_/B vssd1 vssd1 vccd1 vccd1 _4901_/X sky130_fd_sc_hd__a211o_1
XFILLER_45_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5881_ _5707_/A _5124_/X _5880_/X _5707_/Y vssd1 vssd1 vccd1 vccd1 _5881_/X sky130_fd_sc_hd__a31o_1
XFILLER_33_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4832_ _4827_/X _4831_/X _5058_/C vssd1 vssd1 vccd1 vccd1 _4832_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_61_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5718__B _5898_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4763_ _5333_/A _4872_/B _4762_/X _4931_/B vssd1 vssd1 vccd1 vccd1 _4763_/X sky130_fd_sc_hd__o22a_1
XANTENNA__4622__B _4622_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3714_ _5504_/A _3708_/Y _3713_/X _5743_/C vssd1 vssd1 vccd1 vccd1 _3714_/X sky130_fd_sc_hd__o22a_1
X_4694_ _4707_/B _4806_/S _4692_/Y _4693_/X vssd1 vssd1 vccd1 vccd1 _4694_/X sky130_fd_sc_hd__o22a_1
XFILLER_119_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3645_ _3561_/A _3642_/Y _3643_/Y _3608_/A _3644_/X vssd1 vssd1 vccd1 vccd1 _4883_/B
+ sky130_fd_sc_hd__o221a_4
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5734__A _5734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3576_ _3658_/S _3567_/B _3575_/X vssd1 vssd1 vccd1 vccd1 _3618_/B sky130_fd_sc_hd__o21a_1
XANTENNA_fanout107_A _3557_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5544__A1_N _4645_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5315_ _5294_/Y _5309_/X _5312_/X _5314_/Y vssd1 vssd1 vccd1 vccd1 _5315_/X sky130_fd_sc_hd__a31o_1
XFILLER_88_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6295_ _6295_/CLK _6295_/D vssd1 vssd1 vccd1 vccd1 _6295_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_88_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3254__A _5936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5246_ _5075_/A _5245_/X _5080_/B vssd1 vssd1 vccd1 vccd1 _5250_/C sky130_fd_sc_hd__a21oi_1
XFILLER_88_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5177_ _3058_/B _3672_/Y _3121_/X vssd1 vssd1 vccd1 vccd1 _5177_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_68_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4128_ _3819_/B _4069_/B _4072_/C _6083_/Q vssd1 vssd1 vccd1 vccd1 _4128_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_110_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5056__A1 _5090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4059_ _4476_/S _4059_/B vssd1 vssd1 vccd1 vccd1 _4066_/S sky130_fd_sc_hd__nand2_8
XANTENNA__4085__A _4085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3148__B _4577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3790__A1 _4162_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3164__A _3205_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4707__B _4707_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5047__A1 _4625_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_857 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3339__A _5818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3058__B _3058_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3430_ _6261_/Q _5439_/A2 _5924_/B _6030_/Q _3429_/X vssd1 vssd1 vccd1 vccd1 _3430_/X
+ sky130_fd_sc_hd__o221a_2
XANTENNA__4730__B1 _4886_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3361_ _3935_/B _3361_/B vssd1 vssd1 vccd1 vccd1 _3361_/Y sky130_fd_sc_hd__nand2_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5100_ _6009_/Q _3111_/X _5097_/X vssd1 vssd1 vccd1 vccd1 _5100_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_112_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6080_ _6272_/CLK _6080_/D vssd1 vssd1 vccd1 vccd1 _6080_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3292_ _3561_/A _3608_/A vssd1 vssd1 vccd1 vccd1 _3644_/B sky130_fd_sc_hd__nand2_8
XFILLER_112_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5031_ _5031_/A vssd1 vssd1 vccd1 vccd1 _5031_/Y sky130_fd_sc_hd__inv_2
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5286__B2 _5442_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5038__A1 _5567_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5933_ _4657_/A _4586_/Y _5921_/X vssd1 vssd1 vccd1 vccd1 _5940_/S sky130_fd_sc_hd__o21a_1
XFILLER_15_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4261__A2 _4214_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4633__A _5255_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5864_ _6287_/Q _5854_/A _5863_/Y _5866_/B1 vssd1 vssd1 vccd1 vccd1 _6287_/D sky130_fd_sc_hd__o211a_1
XFILLER_21_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4815_ _6188_/Q _4814_/C _6189_/Q vssd1 vssd1 vccd1 vccd1 _4816_/B sky130_fd_sc_hd__a21oi_1
X_5795_ _6261_/Q _3721_/X _5798_/S vssd1 vssd1 vccd1 vccd1 _6261_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4013__A2 _3274_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout224_A _6295_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4746_ _4744_/B _4743_/X _4745_/A _4740_/X _5034_/A vssd1 vssd1 vccd1 vccd1 _4753_/B
+ sky130_fd_sc_hd__a221o_1
X_4677_ _3116_/B _4668_/X _4669_/X _4744_/B _4676_/X vssd1 vssd1 vccd1 vccd1 _4677_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5464__A _5464_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3628_ _3145_/C _3652_/A _3621_/X _3627_/Y _3422_/A vssd1 vssd1 vccd1 vccd1 _3628_/X
+ sky130_fd_sc_hd__a221o_1
Xoutput17 _6191_/Q vssd1 vssd1 vccd1 vccd1 io_out[15] sky130_fd_sc_hd__buf_4
Xoutput28 _6182_/Q vssd1 vssd1 vccd1 vccd1 io_out[25] sky130_fd_sc_hd__buf_4
XFILLER_122_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3559_ _3164_/Y _3443_/Y _3558_/X vssd1 vssd1 vccd1 vccd1 _3559_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_103_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6278_ _6278_/CLK _6278_/D vssd1 vssd1 vccd1 vccd1 _6278_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5229_ _5768_/A0 _5227_/B _5228_/X _5227_/A vssd1 vssd1 vccd1 vccd1 _5229_/X sky130_fd_sc_hd__a211o_1
XANTENNA__4808__A input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3827__A2 _3740_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_640 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_779 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4004__A2 _3030_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5201__A1 _5191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3159__A _3974_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4960__B1 _4648_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5093__B _5093_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5268__A1 _4678_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3279__B1 _5450_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output20_A _6194_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3451__B1 _3450_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4600_ _4963_/A _4654_/A vssd1 vssd1 vccd1 vccd1 _4600_/Y sky130_fd_sc_hd__nor2_1
X_5580_ _5595_/B vssd1 vssd1 vccd1 vccd1 _5580_/Y sky130_fd_sc_hd__inv_2
XFILLER_129_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4531_ _5932_/A _6167_/Q vssd1 vssd1 vccd1 vccd1 _6166_/D sky130_fd_sc_hd__or2_1
XFILLER_7_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5284__A _5512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4462_ _4462_/A _4462_/B _5925_/A vssd1 vssd1 vccd1 vccd1 _4477_/S sky130_fd_sc_hd__or3_4
XANTENNA__3506__A1 _4772_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6201_ _6206_/CLK _6201_/D vssd1 vssd1 vccd1 vccd1 _6201_/Q sky130_fd_sc_hd__dfxtp_1
X_3413_ _3935_/B _3361_/B _3373_/B _3358_/A vssd1 vssd1 vccd1 vccd1 _3414_/B sky130_fd_sc_hd__o22ai_4
X_4393_ _4393_/A _4393_/B _4393_/C vssd1 vssd1 vccd1 vccd1 _4394_/B sky130_fd_sc_hd__or3_1
XFILLER_98_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6132_ _6176_/CLK _6132_/D vssd1 vssd1 vccd1 vccd1 _6132_/Q sky130_fd_sc_hd__dfxtp_1
X_3344_ _3498_/S _3388_/A _3343_/X _3210_/B vssd1 vssd1 vccd1 vccd1 _3344_/X sky130_fd_sc_hd__o211a_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6063_ _6250_/CLK _6063_/D vssd1 vssd1 vccd1 vccd1 _6063_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4628__A _5226_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3275_ _5226_/A _3636_/A _3211_/Y _3269_/Y vssd1 vssd1 vccd1 vccd1 _3275_/X sky130_fd_sc_hd__a211o_1
XFILLER_97_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5014_ _4989_/A _4989_/B _4980_/A vssd1 vssd1 vccd1 vccd1 _5015_/B sky130_fd_sc_hd__a21bo_1
XFILLER_38_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3690__A0 _5935_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout174_A _4214_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5431__A1 _5605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout341_A input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5916_ _4577_/A _5172_/A _3678_/C _5915_/Y vssd1 vssd1 vccd1 vccd1 _5916_/Y sky130_fd_sc_hd__a31oi_1
XFILLER_34_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5847_ _6282_/Q _5854_/A _5846_/Y _5866_/B1 vssd1 vssd1 vccd1 vccd1 _6282_/D sky130_fd_sc_hd__o211a_1
XANTENNA__4082__B _4176_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5778_ _3942_/D _4250_/Y _5776_/X _5777_/Y vssd1 vssd1 vccd1 vccd1 _6253_/D sky130_fd_sc_hd__a22o_1
X_4729_ _4698_/A _4728_/X _4727_/Y vssd1 vssd1 vccd1 vccd1 _4729_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_108_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3707__A _3732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3145__C _3145_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout87_A _5570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3442__A _5818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5670__A1 _5710_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5958__C1 _5960_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5422__A1 _5428_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4273__A _4301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5973__A2 _5503_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5725__A2 _3649_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4161__A1 _4301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4161__B2 _4162_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3055__C _3885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3060_ _3060_/A _3060_/B vssd1 vssd1 vccd1 vccd1 _3060_/Y sky130_fd_sc_hd__nand2_2
XANTENNA__4167__B _4197_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5661__A1 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5413__A1 _5058_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3962_ _3880_/B _5870_/A _3996_/B _5105_/A vssd1 vssd1 vccd1 vccd1 _5645_/A sky130_fd_sc_hd__a31o_2
XANTENNA__5964__A2 _5970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5701_ _3513_/B _3958_/Y _5691_/X _5700_/X vssd1 vssd1 vccd1 vccd1 _5701_/X sky130_fd_sc_hd__a211o_1
XFILLER_50_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3893_ _5124_/S _3893_/B _3893_/C vssd1 vssd1 vccd1 vccd1 _5961_/A sky130_fd_sc_hd__nor3_1
XANTENNA__5177__B1 _3121_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5632_ _5644_/A _5644_/B _5644_/C _5632_/D vssd1 vssd1 vccd1 vccd1 _5632_/X sky130_fd_sc_hd__and4_1
XANTENNA__5716__A2 _3958_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5563_ _4644_/B _5572_/B _5562_/Y _3121_/B _5507_/A vssd1 vssd1 vccd1 vccd1 _5563_/X
+ sky130_fd_sc_hd__a221o_1
X_4514_ _5856_/A _3912_/Y _4512_/X _4513_/Y vssd1 vssd1 vccd1 vccd1 _6153_/D sky130_fd_sc_hd__a22o_1
XFILLER_117_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5494_ _5494_/A _5494_/B _5494_/C vssd1 vssd1 vccd1 vccd1 _5494_/X sky130_fd_sc_hd__and3_1
XFILLER_117_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4445_ _5926_/A0 _3900_/Y _4443_/X _4444_/Y vssd1 vssd1 vccd1 vccd1 _6119_/D sky130_fd_sc_hd__a22o_1
X_4376_ _4376_/A _4376_/B vssd1 vssd1 vccd1 vccd1 _4379_/A sky130_fd_sc_hd__nand2_1
XFILLER_59_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6115_ _6280_/CLK _6115_/D vssd1 vssd1 vccd1 vccd1 _6115_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3327_ _6095_/Q _3589_/A2 _3589_/B1 _6088_/Q vssd1 vssd1 vccd1 vccd1 _3327_/X sky130_fd_sc_hd__o22a_1
XFILLER_98_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout291_A _3105_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3262__A _3885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3338__S0 _4067_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6046_ _6259_/CLK _6046_/D vssd1 vssd1 vccd1 vccd1 _6046_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3258_ _3766_/A _3555_/B vssd1 vssd1 vccd1 vccd1 _3750_/C sky130_fd_sc_hd__nand2_2
XANTENNA__4077__B _4136_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5652__A1 _3251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3189_ _3766_/A _4462_/A vssd1 vssd1 vccd1 vccd1 _3706_/A sky130_fd_sc_hd__or2_4
XFILLER_26_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_54_clk_A _6133_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5404__A1 _4596_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5404__B2 _5463_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4093__A _4162_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3718__A1 _6013_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5128__S _5128_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3156__B _4622_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4694__A2 _4806_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5891__A1 _5653_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3172__A _6200_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3329__S0 _3241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5798__S _5798_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5643__A1 _3103_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3900__A _5767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4851__C1 _3740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5946__A2 _4586_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5159__B1 _4931_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3347__A _3450_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4230_ _4193_/A _4193_/B _4229_/A _4229_/B vssd1 vssd1 vccd1 vccd1 _4230_/X sky130_fd_sc_hd__o211a_2
XFILLER_68_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4161_ _4301_/A _4309_/B _4342_/B _4162_/B vssd1 vssd1 vccd1 vccd1 _4165_/A sky130_fd_sc_hd__a22o_1
XFILLER_122_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3112_ _5065_/A _3112_/B vssd1 vssd1 vccd1 vccd1 _4605_/A sky130_fd_sc_hd__nand2_4
XFILLER_67_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4092_ _4233_/A1 _4090_/X _4091_/X vssd1 vssd1 vccd1 vccd1 _6081_/D sky130_fd_sc_hd__a21o_1
XFILLER_67_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3043_ _3880_/B _5065_/A vssd1 vssd1 vccd1 vccd1 _3043_/Y sky130_fd_sc_hd__nor2_4
XFILLER_55_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4625__B _5093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5398__B1 _5360_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4994_ _5547_/B _4644_/B _4992_/Y _4993_/X vssd1 vssd1 vccd1 vccd1 _4994_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5937__A2 _5934_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3945_ _5634_/B _3945_/B vssd1 vssd1 vccd1 vccd1 _3945_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__4070__B1 _4539_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6084__CLK _6084_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4641__A _5218_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3876_ _5959_/A _5138_/A _5951_/A vssd1 vssd1 vccd1 vccd1 _5911_/D sky130_fd_sc_hd__or3b_1
XANTENNA_fanout137_A _5957_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5615_ _4659_/B _4665_/B _5703_/A vssd1 vssd1 vccd1 vccd1 _5615_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3257__A _3732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5546_ _5538_/Y _5545_/X _5551_/A vssd1 vssd1 vccd1 vccd1 _5546_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout304_A _6067_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3691__S _3902_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5477_ _4974_/A _5476_/Y _3060_/Y vssd1 vssd1 vccd1 vccd1 _5477_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_132_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5322__B1 _5321_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4428_ _4428_/A _4428_/B vssd1 vssd1 vccd1 vccd1 _4429_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__5873__A1 _4003_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3704__B _3704_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4359_ _4383_/S _4359_/B vssd1 vssd1 vccd1 vccd1 _4359_/Y sky130_fd_sc_hd__nor2_1
XFILLER_86_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5086__C1 _5136_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6029_ _6259_/CLK _6029_/D vssd1 vssd1 vccd1 vccd1 _6029_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3939__A1 _5677_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout41 _4072_/Y vssd1 vssd1 vccd1 vccd1 _4437_/A1 sky130_fd_sc_hd__clkbuf_8
Xfanout52 _5871_/C vssd1 vssd1 vccd1 vccd1 _4872_/B sky130_fd_sc_hd__buf_4
Xfanout63 _4642_/Y vssd1 vssd1 vccd1 vccd1 _4645_/B sky130_fd_sc_hd__buf_6
XFILLER_120_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout74 _3195_/X vssd1 vssd1 vccd1 vccd1 _3765_/B sky130_fd_sc_hd__buf_4
XFILLER_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout85 _3090_/Y vssd1 vssd1 vccd1 vccd1 _4946_/A sky130_fd_sc_hd__clkbuf_16
Xfanout96 _3079_/Y vssd1 vssd1 vccd1 vccd1 _5148_/A sky130_fd_sc_hd__buf_8
XANTENNA__5366__B _5367_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4270__B _5109_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3167__A _6009_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4364__A1 _4334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5561__A0 _5567_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4364__B2 _4362_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_331 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5313__B1 _5607_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3614__B _3615_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5616__A1 _5454_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4726__A _5114_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5557__A _5567_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3730_ _6017_/Q _3706_/Y _3729_/X vssd1 vssd1 vccd1 vccd1 _3730_/X sky130_fd_sc_hd__a21o_4
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3661_ _3655_/X _3659_/X _3660_/Y vssd1 vssd1 vccd1 vccd1 _3661_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__3077__A _3105_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5400_ _5498_/A _5397_/X _5399_/X vssd1 vssd1 vccd1 vccd1 _5400_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3592_ _3592_/A _3592_/B vssd1 vssd1 vccd1 vccd1 _3592_/X sky130_fd_sc_hd__or2_1
XFILLER_127_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5331_ _3033_/Y _5330_/B _5330_/Y _3121_/B vssd1 vssd1 vccd1 vccd1 _5331_/X sky130_fd_sc_hd__o211a_1
XFILLER_114_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5292__A _6221_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5262_ _5263_/A _5263_/B vssd1 vssd1 vccd1 vccd1 _5262_/X sky130_fd_sc_hd__and2_2
XFILLER_102_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4213_ _4214_/A _4214_/B vssd1 vssd1 vccd1 vccd1 _4215_/B sky130_fd_sc_hd__nand2_1
XFILLER_130_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5193_ _6215_/Q _5192_/C _5192_/A vssd1 vssd1 vccd1 vccd1 _5193_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_68_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4144_ _4163_/A _4176_/B _4145_/A vssd1 vssd1 vccd1 vccd1 _4144_/X sky130_fd_sc_hd__and3_1
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4075_ _4197_/A _4173_/B vssd1 vssd1 vccd1 vccd1 _4084_/A sky130_fd_sc_hd__nand2_2
XFILLER_37_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3026_ _3312_/A vssd1 vssd1 vccd1 vccd1 _3974_/B sky130_fd_sc_hd__inv_8
XFILLER_36_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout254_A _6237_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3686__S _3902_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4977_ _4745_/A _4975_/X _4992_/B _4744_/B _5034_/A vssd1 vssd1 vccd1 vccd1 _4977_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5240__C1 _4605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3397__A2 _3257_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3928_ _3935_/C _3927_/X _3572_/C vssd1 vssd1 vccd1 vccd1 _3928_/X sky130_fd_sc_hd__o21a_1
XFILLER_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3859_ _6057_/Q _5976_/A vssd1 vssd1 vccd1 vccd1 _3859_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5543__A0 _5344_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4897__A2 _4647_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5529_ _5310_/Y _5522_/Y _5528_/X _5403_/A vssd1 vssd1 vccd1 vccd1 _5531_/A sky130_fd_sc_hd__a211o_1
XFILLER_117_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout220 _3713_/S vssd1 vssd1 vccd1 vccd1 _3709_/S sky130_fd_sc_hd__buf_8
XFILLER_132_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout231 _5625_/A vssd1 vssd1 vccd1 vccd1 _5634_/A sky130_fd_sc_hd__buf_4
XFILLER_120_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout242 _6241_/Q vssd1 vssd1 vccd1 vccd1 _5128_/A0 sky130_fd_sc_hd__buf_6
Xfanout253 _6238_/Q vssd1 vssd1 vccd1 vccd1 _4163_/A sky130_fd_sc_hd__buf_6
Xfanout264 _6235_/Q vssd1 vssd1 vccd1 vccd1 _5109_/A sky130_fd_sc_hd__buf_12
XFILLER_59_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout275 _5480_/B vssd1 vssd1 vccd1 vccd1 _4891_/A sky130_fd_sc_hd__buf_6
Xfanout286 _5768_/A0 vssd1 vssd1 vccd1 vccd1 _5255_/B sky130_fd_sc_hd__buf_8
XFILLER_87_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout297 _6071_/Q vssd1 vssd1 vccd1 vccd1 _3970_/A sky130_fd_sc_hd__buf_12
XFILLER_19_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3450__A _3450_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4265__B _4334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4821__A2 _5367_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4337__A1 _4362_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5837__A1 _5158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5840__A _5840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4175__B _4176_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4900_ _4900_/A _4900_/B vssd1 vssd1 vccd1 vccd1 _4900_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_33_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5880_ _3942_/B _5934_/A _3883_/X vssd1 vssd1 vccd1 vccd1 _5880_/X sky130_fd_sc_hd__a21o_1
XFILLER_34_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4831_ _4990_/A _4829_/Y _4830_/X _4640_/A _4644_/A vssd1 vssd1 vccd1 vccd1 _4831_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3379__A2 _3589_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4762_ _6222_/Q _4587_/B _4761_/X _5239_/A _4753_/Y vssd1 vssd1 vccd1 vccd1 _4762_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_60_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4622__C _5220_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3713_ _6012_/Q _6035_/Q _3713_/S vssd1 vssd1 vccd1 vccd1 _3713_/X sky130_fd_sc_hd__mux2_8
X_4693_ _4692_/A _4692_/B _4842_/B vssd1 vssd1 vccd1 vccd1 _4693_/X sky130_fd_sc_hd__a21o_1
XANTENNA__3238__C _5436_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5525__B1 _5522_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3644_ _3986_/B _3644_/B vssd1 vssd1 vccd1 vccd1 _3644_/X sky130_fd_sc_hd__or2_1
XANTENNA__5734__B _5734_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3575_ _6206_/Q _3575_/B vssd1 vssd1 vccd1 vccd1 _3575_/X sky130_fd_sc_hd__or2_1
X_5314_ _4638_/Y _5302_/B _5313_/Y vssd1 vssd1 vccd1 vccd1 _5314_/Y sky130_fd_sc_hd__a21oi_1
X_6294_ _6295_/CLK _6294_/D vssd1 vssd1 vccd1 vccd1 _6294_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5289__C1 _5948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5828__A1 _5835_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3254__B _3706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5245_ _5911_/A _5244_/A _4648_/Y _5244_/X vssd1 vssd1 vccd1 vccd1 _5245_/X sky130_fd_sc_hd__a31o_1
XFILLER_114_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4500__A1 _4891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5176_ _5191_/A _3092_/B _5071_/A _5175_/X vssd1 vssd1 vccd1 vccd1 _6212_/D sky130_fd_sc_hd__o211a_1
XFILLER_56_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4127_ _4123_/A _4126_/X _4123_/Y vssd1 vssd1 vccd1 vccd1 _4127_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_96_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4366__A _4410_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5056__A2 _4745_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4058_ _5436_/A _4058_/B _5742_/C vssd1 vssd1 vccd1 vccd1 _4059_/B sky130_fd_sc_hd__or3_4
XFILLER_45_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4085__B _4311_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5461__C1 _3122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3009_ _5488_/A vssd1 vssd1 vccd1 vccd1 _3009_/Y sky130_fd_sc_hd__inv_2
XFILLER_43_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_663 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5909__B _5909_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4016__B1 _4850_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5925__A _5925_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3790__A2 _3777_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4040__S _4044_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3180__A _4577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5047__A2 _5093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_54_clk _6133_/CLK vssd1 vssd1 vccd1 vccd1 _6180_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_55_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4007__B1 _3032_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4558__A1 _3942_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3339__B _3555_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3533__A2 _3901_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3360_ _3935_/B _3361_/B vssd1 vssd1 vccd1 vccd1 _3360_/X sky130_fd_sc_hd__or2_1
XFILLER_98_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3291_ _6008_/Q _6009_/Q vssd1 vssd1 vccd1 vccd1 _3608_/A sky130_fd_sc_hd__nand2b_4
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5570__A _5570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5030_ _5547_/A _5547_/B _5504_/A _5488_/A _5029_/B vssd1 vssd1 vccd1 vccd1 _5031_/A
+ sky130_fd_sc_hd__o41a_1
XFILLER_111_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5038__A2 _4645_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5443__C1 _5513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5932_ _5932_/A _5932_/B vssd1 vssd1 vccd1 vccd1 _6293_/D sky130_fd_sc_hd__nor2_1
XANTENNA__4797__A1 _5358_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4914__A _4974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_45_clk _6233_/CLK vssd1 vssd1 vccd1 vccd1 _6232_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_34_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5863_ _3607_/B _5862_/B _5862_/Y _5867_/A1 vssd1 vssd1 vccd1 vccd1 _5863_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_22_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4633__B _4633_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4549__A1 _5926_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4814_ _6189_/Q _6188_/Q _4814_/C vssd1 vssd1 vccd1 vccd1 _4854_/B sky130_fd_sc_hd__and3_1
XFILLER_22_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5794_ _6260_/Q _3718_/X _5798_/S vssd1 vssd1 vccd1 vccd1 _6260_/D sky130_fd_sc_hd__mux2_1
X_4745_ _4745_/A vssd1 vssd1 vccd1 vccd1 _4745_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4676_ _5034_/A _4710_/B _4676_/C vssd1 vssd1 vccd1 vccd1 _4676_/X sky130_fd_sc_hd__and3_1
XFILLER_107_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3627_ _3312_/Y _3623_/Y _3626_/X vssd1 vssd1 vccd1 vccd1 _3627_/Y sky130_fd_sc_hd__a21oi_1
Xoutput18 _6192_/Q vssd1 vssd1 vccd1 vccd1 io_out[16] sky130_fd_sc_hd__buf_4
Xoutput29 _6300_/Q vssd1 vssd1 vccd1 vccd1 io_out[26] sky130_fd_sc_hd__buf_4
X_3558_ _3398_/A _3607_/B _3550_/X _3498_/S vssd1 vssd1 vccd1 vccd1 _3558_/X sky130_fd_sc_hd__o211a_1
XFILLER_1_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6277_ _6279_/CLK _6277_/D vssd1 vssd1 vccd1 vccd1 _6277_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3489_ _6270_/Q _6016_/Q _6084_/Q _6039_/Q _4067_/A _3709_/S vssd1 vssd1 vccd1 vccd1
+ _3490_/C sky130_fd_sc_hd__mux4_1
XANTENNA__5480__A _5488_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5228_ _5225_/Y _5226_/X _5605_/C vssd1 vssd1 vccd1 vccd1 _5228_/X sky130_fd_sc_hd__o21a_1
XFILLER_76_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4808__B _4808_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5682__C1 _3950_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4096__A _4096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5159_ _4589_/Y _5148_/Y _5158_/X _4931_/B _3014_/A vssd1 vssd1 vccd1 vccd1 _5159_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_96_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5434__C1 _5607_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4788__A1 _5367_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4824__A _5509_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_36_clk clkbuf_3_4__f_clk/X vssd1 vssd1 vccd1 vccd1 _6260_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_112_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3460__A1 _3410_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4960__A1 _6193_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4960__B2 _6004_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_556 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5390__A _5392_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4476__A0 _4891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3279__A1 _4216_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3279__B2 _3885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5673__C1 _3974_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_747 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4734__A _5114_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_27_clk _6084_/CLK vssd1 vssd1 vccd1 vccd1 _6280_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5440__A2 _3901_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3451__A1 _3450_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4530_ _4539_/A _6166_/Q vssd1 vssd1 vccd1 vccd1 _6165_/D sky130_fd_sc_hd__and2_1
XFILLER_117_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4461_ _5255_/B _6125_/Q _4476_/S vssd1 vssd1 vccd1 vccd1 _4461_/X sky130_fd_sc_hd__mux2_1
X_6200_ _6302_/CLK _6200_/D vssd1 vssd1 vccd1 vccd1 _6200_/Q sky130_fd_sc_hd__dfxtp_4
X_3412_ _3925_/A vssd1 vssd1 vccd1 vccd1 _3412_/Y sky130_fd_sc_hd__inv_2
X_4392_ _4393_/A _4393_/B _4393_/C vssd1 vssd1 vccd1 vccd1 _4394_/A sky130_fd_sc_hd__o21ai_4
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6131_ _6155_/CLK _6131_/D vssd1 vssd1 vccd1 vccd1 _6131_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3343_ _3211_/Y _3410_/B _3342_/X _3204_/Y vssd1 vssd1 vccd1 vccd1 _3343_/X sky130_fd_sc_hd__a211o_1
XFILLER_112_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4909__A _4945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6062_ _6093_/CLK _6062_/D vssd1 vssd1 vccd1 vccd1 _6062_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4467__A0 _5926_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3274_ _3274_/A _3274_/B vssd1 vssd1 vccd1 vccd1 _3274_/X sky130_fd_sc_hd__or2_4
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4628__B _4806_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5664__C1 _5956_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5013_ _5547_/A _4645_/B _5011_/Y _5012_/X vssd1 vssd1 vccd1 vccd1 _5013_/X sky130_fd_sc_hd__o22a_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4644__A _4644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_18_clk _6084_/CLK vssd1 vssd1 vccd1 vccd1 _6270_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_41_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5915_ _3312_/A _5238_/C _5172_/A vssd1 vssd1 vccd1 vccd1 _5915_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__5719__A0 _4846_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5846_ _5854_/A _5846_/B vssd1 vssd1 vccd1 vccd1 _5846_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_fanout334_A _4846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5777_ _3011_/Y _5788_/B _4250_/Y vssd1 vssd1 vccd1 vccd1 _5777_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__3694__S _3705_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4942__A1 _6192_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4728_ _4697_/A _4697_/B _4660_/A _4660_/B _4657_/X vssd1 vssd1 vccd1 vccd1 _4728_/X
+ sky130_fd_sc_hd__a221o_4
XANTENNA__3707__B _4462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4659_ _5226_/A _4659_/B vssd1 vssd1 vccd1 vccd1 _4660_/B sky130_fd_sc_hd__and2_2
XFILLER_116_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4819__A _5385_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3442__B _3555_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3130__A0 _4707_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5670__A2 _4111_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5958__B1 _5131_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4273__B _4389_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3433__A1 _4301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4630__B1 _4972_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5973__A3 _3883_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5385__A _5385_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4161__A2 _4309_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4167__C _4167_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3100__C_N _3116_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5661__A2 _3179_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3424__A1 _3937_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3961_ _5158_/A _3978_/B vssd1 vssd1 vccd1 vccd1 _5634_/D sky130_fd_sc_hd__nand2_1
X_5700_ _3043_/Y _3495_/B _5698_/X _5699_/Y _5728_/A vssd1 vssd1 vccd1 vccd1 _5700_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3892_ _3893_/B _3892_/B vssd1 vssd1 vccd1 vccd1 _5735_/S sky130_fd_sc_hd__nor2_4
XANTENNA__5177__A1 _3058_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5631_ _5264_/A _3179_/X _5626_/Y _5630_/X _3974_/C vssd1 vssd1 vccd1 vccd1 _5631_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__5295__A _5296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5562_ _3041_/Y _5360_/S _5364_/Y vssd1 vssd1 vccd1 vccd1 _5562_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_129_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4513_ _3010_/Y _4515_/B _3912_/Y vssd1 vssd1 vccd1 vccd1 _4513_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_8_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5493_ _3250_/X _5442_/A _5482_/Y _5943_/C vssd1 vssd1 vccd1 vccd1 _5494_/C sky130_fd_sc_hd__o22a_1
X_4444_ _5305_/A _4458_/B _3900_/Y vssd1 vssd1 vccd1 vccd1 _4444_/Y sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_7_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _6214_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__5742__B _5742_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5885__C1 _5956_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4375_ _4375_/A _4375_/B vssd1 vssd1 vccd1 vccd1 _4376_/B sky130_fd_sc_hd__or2_1
XANTENNA__4639__A _5911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6114_ _6278_/CLK _6114_/D vssd1 vssd1 vccd1 vccd1 _6114_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3326_ _5924_/A _6060_/Q _5436_/C vssd1 vssd1 vccd1 vccd1 _3326_/X sky130_fd_sc_hd__and3_1
XFILLER_98_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3262__B _5264_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6045_ _6293_/CLK _6045_/D vssd1 vssd1 vccd1 vccd1 _6045_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3257_ _3732_/A _3257_/B vssd1 vssd1 vccd1 vccd1 _3749_/C sky130_fd_sc_hd__nor2_1
XANTENNA_fanout284_A _6220_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4077__C _4173_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5652__A2 _5728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3188_ _5730_/A _5617_/B _3940_/A _3215_/B vssd1 vssd1 vccd1 vccd1 _3188_/X sky130_fd_sc_hd__or4_1
XANTENNA__3663__A1 _3511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3689__S _3902_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4093__B _4216_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5168__A1 _3970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5829_ _3529_/X _5819_/B _5828_/X vssd1 vssd1 vccd1 vccd1 _6277_/D sky130_fd_sc_hd__a21o_1
XANTENNA__4915__A1 _5731_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4915__B2 _3101_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5628__C1 _3772_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3329__S1 _3241_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3900__B _3901_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3406__B2 _3541_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_3_7__f_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4906__A1 _4625_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3347__B _3986_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5331__A1 _3033_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4160_ _4202_/A _4173_/B _4146_/B _4144_/X vssd1 vssd1 vccd1 vccd1 _4185_/A sky130_fd_sc_hd__a31o_4
XFILLER_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5619__C1 _4946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3111_ _5075_/B _3111_/B vssd1 vssd1 vccd1 vccd1 _3111_/X sky130_fd_sc_hd__or2_4
XFILLER_56_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4091_ _3795_/B _4069_/B _4072_/C _6081_/Q vssd1 vssd1 vccd1 vccd1 _4091_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_110_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3042_ _6157_/Q vssd1 vssd1 vccd1 vccd1 _3042_/Y sky130_fd_sc_hd__inv_2
XFILLER_82_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5398__A1 _4819_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4993_ _6194_/Q _3671_/Y _5172_/B _6005_/Q _5605_/C vssd1 vssd1 vccd1 vccd1 _4993_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__5398__B2 _6008_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3944_ _3944_/A _3944_/B vssd1 vssd1 vccd1 vccd1 _3945_/B sky130_fd_sc_hd__nand2_1
XANTENNA__4070__A1 _5960_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4641__B _4646_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3875_ _5137_/D _3966_/B vssd1 vssd1 vccd1 vccd1 _5951_/A sky130_fd_sc_hd__nor2_1
XANTENNA__3538__A _3567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5614_ _5653_/A _5889_/B vssd1 vssd1 vccd1 vccd1 _5614_/X sky130_fd_sc_hd__or2_1
XFILLER_118_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3257__B _3257_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5545_ _5072_/B _5551_/B _5544_/X _3060_/B vssd1 vssd1 vccd1 vccd1 _5545_/X sky130_fd_sc_hd__a211o_1
XFILLER_117_354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3581__B1 _3422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5476_ _5476_/A _5476_/B vssd1 vssd1 vccd1 vccd1 _5476_/Y sky130_fd_sc_hd__nor2_2
XFILLER_117_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5858__C1 _5866_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4427_ _4394_/A _4424_/C _4412_/Y vssd1 vssd1 vccd1 vccd1 _4428_/B sky130_fd_sc_hd__o21ai_4
XANTENNA__5322__A1 _5943_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5322__B2 _5442_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3704__C _5767_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4358_ _4358_/A _4358_/B _4358_/C vssd1 vssd1 vccd1 vccd1 _4359_/B sky130_fd_sc_hd__and3_1
XFILLER_99_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3884__A1 _3112_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input4_A io_in[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3309_ _3310_/A _5889_/A vssd1 vssd1 vccd1 vccd1 _3309_/X sky130_fd_sc_hd__and2_1
XFILLER_59_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4289_ _4326_/B _4289_/B _4289_/C vssd1 vssd1 vccd1 vccd1 _4330_/A sky130_fd_sc_hd__nand3_4
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5086__B1 _5158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6028_ _6295_/CLK _6028_/D vssd1 vssd1 vccd1 vccd1 _6028_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3939__A2 _5898_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4061__A1 _3715_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout42 _4072_/Y vssd1 vssd1 vccd1 vccd1 _4233_/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout53 _4654_/Y vssd1 vssd1 vccd1 vccd1 _5871_/C sky130_fd_sc_hd__clkbuf_4
Xfanout64 _4638_/Y vssd1 vssd1 vccd1 vccd1 _5463_/A sky130_fd_sc_hd__buf_6
XFILLER_50_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout75 _5943_/A vssd1 vssd1 vccd1 vccd1 _3832_/A2 sky130_fd_sc_hd__buf_4
Xfanout86 _3090_/Y vssd1 vssd1 vccd1 vccd1 _3740_/A sky130_fd_sc_hd__buf_4
XFILLER_22_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4043__S _4044_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout97 _3058_/Y vssd1 vssd1 vccd1 vccd1 _5227_/A sky130_fd_sc_hd__clkbuf_16
XANTENNA__4270__C _4426_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3167__B _6008_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4364__A2 _4426_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5313__A1 _5464_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3183__A _5870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3627__A1 _3312_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4726__B _4726_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4052__A1 _3880_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4052__B2 _4697_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3660_ _4003_/B _3651_/B _3881_/A vssd1 vssd1 vccd1 vccd1 _3660_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__3077__B _5239_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5552__A1 _5551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3591_ _4410_/B _3832_/A2 _3251_/B _3590_/X _3255_/Y vssd1 vssd1 vccd1 vccd1 _3592_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_127_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5330_ _6006_/Q _5330_/B vssd1 vssd1 vccd1 vccd1 _5330_/Y sky130_fd_sc_hd__nand2_1
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_53_clk_A _6133_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5292__B _5292_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5261_ _5263_/A _5653_/A vssd1 vssd1 vccd1 vccd1 _5261_/Y sky130_fd_sc_hd__nand2_2
XFILLER_126_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4212_ _4165_/A _4165_/C _4165_/B vssd1 vssd1 vccd1 vccd1 _4215_/A sky130_fd_sc_hd__a21bo_1
XFILLER_102_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5192_ _5192_/A _5192_/B _5192_/C vssd1 vssd1 vccd1 vccd1 _6214_/D sky130_fd_sc_hd__nor3_1
X_4143_ _4163_/A _4176_/B vssd1 vssd1 vccd1 vccd1 _4145_/B sky130_fd_sc_hd__nand2_2
XFILLER_110_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5068__B1 _5239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4074_ _6079_/Q _4072_/C _4073_/X vssd1 vssd1 vccd1 vccd1 _6079_/D sky130_fd_sc_hd__a21o_1
XFILLER_37_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4815__B1 _6189_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3025_ _3958_/A vssd1 vssd1 vccd1 vccd1 _3025_/Y sky130_fd_sc_hd__inv_4
XFILLER_64_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4043__A1 _3727_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4976_ _6194_/Q _5002_/C vssd1 vssd1 vccd1 vccd1 _4992_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__5240__B1 _4596_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout247_A _5859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3927_ _3924_/X _3925_/X _3926_/X _3518_/Y vssd1 vssd1 vccd1 vccd1 _3927_/X sky130_fd_sc_hd__o211a_1
XFILLER_137_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3858_ _6058_/Q _3869_/A vssd1 vssd1 vccd1 vccd1 _3858_/X sky130_fd_sc_hd__xor2_1
XFILLER_109_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3789_ _3986_/A _3746_/A _3788_/X _3849_/B vssd1 vssd1 vccd1 vccd1 _3789_/X sky130_fd_sc_hd__a211o_1
X_5528_ _4643_/A _5526_/X _5527_/Y _5291_/Y vssd1 vssd1 vccd1 vccd1 _5528_/X sky130_fd_sc_hd__a22o_1
XFILLER_105_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5459_ _5327_/A _5504_/C _5447_/Y _5458_/Y vssd1 vssd1 vccd1 vccd1 _5459_/X sky130_fd_sc_hd__o31a_1
XFILLER_106_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout210 _5733_/A vssd1 vssd1 vccd1 vccd1 _5239_/A sky130_fd_sc_hd__buf_6
XFILLER_121_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout221 _3713_/S vssd1 vssd1 vccd1 vccd1 _3551_/S sky130_fd_sc_hd__clkbuf_16
Xfanout232 _6290_/Q vssd1 vssd1 vccd1 vccd1 _5625_/A sky130_fd_sc_hd__buf_6
Xfanout243 _5862_/A vssd1 vssd1 vccd1 vccd1 _3942_/A sky130_fd_sc_hd__buf_8
Xfanout254 _6237_/Q vssd1 vssd1 vccd1 vccd1 _3942_/D sky130_fd_sc_hd__buf_8
Xfanout265 _4085_/A vssd1 vssd1 vccd1 vccd1 _3943_/C sky130_fd_sc_hd__buf_6
Xfanout276 _6226_/Q vssd1 vssd1 vccd1 vccd1 _5480_/B sky130_fd_sc_hd__clkbuf_16
XFILLER_47_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5422__S _5456_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout287 _5768_/A0 vssd1 vssd1 vccd1 vccd1 _5256_/B sky130_fd_sc_hd__buf_2
XFILLER_87_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout298 _6070_/Q vssd1 vssd1 vccd1 vccd1 _4622_/B sky130_fd_sc_hd__buf_12
XANTENNA__4806__A0 _5714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3450__B _3986_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4038__S _4044_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4265__C _4309_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_591 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3178__A _3970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5096__C _5096_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4337__A2 _4167_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5534__A1 _5595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5837__A2 _3971_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3848__A1 _3594_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4830_ _6189_/Q _5539_/S vssd1 vssd1 vccd1 vccd1 _4830_/X sky130_fd_sc_hd__and2_1
XFILLER_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4761_ _3011_/Y _4643_/Y _4760_/X _4638_/B vssd1 vssd1 vccd1 vccd1 _4761_/X sky130_fd_sc_hd__o2bb2a_1
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3712_ _6027_/Q _3711_/X _3731_/S vssd1 vssd1 vccd1 vccd1 _6027_/D sky130_fd_sc_hd__mux2_1
X_4692_ _4692_/A _4692_/B vssd1 vssd1 vccd1 vccd1 _4692_/Y sky130_fd_sc_hd__nor2_1
XFILLER_119_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5525__A1 _5498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3643_ _3643_/A _3643_/B vssd1 vssd1 vccd1 vccd1 _3643_/Y sky130_fd_sc_hd__xnor2_2
XANTENNA__5525__B2 _4645_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3816__A _4767_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3574_ _3621_/A _3574_/B _3619_/A vssd1 vssd1 vccd1 vccd1 _3574_/X sky130_fd_sc_hd__or3b_1
XFILLER_115_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5313_ _5464_/A _5312_/A _5607_/B1 vssd1 vssd1 vccd1 vccd1 _5313_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_114_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6293_ _6293_/CLK _6293_/D vssd1 vssd1 vccd1 vccd1 _6293_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__3254__C _4614_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5244_ _5244_/A _5244_/B _5463_/A vssd1 vssd1 vccd1 vccd1 _5244_/X sky130_fd_sc_hd__and3_1
XFILLER_103_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3839__A1 _4846_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4647__A _6184_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5175_ _5050_/C _5166_/Y _5170_/Y _5174_/X _3014_/A vssd1 vssd1 vccd1 vccd1 _5175_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_84_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4126_ _4126_/A _4126_/B vssd1 vssd1 vccd1 vccd1 _4126_/X sky130_fd_sc_hd__or2_1
XFILLER_84_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4366__B _4389_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4057_ _5436_/A _4058_/B _5742_/C vssd1 vssd1 vccd1 vccd1 _4057_/Y sky130_fd_sc_hd__nor3_2
XFILLER_83_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3008_ _5547_/B vssd1 vssd1 vccd1 vccd1 _3008_/Y sky130_fd_sc_hd__inv_2
XFILLER_71_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3697__S _3902_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3472__C1 _3511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5213__A0 _5255_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4016__A1 _6295_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_675 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4016__B2 _6300_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5764__A1 _4891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4959_ _5509_/C _4959_/B vssd1 vssd1 vccd1 vccd1 _4959_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__3775__A0 _5848_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5516__A1 _5607_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5941__A _5948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3164__C _3164_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3180__B _5065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4255__A1 _3718_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5204__B1 _5097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4191__B1 _4072_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3290_ _6009_/Q _6008_/Q vssd1 vssd1 vccd1 vccd1 _3561_/A sky130_fd_sc_hd__nand2b_4
XFILLER_111_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4494__A1 _5385_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4246__A1 _3730_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5931_ _5767_/A _5930_/Y _5931_/S vssd1 vssd1 vccd1 vccd1 _5932_/B sky130_fd_sc_hd__mux2_1
XANTENNA__4797__A2 _4587_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5862_ _5862_/A _5862_/B vssd1 vssd1 vccd1 vccd1 _5862_/Y sky130_fd_sc_hd__nand2_1
XFILLER_61_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4813_ _4972_/A _4806_/X _4812_/X _3740_/A vssd1 vssd1 vccd1 vccd1 _4813_/X sky130_fd_sc_hd__a22o_2
X_5793_ _6259_/Q _3715_/X _5798_/S vssd1 vssd1 vccd1 vccd1 _6259_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4930__A _5034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4744_ _6217_/Q _4744_/B vssd1 vssd1 vccd1 vccd1 _4745_/A sky130_fd_sc_hd__nand2_8
XFILLER_30_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4675_ _4675_/A _4678_/B vssd1 vssd1 vccd1 vccd1 _4676_/C sky130_fd_sc_hd__or2_1
XANTENNA__3546__A _3599_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3626_ _3365_/B _5898_/A _3625_/X _3312_/B _3145_/C vssd1 vssd1 vccd1 vccd1 _3626_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout112_A _3500_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput19 _6193_/Q vssd1 vssd1 vccd1 vccd1 io_out[17] sky130_fd_sc_hd__buf_4
X_3557_ _3557_/A _3557_/B vssd1 vssd1 vccd1 vccd1 _3557_/X sky130_fd_sc_hd__or2_4
X_6276_ _6280_/CLK _6276_/D vssd1 vssd1 vccd1 vccd1 _6276_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3488_ _6016_/Q _6039_/Q _3709_/S vssd1 vssd1 vccd1 vccd1 _3488_/X sky130_fd_sc_hd__mux2_8
XFILLER_103_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5480__B _5480_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5227_ _5227_/A _5227_/B vssd1 vssd1 vccd1 vccd1 _5227_/Y sky130_fd_sc_hd__nor2_4
XFILLER_88_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4485__A1 _5305_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3288__A2 _3287_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5682__B1 _5353_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5158_ _5158_/A _5158_/B _5158_/C _5158_/D vssd1 vssd1 vccd1 vccd1 _5158_/X sky130_fd_sc_hd__or4_1
XANTENNA__4096__B _4136_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4109_ _4163_/A _4173_/B vssd1 vssd1 vccd1 vccd1 _4110_/B sky130_fd_sc_hd__nand2_1
X_5089_ _4644_/A _5088_/X _5086_/X vssd1 vssd1 vccd1 vccd1 _5090_/B sky130_fd_sc_hd__o21ai_1
XFILLER_44_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4788__A2 _5172_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5936__A _5936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4960__A2 _4647_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3175__B _3312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5390__B _5392_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3279__A2 _3257_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3191__A _4622_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4734__B _4734_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_759 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3130__S _3135_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3451__A2 _3986_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5189__C1 _5071_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4460_ _5790_/A1 _3900_/Y _4458_/X _4459_/X vssd1 vssd1 vccd1 vccd1 _6124_/D sky130_fd_sc_hd__a22o_1
XFILLER_7_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3411_ _3465_/A _3926_/A vssd1 vssd1 vccd1 vccd1 _3925_/A sky130_fd_sc_hd__nor2_2
X_4391_ _4391_/A _4391_/B vssd1 vssd1 vccd1 vccd1 _4393_/C sky130_fd_sc_hd__nor2_2
XANTENNA__4703__A2 _6184_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6130_ _6154_/CLK _6130_/D vssd1 vssd1 vccd1 vccd1 _6130_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3342_ _4657_/A _3549_/B _3398_/A _3341_/X vssd1 vssd1 vccd1 vccd1 _3342_/X sky130_fd_sc_hd__o211a_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6061_ _6098_/CLK _6061_/D vssd1 vssd1 vccd1 vccd1 _6061_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4197__A _4197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3273_ _4096_/A _3257_/B _5263_/B _3885_/A vssd1 vssd1 vccd1 vccd1 _3274_/B sky130_fd_sc_hd__a22o_2
XFILLER_98_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5012_ _6195_/Q _4647_/B _4648_/Y _6006_/Q _5227_/B vssd1 vssd1 vccd1 vccd1 _5012_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4628__C _4665_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5020__A1_N _5547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4644__B _4644_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5914_ _3105_/A _5075_/B _5635_/A _3881_/B _5191_/A vssd1 vssd1 vccd1 vccd1 _5914_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__5719__A1 _4837_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5845_ _5845_/A vssd1 vssd1 vccd1 vccd1 _5846_/B sky130_fd_sc_hd__inv_2
XFILLER_22_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout327_A _5072_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5776_ _6253_/Q _5788_/B vssd1 vssd1 vccd1 vccd1 _5776_/X sky130_fd_sc_hd__or2_1
X_4727_ _4727_/A _4727_/B vssd1 vssd1 vccd1 vccd1 _4727_/Y sky130_fd_sc_hd__nor2_1
XFILLER_135_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4658_ _5108_/A _4658_/B vssd1 vssd1 vccd1 vccd1 _4660_/A sky130_fd_sc_hd__xnor2_4
XFILLER_107_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3609_ _3644_/B _3615_/B _3606_/Y _3561_/A _3608_/X vssd1 vssd1 vccd1 vccd1 _4846_/B
+ sky130_fd_sc_hd__o221a_4
XFILLER_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5491__A _5551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4589_ _4589_/A vssd1 vssd1 vccd1 vccd1 _4589_/Y sky130_fd_sc_hd__inv_2
XFILLER_89_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4819__B _4819_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6259_ _6259_/CLK _6259_/D vssd1 vssd1 vccd1 vccd1 _6259_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5958__A1 _3112_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3186__A _3974_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3914__A _4438_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4167__D _4167_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4745__A _4745_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3960_ _5634_/A _3960_/B _3960_/C vssd1 vssd1 vccd1 vccd1 _3978_/B sky130_fd_sc_hd__or3_2
XFILLER_50_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3891_ _4604_/A _4604_/B _5928_/B _5911_/C vssd1 vssd1 vccd1 vccd1 _3953_/A sky130_fd_sc_hd__or4_1
XFILLER_31_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5630_ _3867_/A _3388_/B _5628_/X _5629_/X _3996_/B vssd1 vssd1 vccd1 vccd1 _5630_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5295__B _5296_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5561_ _5567_/A _5040_/Y _5561_/S vssd1 vssd1 vccd1 vccd1 _5561_/X sky130_fd_sc_hd__mux2_2
XFILLER_117_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4512_ _6153_/Q _4515_/B vssd1 vssd1 vccd1 vccd1 _4512_/X sky130_fd_sc_hd__or2_1
X_5492_ _5551_/A _5482_/Y _5491_/Y _3122_/A vssd1 vssd1 vccd1 vccd1 _5494_/B sky130_fd_sc_hd__a211o_1
XFILLER_8_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4443_ _6119_/Q _4458_/B vssd1 vssd1 vccd1 vccd1 _4443_/X sky130_fd_sc_hd__or2_1
XANTENNA__5742__C _5742_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4374_ _4375_/A _4375_/B vssd1 vssd1 vccd1 vccd1 _4376_/A sky130_fd_sc_hd__nand2_1
XANTENNA__4639__B _4643_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3325_ _6011_/Q _3231_/Y _3323_/X vssd1 vssd1 vccd1 vccd1 _6011_/D sky130_fd_sc_hd__o21a_1
X_6113_ _6113_/CLK _6113_/D vssd1 vssd1 vccd1 vccd1 _6113_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6044_ _6295_/CLK _6044_/D vssd1 vssd1 vccd1 vccd1 _6044_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3256_ _3251_/B _3250_/X _3251_/Y _3255_/Y vssd1 vssd1 vccd1 vccd1 _3256_/X sky130_fd_sc_hd__o211a_1
XANTENNA__5101__A2 _5097_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4077__D _4176_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3187_ _5622_/A _5635_/A vssd1 vssd1 vccd1 vccd1 _3215_/B sky130_fd_sc_hd__nand2_1
XANTENNA_fanout277_A _4872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5828_ _5835_/A1 _4405_/Y _5819_/Y _6277_/Q vssd1 vssd1 vccd1 vccd1 _5828_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5168__A2 _5169_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5759_ _5387_/A _5761_/S _5791_/A vssd1 vssd1 vccd1 vccd1 _5759_/X sky130_fd_sc_hd__o21a_1
XFILLER_5_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4128__B1 _4072_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4679__A1 _4678_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3734__A _3734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout92_A _5058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3351__A1 _4658_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4565__A _5238_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4851__A1 _4886_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3900__C _5743_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3406__A2 _3500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4906__A2 _5093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3590__A1 _3590_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3644__A _3986_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5331__A2 _5330_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3342__A1 _4657_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5619__B1 _4648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3110_ _5075_/B _3111_/B vssd1 vssd1 vccd1 vccd1 _4654_/A sky130_fd_sc_hd__nor2_4
XFILLER_68_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4090_ _4103_/A _4090_/B vssd1 vssd1 vccd1 vccd1 _4090_/X sky130_fd_sc_hd__and2_1
XFILLER_95_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3041_ _6007_/Q vssd1 vssd1 vccd1 vccd1 _3041_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5398__A2 _5509_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4992_ _5330_/B _4992_/B vssd1 vssd1 vccd1 vccd1 _4992_/Y sky130_fd_sc_hd__nand2_1
XFILLER_90_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3943_ _3943_/A _5109_/A _3943_/C _3943_/D vssd1 vssd1 vccd1 vccd1 _3944_/B sky130_fd_sc_hd__or4_1
XANTENNA__4070__A2 _4614_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3874_ _3951_/C _3892_/B vssd1 vssd1 vccd1 vccd1 _3966_/B sky130_fd_sc_hd__nor2_2
XFILLER_137_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5613_ _6233_/Q _5250_/X _5612_/X _5948_/A vssd1 vssd1 vccd1 vccd1 _6233_/D sky130_fd_sc_hd__o211a_1
Xclkbuf_3_2__f_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_9_clk/A sky130_fd_sc_hd__clkbuf_16
X_5544_ _4645_/B _5542_/X _5543_/X _3121_/B vssd1 vssd1 vccd1 vccd1 _5544_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_117_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5307__C1 _3060_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3581__A1 _3145_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5475_ _5453_/A _5453_/B _5451_/A vssd1 vssd1 vccd1 vccd1 _5476_/B sky130_fd_sc_hd__o21a_2
XFILLER_105_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5858__B1 _5857_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3318__D1 _4003_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4426_ _4426_/A _4426_/B _4426_/C vssd1 vssd1 vccd1 vccd1 _4428_/A sky130_fd_sc_hd__and3_2
XFILLER_120_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4357_ _4358_/A _4358_/B _4358_/C vssd1 vssd1 vccd1 vccd1 _4383_/S sky130_fd_sc_hd__a21oi_4
XFILLER_59_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3308_ _5889_/A vssd1 vssd1 vccd1 vccd1 _3308_/Y sky130_fd_sc_hd__inv_2
X_4288_ _4225_/A _4225_/B _4225_/C vssd1 vssd1 vccd1 vccd1 _4289_/C sky130_fd_sc_hd__a21bo_2
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5086__A1 _6198_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3239_ _3240_/A _3241_/B vssd1 vssd1 vccd1 vccd1 _3239_/X sky130_fd_sc_hd__or2_4
X_6027_ _6262_/CLK _6027_/D vssd1 vssd1 vccd1 vccd1 _6027_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4833__B2 _5069_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5928__B _5928_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout43 _5867_/A1 vssd1 vssd1 vccd1 vccd1 _5854_/A sky130_fd_sc_hd__buf_4
XFILLER_23_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout54 _3834_/B vssd1 vssd1 vccd1 vccd1 _3845_/B sky130_fd_sc_hd__clkbuf_4
Xfanout65 _4601_/Y vssd1 vssd1 vccd1 vccd1 _5058_/C sky130_fd_sc_hd__buf_6
XFILLER_10_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout76 _3194_/Y vssd1 vssd1 vccd1 vccd1 _5943_/A sky130_fd_sc_hd__clkbuf_4
Xfanout87 _5570_/A vssd1 vssd1 vccd1 vccd1 _4604_/A sky130_fd_sc_hd__buf_6
XANTENNA__3448__B _3450_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout98 _3058_/Y vssd1 vssd1 vccd1 vccd1 _5172_/A sky130_fd_sc_hd__buf_2
XANTENNA__4270__D _4410_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4521__A0 _5790_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3911__B _5766_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3590_ _3590_/A1 _3587_/X _3588_/X _3589_/X vssd1 vssd1 vccd1 vccd1 _3590_/X sky130_fd_sc_hd__a22o_4
XANTENNA__5552__A2 _5542_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3563__A1 _4808_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5260_ _4642_/A _5257_/B _5259_/Y vssd1 vssd1 vccd1 vccd1 _5260_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4211_ _4210_/B _4210_/C _4210_/A vssd1 vssd1 vccd1 vccd1 _4221_/B sky130_fd_sc_hd__o21ai_4
X_5191_ _5191_/A _6214_/Q _5195_/C vssd1 vssd1 vccd1 vccd1 _5192_/C sky130_fd_sc_hd__and3_1
X_4142_ _4270_/A _4111_/B _4114_/B _4112_/X vssd1 vssd1 vccd1 vccd1 _4145_/A sky130_fd_sc_hd__a31o_4
XFILLER_122_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5068__A1 _6197_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4073_ _4136_/A _3709_/X _4233_/A1 _4069_/Y vssd1 vssd1 vccd1 vccd1 _4073_/X sky130_fd_sc_hd__a31o_1
XFILLER_95_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3024_ _3948_/A vssd1 vssd1 vccd1 vccd1 _3024_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4975_ _6005_/Q _4947_/Y _4973_/Y _4974_/X vssd1 vssd1 vccd1 vccd1 _4975_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_51_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3549__A _5392_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3926_ _3926_/A _3926_/B _3926_/C vssd1 vssd1 vccd1 vccd1 _3926_/X sky130_fd_sc_hd__or3_1
XFILLER_32_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3268__B _3388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3857_ _3880_/A _5883_/A _3952_/B vssd1 vssd1 vccd1 vccd1 _3964_/B sky130_fd_sc_hd__nand3_4
XFILLER_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3788_ _3450_/D _3738_/X _3801_/B _3787_/X vssd1 vssd1 vccd1 vccd1 _3788_/X sky130_fd_sc_hd__o211a_1
XANTENNA__4751__B1 _3116_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5527_ _5547_/B _5547_/C vssd1 vssd1 vccd1 vccd1 _5527_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__3263__C_N _4136_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5458_ _5498_/A _5463_/B _5457_/X _5570_/A vssd1 vssd1 vccd1 vccd1 _5458_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_132_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4503__A0 _3943_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4409_ _4410_/B _4426_/B _4410_/D _4426_/A vssd1 vssd1 vccd1 vccd1 _4411_/A sky130_fd_sc_hd__a22oi_4
Xfanout200 _3148_/X vssd1 vssd1 vccd1 vccd1 _3922_/S sky130_fd_sc_hd__buf_6
XFILLER_59_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5700__C1 _5728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5389_ _5420_/B _5389_/B vssd1 vssd1 vccd1 vccd1 _5389_/Y sky130_fd_sc_hd__nor2_4
Xfanout211 _3044_/Y vssd1 vssd1 vccd1 vccd1 _5733_/A sky130_fd_sc_hd__buf_4
XFILLER_114_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout222 _3766_/A vssd1 vssd1 vccd1 vccd1 _3713_/S sky130_fd_sc_hd__buf_6
Xfanout233 _6290_/Q vssd1 vssd1 vccd1 vccd1 _5840_/A sky130_fd_sc_hd__clkbuf_16
Xfanout244 _5862_/A vssd1 vssd1 vccd1 vccd1 _4410_/B sky130_fd_sc_hd__buf_8
XFILLER_113_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout255 _4301_/A vssd1 vssd1 vccd1 vccd1 _4162_/A sky130_fd_sc_hd__buf_8
XFILLER_115_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout266 _4197_/B vssd1 vssd1 vccd1 vccd1 _4136_/A sky130_fd_sc_hd__buf_6
Xfanout277 _4872_/A vssd1 vssd1 vccd1 vccd1 _5446_/B sky130_fd_sc_hd__buf_6
XFILLER_86_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout288 _6219_/Q vssd1 vssd1 vccd1 vccd1 _5768_/A0 sky130_fd_sc_hd__buf_4
XFILLER_46_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout299 _6069_/Q vssd1 vssd1 vccd1 vccd1 _3312_/A sky130_fd_sc_hd__buf_12
XFILLER_101_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3609__A2 _3615_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3450__C _3500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout55_A _5742_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4265__D _4342_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5231__A1 _5075_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3178__B _4577_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3194__A _3960_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6219__CLK _6219_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3133__S _3135_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output36_A _6184_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5849__A _5849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4753__A _4753_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3481__B1 _3589_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5222__A1 _5625_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4760_ _4640_/A _4756_/X _4759_/X vssd1 vssd1 vccd1 vccd1 _4760_/X sky130_fd_sc_hd__o21a_1
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3711_ _6011_/Q _3706_/Y _3710_/X vssd1 vssd1 vccd1 vccd1 _3711_/X sky130_fd_sc_hd__a21o_4
XANTENNA__3784__A1 _4096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4691_ _4691_/A _4691_/B vssd1 vssd1 vccd1 vccd1 _4692_/B sky130_fd_sc_hd__nand2_1
XFILLER_119_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3642_ _3649_/B _3642_/B vssd1 vssd1 vccd1 vccd1 _3642_/Y sky130_fd_sc_hd__xnor2_2
XANTENNA__3536__B2 _3590_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3573_ _3572_/A _3572_/C _3935_/D vssd1 vssd1 vccd1 vccd1 _3619_/A sky130_fd_sc_hd__a21o_1
X_5312_ _5312_/A _5312_/B vssd1 vssd1 vccd1 vccd1 _5312_/X sky130_fd_sc_hd__or2_1
XFILLER_127_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6292_ _6302_/CLK _6292_/D vssd1 vssd1 vccd1 vccd1 _6292_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__5289__A1 _5292_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5243_ _3672_/Y _5097_/B _3118_/Y vssd1 vssd1 vccd1 vccd1 _5250_/B sky130_fd_sc_hd__a21o_1
XFILLER_102_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5523__S _5543_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3839__A2 _3740_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3395__S0 _4067_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5174_ _5171_/X _5172_/Y _5173_/Y _5494_/A vssd1 vssd1 vccd1 vccd1 _5174_/X sky130_fd_sc_hd__o31a_1
XANTENNA__4647__B _4647_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4125_ _4125_/A _4125_/B vssd1 vssd1 vccd1 vccd1 _4126_/B sky130_fd_sc_hd__and2_1
XFILLER_68_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4056_ _5436_/A _4058_/B _5767_/C vssd1 vssd1 vccd1 vccd1 _4476_/S sky130_fd_sc_hd__or3_4
XFILLER_83_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5461__A1 _5507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3007_ _4197_/B vssd1 vssd1 vccd1 vccd1 _3251_/A sky130_fd_sc_hd__inv_2
XFILLER_83_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4663__A _5263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5213__A1 _4634_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4016__A2 _3030_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4958_ _4954_/X _4957_/Y _5050_/B vssd1 vssd1 vccd1 vccd1 _4958_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3909_ _6049_/Q _3730_/X _3909_/S vssd1 vssd1 vccd1 vccd1 _6049_/D sky130_fd_sc_hd__mux2_1
XFILLER_20_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4889_ _4745_/A _4887_/X _4896_/B _3093_/Y _5050_/B vssd1 vssd1 vccd1 vccd1 _4889_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5494__A _5494_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3742__A _3948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3463__B1 _3621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_52_clk_A _6133_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5204__A1 _5136_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4007__A2 _5561_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3189__A _3766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3128__S _3135_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4748__A _5333_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5691__A1 _5730_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3371__B _3575_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5443__A1 _5943_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5930_ _3948_/A _5925_/Y _5929_/X vssd1 vssd1 vccd1 vccd1 _5930_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_18_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5861_ _6286_/Q _5867_/A1 _5860_/Y _5866_/B1 vssd1 vssd1 vccd1 vccd1 _6286_/D sky130_fd_sc_hd__o211a_1
XFILLER_80_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4812_ _5714_/A _4811_/Y _4812_/S vssd1 vssd1 vccd1 vccd1 _4812_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5792_ _6258_/Q _3711_/X _5798_/S vssd1 vssd1 vccd1 vccd1 _6258_/D sky130_fd_sc_hd__mux2_1
XFILLER_22_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3757__A1 _3986_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4743_ _4814_/C _4743_/B vssd1 vssd1 vccd1 vccd1 _4743_/X sky130_fd_sc_hd__or2_1
XFILLER_119_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4674_ _4675_/A _4678_/B vssd1 vssd1 vccd1 vccd1 _4710_/B sky130_fd_sc_hd__nand2_1
XANTENNA__3509__A1 _5707_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3546__B _5707_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3625_ _6207_/Q _3615_/B _3658_/S vssd1 vssd1 vccd1 vccd1 _3625_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3556_ _3557_/A _3557_/B vssd1 vssd1 vccd1 vccd1 _3607_/B sky130_fd_sc_hd__nor2_8
XFILLER_115_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6275_ _6280_/CLK _6275_/D vssd1 vssd1 vccd1 vccd1 _6275_/Q sky130_fd_sc_hd__dfxtp_1
X_3487_ _4202_/A _3136_/Y _5392_/B _3053_/X vssd1 vssd1 vccd1 vccd1 _3492_/A sky130_fd_sc_hd__a22o_4
XFILLER_102_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5226_ _5226_/A _5454_/B _5264_/B vssd1 vssd1 vccd1 vccd1 _5226_/X sky130_fd_sc_hd__and3_1
XFILLER_102_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5682__A1 _5710_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5682__B2 _5734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3693__A0 _5333_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5157_ _4593_/Y _5144_/X _3116_/X vssd1 vssd1 vccd1 vccd1 _5158_/D sky130_fd_sc_hd__o21a_1
XFILLER_29_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4096__C _4311_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4108_ _4108_/A _4108_/B vssd1 vssd1 vccd1 vccd1 _4110_/A sky130_fd_sc_hd__nor2_2
XFILLER_110_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5088_ _6198_/Q _4646_/Y _5087_/X _5072_/A _5403_/A vssd1 vssd1 vccd1 vccd1 _5088_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__5434__A1 _4644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5434__B2 _5464_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4039_ _6060_/Q _3715_/X _4044_/S vssd1 vssd1 vccd1 vccd1 _6060_/D sky130_fd_sc_hd__mux2_1
XFILLER_37_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5936__B _5943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3456__B _3458_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3920__A1 _3727_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4568__A _5244_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5673__A1 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3191__B _6071_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4242__S _4246_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5862__A _5862_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3085__C _5058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3410_ _6203_/Q _3410_/B vssd1 vssd1 vccd1 vccd1 _3926_/A sky130_fd_sc_hd__nor2_2
X_4390_ _4426_/A _4389_/B _4389_/C vssd1 vssd1 vccd1 vccd1 _4391_/B sky130_fd_sc_hd__a21oi_1
X_3341_ _3636_/A _4619_/A vssd1 vssd1 vccd1 vccd1 _3341_/X sky130_fd_sc_hd__or2_1
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6060_ _6248_/CLK _6060_/D vssd1 vssd1 vccd1 vccd1 _6060_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4197__B _4197_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3272_ _6274_/Q _6110_/Q _3551_/S vssd1 vssd1 vccd1 vccd1 _5263_/B sky130_fd_sc_hd__mux2_8
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5664__A1 _4096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5011_ _5509_/C _5011_/B vssd1 vssd1 vccd1 vccd1 _5011_/Y sky130_fd_sc_hd__nor2_1
XFILLER_87_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3427__B1 _3589_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3321__S _3511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5913_ _3880_/B _4604_/C _3877_/B _5959_/A vssd1 vssd1 vccd1 vccd1 _5919_/B sky130_fd_sc_hd__a31o_1
XFILLER_34_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5844_ _3274_/X _5935_/A0 _5862_/B vssd1 vssd1 vccd1 vccd1 _5845_/A sky130_fd_sc_hd__mux2_8
XFILLER_34_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5775_ _5926_/A0 _4250_/Y _5773_/X _5774_/Y vssd1 vssd1 vccd1 vccd1 _6252_/D sky130_fd_sc_hd__a22o_1
XANTENNA_fanout222_A _3766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4726_ _5114_/A _4726_/B vssd1 vssd1 vccd1 vccd1 _4727_/B sky130_fd_sc_hd__and2_2
X_4657_ _4657_/A _4658_/B vssd1 vssd1 vccd1 vccd1 _4657_/X sky130_fd_sc_hd__and2_1
XFILLER_107_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3608_ _3608_/A _3611_/B vssd1 vssd1 vccd1 vccd1 _3608_/X sky130_fd_sc_hd__or2_1
X_4588_ _5090_/A _5095_/A vssd1 vssd1 vccd1 vccd1 _4589_/A sky130_fd_sc_hd__or2_4
XFILLER_122_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3539_ _3567_/B _3593_/B vssd1 vssd1 vccd1 vccd1 _3540_/B sky130_fd_sc_hd__nor2_1
XFILLER_115_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6258_ _6258_/CLK _6258_/D vssd1 vssd1 vccd1 vccd1 _6258_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5655__A1 _5454_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5209_ _5206_/B _5207_/X _5208_/X vssd1 vssd1 vccd1 vccd1 _5209_/X sky130_fd_sc_hd__o21a_1
X_6189_ _6288_/CLK _6189_/D vssd1 vssd1 vccd1 vccd1 _6189_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_69_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4863__C1 _4852_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5407__B2 _3236_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5958__A2 _3975_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4091__B1 _4072_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5460__B1_N _5227_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4062__S _4066_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5646__A1 _4577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3890_ _5138_/A _5137_/D _3966_/B vssd1 vssd1 vccd1 vccd1 _5959_/B sky130_fd_sc_hd__or3_2
XANTENNA__4385__B2 _4437_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5560_ _6007_/Q _5560_/B vssd1 vssd1 vccd1 vccd1 _5560_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3096__B _4744_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4511_ _3942_/D _3912_/Y _4509_/X _4510_/Y vssd1 vssd1 vccd1 vccd1 _6152_/D sky130_fd_sc_hd__a22o_1
X_5491_ _5551_/A _5491_/B vssd1 vssd1 vccd1 vccd1 _5491_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__4700__S _4812_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4442_ _5935_/A0 _3900_/Y _4440_/X _4441_/X vssd1 vssd1 vccd1 vccd1 _6118_/D sky130_fd_sc_hd__a22o_1
X_4373_ _4373_/A _4373_/B vssd1 vssd1 vccd1 vccd1 _4375_/B sky130_fd_sc_hd__xor2_1
XANTENNA__3896__A0 _5859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6112_ _6113_/CLK _6112_/D vssd1 vssd1 vccd1 vccd1 _6112_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3324_ _3324_/A _4614_/B vssd1 vssd1 vccd1 vccd1 _5138_/A sky130_fd_sc_hd__nand2_4
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6043_ _6262_/CLK _6043_/D vssd1 vssd1 vccd1 vccd1 _6043_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3255_ _3255_/A _5799_/B vssd1 vssd1 vccd1 vccd1 _3255_/Y sky130_fd_sc_hd__nand2_4
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3186_ _3974_/B _3677_/B vssd1 vssd1 vccd1 vccd1 _3940_/A sky130_fd_sc_hd__nor2_4
XFILLER_66_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout172_A _5638_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5767__A _5767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4671__A _4672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3820__B1 _3484_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5827_ _3477_/Y _5819_/B _5826_/X vssd1 vssd1 vccd1 vccd1 _6276_/D sky130_fd_sc_hd__a21o_1
XANTENNA__5168__A3 _4604_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3287__A _3287_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5758_ _6247_/Q _5763_/B vssd1 vssd1 vccd1 vccd1 _5758_/X sky130_fd_sc_hd__or2_1
XFILLER_136_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4709_ _4710_/A _4710_/B _4713_/A vssd1 vssd1 vccd1 vccd1 _4750_/B sky130_fd_sc_hd__a21o_1
XFILLER_108_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5689_ _4772_/B _4767_/B _5703_/A vssd1 vssd1 vccd1 vccd1 _5690_/B sky130_fd_sc_hd__mux2_1
XFILLER_1_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5628__A1 _6295_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout85_A _3090_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4846__A _4846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3750__A _5617_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4565__B _4753_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_866 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3896__S _4643_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3811__A0 _3593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3197__A _3873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4367__A1 _4410_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5867__A1 _5867_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5619__A1 _5622_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3040_ _6004_/Q vssd1 vssd1 vccd1 vccd1 _4943_/B sky130_fd_sc_hd__inv_2
XFILLER_48_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4991_ _6194_/Q _4990_/A _4640_/Y _4990_/Y vssd1 vssd1 vccd1 vccd1 _4991_/X sky130_fd_sc_hd__o211a_1
XFILLER_16_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3942_ _3942_/A _3942_/B _5856_/A _3942_/D vssd1 vssd1 vccd1 vccd1 _3943_/D sky130_fd_sc_hd__or4_1
XANTENNA__3802__B1 _3777_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3819__B _3819_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3873_ _3873_/A _3893_/C vssd1 vssd1 vccd1 vccd1 _3892_/B sky130_fd_sc_hd__or2_2
X_5612_ _5412_/A _5598_/Y _5607_/X _5611_/X _5251_/Y vssd1 vssd1 vccd1 vccd1 _5612_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5555__B1 _5556_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5543_ _5344_/A _6006_/Q _5543_/S vssd1 vssd1 vccd1 vccd1 _5543_/X sky130_fd_sc_hd__mux2_1
X_5474_ _4891_/A _5251_/A _5473_/Y _5948_/A vssd1 vssd1 vccd1 vccd1 _6226_/D sky130_fd_sc_hd__o211a_1
XANTENNA__3318__C1 _4003_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4425_ _4426_/A _4426_/B vssd1 vssd1 vccd1 vccd1 _4425_/Y sky130_fd_sc_hd__nand2_1
XFILLER_99_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4356_ _4382_/B _4356_/B vssd1 vssd1 vccd1 vccd1 _4358_/C sky130_fd_sc_hd__or2_2
XFILLER_98_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3307_ _3575_/B _3267_/A _3267_/B _3306_/Y vssd1 vssd1 vccd1 vccd1 _5889_/A sky130_fd_sc_hd__a31o_4
XFILLER_98_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4287_ _4326_/A _4285_/Y _4214_/X _4218_/A vssd1 vssd1 vccd1 vccd1 _4289_/B sky130_fd_sc_hd__a211o_2
XFILLER_98_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5086__A2 _5870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6026_ _6257_/CLK _6026_/D vssd1 vssd1 vccd1 vccd1 _6026_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3238_ _5924_/A _6059_/Q _5436_/C vssd1 vssd1 vccd1 vccd1 _3238_/X sky130_fd_sc_hd__and3_1
XFILLER_74_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3169_ _6217_/Q _5143_/A vssd1 vssd1 vccd1 vccd1 _4592_/B sky130_fd_sc_hd__nor2_4
XTAP_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout44 _5839_/X vssd1 vssd1 vccd1 vccd1 _5867_/A1 sky130_fd_sc_hd__buf_8
XFILLER_22_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout55 _5742_/C vssd1 vssd1 vccd1 vccd1 _5743_/C sky130_fd_sc_hd__buf_8
Xfanout66 _4601_/Y vssd1 vssd1 vccd1 vccd1 _5412_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_80_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout77 _3121_/X vssd1 vssd1 vccd1 vccd1 _5498_/A sky130_fd_sc_hd__buf_6
Xfanout88 _5570_/A vssd1 vssd1 vccd1 vccd1 _5959_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__5546__B1 _5551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout99 _3060_/B vssd1 vssd1 vccd1 vccd1 _5507_/A sky130_fd_sc_hd__buf_6
XFILLER_10_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3745__A _5503_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4576__A _4576_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3480__A _5924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4760__A1 _4640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5870__A _5870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4210_ _4210_/A _4210_/B _4210_/C vssd1 vssd1 vccd1 vccd1 _4221_/A sky130_fd_sc_hd__or3_4
XANTENNA__5170__D1 _3880_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5190_ _5191_/A _5195_/C _6214_/Q vssd1 vssd1 vccd1 vccd1 _5192_/B sky130_fd_sc_hd__a21oi_1
XFILLER_96_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4141_ _4202_/A _4173_/B vssd1 vssd1 vccd1 vccd1 _4146_/A sky130_fd_sc_hd__nand2_2
XFILLER_68_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5068__A2 _5238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4072_ _5936_/A _4072_/B _4072_/C _5138_/A vssd1 vssd1 vccd1 vccd1 _4072_/Y sky130_fd_sc_hd__nor4b_4
XFILLER_110_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5473__C1 _5251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3023_ _3869_/A vssd1 vssd1 vccd1 vccd1 _3197_/B sky130_fd_sc_hd__inv_2
XFILLER_83_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4974_ _4974_/A _6004_/Q _6005_/Q vssd1 vssd1 vccd1 vccd1 _4974_/X sky130_fd_sc_hd__and3_2
XFILLER_52_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5110__A _5110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3925_ _3925_/A _3926_/C vssd1 vssd1 vccd1 vccd1 _3925_/X sky130_fd_sc_hd__or2_2
XFILLER_32_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3856_ _4642_/A _5883_/A _3952_/B vssd1 vssd1 vccd1 vccd1 _3856_/X sky130_fd_sc_hd__and3_2
XFILLER_20_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout135_A _3084_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3787_ _4697_/A _3845_/B _3737_/Y _3786_/Y vssd1 vssd1 vccd1 vccd1 _3787_/X sky130_fd_sc_hd__a211o_1
XFILLER_118_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5526_ _3059_/Y _5520_/X _5525_/X vssd1 vssd1 vccd1 vccd1 _5526_/X sky130_fd_sc_hd__a21o_1
XFILLER_106_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout302_A _4642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5457_ _4644_/B _5464_/B _5456_/X _4646_/A vssd1 vssd1 vccd1 vccd1 _5457_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_59_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4408_ _4388_/A _4426_/C _4391_/A vssd1 vssd1 vccd1 vccd1 _4413_/A sky130_fd_sc_hd__o21bai_4
X_5388_ _5387_/B _5387_/C _5387_/A vssd1 vssd1 vccd1 vccd1 _5389_/B sky130_fd_sc_hd__a21oi_2
Xfanout201 _3869_/B vssd1 vssd1 vccd1 vccd1 _3658_/S sky130_fd_sc_hd__buf_6
XFILLER_120_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout212 _3025_/Y vssd1 vssd1 vccd1 vccd1 _4963_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_59_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout223 _6297_/Q vssd1 vssd1 vccd1 vccd1 _3766_/A sky130_fd_sc_hd__buf_8
XFILLER_132_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4339_ _4302_/A _4302_/B _4305_/A vssd1 vssd1 vccd1 vccd1 _4340_/B sky130_fd_sc_hd__o21bai_2
XFILLER_86_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout234 _6290_/Q vssd1 vssd1 vccd1 vccd1 _5883_/A sky130_fd_sc_hd__buf_6
Xfanout245 _5862_/A vssd1 vssd1 vccd1 vccd1 _4214_/A sky130_fd_sc_hd__buf_6
Xfanout256 _6237_/Q vssd1 vssd1 vccd1 vccd1 _4301_/A sky130_fd_sc_hd__buf_12
Xfanout267 _4085_/A vssd1 vssd1 vccd1 vccd1 _4197_/B sky130_fd_sc_hd__buf_8
Xfanout278 _6225_/Q vssd1 vssd1 vccd1 vccd1 _4872_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_75_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout289 _6213_/Q vssd1 vssd1 vccd1 vccd1 _5179_/A sky130_fd_sc_hd__buf_4
XFILLER_28_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6009_ _6209_/CLK _6009_/D vssd1 vssd1 vccd1 vccd1 _6009_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__3450__D _3450_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4019__B1 _3032_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5216__C1 _4646_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3545__A2 _3567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_608 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output29_A _6300_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4245__S _4246_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5222__A2 _4622_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3710_ _5488_/A _3708_/Y _3709_/X _5743_/C vssd1 vssd1 vccd1 vccd1 _3710_/X sky130_fd_sc_hd__o22a_1
XFILLER_81_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3784__A2 _5943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4690_ _4707_/B _4690_/B vssd1 vssd1 vccd1 vccd1 _4691_/B sky130_fd_sc_hd__nand2_1
XFILLER_119_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3641_ _4216_/A _3210_/B _3640_/X vssd1 vssd1 vccd1 vccd1 _3641_/X sky130_fd_sc_hd__o21a_1
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3572_ _3572_/A _3935_/D _3572_/C vssd1 vssd1 vccd1 vccd1 _3574_/B sky130_fd_sc_hd__and3_1
XFILLER_127_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5311_ _5605_/C _5311_/B vssd1 vssd1 vccd1 vccd1 _5312_/B sky130_fd_sc_hd__or2_4
X_6291_ _6299_/CLK _6291_/D vssd1 vssd1 vccd1 vccd1 _6291_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5289__A2 _5251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5242_ _5242_/A vssd1 vssd1 vccd1 vccd1 _5248_/C sky130_fd_sc_hd__inv_2
XANTENNA__5694__C1 _5710_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3395__S1 _3709_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5173_ _3126_/A _5075_/C _5136_/C vssd1 vssd1 vccd1 vccd1 _5173_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_96_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4124_ _4125_/A _4125_/B vssd1 vssd1 vccd1 vccd1 _4126_/A sky130_fd_sc_hd__nor2_1
XFILLER_96_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput1 io_in[0] vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_2
XFILLER_84_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4055_ _3970_/A _4051_/S _5869_/S _5072_/A vssd1 vssd1 vccd1 vccd1 _6071_/D sky130_fd_sc_hd__a22o_1
XFILLER_110_395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_48_clk _6230_/CLK vssd1 vssd1 vccd1 vccd1 _6257_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_37_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3006_ _4216_/A vssd1 vssd1 vccd1 vccd1 _3944_/A sky130_fd_sc_hd__inv_2
XANTENNA__4663__B _4663_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3472__A1 _3960_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_611 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout252_A _6238_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4957_ _4987_/B _4957_/B vssd1 vssd1 vccd1 vccd1 _4957_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_52_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3908_ _6048_/Q _3727_/X _3909_/S vssd1 vssd1 vccd1 vccd1 _6048_/D sky130_fd_sc_hd__mux2_1
X_4888_ _6191_/Q _4916_/C vssd1 vssd1 vccd1 vccd1 _4896_/B sky130_fd_sc_hd__xnor2_1
XFILLER_20_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3839_ _4846_/B _3740_/X _3749_/X _3838_/X vssd1 vssd1 vccd1 vccd1 _3839_/X sky130_fd_sc_hd__a211o_1
XFILLER_137_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3295__A _6200_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3527__A2 _4767_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5509_ _5476_/B _5509_/B _5509_/C vssd1 vssd1 vccd1 vccd1 _5537_/B sky130_fd_sc_hd__and3b_1
XFILLER_106_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3742__B _5124_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4854__A _6190_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_39_clk clkbuf_3_4__f_clk/X vssd1 vssd1 vccd1 vccd1 _6256_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_74_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4065__S _4066_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3189__B _4462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5204__A2 _5203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_443 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4748__B _5344_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5676__C1 _5956_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5140__A1 _5131_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5691__A2 _3937_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4651__B1 _4640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5860_ _3597_/B _5862_/B _5859_/Y _5867_/A1 vssd1 vssd1 vccd1 vccd1 _5860_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_33_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4811_ _4811_/A _4811_/B vssd1 vssd1 vccd1 vccd1 _4811_/Y sky130_fd_sc_hd__xnor2_1
XTAP_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5791_ _5791_/A _5791_/B vssd1 vssd1 vccd1 vccd1 _5798_/S sky130_fd_sc_hd__nand2_8
XFILLER_33_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5595__A _5595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5600__C1 _5169_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4742_ _6187_/Q _4742_/B vssd1 vssd1 vccd1 vccd1 _4743_/B sky130_fd_sc_hd__nor2_1
XFILLER_14_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4954__B2 _4745_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4673_ _4673_/A _4673_/B vssd1 vssd1 vccd1 vccd1 _4678_/B sky130_fd_sc_hd__nor2_2
XFILLER_119_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3624_ _6207_/Q _3615_/B _5635_/A vssd1 vssd1 vccd1 vccd1 _5898_/A sky130_fd_sc_hd__mux2_2
XFILLER_128_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3555_ _5818_/A _3555_/B _3555_/C vssd1 vssd1 vccd1 vccd1 _3557_/B sky130_fd_sc_hd__and3_4
XFILLER_127_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6274_ _6274_/CLK _6274_/D vssd1 vssd1 vccd1 vccd1 _6274_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3486_ _6278_/Q _6114_/Q _3709_/S vssd1 vssd1 vccd1 vccd1 _5392_/B sky130_fd_sc_hd__mux2_4
XFILLER_89_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4658__B _4658_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5225_ _5454_/B _5264_/B _5226_/A vssd1 vssd1 vccd1 vccd1 _5225_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_88_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5682__A2 _4112_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5156_ _5058_/D _5133_/X _5155_/X vssd1 vssd1 vccd1 vccd1 _5156_/X sky130_fd_sc_hd__o21a_1
XFILLER_69_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4096__D _4309_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4107_ _4162_/A _4176_/B _4107_/C vssd1 vssd1 vccd1 vccd1 _4108_/B sky130_fd_sc_hd__and3_1
XFILLER_84_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5087_ _5227_/A _3672_/Y _4648_/Y vssd1 vssd1 vccd1 vccd1 _5087_/X sky130_fd_sc_hd__a21o_1
XFILLER_84_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5434__A2 _5418_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4038_ _6059_/Q _3711_/X _4044_/S vssd1 vssd1 vccd1 vccd1 _6059_/D sky130_fd_sc_hd__mux2_1
XFILLER_37_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5198__A1 _3116_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5989_ _6103_/Q vssd1 vssd1 vccd1 vccd1 _6103_/D sky130_fd_sc_hd__clkbuf_2
XANTENNA__5709__S _5734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4568__B _5165_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3133__A0 _4819_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5673__A2 _3179_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4881__B1 _3029_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5189__A1 _5191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4936__A1 _4990_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3340_ _4162_/B _3257_/B _5296_/B _3885_/A _3339_/X vssd1 vssd1 vccd1 vccd1 _3340_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_124_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3271_ _4022_/C _5622_/A _3271_/C vssd1 vssd1 vccd1 vccd1 _3274_/A sky130_fd_sc_hd__and3_1
XFILLER_97_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4197__C _4426_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5010_ _5005_/X _5009_/Y _5034_/A vssd1 vssd1 vccd1 vccd1 _5010_/X sky130_fd_sc_hd__mux2_1
XFILLER_85_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5664__A2 _5649_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5912_ _5244_/A _3081_/Y _3886_/X _4586_/Y vssd1 vssd1 vccd1 vccd1 _5920_/C sky130_fd_sc_hd__o22a_1
XFILLER_81_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5843_ _5854_/A _5841_/X _5842_/Y vssd1 vssd1 vccd1 vccd1 _6281_/D sky130_fd_sc_hd__a21oi_1
XFILLER_34_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5774_ _5305_/A _5788_/B _4250_/Y vssd1 vssd1 vccd1 vccd1 _5774_/Y sky130_fd_sc_hd__a21oi_1
X_4725_ _5114_/A _4726_/B vssd1 vssd1 vccd1 vccd1 _4725_/X sky130_fd_sc_hd__or2_2
XFILLER_135_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4656_ _6184_/Q _4970_/B _4653_/X _4655_/Y _5071_/A vssd1 vssd1 vccd1 vccd1 _6184_/D
+ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout215_A _3024_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3607_ _3607_/A _3607_/B vssd1 vssd1 vccd1 vccd1 _3611_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__5352__B2 _5470_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4587_ _5241_/A _4587_/B _5911_/B _5911_/C vssd1 vssd1 vccd1 vccd1 _5870_/B sky130_fd_sc_hd__or4_4
XFILLER_89_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3538_ _3567_/B _3593_/B vssd1 vssd1 vccd1 vccd1 _3594_/A sky130_fd_sc_hd__and2_2
XANTENNA_clkbuf_leaf_51_clk_A _6133_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6257_ _6257_/CLK _6257_/D vssd1 vssd1 vccd1 vccd1 _6257_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3469_ _3365_/B _3518_/B _3468_/X _3312_/B _3145_/C vssd1 vssd1 vccd1 vccd1 _3469_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_67_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5208_ _5790_/A1 _5206_/A _5206_/Y _6162_/Q vssd1 vssd1 vccd1 vccd1 _5208_/X sky130_fd_sc_hd__o22a_1
XFILLER_130_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6188_ _6193_/CLK _6188_/D vssd1 vssd1 vccd1 vccd1 _6188_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_57_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5139_ _5360_/S _3971_/B _5131_/Y _5138_/X vssd1 vssd1 vccd1 vccd1 _5139_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_29_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5407__A2 _5767_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3418__B2 _4003_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5591__A1 _6232_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5591__B2 _3948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5963__A _5970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5139__A2_N _3971_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4579__A _5071_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5894__A2 _5677_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_19_clk_A _6084_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5646__A2 _5128_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5203__A _5203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4606__B1 _5048_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4510_ _3011_/Y _4515_/B _3912_/Y vssd1 vssd1 vccd1 vccd1 _4510_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_117_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5490_ _5310_/Y _5482_/Y _5486_/Y _5489_/X vssd1 vssd1 vccd1 vccd1 _5490_/X sky130_fd_sc_hd__a211o_1
X_4441_ _5292_/B _4438_/S _4439_/S vssd1 vssd1 vccd1 vccd1 _4441_/X sky130_fd_sc_hd__o21a_1
X_4372_ _4340_/A _4340_/B _4345_/A _4345_/B vssd1 vssd1 vccd1 vccd1 _4373_/B sky130_fd_sc_hd__o2bb2a_1
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6111_ _6113_/CLK _6111_/D vssd1 vssd1 vccd1 vccd1 _6111_/Q sky130_fd_sc_hd__dfxtp_1
X_3323_ _3631_/A _3322_/X _3256_/X _3592_/A vssd1 vssd1 vccd1 vccd1 _3323_/X sky130_fd_sc_hd__a211o_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5098__B1 _5097_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6042_ _6218_/CLK _6042_/D vssd1 vssd1 vccd1 vccd1 _6042_/Q sky130_fd_sc_hd__dfxtp_1
X_3254_ _5936_/A _3706_/A _4614_/B vssd1 vssd1 vccd1 vccd1 _5799_/B sky130_fd_sc_hd__or3_4
XFILLER_85_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3185_ _3212_/A _3736_/A vssd1 vssd1 vccd1 vccd1 _3549_/B sky130_fd_sc_hd__or2_4
XFILLER_54_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4952__A _6193_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout165_A _3704_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4073__A1 _4136_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5767__B _5767_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4671__B _5263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3820__A1 _4334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout332_A _5029_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5826_ _5835_/A1 _4384_/Y _5819_/Y _6276_/Q vssd1 vssd1 vccd1 vccd1 _5826_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3259__S0 _4067_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5573__A1 _5412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5757_ _5856_/A _5742_/Y _5755_/X _5756_/Y vssd1 vssd1 vccd1 vccd1 _6246_/D sky130_fd_sc_hd__a22o_1
XFILLER_136_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4708_ _4750_/A _4708_/B vssd1 vssd1 vccd1 vccd1 _4713_/A sky130_fd_sc_hd__nand2_2
XFILLER_5_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5688_ _4162_/A _5649_/X _5687_/X _5956_/A vssd1 vssd1 vccd1 vccd1 _6237_/D sky130_fd_sc_hd__o211a_1
XFILLER_135_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4639_ _5911_/A _4643_/A vssd1 vssd1 vccd1 vccd1 _4644_/A sky130_fd_sc_hd__nand2_8
XFILLER_104_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5628__A2 _4615_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4846__B _4846_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout78_A _3115_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_878 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5677__B _5677_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_466 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4367__A2 _4389_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5564__A1 _5072_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3417__S _3658_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3327__B1 _3589_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5867__A2 _5865_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3952__D_N _4614_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3941__A _3941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4772__A _5119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4055__A1 _3970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4990_ _4990_/A _4990_/B vssd1 vssd1 vccd1 vccd1 _4990_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__3489__S0 _4067_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4055__B2 _5072_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3941_ _3941_/A _3974_/B _3952_/B vssd1 vssd1 vccd1 vccd1 _5634_/B sky130_fd_sc_hd__and3_4
XFILLER_16_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3388__A _3388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3872_ _5943_/B _4608_/C vssd1 vssd1 vccd1 vccd1 _5137_/D sky130_fd_sc_hd__or2_1
X_5611_ _5611_/A _5611_/B vssd1 vssd1 vccd1 vccd1 _5611_/X sky130_fd_sc_hd__and2_1
XANTENNA__5555__A1 _5494_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5542_ _5558_/B _5542_/B vssd1 vssd1 vccd1 vccd1 _5542_/X sky130_fd_sc_hd__or2_4
XFILLER_117_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5307__A1 _3121_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5473_ _5513_/A _5464_/B _5472_/X _5251_/A vssd1 vssd1 vccd1 vccd1 _5473_/Y sky130_fd_sc_hd__o211ai_1
XANTENNA__5307__B2 _4644_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4424_ _4424_/A _4424_/B _4424_/C vssd1 vssd1 vccd1 vccd1 _4429_/A sky130_fd_sc_hd__or3_4
XFILLER_133_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4355_ _4355_/A _4355_/B _4355_/C vssd1 vssd1 vccd1 vccd1 _4356_/B sky130_fd_sc_hd__nor3_1
XFILLER_99_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3306_ _6201_/Q _3575_/B vssd1 vssd1 vccd1 vccd1 _3306_/Y sky130_fd_sc_hd__nor2_1
XFILLER_99_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4286_ _4214_/X _4218_/A _4326_/A _4285_/Y vssd1 vssd1 vccd1 vccd1 _4326_/B sky130_fd_sc_hd__o211ai_4
XFILLER_58_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5086__A3 _3971_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6025_ _6248_/CLK _6025_/D vssd1 vssd1 vccd1 vccd1 _6025_/Q sky130_fd_sc_hd__dfxtp_1
X_3237_ _5436_/A _5436_/C vssd1 vssd1 vccd1 vccd1 _3913_/A sky130_fd_sc_hd__nand2_8
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3168_ _4648_/A _4946_/A vssd1 vssd1 vccd1 vccd1 _3168_/Y sky130_fd_sc_hd__nand2_1
XFILLER_104_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3099_ _3170_/A _6215_/Q _6214_/Q _5051_/C vssd1 vssd1 vccd1 vccd1 _3116_/B sky130_fd_sc_hd__or4_4
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5794__A1 _3718_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3298__A _3541_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout45 _5556_/A2 vssd1 vssd1 vccd1 vccd1 _5251_/A sky130_fd_sc_hd__buf_6
Xfanout56 _3684_/X vssd1 vssd1 vccd1 vccd1 _5742_/C sky130_fd_sc_hd__clkbuf_16
Xfanout67 _5513_/A vssd1 vssd1 vccd1 vccd1 _5595_/A sky130_fd_sc_hd__buf_4
XFILLER_23_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout78 _3115_/Y vssd1 vssd1 vccd1 vccd1 _5034_/A sky130_fd_sc_hd__clkbuf_8
X_5809_ _5835_/A1 _4103_/X _5808_/X vssd1 vssd1 vccd1 vccd1 _6268_/D sky130_fd_sc_hd__a21o_1
XFILLER_22_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout89 _3205_/A vssd1 vssd1 vccd1 vccd1 _5570_/A sky130_fd_sc_hd__buf_8
XFILLER_129_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4857__A _4872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3700__S _3705_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3796__B1 _3382_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4993__C1 _5605_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4767__A _4767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3671__A _4648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4140_ _4171_/A _4140_/B vssd1 vssd1 vccd1 vccd1 _4148_/A sky130_fd_sc_hd__or2_4
XFILLER_96_723 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5068__A3 _5128_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4071_ _4071_/A _4296_/A vssd1 vssd1 vccd1 vccd1 _4072_/C sky130_fd_sc_hd__nor2_8
XFILLER_95_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3022_ _3873_/A vssd1 vssd1 vccd1 vccd1 _3878_/A sky130_fd_sc_hd__inv_2
XANTENNA__5598__A _6233_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_867 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4028__A1 _3940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5225__B1 _5226_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4973_ _5731_/S _4945_/A _4945_/B _4972_/Y vssd1 vssd1 vccd1 vccd1 _4973_/Y sky130_fd_sc_hd__o31ai_4
XANTENNA__5240__A3 _5090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3924_ _3309_/X _3935_/B _3373_/B _3358_/A vssd1 vssd1 vccd1 vccd1 _3924_/X sky130_fd_sc_hd__o22a_1
XFILLER_20_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5528__A1 _4643_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3855_ _3853_/X _3854_/X _3855_/S vssd1 vssd1 vccd1 vccd1 _6041_/D sky130_fd_sc_hd__mux2_1
X_3786_ _4620_/B _3845_/B vssd1 vssd1 vccd1 vccd1 _3786_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__3565__B _3567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5525_ _5498_/A _5521_/X _5522_/Y _4645_/B _5524_/Y vssd1 vssd1 vccd1 vccd1 _5525_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_118_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5456_ _6010_/Q _5454_/A _5456_/S vssd1 vssd1 vccd1 vccd1 _5456_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4407_ _3819_/B _4295_/A _4406_/Y vssd1 vssd1 vccd1 vccd1 _6113_/D sky130_fd_sc_hd__o21ai_1
XFILLER_121_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5700__A1 _3043_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5387_ _5387_/A _5387_/B _5387_/C vssd1 vssd1 vccd1 vccd1 _5420_/B sky130_fd_sc_hd__and3_2
XFILLER_114_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout202 _3147_/Y vssd1 vssd1 vccd1 vccd1 _3869_/B sky130_fd_sc_hd__buf_6
Xfanout213 _3025_/Y vssd1 vssd1 vccd1 vccd1 _5065_/A sky130_fd_sc_hd__buf_8
Xfanout224 _6295_/Q vssd1 vssd1 vccd1 vccd1 _3241_/A sky130_fd_sc_hd__buf_12
X_4338_ _4338_/A _4338_/B vssd1 vssd1 vccd1 vccd1 _4340_/A sky130_fd_sc_hd__nor2_1
Xfanout235 _4577_/A vssd1 vssd1 vccd1 vccd1 _5136_/C sky130_fd_sc_hd__buf_6
XFILLER_87_745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout246 _6240_/Q vssd1 vssd1 vccd1 vccd1 _5862_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_86_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input2_A io_in[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout257 _3943_/A vssd1 vssd1 vccd1 vccd1 _5926_/A0 sky130_fd_sc_hd__buf_6
XFILLER_86_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout268 _6234_/Q vssd1 vssd1 vccd1 vccd1 _4085_/A sky130_fd_sc_hd__buf_4
XFILLER_115_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4269_ _4270_/A _4426_/B vssd1 vssd1 vccd1 vccd1 _4302_/A sky130_fd_sc_hd__nand2_2
Xfanout279 _6224_/Q vssd1 vssd1 vccd1 vccd1 _5385_/A sky130_fd_sc_hd__buf_6
XFILLER_86_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6008_ _6209_/CLK _6008_/D vssd1 vssd1 vccd1 vccd1 _6008_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_28_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_804 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4019__A1 _5940_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4019__B2 _6293_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4587__A _5241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3702__A0 _5790_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4258__A1 _3727_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5455__A0 _5480_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3481__A2 _3589_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4966__C1 _4638_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_550 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3640_ _3164_/Y _3594_/B _3639_/X _3560_/S vssd1 vssd1 vccd1 vccd1 _3640_/X sky130_fd_sc_hd__a211o_1
X_3571_ _3571_/A _3571_/B vssd1 vssd1 vccd1 vccd1 _3572_/C sky130_fd_sc_hd__or2_1
XANTENNA__5930__A1 _3948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5310_ _5605_/C _5311_/B vssd1 vssd1 vccd1 vccd1 _5310_/Y sky130_fd_sc_hd__nor2_4
XFILLER_115_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6290_ _6290_/CLK _6290_/D vssd1 vssd1 vccd1 vccd1 _6290_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5241_ _5241_/A _5241_/B _5241_/C vssd1 vssd1 vccd1 vccd1 _5242_/A sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_3_0__f_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4497__A1 _4872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5172_ _5172_/A _5172_/B vssd1 vssd1 vccd1 vccd1 _5172_/Y sky130_fd_sc_hd__nor2_1
X_4123_ _4123_/A _4125_/B vssd1 vssd1 vccd1 vccd1 _4123_/Y sky130_fd_sc_hd__nor2_1
XFILLER_111_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput2 io_in[1] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__buf_6
X_4054_ _6070_/Q _4051_/S _5869_/S _4846_/A vssd1 vssd1 vccd1 vccd1 _6070_/D sky130_fd_sc_hd__a22o_1
XFILLER_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3005_ _5924_/A vssd1 vssd1 vccd1 vccd1 _5742_/A sky130_fd_sc_hd__clkinv_4
XFILLER_37_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4956_ _4964_/A _4983_/A vssd1 vssd1 vccd1 vccd1 _4957_/B sky130_fd_sc_hd__nand2_1
XFILLER_51_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout245_A _5862_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4421__B2 _4437_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3907_ _6047_/Q _3724_/X _3909_/S vssd1 vssd1 vccd1 vccd1 _6047_/D sky130_fd_sc_hd__mux2_1
X_4887_ _3740_/A _4885_/Y _4886_/Y _4972_/A _4881_/X vssd1 vssd1 vccd1 vccd1 _4887_/X
+ sky130_fd_sc_hd__a32o_2
XFILLER_137_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3838_ _4214_/A _3777_/S _3837_/X _3751_/A vssd1 vssd1 vccd1 vccd1 _3838_/X sky130_fd_sc_hd__o211a_1
XFILLER_20_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3295__B _3297_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3769_ _5210_/B _4539_/A _3772_/B _3769_/D vssd1 vssd1 vccd1 vccd1 _3769_/X sky130_fd_sc_hd__and4_1
XFILLER_118_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5508_ _6003_/Q _5476_/Y _6004_/Q vssd1 vssd1 vccd1 vccd1 _5510_/A sky130_fd_sc_hd__a21oi_1
XFILLER_105_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5134__C1 _5638_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5439_ _6256_/Q _5439_/A2 _5743_/B _6248_/Q vssd1 vssd1 vccd1 vccd1 _5439_/X sky130_fd_sc_hd__o22a_1
XANTENNA__4488__A1 _3011_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5685__B1 _3974_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3742__C _5712_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5437__B1 _4058_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5966__A _5970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4715__A2 _5041_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5912__A1 _5244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5912__B2 _4586_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4479__A1 _5221_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5676__B1 _5675_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5140__A2 _4594_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5979__B2 _5862_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_612 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4780__A _5358_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4810_ _4774_/A _4774_/B _4771_/Y vssd1 vssd1 vccd1 vccd1 _4811_/B sky130_fd_sc_hd__o21ai_2
XTAP_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4939__C1 _5494_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5790_ _5790_/A1 _4250_/Y _5788_/X _5789_/X vssd1 vssd1 vccd1 vccd1 _6257_/D sky130_fd_sc_hd__a22o_1
XANTENNA__5600__B1 _3121_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4741_ _6187_/Q _4742_/B vssd1 vssd1 vccd1 vccd1 _4814_/C sky130_fd_sc_hd__and2_1
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3396__A _5818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4672_ _4672_/A _5263_/A vssd1 vssd1 vccd1 vccd1 _4673_/B sky130_fd_sc_hd__nor2_1
XFILLER_119_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3623_ _3923_/A _3623_/B vssd1 vssd1 vccd1 vccd1 _3623_/Y sky130_fd_sc_hd__xnor2_1
X_3554_ _6271_/Q _6017_/Q _6085_/Q _6040_/Q _4067_/A _3713_/S vssd1 vssd1 vccd1 vccd1
+ _3555_/C sky130_fd_sc_hd__mux4_1
XFILLER_127_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3485_ _4334_/A _3832_/A2 _3251_/B _3484_/X _3255_/Y vssd1 vssd1 vccd1 vccd1 _3485_/X
+ sky130_fd_sc_hd__o221a_1
X_6273_ _6280_/CLK _6273_/D vssd1 vssd1 vccd1 vccd1 _6273_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5224_ _4643_/A _5217_/Y _5223_/X _3060_/B vssd1 vssd1 vccd1 vccd1 _5224_/X sky130_fd_sc_hd__a211o_1
XANTENNA__4020__A _5976_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4955__A _5504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5155_ _4614_/A _5138_/X _5153_/Y _4593_/Y _5154_/Y vssd1 vssd1 vccd1 vccd1 _5155_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_69_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4106_ _4162_/A _4176_/B _4107_/C vssd1 vssd1 vccd1 vccd1 _4108_/A sky130_fd_sc_hd__a21oi_1
X_5086_ _6198_/Q _5870_/A _3971_/B _5158_/A _5136_/C vssd1 vssd1 vccd1 vccd1 _5086_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_110_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4037_ _4475_/S _4520_/S vssd1 vssd1 vccd1 vccd1 _4044_/S sky130_fd_sc_hd__nand2_8
XFILLER_84_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3445__A2 _5707_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4690__A _4707_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5988_ _6102_/Q vssd1 vssd1 vccd1 vccd1 _6102_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_40_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4939_ _3009_/Y _4644_/Y _4826_/Y _4938_/Y _5494_/A vssd1 vssd1 vccd1 vccd1 _4939_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_21_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4158__B1 _4072_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3753__B _3777_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5658__B1 _3950_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4568__C _5241_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3133__A1 _6008_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4881__B2 _4806_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_751 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3944__A _3944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3372__A1 _3658_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3270_ _6266_/Q _6012_/Q _6080_/Q _6035_/Q _4067_/A _3713_/S vssd1 vssd1 vccd1 vccd1
+ _3271_/C sky130_fd_sc_hd__mux4_2
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4197__D _4410_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_862 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_748 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3427__A2 _5439_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5911_ _5911_/A _5911_/B _5911_/C _5911_/D vssd1 vssd1 vccd1 vccd1 _5921_/B sky130_fd_sc_hd__or4_1
XFILLER_19_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5842_ _6281_/Q _5854_/A _5866_/B1 vssd1 vssd1 vccd1 vccd1 _5842_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_34_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5773_ _6252_/Q _5788_/B vssd1 vssd1 vccd1 vccd1 _5773_/X sky130_fd_sc_hd__or2_1
XFILLER_21_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4724_ _5114_/A _4726_/B vssd1 vssd1 vccd1 vccd1 _4727_/A sky130_fd_sc_hd__nor2_1
XANTENNA__5337__C1 _5244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4655_ _5221_/A _4872_/B _4970_/B vssd1 vssd1 vccd1 vccd1 _4655_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_135_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout110_A _3443_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3606_ _3642_/B _3606_/B vssd1 vssd1 vccd1 vccd1 _3606_/Y sky130_fd_sc_hd__nor2_2
XANTENNA__4669__B _6184_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4586_ _4643_/A _4586_/B vssd1 vssd1 vccd1 vccd1 _4586_/Y sky130_fd_sc_hd__nand2_4
X_3537_ _4362_/A _3832_/A2 _3251_/B _3536_/X _3255_/Y vssd1 vssd1 vccd1 vccd1 _3537_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_89_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6256_ _6256_/CLK _6256_/D vssd1 vssd1 vccd1 vccd1 _6256_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3468_ _6204_/Q _3458_/B _3658_/S vssd1 vssd1 vccd1 vccd1 _3468_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5207_ _6218_/Q _5934_/B _5207_/S vssd1 vssd1 vccd1 vccd1 _5207_/X sky130_fd_sc_hd__mux2_1
XFILLER_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6187_ _6193_/CLK _6187_/D vssd1 vssd1 vccd1 vccd1 _6187_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_130_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4863__A1 _5034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3666__A2 _5900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3399_ _3388_/A _3388_/B _3500_/A vssd1 vssd1 vccd1 vccd1 _3405_/C sky130_fd_sc_hd__o21a_1
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5138_ _5138_/A _5138_/B vssd1 vssd1 vccd1 vccd1 _5138_/X sky130_fd_sc_hd__or2_2
XFILLER_85_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5069_ _5069_/A _5069_/B _5069_/C _5069_/D vssd1 vssd1 vccd1 vccd1 _5069_/X sky130_fd_sc_hd__and4_1
XFILLER_84_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5576__C1 _5948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5591__A2 _5454_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5455__S _5539_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5646__A3 _4614_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4606__A1 _5976_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3004__A _3241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4440_ _6118_/Q _4458_/B vssd1 vssd1 vccd1 vccd1 _4440_/X sky130_fd_sc_hd__or2_1
XFILLER_7_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3345__A1 _4096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4371_ _4371_/A _4371_/B vssd1 vssd1 vccd1 vccd1 _4373_/A sky130_fd_sc_hd__xnor2_2
XFILLER_125_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6110_ _6274_/CLK _6110_/D vssd1 vssd1 vccd1 vccd1 _6110_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3322_ _3300_/X _5889_/B _3583_/S vssd1 vssd1 vccd1 vccd1 _3322_/X sky130_fd_sc_hd__mux2_4
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5098__A1 _6008_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6041_ _6041_/CLK _6041_/D vssd1 vssd1 vccd1 vccd1 _6041_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3253_ _5936_/A _3706_/A _4614_/B vssd1 vssd1 vccd1 vccd1 _3253_/Y sky130_fd_sc_hd__nor3_2
XFILLER_100_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3184_ _3212_/A _3736_/A vssd1 vssd1 vccd1 vccd1 _3495_/A sky130_fd_sc_hd__nor2_1
XFILLER_66_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4073__A2 _3709_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3849__A _3944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5270__B2 _3121_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5767__C _5767_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout158_A _3060_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5825_ _3425_/B _5819_/B _5824_/X vssd1 vssd1 vccd1 vccd1 _6275_/D sky130_fd_sc_hd__a21o_1
XFILLER_50_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5022__A1 _6195_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3259__S1 _3709_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5756_ _3010_/Y _5763_/B _5742_/Y vssd1 vssd1 vccd1 vccd1 _5756_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_22_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout325_A input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4707_ _6221_/Q _4707_/B vssd1 vssd1 vccd1 vccd1 _4708_/B sky130_fd_sc_hd__or2_1
X_5687_ _5728_/A _5687_/B _5687_/C vssd1 vssd1 vccd1 vccd1 _5687_/X sky130_fd_sc_hd__or3_2
XFILLER_136_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4638_ _4638_/A _4638_/B vssd1 vssd1 vccd1 vccd1 _4638_/Y sky130_fd_sc_hd__nor2_4
XFILLER_123_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4569_ _5928_/B _5147_/C _5876_/A vssd1 vssd1 vccd1 vccd1 _4569_/X sky130_fd_sc_hd__or3b_1
XFILLER_89_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5089__A1 _4644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6239_ _6270_/CLK _6239_/D vssd1 vssd1 vccd1 vccd1 _6239_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3639__A2 _3987_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5304__A _5305_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3052__A_N _4622_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5013__A1 _5547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3494__A _5707_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3941__B _3974_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4827__A1 _5385_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4827__B2 _4826_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4772__B _4772_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3489__S1 _3709_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3940_ _3940_/A _3940_/B vssd1 vssd1 vccd1 vccd1 _3940_/Y sky130_fd_sc_hd__nor2_1
XFILLER_72_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3388__B _3388_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_50_clk_A _6230_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3871_ _3893_/B _3893_/C vssd1 vssd1 vccd1 vccd1 _3877_/B sky130_fd_sc_hd__or2_2
X_5610_ _3590_/X _5442_/A _5598_/Y _5943_/C _5513_/A vssd1 vssd1 vccd1 vccd1 _5611_/B
+ sky130_fd_sc_hd__o221a_1
XANTENNA__5555__A2 _5542_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5541_ _5540_/B _5540_/C _5547_/A vssd1 vssd1 vccd1 vccd1 _5542_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__5960__C1 _5960_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5472_ _5465_/X _5471_/X _5058_/C vssd1 vssd1 vccd1 vccd1 _5472_/X sky130_fd_sc_hd__a21o_1
X_4423_ _3842_/B _4295_/A _4296_/Y _6115_/Q vssd1 vssd1 vccd1 vccd1 _4423_/X sky130_fd_sc_hd__a2bb2o_1
XANTENNA__5108__B _5108_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4354_ _4355_/A _4355_/B _4355_/C vssd1 vssd1 vccd1 vccd1 _4382_/B sky130_fd_sc_hd__o21a_2
XFILLER_99_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3305_ _3575_/B _3266_/A _3266_/B _3304_/X vssd1 vssd1 vccd1 vccd1 _3310_/A sky130_fd_sc_hd__o31a_4
X_4285_ _4321_/B _4283_/Y _4221_/A _4221_/Y vssd1 vssd1 vccd1 vccd1 _4285_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_98_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6024_ _6293_/CLK _6024_/D vssd1 vssd1 vccd1 vccd1 _6024_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3236_ _5924_/A _3236_/B vssd1 vssd1 vccd1 vccd1 _3236_/Y sky130_fd_sc_hd__nor2_8
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4963__A _4963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3167_ _6009_/Q _6008_/Q vssd1 vssd1 vccd1 vccd1 _5840_/B sky130_fd_sc_hd__nor2_8
XFILLER_94_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout275_A _5480_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3098_ _5731_/S _5049_/A vssd1 vssd1 vccd1 vccd1 _3101_/A sky130_fd_sc_hd__nand2_4
XFILLER_82_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_18_clk_A _6084_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout46 _5250_/X vssd1 vssd1 vccd1 vccd1 _5556_/A2 sky130_fd_sc_hd__buf_6
XFILLER_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout57 _3203_/X vssd1 vssd1 vccd1 vccd1 _3498_/S sky130_fd_sc_hd__buf_4
XFILLER_22_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5808_ _3477_/Y _5801_/B _5801_/Y _6268_/Q vssd1 vssd1 vccd1 vccd1 _5808_/X sky130_fd_sc_hd__a22o_1
Xfanout68 _5494_/A vssd1 vssd1 vccd1 vccd1 _5513_/A sky130_fd_sc_hd__buf_4
Xfanout79 _3115_/Y vssd1 vssd1 vccd1 vccd1 _5050_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_13_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5739_ _3986_/B _3958_/Y _5738_/Y _3180_/Y _5728_/A vssd1 vssd1 vccd1 vccd1 _5740_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_135_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout90_A _3205_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4857__B _4979_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5034__A _5034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3480__C _5436_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4592__B _4592_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3796__A1 _4270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4993__B1 _5172_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4812__S _4812_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3952__A _4587_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4767__B _4767_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3720__A1 _4112_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3671__B _5509_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3720__B2 _6230_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4070_ _5960_/C1 _4614_/B _3766_/Y _4539_/A vssd1 vssd1 vccd1 vccd1 _4296_/A sky130_fd_sc_hd__o31ai_4
XANTENNA__5473__A1 _5513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3021_ _6057_/Q vssd1 vssd1 vccd1 vccd1 _3021_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5225__A1 _5454_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4028__A2 _5900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4972_ _4972_/A _4972_/B _4972_/C vssd1 vssd1 vccd1 vccd1 _4972_/Y sky130_fd_sc_hd__nand3_2
XFILLER_63_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3787__A1 _4697_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3923_ _3923_/A _3923_/B vssd1 vssd1 vccd1 vccd1 _3923_/Y sky130_fd_sc_hd__nand2_1
X_3854_ _5128_/A0 _3765_/X _3772_/X _3771_/B _6041_/Q vssd1 vssd1 vccd1 vccd1 _3854_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_20_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3785_ _6035_/Q _3771_/X _3783_/Y _3784_/X vssd1 vssd1 vccd1 vccd1 _6035_/D sky130_fd_sc_hd__a211o_1
XANTENNA__5119__A _5119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5524_ _3121_/B _5523_/X _3060_/B vssd1 vssd1 vccd1 vccd1 _5524_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_117_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5455_ _5480_/B _4900_/Y _5539_/S vssd1 vssd1 vccd1 vccd1 _5463_/B sky130_fd_sc_hd__mux2_2
XANTENNA__3862__A _3885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4406_ _6113_/Q _4296_/Y _4405_/Y _4437_/A1 vssd1 vssd1 vccd1 vccd1 _4406_/Y sky130_fd_sc_hd__a22oi_1
X_5386_ _5387_/B _5385_/C _5387_/A vssd1 vssd1 vccd1 vccd1 _5386_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__5700__A2 _3495_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout203 _5622_/A vssd1 vssd1 vccd1 vccd1 _3555_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_120_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3711__A1 _6011_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout214 _3025_/Y vssd1 vssd1 vccd1 vccd1 _3941_/A sky130_fd_sc_hd__buf_6
X_4337_ _4362_/A _4167_/C _4336_/C vssd1 vssd1 vccd1 vccd1 _4338_/B sky130_fd_sc_hd__a21oi_1
XFILLER_87_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout225 _5940_/A0 vssd1 vssd1 vccd1 vccd1 _3241_/B sky130_fd_sc_hd__buf_8
XFILLER_86_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout236 _5911_/A vssd1 vssd1 vccd1 vccd1 _4577_/A sky130_fd_sc_hd__buf_6
XFILLER_59_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout247 _5859_/A vssd1 vssd1 vccd1 vccd1 _3942_/B sky130_fd_sc_hd__buf_8
XFILLER_113_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout258 _4270_/A vssd1 vssd1 vccd1 vccd1 _4162_/B sky130_fd_sc_hd__buf_8
XFILLER_87_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout269 _6231_/Q vssd1 vssd1 vccd1 vccd1 _5567_/A sky130_fd_sc_hd__buf_8
X_4268_ _4268_/A _4268_/B vssd1 vssd1 vccd1 vccd1 _4278_/A sky130_fd_sc_hd__xnor2_4
XFILLER_115_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6007_ _6007_/CLK _6007_/D vssd1 vssd1 vccd1 vccd1 _6007_/Q sky130_fd_sc_hd__dfxtp_4
X_3219_ _3869_/A _5818_/B vssd1 vssd1 vccd1 vccd1 _3231_/C sky130_fd_sc_hd__or2_4
XANTENNA__3475__A0 _4734_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4199_ _4195_/Y _4199_/B _4275_/A vssd1 vssd1 vccd1 vccd1 _4275_/B sky130_fd_sc_hd__nand3b_4
XFILLER_55_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5216__A1 _5218_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3102__A _5090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3778__A1 _4658_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5029__A _5567_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5152__B1 _5136_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4587__B _4587_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5455__A1 _4900_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5207__A1 _5934_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3012__A _6221_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4966__B1 _4640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4194__A1 _4214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3570_ _3935_/D _3570_/B vssd1 vssd1 vccd1 vccd1 _3570_/X sky130_fd_sc_hd__xor2_1
XFILLER_6_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3682__A _5635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5240_ _3170_/A _6216_/Q _5090_/A _4596_/B _4605_/A vssd1 vssd1 vccd1 vccd1 _5249_/B
+ sky130_fd_sc_hd__o311a_1
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5694__A1 _3765_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5171_ _5172_/A _3072_/A _3084_/B _5498_/A _5164_/Y vssd1 vssd1 vccd1 vccd1 _5171_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_111_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4122_ _4122_/A _4122_/B vssd1 vssd1 vccd1 vccd1 _4125_/B sky130_fd_sc_hd__or2_1
XFILLER_84_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4053_ _3312_/A _4819_/B _5869_/S vssd1 vssd1 vccd1 vccd1 _6069_/D sky130_fd_sc_hd__mux2_1
Xinput3 io_in[2] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__buf_8
X_3004_ _3241_/A vssd1 vssd1 vccd1 vccd1 _3240_/A sky130_fd_sc_hd__inv_2
XFILLER_37_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4955_ _5504_/A _4979_/B vssd1 vssd1 vccd1 vccd1 _4987_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__3857__A _3880_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3906_ _6046_/Q _3721_/X _3909_/S vssd1 vssd1 vccd1 vccd1 _6046_/D sky130_fd_sc_hd__mux2_1
X_4886_ _5454_/A _4886_/B vssd1 vssd1 vccd1 vccd1 _4886_/Y sky130_fd_sc_hd__nand2_1
XFILLER_138_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3837_ _3593_/A _3746_/A _3836_/X _3849_/B vssd1 vssd1 vccd1 vccd1 _3837_/X sky130_fd_sc_hd__a211o_1
XFILLER_137_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3768_ _3768_/A vssd1 vssd1 vccd1 vccd1 _3771_/B sky130_fd_sc_hd__inv_2
X_5507_ _5507_/A _5507_/B vssd1 vssd1 vccd1 vccd1 _5507_/X sky130_fd_sc_hd__or2_1
X_3699_ _5446_/B _6025_/Q _3902_/A vssd1 vssd1 vccd1 vccd1 _3699_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5134__B1 _5133_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5438_ _6131_/Q _5767_/B _5436_/X _3236_/Y _5437_/X vssd1 vssd1 vccd1 vccd1 _5438_/X
+ sky130_fd_sc_hd__o221a_2
XANTENNA__5685__A1 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3696__A0 _5856_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5369_ _5340_/X _5343_/Y _5366_/Y _5367_/X vssd1 vssd1 vccd1 vccd1 _5370_/A sky130_fd_sc_hd__o211a_1
XFILLER_59_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4948__B1 _6004_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5676__A1 _4270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5206__B _5206_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3007__A _4197_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3439__B1 _5367_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4939__B1 _4826_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4780__B _5367_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5600__A1 _6009_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4740_ _5703_/A _4731_/X _4739_/X _4972_/A vssd1 vssd1 vccd1 vccd1 _4740_/X sky130_fd_sc_hd__a2bb2o_4
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3396__B _3555_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4671_ _4672_/A _5263_/A vssd1 vssd1 vccd1 vccd1 _4710_/A sky130_fd_sc_hd__nand2_1
XFILLER_119_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3622_ _3568_/B _3570_/B _3618_/A vssd1 vssd1 vccd1 vccd1 _3623_/B sky130_fd_sc_hd__o21ai_2
XFILLER_134_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3553_ _6017_/Q _6040_/Q _3709_/S vssd1 vssd1 vccd1 vccd1 _3553_/X sky130_fd_sc_hd__mux2_2
XFILLER_115_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4301__A _4301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6272_ _6272_/CLK _6272_/D vssd1 vssd1 vccd1 vccd1 _6272_/Q sky130_fd_sc_hd__dfxtp_1
X_3484_ _3590_/A1 _3483_/X _3482_/X vssd1 vssd1 vccd1 vccd1 _3484_/X sky130_fd_sc_hd__a21o_2
XFILLER_115_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5667__A1 _5730_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5223_ _3156_/Y _5220_/X _5222_/X _4638_/B vssd1 vssd1 vccd1 vccd1 _5223_/X sky130_fd_sc_hd__o211a_1
XFILLER_97_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5154_ _3863_/X _5909_/B _5065_/A _5095_/A vssd1 vssd1 vccd1 vccd1 _5154_/Y sky130_fd_sc_hd__a211oi_1
XFILLER_69_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4955__B _4979_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4105_ _4437_/A1 _4103_/X _4104_/X vssd1 vssd1 vccd1 vccd1 _6082_/D sky130_fd_sc_hd__a21o_1
XFILLER_110_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5085_ _5093_/A _5093_/B vssd1 vssd1 vccd1 vccd1 _5085_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_fanout188_A _3280_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4036_ _5767_/C _5925_/A vssd1 vssd1 vccd1 vccd1 _4520_/S sky130_fd_sc_hd__or2_4
XFILLER_56_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3850__B1 _3740_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4690__B _4690_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5987_ _6101_/Q vssd1 vssd1 vccd1 vccd1 _6101_/D sky130_fd_sc_hd__clkbuf_2
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5198__A3 _5617_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4938_ _5543_/S _4918_/Y _4937_/X vssd1 vssd1 vccd1 vccd1 _4938_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_21_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4869_ _4864_/Y _4865_/X _4868_/X _3122_/Y vssd1 vssd1 vccd1 vccd1 _4869_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3905__A1 _3718_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5658__A1 _5710_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5830__A1 _5835_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3841__A0 _5898_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5346__B1 _5345_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3372__A2 _3388_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_616 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5821__A1 _3322_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5910_ _4826_/Y _5239_/D _5909_/Y _5551_/A _5074_/Y vssd1 vssd1 vccd1 vccd1 _5921_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_81_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3832__B1 _3536_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5841_ _4010_/B _3251_/A _5862_/B vssd1 vssd1 vccd1 vccd1 _5841_/X sky130_fd_sc_hd__mux2_8
X_5772_ _5935_/A0 _4250_/Y _5770_/X _5771_/X vssd1 vssd1 vccd1 vccd1 _6251_/D sky130_fd_sc_hd__a22o_1
XFILLER_21_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3200__A _3765_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4723_ _4625_/A _5093_/A _4722_/X _4721_/X _5866_/B1 vssd1 vssd1 vccd1 vccd1 _6186_/D
+ sky130_fd_sc_hd__o311a_1
X_4654_ _4654_/A _5203_/A vssd1 vssd1 vccd1 vccd1 _4654_/Y sky130_fd_sc_hd__nor2_1
XFILLER_135_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3605_ _4214_/A _3210_/B _3210_/C _3604_/X vssd1 vssd1 vccd1 vccd1 _3605_/X sky130_fd_sc_hd__o211a_1
XFILLER_128_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4585_ _3084_/B _3979_/B _4583_/X _4584_/Y _5192_/A vssd1 vssd1 vccd1 vccd1 _6183_/D
+ sky130_fd_sc_hd__a311o_1
X_3536_ _3532_/X _3533_/X _3535_/X _3590_/A1 vssd1 vssd1 vccd1 vccd1 _3536_/X sky130_fd_sc_hd__a22o_4
XANTENNA__4560__A1 _4872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6255_ _6256_/CLK _6255_/D vssd1 vssd1 vccd1 vccd1 _6255_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3467_ _6204_/Q _3458_/B _3575_/B vssd1 vssd1 vccd1 vccd1 _3518_/B sky130_fd_sc_hd__mux2_4
XANTENNA__5561__S _5561_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4312__A1 _4426_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5206_ _5206_/A _5206_/B vssd1 vssd1 vccd1 vccd1 _5206_/Y sky130_fd_sc_hd__nand2_1
XFILLER_130_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6186_ _6196_/CLK _6186_/D vssd1 vssd1 vccd1 vccd1 _6186_/Q sky130_fd_sc_hd__dfxtp_2
X_3398_ _3398_/A _3500_/C vssd1 vssd1 vccd1 vccd1 _3398_/X sky130_fd_sc_hd__or2_1
XFILLER_97_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4685__A2_N _4872_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5137_ _5258_/A _5928_/B _5911_/C _5137_/D vssd1 vssd1 vccd1 vccd1 _5138_/B sky130_fd_sc_hd__or4_1
XFILLER_84_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5068_ _6197_/Q _5238_/A _5128_/S _5239_/A vssd1 vssd1 vccd1 vccd1 _5069_/D sky130_fd_sc_hd__a31o_1
XFILLER_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5812__A1 _3583_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4019_ _5940_/A0 _5108_/A _3032_/Y _6293_/Q _4018_/X vssd1 vssd1 vccd1 vccd1 _4020_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_84_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4206__A _4362_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3110__A _5075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5591__A3 _4638_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5328__A0 _6222_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5879__A1 _4819_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4000__B1 _5932_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4551__A1 _3011_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3354__A2 _4663_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4876__A _5454_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3955__A _5128_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5319__B1 _5742_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4542__A1 _5221_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4370_ _4370_/A _4370_/B vssd1 vssd1 vccd1 vccd1 _4371_/B sky130_fd_sc_hd__xnor2_4
XFILLER_125_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3321_ _3311_/Y _3320_/X _3511_/A vssd1 vssd1 vccd1 vccd1 _5889_/B sky130_fd_sc_hd__mux2_8
XFILLER_4_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5098__A2 _3111_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6040_ _6079_/CLK _6040_/D vssd1 vssd1 vccd1 vccd1 _6040_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3252_ _3960_/C _3951_/C vssd1 vssd1 vccd1 vccd1 _4614_/B sky130_fd_sc_hd__or2_4
XFILLER_86_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3183_ _5870_/A _4566_/B vssd1 vssd1 vccd1 vccd1 _3736_/A sky130_fd_sc_hd__or2_4
XFILLER_27_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5824_ _5835_/A1 _4359_/Y _5819_/Y _6275_/Q vssd1 vssd1 vccd1 vccd1 _5824_/X sky130_fd_sc_hd__a22o_1
XFILLER_34_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5755_ _6246_/Q _5763_/B vssd1 vssd1 vccd1 vccd1 _5755_/X sky130_fd_sc_hd__or2_1
XANTENNA__3865__A _4604_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4706_ _6221_/Q _4707_/B vssd1 vssd1 vccd1 vccd1 _4750_/A sky130_fd_sc_hd__nand2_2
XANTENNA__3584__A2 _3583_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5686_ _5075_/A _4619_/B _5203_/A _3458_/B _5685_/X vssd1 vssd1 vccd1 vccd1 _5687_/C
+ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout318_A _5799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4637_ _6184_/Q _4634_/X _5041_/S vssd1 vssd1 vccd1 vccd1 _4637_/X sky130_fd_sc_hd__mux2_1
XFILLER_135_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4568_ _5244_/B _5165_/B _5241_/B vssd1 vssd1 vccd1 vccd1 _5147_/C sky130_fd_sc_hd__and3_1
XFILLER_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3519_ _3462_/X _3518_/Y _3935_/C vssd1 vssd1 vccd1 vccd1 _3572_/A sky130_fd_sc_hd__a21o_1
XANTENNA__4696__A _4697_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4499_ _6140_/Q _4499_/B vssd1 vssd1 vccd1 vccd1 _4499_/X sky130_fd_sc_hd__or2_1
XFILLER_89_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6238_ _6270_/CLK _6238_/D vssd1 vssd1 vccd1 vccd1 _6238_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_89_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6169_ _6170_/CLK _6169_/D vssd1 vssd1 vccd1 vccd1 _6169_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3105__A _3105_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5013__A2 _4645_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_20_clk _6084_/CLK vssd1 vssd1 vccd1 vccd1 _6274_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_5_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3327__A2 _3589_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3941__C _3952_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4827__A2 _4644_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3388__C _3500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3870_ _3893_/B _3893_/C vssd1 vssd1 vccd1 vccd1 _4608_/C sky130_fd_sc_hd__nor2_4
XANTENNA__3685__A _5767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5540_ _6230_/Q _5540_/B _5540_/C vssd1 vssd1 vccd1 vccd1 _5558_/B sky130_fd_sc_hd__and3_1
XANTENNA__4763__A1 _5333_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4763__B2 _4931_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5960__B1 _5131_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_11_clk _6219_/CLK vssd1 vssd1 vccd1 vccd1 _6301_/CLK sky130_fd_sc_hd__clkbuf_16
X_5471_ _5909_/B _5734_/B _5464_/B _5943_/C vssd1 vssd1 vccd1 vccd1 _5471_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_118_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4422_ _3831_/B _4295_/A _4421_/Y vssd1 vssd1 vccd1 vccd1 _6114_/D sky130_fd_sc_hd__o21ai_1
XANTENNA__5712__A0 _3615_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4353_ _4353_/A _4353_/B vssd1 vssd1 vccd1 vccd1 _4355_/C sky130_fd_sc_hd__xnor2_1
XFILLER_98_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3624__S _5635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5405__A _5436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3304_ _6201_/Q _3869_/B vssd1 vssd1 vccd1 vccd1 _3304_/X sky130_fd_sc_hd__or2_1
XFILLER_101_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4284_ _4221_/A _4221_/Y _4321_/B _4283_/Y vssd1 vssd1 vccd1 vccd1 _4326_/A sky130_fd_sc_hd__a211o_2
XFILLER_113_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6023_ _6254_/CLK _6023_/D vssd1 vssd1 vccd1 vccd1 _6023_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3235_ _3241_/A _3241_/B vssd1 vssd1 vccd1 vccd1 _3235_/X sky130_fd_sc_hd__or2_2
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3166_ _5840_/A _4462_/A vssd1 vssd1 vccd1 vccd1 _3741_/B sky130_fd_sc_hd__or2_4
XFILLER_104_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout170_A _3239_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3097_ _4946_/A _4999_/B vssd1 vssd1 vccd1 vccd1 _4972_/A sky130_fd_sc_hd__nor2_8
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout47 _4553_/B vssd1 vssd1 vccd1 vccd1 _4562_/B sky130_fd_sc_hd__clkbuf_4
Xfanout58 _3495_/A vssd1 vssd1 vccd1 vccd1 _3636_/A sky130_fd_sc_hd__clkbuf_4
X_5807_ _5835_/A1 _4090_/X _5806_/X vssd1 vssd1 vccd1 vccd1 _6267_/D sky130_fd_sc_hd__a21o_1
XANTENNA__4203__B1 _4342_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout69 _4600_/Y vssd1 vssd1 vccd1 vccd1 _5494_/A sky130_fd_sc_hd__clkbuf_8
X_3999_ _3995_/Y _3999_/B _3999_/C vssd1 vssd1 vccd1 vccd1 _3999_/X sky130_fd_sc_hd__and3b_1
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5738_ _5738_/A _5738_/B vssd1 vssd1 vccd1 vccd1 _5738_/Y sky130_fd_sc_hd__nand2_1
XFILLER_6_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5669_ _6293_/Q _4615_/A _3772_/B vssd1 vssd1 vccd1 vccd1 _5669_/X sky130_fd_sc_hd__a21o_1
XFILLER_136_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout83_A _5731_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3493__B2 _3599_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5050__A _5072_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4993__A1 _6194_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3709__S _3709_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5942__B1 _5921_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3952__B _3952_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3720__A2 _5743_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5458__C1 _5570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3020_ _6058_/Q vssd1 vssd1 vccd1 vccd1 _3020_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_0_clk _6133_/CLK vssd1 vssd1 vccd1 vccd1 _6288_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__3484__A1 _3590_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5225__A2 _5264_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4971_ _4625_/A _5093_/A _4969_/X _4970_/X _5071_/A vssd1 vssd1 vccd1 vccd1 _6193_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_64_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5630__C1 _3996_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3922_ _3649_/A _3649_/B _3922_/S vssd1 vssd1 vccd1 vccd1 _5900_/B sky130_fd_sc_hd__mux2_1
XFILLER_32_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3853_ _5900_/A _3841_/S _3852_/X vssd1 vssd1 vccd1 vccd1 _3853_/X sky130_fd_sc_hd__o21a_2
XFILLER_20_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4736__A1 _5296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5933__B1 _5921_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3784_ _4096_/A _5943_/A _3331_/Y _3765_/X _3772_/X vssd1 vssd1 vccd1 vccd1 _3784_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_118_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5119__B _5934_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5523_ _4707_/B _6005_/Q _5543_/S vssd1 vssd1 vccd1 vccd1 _5523_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5454_ _5454_/A _5454_/B vssd1 vssd1 vccd1 vccd1 _5454_/Y sky130_fd_sc_hd__nor2_1
XFILLER_117_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4405_ _4405_/A _4405_/B vssd1 vssd1 vccd1 vccd1 _4405_/Y sky130_fd_sc_hd__xnor2_1
X_5385_ _5385_/A _5387_/B _5385_/C vssd1 vssd1 vccd1 vccd1 _5446_/C sky130_fd_sc_hd__and3_2
XFILLER_99_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4336_ _4362_/A _4389_/B _4336_/C vssd1 vssd1 vccd1 vccd1 _4338_/A sky130_fd_sc_hd__and3_1
XFILLER_5_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout204 _3137_/X vssd1 vssd1 vccd1 vccd1 _5622_/A sky130_fd_sc_hd__buf_8
Xfanout215 _3024_/Y vssd1 vssd1 vccd1 vccd1 _4638_/A sky130_fd_sc_hd__buf_12
Xfanout226 _6294_/Q vssd1 vssd1 vccd1 vccd1 _5940_/A0 sky130_fd_sc_hd__buf_4
XFILLER_113_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout237 _5911_/A vssd1 vssd1 vccd1 vccd1 _3948_/A sky130_fd_sc_hd__buf_12
Xfanout248 _4362_/A vssd1 vssd1 vccd1 vccd1 _4202_/A sky130_fd_sc_hd__buf_8
X_4267_ _4410_/B _4311_/B vssd1 vssd1 vccd1 vccd1 _4268_/B sky130_fd_sc_hd__nand2_4
XANTENNA__4974__A _4974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout259 _3943_/A vssd1 vssd1 vccd1 vccd1 _4270_/A sky130_fd_sc_hd__buf_12
XFILLER_87_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6006_ _6007_/CLK _6006_/D vssd1 vssd1 vccd1 vccd1 _6006_/Q sky130_fd_sc_hd__dfxtp_4
X_3218_ _3498_/S _3218_/B _3398_/A _3218_/D vssd1 vssd1 vccd1 vccd1 _5818_/B sky130_fd_sc_hd__and4_4
XFILLER_74_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4198_ _4199_/B _4275_/A _4195_/Y vssd1 vssd1 vccd1 vccd1 _4200_/B sky130_fd_sc_hd__a21bo_2
XFILLER_67_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3149_ _3948_/A _5936_/A _5712_/S vssd1 vssd1 vccd1 vccd1 _3738_/A sky130_fd_sc_hd__or3_4
XFILLER_28_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3102__B _4638_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3778__A2 _3740_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_747 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4214__A _4214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5029__B _5029_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3772__B _3772_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5688__C1 _5956_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5152__A1 _5238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5860__C1 _5867_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5612__C1 _5251_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4966__A1 _4990_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5915__B1 _5172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4194__A2 _4173_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5654__S _5703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3963__A _4604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_784 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5694__A2 _5380_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5170_ _3050_/B _3964_/B _5168_/X _5169_/Y _3880_/B vssd1 vssd1 vccd1 vccd1 _5170_/Y
+ sky130_fd_sc_hd__o2111ai_2
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_17_clk_A _6084_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4121_ _4121_/A _4121_/B vssd1 vssd1 vccd1 vccd1 _4122_/B sky130_fd_sc_hd__nor2_1
XFILLER_96_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4052_ _3880_/A _4051_/S _5869_/S _4697_/A vssd1 vssd1 vccd1 vccd1 _6068_/D sky130_fd_sc_hd__a22o_1
XFILLER_110_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput4 io_in[3] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__buf_6
XFILLER_77_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5851__C1 _5866_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3003_ _6296_/Q vssd1 vssd1 vccd1 vccd1 _5955_/A sky130_fd_sc_hd__inv_2
XFILLER_36_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4954_ _4705_/A _4959_/B _4950_/X _4745_/A vssd1 vssd1 vccd1 vccd1 _4954_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_51_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3857__B _5883_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3905_ _6045_/Q _3718_/X _3909_/S vssd1 vssd1 vccd1 vccd1 _6045_/D sky130_fd_sc_hd__mux2_1
XFILLER_33_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4885_ _4882_/Y _4883_/Y _4884_/Y vssd1 vssd1 vccd1 vccd1 _4885_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_32_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4034__A _5742_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3836_ _3643_/A _3738_/X _3801_/B _3835_/X vssd1 vssd1 vccd1 vccd1 _3836_/X sky130_fd_sc_hd__o211a_1
XANTENNA_fanout133_A _3084_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5382__A1 _5412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3767_ _5210_/B _3772_/B _3769_/D _5932_/A vssd1 vssd1 vccd1 vccd1 _3768_/A sky130_fd_sc_hd__a31o_1
XANTENNA__3873__A _3873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5506_ _5327_/A _5547_/C _5505_/Y _5503_/X vssd1 vssd1 vccd1 vccd1 _5507_/B sky130_fd_sc_hd__o31a_1
XANTENNA_fanout300_A _6069_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4072__D_N _5138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3698_ _3942_/B _3697_/X _3705_/A vssd1 vssd1 vccd1 vccd1 _6024_/D sky130_fd_sc_hd__mux2_1
XFILLER_106_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5437_ _6179_/Q _4234_/B _4058_/B _6139_/Q vssd1 vssd1 vccd1 vccd1 _5437_/X sky130_fd_sc_hd__o22a_1
XANTENNA__5685__A2 _3179_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5368_ _5366_/Y _5367_/X _5340_/X _5343_/Y vssd1 vssd1 vccd1 vccd1 _5368_/X sky130_fd_sc_hd__a211o_1
XFILLER_87_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4319_ _4320_/A _4320_/B vssd1 vssd1 vccd1 vccd1 _4351_/B sky130_fd_sc_hd__and2b_1
X_5299_ _5297_/Y _5298_/X _5653_/A vssd1 vssd1 vccd1 vccd1 _5299_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__5437__A2 _4234_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3113__A _5069_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout46_A _5250_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4948__A1 _4974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5070__A0 _6197_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_499 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5676__A2 _5649_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4884__B1 _4886_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3722__S _3731_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5503__A _5503_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3439__A1 _4163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3439__B2 _3885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3023__A _3869_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3958__A _3958_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output27_A _6183_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5600__A2 _4646_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_820 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4670_ _4672_/A _5263_/A vssd1 vssd1 vccd1 vccd1 _4673_/A sky130_fd_sc_hd__and2_1
X_3621_ _3621_/A _3621_/B _3653_/A vssd1 vssd1 vccd1 vccd1 _3621_/X sky130_fd_sc_hd__or3_1
X_3552_ _4214_/A _3136_/Y _5428_/B _3053_/X vssd1 vssd1 vccd1 vccd1 _3557_/A sky130_fd_sc_hd__a22o_4
XFILLER_115_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6271_ _6274_/CLK _6271_/D vssd1 vssd1 vccd1 vccd1 _6271_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5116__A1 _3033_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3483_ _6262_/Q _6054_/Q _6047_/Q _6031_/Q _3241_/A _5940_/A0 vssd1 vssd1 vccd1 vccd1
+ _3483_/X sky130_fd_sc_hd__mux4_1
XANTENNA__4301__B _4410_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5222_ _5625_/A _4622_/B _5221_/B _5219_/X _5221_/Y vssd1 vssd1 vccd1 vccd1 _5222_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5667__A2 _3937_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5153_ _5131_/B _5152_/Y _5077_/C _3123_/A vssd1 vssd1 vccd1 vccd1 _5153_/Y sky130_fd_sc_hd__a211oi_1
XFILLER_69_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4104_ _3807_/B _4069_/B _4072_/C _6082_/Q vssd1 vssd1 vccd1 vccd1 _4104_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_84_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5084_ _5090_/A _5074_/A _5080_/X _5083_/Y vssd1 vssd1 vccd1 vccd1 _5093_/B sky130_fd_sc_hd__a211o_2
XFILLER_110_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4627__B1 _5703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4035_ _5767_/C _5925_/A vssd1 vssd1 vccd1 vccd1 _4515_/B sky130_fd_sc_hd__nor2_2
XFILLER_72_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3868__A _5712_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout348_A _4633_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5986_ _5984_/Y _5985_/X _5986_/B1 vssd1 vssd1 vccd1 vccd1 _6302_/D sky130_fd_sc_hd__a21oi_1
XFILLER_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4937_ _6192_/Q _3671_/Y _5172_/B _4974_/A vssd1 vssd1 vccd1 vccd1 _4937_/X sky130_fd_sc_hd__o22a_1
XANTENNA__3602__A1 _5428_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4868_ _6190_/Q _4867_/X _4990_/A vssd1 vssd1 vccd1 vccd1 _4868_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5355__A1 _5943_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5355__B2 _5442_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3819_ _3855_/S _3819_/B vssd1 vssd1 vccd1 vccd1 _3819_/Y sky130_fd_sc_hd__nor2_1
XFILLER_119_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4799_ _6188_/Q _4970_/B vssd1 vssd1 vccd1 vccd1 _4799_/X sky130_fd_sc_hd__or2_1
XFILLER_118_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3108__A _3958_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5658__A2 _3713_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5346__A1 _5507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3960__B _3960_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5887__B _5888_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3832__A1 _4202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5840_ _5840_/A _5840_/B vssd1 vssd1 vccd1 vccd1 _5865_/S sky130_fd_sc_hd__nor2_4
XFILLER_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5771_ _5292_/B _5791_/B _5769_/S vssd1 vssd1 vccd1 vccd1 _5771_/X sky130_fd_sc_hd__o21a_1
XANTENNA__3200__B _4604_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4722_ _6221_/Q _4872_/B _4720_/X _4931_/B vssd1 vssd1 vccd1 vccd1 _4722_/X sky130_fd_sc_hd__o22a_1
XANTENNA__5337__A1 _5133_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4653_ _4636_/Y _4652_/X _5069_/A vssd1 vssd1 vccd1 vccd1 _4653_/X sky130_fd_sc_hd__o21a_1
X_3604_ _3225_/X _3593_/A _3603_/X _3560_/S vssd1 vssd1 vccd1 vccd1 _3604_/X sky130_fd_sc_hd__a211o_1
X_4584_ _3979_/B _4583_/X _6183_/Q vssd1 vssd1 vccd1 vccd1 _4584_/Y sky130_fd_sc_hd__a21boi_1
X_3535_ _6055_/Q _3589_/A2 _3589_/B1 _6048_/Q _3534_/X vssd1 vssd1 vccd1 vccd1 _3535_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__4560__A2 _4252_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3466_ _3926_/C _3466_/B vssd1 vssd1 vccd1 vccd1 _3466_/Y sky130_fd_sc_hd__xnor2_1
X_6254_ _6254_/CLK _6254_/D vssd1 vssd1 vccd1 vccd1 _6254_/Q sky130_fd_sc_hd__dfxtp_1
X_5205_ _5097_/A _3170_/A _5203_/X _5204_/Y _5192_/A vssd1 vssd1 vccd1 vccd1 _6217_/D
+ sky130_fd_sc_hd__a221oi_2
XFILLER_103_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4312__A2 _4311_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6185_ _6288_/CLK _6185_/D vssd1 vssd1 vccd1 vccd1 _6185_/Q sky130_fd_sc_hd__dfxtp_4
X_3397_ _4162_/A _3257_/B _5341_/B _3885_/A _3396_/X vssd1 vssd1 vccd1 vccd1 _3397_/X
+ sky130_fd_sc_hd__a221o_2
XANTENNA_fanout298_A _6070_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3520__B1 _3621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5136_ _5134_/X _5136_/B _5136_/C vssd1 vssd1 vccd1 vccd1 _5136_/X sky130_fd_sc_hd__and3b_1
XFILLER_123_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5067_ _6197_/Q _4604_/A _3996_/B _5066_/Y vssd1 vssd1 vccd1 vccd1 _5069_/C sky130_fd_sc_hd__a31o_1
XANTENNA__5273__B1 _5227_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4018_ _6218_/Q _3029_/Y _5714_/A _6042_/Q _4017_/X vssd1 vssd1 vccd1 vccd1 _4018_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_38_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3823__A1 _5392_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5576__A1 _5567_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4206__B _4311_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5969_ _3033_/Y _5158_/A _4023_/A _5115_/Y vssd1 vssd1 vccd1 vccd1 _5970_/B sky130_fd_sc_hd__o31a_1
XANTENNA__3587__B1 _3589_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4876__B _4877_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3272__S _3551_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5053__A _5090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5510__C_N _5227_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3814__A1 _4163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5016__A0 _6195_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3301__A _3312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3971__A _4577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3320_ _3315_/Y _3318_/X _3319_/X _3303_/X _3960_/B vssd1 vssd1 vccd1 vccd1 _3320_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_125_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3251_ _3251_/A _3251_/B vssd1 vssd1 vccd1 vccd1 _3251_/Y sky130_fd_sc_hd__nand2_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3182_ _3880_/B _3996_/B vssd1 vssd1 vccd1 vccd1 _4566_/B sky130_fd_sc_hd__nand2_1
XFILLER_67_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3805__A1 _4734_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5823_ _3375_/X _5819_/B _5822_/X vssd1 vssd1 vccd1 vccd1 _6274_/D sky130_fd_sc_hd__a21o_1
XFILLER_62_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5754_ _3942_/D _5742_/Y _5752_/X _5753_/Y vssd1 vssd1 vccd1 vccd1 _6245_/D sky130_fd_sc_hd__a22o_1
XANTENNA__3865__B _5928_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4705_ _4705_/A _4716_/B vssd1 vssd1 vccd1 vccd1 _4705_/Y sky130_fd_sc_hd__nor2_1
X_5685_ input4/X _3179_/X _3974_/C _5684_/X vssd1 vssd1 vccd1 vccd1 _5685_/X sky130_fd_sc_hd__o211a_1
XANTENNA__5138__A _5138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4636_ _3116_/B _4631_/Y _4635_/X vssd1 vssd1 vccd1 vccd1 _4636_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout213_A _3025_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4567_ _5097_/A _5075_/A vssd1 vssd1 vccd1 vccd1 _5876_/A sky130_fd_sc_hd__nor2_2
XANTENNA__3881__A _3881_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3518_ _3518_/A _3518_/B vssd1 vssd1 vccd1 vccd1 _3518_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__4696__B _4697_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4498_ _3942_/A _4501_/A2 _4496_/X _4497_/X vssd1 vssd1 vccd1 vccd1 _6139_/D sky130_fd_sc_hd__a22o_1
X_6237_ _6241_/CLK _6237_/D vssd1 vssd1 vccd1 vccd1 _6237_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_104_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3449_ _3500_/A _3458_/B vssd1 vssd1 vccd1 vccd1 _3986_/C sky130_fd_sc_hd__or2_1
XANTENNA__4297__A1 _4437_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6168_ _6170_/CLK _6168_/D vssd1 vssd1 vccd1 vccd1 _6168_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3105__B _5075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5119_ _5119_/A _5934_/A vssd1 vssd1 vccd1 vccd1 _5119_/Y sky130_fd_sc_hd__nor2_1
XFILLER_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4049__A1 _3873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6099_ _6260_/CLK _6099_/D vssd1 vssd1 vccd1 vccd1 _6099_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4049__B2 _4633_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5797__A1 _3727_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_775 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3121__A _5218_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5182__C1 _5731_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5237__B1 _5638_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4460__A1 _5790_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3031__A _4657_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3966__A _5934_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3685__B _3704_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4763__A2 _4872_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5960__A1 _3112_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3420__C1 _3960_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5470_ _5467_/X _5469_/X _5470_/S vssd1 vssd1 vccd1 vccd1 _5734_/B sky130_fd_sc_hd__mux2_4
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4421_ _6114_/Q _4296_/Y _4420_/X _4437_/A1 vssd1 vssd1 vccd1 vccd1 _4421_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_126_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4352_ _4353_/B _4353_/A vssd1 vssd1 vccd1 vccd1 _4382_/A sky130_fd_sc_hd__and2b_2
XFILLER_125_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3303_ _6201_/Q _3388_/A vssd1 vssd1 vccd1 vccd1 _3303_/X sky130_fd_sc_hd__and2_1
X_4283_ _4283_/A _4283_/B vssd1 vssd1 vccd1 vccd1 _4283_/Y sky130_fd_sc_hd__nor2_2
XFILLER_59_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3206__A _5054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3234_ _3241_/A _3241_/B vssd1 vssd1 vccd1 vccd1 _3236_/B sky130_fd_sc_hd__nor2_4
X_6022_ _6154_/CLK _6022_/D vssd1 vssd1 vccd1 vccd1 _6022_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3165_ _5840_/A _4462_/A vssd1 vssd1 vccd1 vccd1 _3740_/B sky130_fd_sc_hd__nor2_1
XFILLER_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5228__B1 _5605_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3096_ _3170_/A _4744_/B vssd1 vssd1 vccd1 vccd1 _5049_/A sky130_fd_sc_hd__nand2_2
XFILLER_81_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4451__A1 _5856_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout48 _4490_/B vssd1 vssd1 vccd1 vccd1 _4499_/B sky130_fd_sc_hd__buf_4
X_5806_ _3425_/B _5801_/B _5801_/Y _6267_/Q vssd1 vssd1 vccd1 vccd1 _5806_/X sky130_fd_sc_hd__a22o_1
XANTENNA_fanout330_A _5207_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout59 _3958_/Y vssd1 vssd1 vccd1 vccd1 _5203_/A sky130_fd_sc_hd__buf_6
XFILLER_10_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4203__A1 _4334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4203__B2 _4162_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3998_ _5226_/A _4657_/A _3998_/C _3998_/D vssd1 vssd1 vccd1 vccd1 _3999_/B sky130_fd_sc_hd__or4_1
XFILLER_50_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5737_ _3868_/Y _5736_/X _4002_/X vssd1 vssd1 vccd1 vccd1 _5738_/B sky130_fd_sc_hd__o21ai_1
XFILLER_109_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5668_ _5955_/A _5735_/S vssd1 vssd1 vccd1 vccd1 _5668_/Y sky130_fd_sc_hd__nor2_1
XFILLER_129_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4619_ _4619_/A _4619_/B vssd1 vssd1 vccd1 vccd1 _4620_/D sky130_fd_sc_hd__nor2_1
X_5599_ _6233_/Q _5599_/B vssd1 vssd1 vccd1 vccd1 _5599_/X sky130_fd_sc_hd__and2_1
XANTENNA__3714__B1 _3713_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5467__B1 _3704_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout76_A _3194_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3493__A2 _3450_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_807 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5050__B _5050_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4442__A1 _5935_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5942__A1 _5264_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3725__S _3731_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4410__A _4426_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5170__A2 _3964_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3026__A _3312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3469__C1 _3145_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3460__S _3575_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5241__A _5241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4970_ _6193_/Q _4970_/B vssd1 vssd1 vccd1 vccd1 _4970_/X sky130_fd_sc_hd__or2_1
XFILLER_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4433__A1 _4437_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3921_ _6056_/Q _3730_/X _3921_/S vssd1 vssd1 vccd1 vccd1 _6056_/D sky130_fd_sc_hd__mux2_1
XFILLER_32_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3852_ _4877_/B _3749_/X _3851_/X _3748_/Y vssd1 vssd1 vccd1 vccd1 _3852_/X sky130_fd_sc_hd__a211o_1
XFILLER_32_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5933__A1 _4657_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4736__A2 _4690_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3783_ _3855_/S _3783_/B vssd1 vssd1 vccd1 vccd1 _3783_/Y sky130_fd_sc_hd__nor2_1
X_5522_ _5540_/B _5540_/C vssd1 vssd1 vccd1 vccd1 _5522_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_118_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5453_ _5453_/A _5453_/B vssd1 vssd1 vccd1 vccd1 _5453_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_133_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5697__A0 _3593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5416__A _5446_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4404_ _4382_/A _4382_/B _4383_/S _4384_/A _4405_/A vssd1 vssd1 vccd1 vccd1 _4419_/B
+ sky130_fd_sc_hd__o311a_1
X_5384_ _5387_/B _5251_/A _5382_/Y _5383_/Y _5556_/C1 vssd1 vssd1 vccd1 vccd1 _6223_/D
+ sky130_fd_sc_hd__o221a_1
X_4335_ _4335_/A _4363_/A vssd1 vssd1 vccd1 vccd1 _4336_/C sky130_fd_sc_hd__xor2_1
Xfanout205 _3136_/Y vssd1 vssd1 vccd1 vccd1 _3257_/B sky130_fd_sc_hd__buf_8
Xfanout216 _3024_/Y vssd1 vssd1 vccd1 vccd1 _3880_/B sky130_fd_sc_hd__buf_6
Xfanout227 _6293_/Q vssd1 vssd1 vccd1 vccd1 _5436_/A sky130_fd_sc_hd__buf_6
Xfanout238 _6289_/Q vssd1 vssd1 vccd1 vccd1 _5911_/A sky130_fd_sc_hd__buf_12
XFILLER_113_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout249 _5859_/A vssd1 vssd1 vccd1 vccd1 _4362_/A sky130_fd_sc_hd__buf_12
X_4266_ _4266_/A _4266_/B vssd1 vssd1 vccd1 vccd1 _4268_/A sky130_fd_sc_hd__or2_4
XANTENNA__4974__B _6004_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6005_ _6007_/CLK _6005_/D vssd1 vssd1 vccd1 vccd1 _6005_/Q sky130_fd_sc_hd__dfxtp_4
X_3217_ _3212_/A _3156_/Y _5464_/A _3216_/X _3706_/A vssd1 vssd1 vccd1 vccd1 _3218_/D
+ sky130_fd_sc_hd__o32a_1
X_4197_ _4197_/A _4197_/B _4426_/B _4410_/D vssd1 vssd1 vccd1 vccd1 _4275_/A sky130_fd_sc_hd__nand4_4
XFILLER_55_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5151__A _5192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3148_ _3880_/A _4577_/A vssd1 vssd1 vccd1 vccd1 _3148_/X sky130_fd_sc_hd__or2_1
XFILLER_39_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4990__A _4990_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3079_ _5258_/A _5605_/C vssd1 vssd1 vccd1 vccd1 _3079_/Y sky130_fd_sc_hd__nor2_2
XFILLER_42_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5621__B1 _3736_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_759 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4214__B _4214_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5326__A _6222_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3772__C _4539_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5152__A2 _5158_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3280__S _3709_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5915__A1 _3312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5935__S _5943_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5236__A _5236_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4120_ _4154_/A vssd1 vssd1 vccd1 vccd1 _4122_/A sky130_fd_sc_hd__inv_2
XFILLER_96_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4794__B _5041_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4051_ _4050_/X _3869_/A _4051_/S vssd1 vssd1 vccd1 vccd1 _6067_/D sky130_fd_sc_hd__mux2_1
XFILLER_111_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput5 io_in[4] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__buf_4
XFILLER_77_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3002_ _3766_/A vssd1 vssd1 vccd1 vccd1 _3732_/A sky130_fd_sc_hd__clkinv_4
XFILLER_49_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4406__B2 _4437_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4953_ _5002_/C _4953_/B vssd1 vssd1 vccd1 vccd1 _4959_/B sky130_fd_sc_hd__or2_1
XFILLER_33_862 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3904_ _6044_/Q _3715_/X _3909_/S vssd1 vssd1 vccd1 vccd1 _6044_/D sky130_fd_sc_hd__mux2_1
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3857__C _3952_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4884_ _4882_/Y _4883_/Y _4886_/B vssd1 vssd1 vccd1 vccd1 _4884_/Y sky130_fd_sc_hd__a21oi_1
X_3835_ _5428_/A _3834_/B _3737_/Y _3834_/Y vssd1 vssd1 vccd1 vccd1 _3835_/X sky130_fd_sc_hd__a211o_1
XANTENNA__5906__A1 _5883_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4034__B _5925_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3766_ _3766_/A _5503_/A vssd1 vssd1 vccd1 vccd1 _3766_/Y sky130_fd_sc_hd__nand2_2
XANTENNA_fanout126_A _5714_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5505_ _6227_/Q _5504_/C _5504_/A vssd1 vssd1 vccd1 vccd1 _5505_/Y sky130_fd_sc_hd__a21oi_1
X_3697_ _5387_/A _6024_/Q _3902_/A vssd1 vssd1 vccd1 vccd1 _3697_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5436_ _5436_/A _6155_/Q _5436_/C vssd1 vssd1 vccd1 vccd1 _5436_/X sky130_fd_sc_hd__and3_1
XFILLER_133_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5367_ _5367_/A _5367_/B vssd1 vssd1 vccd1 vccd1 _5367_/X sky130_fd_sc_hd__or2_1
XFILLER_59_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4318_ _4318_/A _4318_/B vssd1 vssd1 vccd1 vccd1 _4320_/B sky130_fd_sc_hd__xnor2_4
XFILLER_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5298_ _5295_/Y _5296_/X _5262_/X _5265_/Y vssd1 vssd1 vccd1 vccd1 _5298_/X sky130_fd_sc_hd__a211o_1
XFILLER_59_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4249_ _5767_/C _4251_/B vssd1 vssd1 vccd1 vccd1 _4252_/A sky130_fd_sc_hd__or2_4
XFILLER_75_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5842__B1 _5866_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3113__B _4605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4948__A2 _4972_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4030__C1 _5883_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3783__B _3783_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4636__A1 _3116_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3439__A2 _3257_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3958__B _4604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4939__A2 _4644_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5597__C1 _5948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5061__A1 _4604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_832 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5349__C1 _5929_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5665__S _5703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3620_ _3619_/A _3619_/C _3619_/B vssd1 vssd1 vccd1 vccd1 _3653_/A sky130_fd_sc_hd__a21oi_2
X_3551_ _6279_/Q _6115_/Q _3551_/S vssd1 vssd1 vccd1 vccd1 _5428_/B sky130_fd_sc_hd__mux2_4
XFILLER_6_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6270_ _6270_/CLK _6270_/D vssd1 vssd1 vccd1 vccd1 _6270_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5116__A2 _5241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3482_ _6076_/Q _5743_/B _3480_/X _3236_/Y _3481_/X vssd1 vssd1 vccd1 vccd1 _3482_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_115_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5221_ _5221_/A _5221_/B vssd1 vssd1 vccd1 vccd1 _5221_/Y sky130_fd_sc_hd__nor2_1
XFILLER_88_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5152_ _5238_/A _5158_/B _5136_/C vssd1 vssd1 vccd1 vccd1 _5152_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_96_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4103_ _4103_/A _4103_/B vssd1 vssd1 vccd1 vccd1 _4103_/X sky130_fd_sc_hd__xor2_2
XFILLER_110_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5083_ _5083_/A _5083_/B vssd1 vssd1 vccd1 vccd1 _5083_/Y sky130_fd_sc_hd__nand2_1
XFILLER_56_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4627__A1 _3030_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3214__A _3948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4034_ _5742_/C _5925_/A vssd1 vssd1 vccd1 vccd1 _4475_/S sky130_fd_sc_hd__or2_4
XFILLER_110_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5985_ _5985_/A _5985_/B _5985_/C vssd1 vssd1 vccd1 vccd1 _5985_/X sky130_fd_sc_hd__or3_1
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4936_ _4990_/A _4934_/X _4935_/Y vssd1 vssd1 vccd1 vccd1 _4936_/X sky130_fd_sc_hd__a21o_1
XFILLER_52_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout243_A _5862_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4260__C1 _4214_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4867_ _4867_/A _4867_/B vssd1 vssd1 vccd1 vccd1 _4867_/X sky130_fd_sc_hd__xor2_2
XFILLER_138_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3818_ _3937_/D _3841_/S _3817_/X vssd1 vssd1 vccd1 vccd1 _3819_/B sky130_fd_sc_hd__o21ai_4
X_4798_ _5358_/A _5871_/C _4797_/X _4931_/B vssd1 vssd1 vccd1 vccd1 _4798_/X sky130_fd_sc_hd__o22a_1
XFILLER_21_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3366__A1 _3388_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3749_ _4592_/B _3749_/B _3749_/C vssd1 vssd1 vccd1 vccd1 _3749_/X sky130_fd_sc_hd__and3_4
XFILLER_106_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5419_ _5446_/B _5420_/B vssd1 vssd1 vccd1 vccd1 _5480_/C sky130_fd_sc_hd__and2_4
XFILLER_114_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3124__A _5097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5043__A1 _5567_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5043__B2 _4638_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_16_clk_A _6233_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5346__A2 _5227_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3960__C _3960_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4609__A1 _5241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3034__A _5119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5282__A1 _5929_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3969__A _4596_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5770_ _6251_/Q _5788_/B vssd1 vssd1 vccd1 vccd1 _5770_/X sky130_fd_sc_hd__or2_1
XTAP_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3596__A1 _3599_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4721_ _6186_/Q _4721_/B vssd1 vssd1 vccd1 vccd1 _4721_/X sky130_fd_sc_hd__or2_1
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3596__B2 _3387_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4652_ _5255_/B _4644_/Y _4651_/X _4644_/A _5090_/A vssd1 vssd1 vccd1 vccd1 _4652_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_30_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3603_ _3398_/A _3643_/A _3602_/X _3498_/S vssd1 vssd1 vccd1 vccd1 _3603_/X sky130_fd_sc_hd__o211a_1
X_4583_ _5911_/B _3879_/X _4582_/Y _4654_/A _4581_/X vssd1 vssd1 vccd1 vccd1 _4583_/X
+ sky130_fd_sc_hd__o221a_2
XFILLER_116_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3534_ _6263_/Q _5439_/A2 _5924_/B _6032_/Q vssd1 vssd1 vccd1 vccd1 _3534_/X sky130_fd_sc_hd__o22a_1
X_6253_ _6257_/CLK _6253_/D vssd1 vssd1 vccd1 vccd1 _6253_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3465_ _3465_/A _3465_/B vssd1 vssd1 vccd1 vccd1 _3466_/B sky130_fd_sc_hd__nor2_1
XFILLER_88_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5204_ _5136_/C _5203_/A _5097_/A vssd1 vssd1 vccd1 vccd1 _5204_/Y sky130_fd_sc_hd__a21oi_1
X_6184_ _6193_/CLK _6184_/D vssd1 vssd1 vccd1 vccd1 _6184_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_69_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3396_ _5818_/A _3555_/B _3396_/C vssd1 vssd1 vccd1 vccd1 _3396_/X sky130_fd_sc_hd__and3_1
XANTENNA__5143__B _5143_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5135_ _4046_/A _3072_/A _4648_/Y _5227_/A vssd1 vssd1 vccd1 vccd1 _5136_/B sky130_fd_sc_hd__a211o_1
XFILLER_97_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5066_ _4604_/A _3971_/B _3974_/C vssd1 vssd1 vccd1 vccd1 _5066_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__5273__A1 _5258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4017_ _6302_/Q _3033_/Y _4767_/A _6301_/Q _4016_/X vssd1 vssd1 vccd1 vccd1 _4017_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_37_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5576__A2 _5250_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5968_ _5114_/Y _5970_/A _6298_/Q vssd1 vssd1 vccd1 vccd1 _5968_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_40_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4784__B1 _3116_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4919_ _4745_/Y _4915_/X _4918_/Y _4705_/A _3116_/X vssd1 vssd1 vccd1 vccd1 _4931_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_21_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5899_ _5900_/A _5900_/B _5896_/Y _5897_/Y _5898_/Y vssd1 vssd1 vccd1 vccd1 _5899_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_21_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3119__A _5050_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4423__A1_N _3842_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3553__S _3709_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4839__A1 _5392_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5060__A2_N _5244_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5053__B _5731_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3814__A2 _3777_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3301__B _3952_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4775__A0 _5119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3578__A1 _3567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3728__S _3731_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5319__A2 _5349_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3029__A _4990_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3971__B _3971_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5244__A _5244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3250_ _3590_/A1 _3248_/X _3249_/X _3247_/X vssd1 vssd1 vccd1 vccd1 _3250_/X sky130_fd_sc_hd__a31o_4
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3181_ _4638_/A _5840_/A vssd1 vssd1 vccd1 vccd1 _4587_/B sky130_fd_sc_hd__nand2_8
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5898__B _5898_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5822_ _5835_/A1 _4331_/X _5819_/Y _6274_/Q vssd1 vssd1 vccd1 vccd1 _5822_/X sky130_fd_sc_hd__a22o_1
XFILLER_90_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5753_ _3011_/Y _5763_/B _5742_/Y vssd1 vssd1 vccd1 vccd1 _5753_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_50_779 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5419__A _5446_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4704_ _4742_/B _4704_/B vssd1 vssd1 vccd1 vccd1 _4716_/B sky130_fd_sc_hd__or2_1
X_5684_ _5681_/X _5682_/X _5683_/X vssd1 vssd1 vccd1 vccd1 _5684_/X sky130_fd_sc_hd__a21o_1
XANTENNA__4518__A0 _5446_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4635_ _6184_/Q _4744_/B _5050_/B _4634_/X _5051_/D vssd1 vssd1 vccd1 vccd1 _4635_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_135_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout206_A _3734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4566_ _3114_/C _4566_/B _4605_/B vssd1 vssd1 vccd1 vccd1 _5839_/A sky130_fd_sc_hd__and3b_1
XANTENNA__4469__S _4477_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3517_ _3935_/C _3516_/B _3312_/Y vssd1 vssd1 vccd1 vccd1 _3517_/X sky130_fd_sc_hd__o21a_1
XFILLER_116_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4497_ _4872_/A _4239_/A _4059_/B vssd1 vssd1 vccd1 vccd1 _4497_/X sky130_fd_sc_hd__o21a_1
XFILLER_103_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6236_ _6241_/CLK _6236_/D vssd1 vssd1 vccd1 vccd1 _6236_/Q sky130_fd_sc_hd__dfxtp_1
X_3448_ _3448_/A _3450_/D vssd1 vssd1 vccd1 vccd1 _3448_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_134_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6167_ _6170_/CLK _6167_/D vssd1 vssd1 vccd1 vccd1 _6167_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3379_ _6096_/Q _3589_/A2 _3589_/B1 _6089_/Q vssd1 vssd1 vccd1 vccd1 _3379_/X sky130_fd_sc_hd__o22a_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5118_ _5117_/Y _6204_/Q _5129_/S vssd1 vssd1 vccd1 vccd1 _6204_/D sky130_fd_sc_hd__mux2_1
X_6098_ _6098_/CLK _6098_/D vssd1 vssd1 vccd1 vccd1 _6098_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5246__A1 _5075_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5049_ _5049_/A _5051_/D vssd1 vssd1 vccd1 vccd1 _5052_/A sky130_fd_sc_hd__nor2_1
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3121__B _3121_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_787 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5485__A1 _5072_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5237__B2 _5236_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3248__B1 _5924_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3312__A _3312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3799__A1 _3033_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4460__A2 _3900_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5239__A _5239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3685__C _5743_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4143__A _4163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5960__A2 _3975_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3982__A _5239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4420_ _4431_/B _4420_/B vssd1 vssd1 vccd1 vccd1 _4420_/X sky130_fd_sc_hd__and2_1
XANTENNA__5173__B1 _5136_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3723__A1 _4112_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3723__B2 _5567_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4351_ _4351_/A _4351_/B vssd1 vssd1 vccd1 vccd1 _4353_/B sky130_fd_sc_hd__nor2_1
X_3302_ _3312_/A _3952_/B vssd1 vssd1 vccd1 vccd1 _3511_/A sky130_fd_sc_hd__nand2_8
XFILLER_113_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5405__C _5436_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4282_ _4283_/A _4283_/B vssd1 vssd1 vccd1 vccd1 _4321_/B sky130_fd_sc_hd__and2_2
XFILLER_98_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6021_ _6254_/CLK _6021_/D vssd1 vssd1 vccd1 vccd1 _6021_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3233_ _5936_/A _3706_/A _5734_/A vssd1 vssd1 vccd1 vccd1 _3251_/B sky130_fd_sc_hd__or3_4
XANTENNA_clkbuf_3_3__f_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3921__S _3921_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3487__B1 _5392_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3164_ _3205_/A _3212_/A _3164_/C vssd1 vssd1 vccd1 vccd1 _3164_/Y sky130_fd_sc_hd__nor3_2
XFILLER_104_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3095_ _6217_/Q _4705_/A vssd1 vssd1 vccd1 vccd1 _4999_/B sky130_fd_sc_hd__nor2_8
XANTENNA__3222__A _3706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4451__A2 _3900_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout156_A _3069_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout38 _4721_/B vssd1 vssd1 vccd1 vccd1 _5046_/B sky130_fd_sc_hd__buf_4
XANTENNA__3876__B _5138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout49 _5766_/C vssd1 vssd1 vccd1 vccd1 _5767_/C sky130_fd_sc_hd__buf_6
X_5805_ _5817_/A1 _4078_/Y _5804_/X vssd1 vssd1 vccd1 vccd1 _6266_/D sky130_fd_sc_hd__a21o_1
XANTENNA__5400__A1 _5498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4203__A2 _4309_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3997_ _4697_/A _5114_/A _5119_/A _5392_/A vssd1 vssd1 vccd1 vccd1 _3998_/D sky130_fd_sc_hd__or4_1
XFILLER_10_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5736_ _5710_/S _3280_/X _5735_/X _3772_/B _5734_/X vssd1 vssd1 vccd1 vccd1 _5736_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout323_A input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3962__A1 _3880_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5667_ _5730_/A _3937_/C _5666_/X vssd1 vssd1 vccd1 vccd1 _5675_/A sky130_fd_sc_hd__o21a_1
XFILLER_136_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4618_ _4618_/A _4618_/B _4618_/C _5062_/B vssd1 vssd1 vccd1 vccd1 _4625_/A sky130_fd_sc_hd__or4b_4
X_5598_ _6233_/Q _5598_/B vssd1 vssd1 vccd1 vccd1 _5598_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_135_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_606 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3714__A1 _5504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3714__B2 _5743_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4549_ _5926_/A0 _4564_/A2 _4547_/X _4548_/Y vssd1 vssd1 vccd1 vccd1 _6175_/D sky130_fd_sc_hd__a22o_1
XFILLER_104_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3116__B _3116_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6219_ _6219_/CLK _6219_/D vssd1 vssd1 vccd1 vccd1 _6219_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4442__A2 _3900_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3278__S _3551_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5942__A2 _4586_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4902__B1 _5239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4410__B _4410_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5458__A1 _5498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5522__A _5540_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4130__A1 _4163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5241__B _5241_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3977__A _5191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3920_ _6055_/Q _3727_/X _3921_/S vssd1 vssd1 vccd1 vccd1 _6055_/D sky130_fd_sc_hd__mux2_1
XFILLER_44_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3851_ _4883_/B _3751_/A _3816_/B _3850_/X vssd1 vssd1 vccd1 vccd1 _3851_/X sky130_fd_sc_hd__o211a_1
XFILLER_32_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3782_ _3748_/Y _3780_/X _3781_/X vssd1 vssd1 vccd1 vccd1 _3783_/B sky130_fd_sc_hd__o21ai_4
XANTENNA__5933__A2 _4586_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5521_ _3008_/Y _4990_/B _5539_/S vssd1 vssd1 vccd1 vccd1 _5521_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3916__S _3921_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5452_ _5452_/A _5452_/B vssd1 vssd1 vccd1 vccd1 _5453_/B sky130_fd_sc_hd__nor2_1
XANTENNA__4601__A _5090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4403_ _4382_/A _4382_/B _4383_/S _4384_/A vssd1 vssd1 vccd1 vccd1 _4405_/B sky130_fd_sc_hd__o31ai_2
XFILLER_117_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5383_ _5943_/C _5358_/Y _5251_/A vssd1 vssd1 vccd1 vccd1 _5383_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_99_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4334_ _4334_/A _4410_/D vssd1 vssd1 vccd1 vccd1 _4363_/A sky130_fd_sc_hd__nand2_2
XFILLER_113_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout206 _3734_/A vssd1 vssd1 vccd1 vccd1 _4462_/A sky130_fd_sc_hd__buf_12
XFILLER_87_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout217 _5131_/A vssd1 vssd1 vccd1 vccd1 _4046_/A sky130_fd_sc_hd__buf_6
Xfanout228 _6293_/Q vssd1 vssd1 vccd1 vccd1 _5924_/A sky130_fd_sc_hd__buf_6
XFILLER_86_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4265_ _4362_/A _4334_/A _4309_/B _4342_/B vssd1 vssd1 vccd1 vccd1 _4266_/B sky130_fd_sc_hd__and4_1
Xfanout239 _5128_/A0 vssd1 vssd1 vccd1 vccd1 _5790_/A1 sky130_fd_sc_hd__buf_8
XFILLER_115_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6004_ _6007_/CLK _6004_/D vssd1 vssd1 vccd1 vccd1 _6004_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_39_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3216_ _5840_/A _5653_/A _4806_/S _3221_/D vssd1 vssd1 vccd1 vccd1 _3216_/X sky130_fd_sc_hd__or4_1
X_4196_ _4197_/B _3280_/X _4167_/D _4197_/A vssd1 vssd1 vccd1 vccd1 _4199_/B sky130_fd_sc_hd__a22o_2
XFILLER_54_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4048__A _5733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3147_ _3880_/A _3948_/A vssd1 vssd1 vccd1 vccd1 _3147_/Y sky130_fd_sc_hd__nor2_1
XFILLER_28_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3078_ _3105_/A _5239_/B vssd1 vssd1 vccd1 vccd1 _3078_/Y sky130_fd_sc_hd__nand2_2
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5621__A1 _4614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3887__A _5097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_863 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5719_ _4846_/B _4837_/B _5731_/S vssd1 vssd1 vccd1 vccd1 _5719_/X sky130_fd_sc_hd__mux2_1
XFILLER_108_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5688__A1 _4162_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3699__A0 _5446_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3772__D _5191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4360__B2 _4437_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5860__A1 _3597_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5612__A1 _5412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5915__A2 _5238_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5128__A0 _5128_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3037__A _5428_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4050_ _4657_/A _5075_/A _4596_/B vssd1 vssd1 vccd1 vccd1 _4050_/X sky130_fd_sc_hd__mux2_1
X_3001_ _6299_/Q vssd1 vssd1 vccd1 vccd1 _5656_/A sky130_fd_sc_hd__clkinv_2
Xinput6 io_in[5] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__buf_4
XFILLER_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3203__C _4614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5064__C1 _5148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4952_ _6193_/Q _4952_/B vssd1 vssd1 vccd1 vccd1 _4953_/B sky130_fd_sc_hd__nor2_1
XFILLER_33_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3500__A _3500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3903_ _6043_/Q _3711_/X _3909_/S vssd1 vssd1 vccd1 vccd1 _6043_/D sky130_fd_sc_hd__mux2_1
XFILLER_33_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4883_ _5454_/A _4883_/B vssd1 vssd1 vccd1 vccd1 _4883_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_32_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3834_ _5721_/B _3834_/B vssd1 vssd1 vccd1 vccd1 _3834_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__3917__A1 _3718_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3765_ _5108_/B _3765_/B _4072_/B vssd1 vssd1 vccd1 vccd1 _3765_/X sky130_fd_sc_hd__or3_4
XFILLER_118_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5504_ _5504_/A _6227_/Q _5504_/C vssd1 vssd1 vccd1 vccd1 _5547_/C sky130_fd_sc_hd__and3_2
X_3696_ _5856_/A _3695_/X _3705_/A vssd1 vssd1 vccd1 vccd1 _6023_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4761__A1_N _3011_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout119_A _3388_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5435_ _5432_/Y _5433_/X _5434_/X vssd1 vssd1 vccd1 vccd1 _5435_/X sky130_fd_sc_hd__a21o_1
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5366_ _5367_/A _5367_/B vssd1 vssd1 vccd1 vccd1 _5366_/Y sky130_fd_sc_hd__nand2_1
XFILLER_102_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4477__S _4477_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4317_ _4318_/B _4318_/A vssd1 vssd1 vccd1 vccd1 _4351_/A sky130_fd_sc_hd__and2b_1
XANTENNA__4776__A1_N _3101_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5297_ _5262_/X _5265_/Y _5295_/Y _5296_/X vssd1 vssd1 vccd1 vccd1 _5297_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_87_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4248_ _5767_/C _4251_/B vssd1 vssd1 vccd1 vccd1 _4553_/B sky130_fd_sc_hd__nor2_1
XFILLER_87_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4179_ _4180_/A _4180_/B _4180_/C vssd1 vssd1 vccd1 vccd1 _4181_/B sky130_fd_sc_hd__a21o_2
XFILLER_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_3__f_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _6219_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_128_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3908__A1 _3727_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4581__B2 _3060_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4333__A1 _3783_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5530__B1 _5522_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5072__A _5072_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4097__B1 _4112_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5833__A1 _5835_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4636__A2 _4631_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3304__B _3869_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5800__A _5800_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5349__B1 _5349_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_844 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3974__B _3974_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3375__A2 _5653_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3550_ _3549_/B _5706_/B _3549_/Y _3211_/Y vssd1 vssd1 vccd1 vccd1 _3550_/X sky130_fd_sc_hd__a211o_1
XFILLER_6_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3481_ _6098_/Q _3589_/A2 _3589_/B1 _6091_/Q vssd1 vssd1 vccd1 vccd1 _3481_/X sky130_fd_sc_hd__o22a_1
XFILLER_115_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5220_ _5256_/B _5219_/X _5220_/S vssd1 vssd1 vccd1 vccd1 _5220_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5151_ _5192_/A _5151_/B vssd1 vssd1 vccd1 vccd1 _6210_/D sky130_fd_sc_hd__nor2_1
XFILLER_97_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4102_ _4103_/A _4103_/B vssd1 vssd1 vccd1 vccd1 _4125_/A sky130_fd_sc_hd__or2_2
XFILLER_97_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5082_ _4589_/A _5104_/B _4597_/Y _5081_/X vssd1 vssd1 vccd1 vccd1 _5083_/B sky130_fd_sc_hd__o211a_1
XFILLER_96_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5285__C1 _3122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3214__B _5512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5824__A1 _5835_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4627__A2 _4812_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4033_ _5436_/A _5742_/B vssd1 vssd1 vccd1 vccd1 _5925_/A sky130_fd_sc_hd__or2_4
XFILLER_56_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5037__C1 _5227_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3230__A _4539_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5984_ _5114_/Y _5985_/C _6302_/Q vssd1 vssd1 vccd1 vccd1 _5984_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_24_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4935_ _6192_/Q _4990_/A _4640_/Y vssd1 vssd1 vccd1 vccd1 _4935_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__4260__B1 _4216_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4866_ _4820_/B _4829_/B _4860_/B vssd1 vssd1 vccd1 vccd1 _4867_/B sky130_fd_sc_hd__a21bo_4
XANTENNA_fanout236_A _5911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3817_ _3815_/X _3816_/X _3748_/Y vssd1 vssd1 vccd1 vccd1 _3817_/X sky130_fd_sc_hd__a21o_1
XFILLER_119_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4797_ _5358_/A _4587_/B _4786_/X _4796_/X vssd1 vssd1 vccd1 vccd1 _4797_/X sky130_fd_sc_hd__o211a_1
XANTENNA__4012__B1 _3513_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4563__A1 _4891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3748_ _3841_/S vssd1 vssd1 vccd1 vccd1 _3748_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_119_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3679_ _3974_/B _5172_/A _5330_/B vssd1 vssd1 vccd1 vccd1 _3679_/X sky130_fd_sc_hd__or3_1
XFILLER_133_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5418_ _4872_/A _4867_/X _5539_/S vssd1 vssd1 vccd1 vccd1 _5418_/X sky130_fd_sc_hd__mux2_4
XFILLER_121_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3523__C1 _3145_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5349_ _6120_/Q _4234_/B _5349_/B1 _6022_/Q _5929_/B2 vssd1 vssd1 vccd1 vccd1 _5349_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_102_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4079__B1 _4072_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5276__C1 _5607_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3124__B _5192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4236__A _5767_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3140__A _4462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5043__A2 _5463_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_50_clk _6230_/CLK vssd1 vssd1 vccd1 vccd1 _6154_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_129_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5200__C1 _5097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4554__A1 _3010_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4306__A1 _4301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5806__A1 _3425_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3969__B _4605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4720_ _5051_/D _4705_/Y _4711_/X _4719_/X vssd1 vssd1 vccd1 vccd1 _4720_/X sky130_fd_sc_hd__o31a_1
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_41_clk clkbuf_3_4__f_clk/X vssd1 vssd1 vccd1 vccd1 _6293_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_30_663 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4651_ _4647_/Y _4650_/X _4640_/A _4637_/X vssd1 vssd1 vccd1 vccd1 _4651_/X sky130_fd_sc_hd__o2bb2a_1
X_3602_ _5428_/A _3495_/A _3211_/Y _3601_/Y vssd1 vssd1 vccd1 vccd1 _3602_/X sky130_fd_sc_hd__a211o_1
XANTENNA__4545__A1 _4672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4582_ _5605_/C _3996_/B _4587_/B vssd1 vssd1 vccd1 vccd1 _4582_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_116_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3533_ _6099_/Q _3901_/B _3704_/B _6092_/Q _5470_/S vssd1 vssd1 vccd1 vccd1 _3533_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__3209__B _5617_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6252_ _6257_/CLK _6252_/D vssd1 vssd1 vccd1 vccd1 _6252_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3464_ _3926_/A _3464_/B vssd1 vssd1 vccd1 vccd1 _3465_/B sky130_fd_sc_hd__nor2_1
XFILLER_115_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5203_ _5203_/A _5203_/B _5203_/C _5647_/B vssd1 vssd1 vccd1 vccd1 _5203_/X sky130_fd_sc_hd__or4b_1
X_6183_ _6290_/CLK _6183_/D vssd1 vssd1 vccd1 vccd1 _6183_/Q sky130_fd_sc_hd__dfxtp_1
X_3395_ _6268_/Q _6014_/Q _6082_/Q _6037_/Q _4067_/A _3709_/S vssd1 vssd1 vccd1 vccd1
+ _3396_/C sky130_fd_sc_hd__mux4_1
XANTENNA__3225__A _3555_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5134_ _3062_/Y _5131_/Y _5133_/X _5638_/A vssd1 vssd1 vccd1 vccd1 _5134_/X sky130_fd_sc_hd__o211a_1
XFILLER_85_803 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5065_ _5065_/A _5065_/B vssd1 vssd1 vccd1 vccd1 _5069_/B sky130_fd_sc_hd__nand2_1
XFILLER_123_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout186_A _4111_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4016_ _6295_/Q _3030_/Y _4850_/A _6300_/Q vssd1 vssd1 vccd1 vccd1 _4016_/X sky130_fd_sc_hd__o22a_1
XANTENNA__3879__B _4587_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4056__A _5436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5967_ _5964_/Y _5966_/X _5986_/B1 vssd1 vssd1 vccd1 vccd1 _6297_/D sky130_fd_sc_hd__a21oi_1
XANTENNA__3587__A2 _3589_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4918_ _4952_/B _4918_/B vssd1 vssd1 vccd1 vccd1 _4918_/Y sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_32_clk clkbuf_3_5__f_clk/X vssd1 vssd1 vccd1 vccd1 _6143_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__5981__B1 _6301_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5898_ _5898_/A _5898_/B vssd1 vssd1 vccd1 vccd1 _5898_/Y sky130_fd_sc_hd__nand2_1
XFILLER_32_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5408__S0 _3241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3992__C1 _3179_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4849_ _4849_/A _4849_/B vssd1 vssd1 vccd1 vccd1 _4849_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_4_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout99_A _3060_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4839__A2 _5703_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4472__A0 _5387_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3275__A1 _5226_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5185__D1 _3958_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5244__B _5244_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3180_ _4577_/A _5065_/A vssd1 vssd1 vccd1 vccd1 _3180_/Y sky130_fd_sc_hd__nor2_2
XFILLER_39_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4575__S _4575_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4463__A0 _3943_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5660__C1 _3996_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5821_ _3322_/X _5819_/B _5820_/X vssd1 vssd1 vccd1 vccd1 _6273_/D sky130_fd_sc_hd__a21o_1
XANTENNA__3919__S _3921_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5752_ _6245_/Q _5763_/B vssd1 vssd1 vccd1 vccd1 _5752_/X sky130_fd_sc_hd__or2_1
XANTENNA__4604__A _4604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_14_clk _6233_/CLK vssd1 vssd1 vccd1 vccd1 _6299_/CLK sky130_fd_sc_hd__clkbuf_16
X_4703_ _6185_/Q _6184_/Q _6186_/Q vssd1 vssd1 vccd1 vccd1 _4704_/B sky130_fd_sc_hd__a21oi_1
XFILLER_30_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5683_ _3867_/B _5848_/A0 _3513_/B _3867_/A _3996_/B vssd1 vssd1 vccd1 vccd1 _5683_/X
+ sky130_fd_sc_hd__a221o_1
X_4634_ _4678_/A _4675_/A vssd1 vssd1 vccd1 vccd1 _4634_/X sky130_fd_sc_hd__and2_2
XFILLER_8_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5715__B1 _5728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4565_ _5238_/C _4753_/A vssd1 vssd1 vccd1 vccd1 _4605_/B sky130_fd_sc_hd__nand2_2
XFILLER_104_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3516_ _3935_/C _3516_/B vssd1 vssd1 vccd1 vccd1 _3516_/Y sky130_fd_sc_hd__nand2_1
X_4496_ _6139_/Q _4499_/B vssd1 vssd1 vccd1 vccd1 _4496_/X sky130_fd_sc_hd__or2_1
XFILLER_116_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6235_ _6270_/CLK _6235_/D vssd1 vssd1 vccd1 vccd1 _6235_/Q sky130_fd_sc_hd__dfxtp_1
X_3447_ _3446_/X _4162_/A _3560_/S vssd1 vssd1 vccd1 vccd1 _3447_/X sky130_fd_sc_hd__mux2_1
XFILLER_103_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6166_ _6170_/CLK _6166_/D vssd1 vssd1 vccd1 vccd1 _6166_/Q sky130_fd_sc_hd__dfxtp_1
X_3378_ _5924_/A _6061_/Q _5436_/C vssd1 vssd1 vccd1 vccd1 _3378_/X sky130_fd_sc_hd__and3_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_15_clk_A _6233_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5117_ _5985_/A vssd1 vssd1 vccd1 vccd1 _5117_/Y sky130_fd_sc_hd__inv_2
X_6097_ _6098_/CLK _6097_/D vssd1 vssd1 vccd1 vccd1 _6097_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5048_ _4618_/A _5048_/B _5048_/C vssd1 vssd1 vccd1 vccd1 _5250_/A sky130_fd_sc_hd__and3b_1
XFILLER_84_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4757__A1 _5543_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5048__C _5048_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5182__A1 _5143_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3496__A1 _4767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4693__B1 _4842_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3312__B _3312_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4996__A1 _5547_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5945__B1 _5944_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5239__B _5239_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4143__B _4176_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5255__A _5292_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4350_ _4350_/A _4350_/B vssd1 vssd1 vccd1 vccd1 _4353_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__3723__A2 _5742_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3301_ _3312_/A _3952_/B vssd1 vssd1 vccd1 vccd1 _3422_/A sky130_fd_sc_hd__and2_4
XFILLER_113_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4281_ _4281_/A _4281_/B vssd1 vssd1 vccd1 vccd1 _4283_/B sky130_fd_sc_hd__xnor2_2
X_6020_ _6257_/CLK _6020_/D vssd1 vssd1 vccd1 vccd1 _6020_/Q sky130_fd_sc_hd__dfxtp_1
X_3232_ _5570_/A _5734_/A vssd1 vssd1 vccd1 vccd1 _5928_/A sky130_fd_sc_hd__nor2_2
XFILLER_67_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3487__A1 _4202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3487__B2 _3053_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3163_ _3575_/B _3163_/B vssd1 vssd1 vccd1 vccd1 _3164_/C sky130_fd_sc_hd__or2_4
XFILLER_94_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3094_ _5051_/B _5051_/C vssd1 vssd1 vccd1 vccd1 _4705_/A sky130_fd_sc_hd__or2_4
XFILLER_48_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4739__A1 _3033_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5804_ _3375_/X _5801_/B _5801_/Y _6266_/Q vssd1 vssd1 vccd1 vccd1 _5804_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4334__A _4334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout39 _4970_/B vssd1 vssd1 vccd1 vccd1 _4721_/B sky130_fd_sc_hd__buf_2
XANTENNA_fanout149_A _5476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3996_ _4850_/A _3996_/B vssd1 vssd1 vccd1 vccd1 _3998_/C sky130_fd_sc_hd__nand2_1
XANTENNA__3947__C1 _3941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5735_ _6058_/Q _6218_/Q _5735_/S vssd1 vssd1 vccd1 vccd1 _5735_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3962__A2 _5870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout316_A _4576_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5666_ _5718_/A _5665_/X _5732_/C1 vssd1 vssd1 vccd1 vccd1 _5666_/X sky130_fd_sc_hd__o21a_1
XFILLER_108_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4617_ _5062_/A _5083_/A _4617_/C vssd1 vssd1 vccd1 vccd1 _4618_/C sky130_fd_sc_hd__nand3_1
XFILLER_135_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5597_ _6232_/Q _5250_/X _5595_/Y _5596_/X _5948_/A vssd1 vssd1 vccd1 vccd1 _6232_/D
+ sky130_fd_sc_hd__o221a_1
XANTENNA__5165__A _5635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4548_ _5305_/A _4562_/B _4564_/A2 vssd1 vssd1 vccd1 vccd1 _4548_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_2_618 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3270__S0 _4067_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4479_ _5221_/A _4499_/B _4057_/Y vssd1 vssd1 vccd1 vccd1 _4479_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_89_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5467__A2 _3901_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6218_ _6218_/CLK _6218_/D vssd1 vssd1 vccd1 vccd1 _6218_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5872__C1 _5206_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6149_ _6154_/CLK _6149_/D vssd1 vssd1 vccd1 vccd1 _6149_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_412 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5155__A1 _4614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5075__A _5075_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4410__C _4426_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5458__A2 _5463_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3469__B2 _3312_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5863__C1 _5867_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4130__A2 _4173_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4969__A1 _5504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4969__B2 _4931_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5091__B1 _5051_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5630__A2 _3388_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3977__B _4596_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3641__A1 _4216_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3850_ _3848_/X _3849_/Y _3740_/X vssd1 vssd1 vccd1 vccd1 _3850_/X sky130_fd_sc_hd__a21o_1
X_3781_ _5653_/B _3841_/S vssd1 vssd1 vccd1 vccd1 _3781_/X sky130_fd_sc_hd__or2_2
X_5520_ _4974_/X _5476_/Y _5519_/Y vssd1 vssd1 vccd1 vccd1 _5520_/X sky130_fd_sc_hd__a21o_1
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5146__A1 _5258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5451_ _5451_/A _5451_/B vssd1 vssd1 vccd1 vccd1 _5453_/A sky130_fd_sc_hd__nand2_1
XANTENNA__4601__B _5069_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4402_ _4419_/A _4402_/B vssd1 vssd1 vccd1 vccd1 _4405_/A sky130_fd_sc_hd__nor2_1
X_5382_ _5412_/A _5358_/Y _5381_/X vssd1 vssd1 vccd1 vccd1 _5382_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_114_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4333_ _3783_/B _4295_/A _4332_/Y vssd1 vssd1 vccd1 vccd1 _6110_/D sky130_fd_sc_hd__o21ai_1
XFILLER_125_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5713__A _5714_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout207 _4022_/C vssd1 vssd1 vccd1 vccd1 _5818_/A sky130_fd_sc_hd__buf_8
Xfanout218 _5210_/B vssd1 vssd1 vccd1 vccd1 _5191_/A sky130_fd_sc_hd__buf_8
XFILLER_99_577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4264_ _4362_/A _4342_/B vssd1 vssd1 vccd1 vccd1 _4310_/A sky130_fd_sc_hd__nand2_1
XFILLER_59_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout229 _5625_/A vssd1 vssd1 vccd1 vccd1 _5090_/A sky130_fd_sc_hd__buf_8
XFILLER_101_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6003_ _6217_/CLK _6003_/D vssd1 vssd1 vccd1 vccd1 _6003_/Q sky130_fd_sc_hd__dfxtp_2
X_3215_ _3940_/A _3215_/B vssd1 vssd1 vccd1 vccd1 _3221_/D sky130_fd_sc_hd__or2_2
XFILLER_86_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4195_ _4270_/A _4389_/B vssd1 vssd1 vccd1 vccd1 _4195_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__3233__A _5936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3146_ _3880_/A _5065_/A _3960_/B vssd1 vssd1 vccd1 vccd1 _5882_/S sky130_fd_sc_hd__or3_4
XFILLER_95_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4409__B1 _4410_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4048__B _5096_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5606__C1 _5227_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3077_ _3105_/A _5239_/B vssd1 vssd1 vccd1 vccd1 _5625_/B sky130_fd_sc_hd__and2_2
XANTENNA_fanout266_A _4197_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5621__A2 _3950_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3887__B _5131_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3979_ _5638_/B _3979_/B _5647_/C vssd1 vssd1 vccd1 vccd1 _3982_/B sky130_fd_sc_hd__and3_1
X_5718_ _5718_/A _5898_/B vssd1 vssd1 vccd1 vccd1 _5718_/Y sky130_fd_sc_hd__nand2_1
XFILLER_136_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5649_ _5649_/A _5649_/B _5649_/C vssd1 vssd1 vccd1 vccd1 _5649_/X sky130_fd_sc_hd__and3_4
XFILLER_108_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5688__A2 _5649_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3127__B _4462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout81_A _3102_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3143__A _4003_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5376__B2 _5595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5128__A1 _5072_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4887__B1 _4972_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5300__A1 _3032_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3053__A _5800_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput7 io_in[6] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__clkbuf_4
XFILLER_25_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5064__B1 _5158_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4951_ _6193_/Q _4952_/B vssd1 vssd1 vccd1 vccd1 _5002_/C sky130_fd_sc_hd__and2_2
XFILLER_33_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3500__B _3500_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3902_ _3902_/A _4439_/S vssd1 vssd1 vccd1 vccd1 _3909_/S sky130_fd_sc_hd__nand2_8
XFILLER_32_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4882_ _4847_/B _4849_/B _4845_/Y vssd1 vssd1 vccd1 vccd1 _4882_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_33_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3833_ _6039_/Q _3771_/X _3831_/Y _3832_/X vssd1 vssd1 vccd1 vccd1 _6039_/D sky130_fd_sc_hd__a211o_1
XANTENNA__4612__A _5239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3764_ _3855_/S _4069_/A vssd1 vssd1 vccd1 vccd1 _3764_/Y sky130_fd_sc_hd__nor2_1
X_5503_ _5503_/A _5503_/B _5503_/C vssd1 vssd1 vccd1 vccd1 _5503_/X sky130_fd_sc_hd__or3_1
XFILLER_9_592 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3695_ _5358_/A _6023_/Q _3902_/A vssd1 vssd1 vccd1 vccd1 _3695_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5434_ _4644_/A _5418_/X _5421_/Y _5464_/A _5607_/B1 vssd1 vssd1 vccd1 vccd1 _5434_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_133_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5365_ _5367_/A _5367_/B vssd1 vssd1 vccd1 vccd1 _5365_/X sky130_fd_sc_hd__and2_1
X_4316_ _4278_/A _4278_/B _4276_/Y vssd1 vssd1 vccd1 vccd1 _4318_/B sky130_fd_sc_hd__o21a_2
XFILLER_59_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5296_ _5296_/A _5296_/B vssd1 vssd1 vccd1 vccd1 _5296_/X sky130_fd_sc_hd__or2_2
XFILLER_113_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4247_ _5767_/A _5436_/C vssd1 vssd1 vccd1 vccd1 _4251_/B sky130_fd_sc_hd__nand2_8
XFILLER_102_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4178_ _4178_/A _4178_/B vssd1 vssd1 vccd1 vccd1 _4180_/C sky130_fd_sc_hd__xnor2_4
XANTENNA__3853__A1 _5900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3129_ _4657_/A _6004_/Q _3135_/S vssd1 vssd1 vccd1 vccd1 _6004_/D sky130_fd_sc_hd__mux2_1
XANTENNA__5055__B1 _4596_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3605__A1 _4214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3410__B _3410_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4522__A _4539_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4030__A1 _5934_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4581__A2 _5638_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3138__A _3766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5530__A1 _5463_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5530__B2 _4596_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5353__A _5353_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5072__B _5072_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4097__A1 _4096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4097__B2 _4197_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5800__B _5818_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5597__A1 _6232_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3974__C _3974_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4021__A1 _4022_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3480_ _5924_/A _6063_/Q _5436_/C vssd1 vssd1 vccd1 vccd1 _3480_/X sky130_fd_sc_hd__and3_1
XFILLER_115_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5263__A _5263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3532__B1 _5743_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5150_ _5191_/A _4046_/A _4577_/D _5149_/X vssd1 vssd1 vccd1 vccd1 _5151_/B sky130_fd_sc_hd__o22a_1
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4101_ _4083_/Y _4087_/A _4099_/X _4123_/A vssd1 vssd1 vccd1 vccd1 _4103_/B sky130_fd_sc_hd__o31ai_4
X_5081_ _5570_/A _4604_/C _4642_/Y _5244_/A _4581_/X vssd1 vssd1 vccd1 vccd1 _5081_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_110_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4627__A3 _4659_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4032_ _3020_/Y _3984_/X _4031_/Y _5932_/A vssd1 vssd1 vccd1 vccd1 _6058_/D sky130_fd_sc_hd__a211oi_1
XFILLER_84_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3835__A1 _5428_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5037__B1 _4648_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3511__A _3511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5588__A1 _6232_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5983_ _5981_/Y _5982_/X _5986_/B1 vssd1 vssd1 vccd1 vccd1 _6301_/D sky130_fd_sc_hd__a21oi_1
XFILLER_18_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4934_ _4934_/A _4934_/B vssd1 vssd1 vccd1 vccd1 _4934_/X sky130_fd_sc_hd__xor2_2
XANTENNA__4796__C1 _5239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4865_ _6190_/Q _3671_/Y _5172_/B _5029_/B _4646_/Y vssd1 vssd1 vccd1 vccd1 _4865_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__4342__A _4426_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3816_ _4767_/B _3816_/B vssd1 vssd1 vccd1 vccd1 _3816_/X sky130_fd_sc_hd__or2_1
XANTENNA__4012__A1 _3032_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4796_ _5358_/A _4643_/Y _4795_/X _4643_/A _5239_/A vssd1 vssd1 vccd1 vccd1 _4796_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4012__B2 _4767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout229_A _5625_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5760__A1 _3942_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4563__A2 _4252_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3747_ _3747_/A _4072_/B vssd1 vssd1 vccd1 vccd1 _3793_/B sky130_fd_sc_hd__or2_4
XFILLER_119_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3678_ _3678_/A _3678_/B _3678_/C vssd1 vssd1 vccd1 vccd1 _3678_/X sky130_fd_sc_hd__or3_1
XFILLER_134_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5417_ _5415_/Y _5416_/X _5507_/A _5327_/A vssd1 vssd1 vccd1 vccd1 _5417_/X sky130_fd_sc_hd__a211o_1
XFILLER_133_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5348_ _6253_/Q _3243_/A _5742_/B _6245_/Q vssd1 vssd1 vccd1 vccd1 _5348_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5279_ _6126_/Q _5767_/B _5277_/X _3236_/Y _5278_/X vssd1 vssd1 vccd1 vccd1 _5279_/X
+ sky130_fd_sc_hd__o221a_2
XFILLER_87_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3826__A1 _4202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5112__S _5124_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3421__A _3960_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout44_A _5839_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4252__A _4252_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5751__A1 _5926_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4306__A2 _4389_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5267__B1 _3059_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3331__A _3331_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output25_A _6198_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4242__A1 _3718_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5258__A _5258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4162__A _4162_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4650_ _6184_/Q _5543_/S _5172_/B _3030_/Y _4646_/Y vssd1 vssd1 vccd1 vccd1 _4650_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_30_675 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3601_ _3636_/A _5721_/B vssd1 vssd1 vccd1 vccd1 _3601_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__4545__A2 _4252_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4581_ _5095_/A _5638_/B _4580_/C _3060_/A _4580_/X vssd1 vssd1 vccd1 vccd1 _4581_/X
+ sky130_fd_sc_hd__o221a_2
X_3532_ _6064_/Q _5439_/A2 _5743_/B _6077_/Q vssd1 vssd1 vccd1 vccd1 _3532_/X sky130_fd_sc_hd__o22a_1
XFILLER_116_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6251_ _6256_/CLK _6251_/D vssd1 vssd1 vccd1 vccd1 _6251_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3463_ _3926_/C _3462_/B _3621_/A vssd1 vssd1 vccd1 vccd1 _3463_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_103_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5202_ _6217_/Q _5202_/B vssd1 vssd1 vccd1 vccd1 _5203_/B sky130_fd_sc_hd__xnor2_1
X_6182_ _6290_/CLK _6182_/D vssd1 vssd1 vccd1 vccd1 _6182_/Q sky130_fd_sc_hd__dfxtp_1
X_3394_ _6014_/Q _6037_/Q _3709_/S vssd1 vssd1 vccd1 vccd1 _3394_/X sky130_fd_sc_hd__mux2_2
X_5133_ _5570_/A _5603_/S vssd1 vssd1 vccd1 vccd1 _5133_/X sky130_fd_sc_hd__or2_4
XFILLER_97_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_815 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5721__A _5733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5064_ _3019_/Y _5143_/B _5158_/B _5148_/A vssd1 vssd1 vccd1 vccd1 _5065_/B sky130_fd_sc_hd__a211o_1
XANTENNA__3808__A1 _4301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4015_ _3878_/A _4009_/B _4009_/X _4014_/X vssd1 vssd1 vccd1 vccd1 _4015_/X sky130_fd_sc_hd__a211o_1
XFILLER_72_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3241__A _3241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout179_A _3553_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4056__B _4058_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5966_ _5970_/A _5966_/B vssd1 vssd1 vccd1 vccd1 _5966_/X sky130_fd_sc_hd__or2_1
XANTENNA_fanout346_A input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4917_ _6191_/Q _4916_/C _6192_/Q vssd1 vssd1 vccd1 vccd1 _4918_/B sky130_fd_sc_hd__a21oi_1
X_5897_ _5898_/A _5898_/B vssd1 vssd1 vccd1 vccd1 _5897_/Y sky130_fd_sc_hd__nor2_1
XFILLER_138_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5408__S1 _3241_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4072__A _5936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4848_ _4809_/B _4811_/B _4807_/X vssd1 vssd1 vccd1 vccd1 _4849_/B sky130_fd_sc_hd__a21o_2
XFILLER_20_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4779_ _5358_/A _5367_/A vssd1 vssd1 vccd1 vccd1 _4860_/A sky130_fd_sc_hd__nand2_2
XFILLER_107_703 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5497__A0 _5504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5107__S _5129_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4247__A _5767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3151__A _3312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4681__S _5543_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5972__A1 _5110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5509__C _5509_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5724__A1 _3772_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3326__A _5924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5244__C _5463_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5660__B1 _3410_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3996__A _4850_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5820_ _5835_/A1 _4293_/X _5819_/Y _6273_/Q vssd1 vssd1 vccd1 vccd1 _5820_/X sky130_fd_sc_hd__a22o_1
XFILLER_34_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5751_ _5926_/A0 _5742_/Y _5749_/X _5750_/Y vssd1 vssd1 vccd1 vccd1 _6244_/D sky130_fd_sc_hd__a22o_1
XANTENNA__4604__B _4604_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4702_ _6186_/Q _6185_/Q _6184_/Q vssd1 vssd1 vccd1 vccd1 _4742_/B sky130_fd_sc_hd__and3_1
X_5682_ _5710_/S _4112_/C _5353_/A _5734_/A _3950_/C vssd1 vssd1 vccd1 vccd1 _5682_/X
+ sky130_fd_sc_hd__o221a_1
X_4633_ _5255_/B _4633_/B vssd1 vssd1 vccd1 vccd1 _4675_/A sky130_fd_sc_hd__or2_1
XANTENNA__5715__A1 _3974_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4564_ _5790_/A1 _4564_/A2 _4562_/X _4563_/X vssd1 vssd1 vccd1 vccd1 _6180_/D sky130_fd_sc_hd__a22o_1
XFILLER_118_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3515_ _3465_/A _3456_/X _3465_/B _3459_/B vssd1 vssd1 vccd1 vccd1 _3516_/B sky130_fd_sc_hd__o31a_2
X_4495_ _3942_/B _4501_/A2 _4493_/X _4494_/X vssd1 vssd1 vccd1 vccd1 _6138_/D sky130_fd_sc_hd__a22o_1
XFILLER_131_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3236__A _5924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6234_ _6234_/CLK _6234_/D vssd1 vssd1 vccd1 vccd1 _6234_/Q sky130_fd_sc_hd__dfxtp_1
X_3446_ _3203_/X _3801_/A _3437_/X _3445_/Y vssd1 vssd1 vccd1 vccd1 _3446_/X sky130_fd_sc_hd__o22a_1
XFILLER_103_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6165_ _6263_/CLK _6165_/D vssd1 vssd1 vccd1 vccd1 _6165_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3377_ _6012_/Q _3231_/Y _3376_/X vssd1 vssd1 vccd1 vccd1 _6012_/D sky130_fd_sc_hd__o21a_1
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5116_ _3033_/Y _5241_/A _5115_/Y vssd1 vssd1 vccd1 vccd1 _5985_/A sky130_fd_sc_hd__o21a_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6096_ _6098_/CLK _6096_/D vssd1 vssd1 vccd1 vccd1 _6096_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5047_ _4625_/A _5093_/A _5045_/X _5046_/X _5047_/C1 vssd1 vssd1 vccd1 vccd1 _6196_/D
+ sky130_fd_sc_hd__o311a_1
XANTENNA__4067__A _4067_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4454__A1 _3942_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_862 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5954__A1 _3941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5949_ _5949_/A _5949_/B vssd1 vssd1 vccd1 vccd1 _5949_/X sky130_fd_sc_hd__or2_1
XFILLER_40_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4530__A _4539_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5182__A2 _5617_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3146__A _3880_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3248__A2 _5439_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4445__A1 _5926_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4996__A2 _4872_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4705__A _4705_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5945__A1 _5264_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5239__C _5403_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5173__A2 _5075_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5255__B _5255_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3056__A _5239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3300_ _3564_/S _4665_/B _3294_/X vssd1 vssd1 vccd1 vccd1 _3300_/X sky130_fd_sc_hd__o21a_1
X_4280_ _4281_/B _4281_/A vssd1 vssd1 vccd1 vccd1 _4321_/A sky130_fd_sc_hd__and2b_1
XFILLER_4_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3231_ _5799_/A _3255_/A _3231_/C vssd1 vssd1 vccd1 vccd1 _3231_/Y sky130_fd_sc_hd__nand3_4
XFILLER_98_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4684__A1 _5051_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3162_ _3575_/B _3163_/B vssd1 vssd1 vccd1 vccd1 _3745_/B sky130_fd_sc_hd__nor2_1
XFILLER_67_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3093_ _5051_/B _5051_/C vssd1 vssd1 vccd1 vccd1 _3093_/Y sky130_fd_sc_hd__nor2_2
XFILLER_82_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5633__B1 _5097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4615__A _4615_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5803_ _6265_/Q _5801_/Y _5802_/X vssd1 vssd1 vccd1 vccd1 _6265_/D sky130_fd_sc_hd__a21o_1
XFILLER_62_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4334__B _4410_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4739__A2 _4806_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3995_ _5883_/A _5738_/A vssd1 vssd1 vccd1 vccd1 _3995_/Y sky130_fd_sc_hd__nand2_1
XFILLER_50_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5734_ _5734_/A _5734_/B vssd1 vssd1 vccd1 vccd1 _5734_/X sky130_fd_sc_hd__or2_1
XFILLER_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5665_ _4697_/B _4690_/B _5703_/A vssd1 vssd1 vccd1 vccd1 _5665_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3962__A3 _3996_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5446__A _5480_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4616_ _4604_/A _4615_/Y _5919_/A _4613_/X _5048_/C vssd1 vssd1 vccd1 vccd1 _4617_/C
+ sky130_fd_sc_hd__o2111a_1
X_5596_ _5595_/A _5594_/X _5251_/Y vssd1 vssd1 vccd1 vccd1 _5596_/X sky130_fd_sc_hd__a21o_1
XANTENNA_fanout309_A _6010_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5165__B _5165_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4547_ _6175_/Q _4562_/B vssd1 vssd1 vccd1 vccd1 _4547_/X sky130_fd_sc_hd__or2_1
XFILLER_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4478_ _6133_/Q _4490_/B vssd1 vssd1 vccd1 vccd1 _4478_/X sky130_fd_sc_hd__or2_1
XFILLER_132_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6217_ _6217_/CLK _6217_/D vssd1 vssd1 vccd1 vccd1 _6217_/Q sky130_fd_sc_hd__dfxtp_4
X_3429_ _6053_/Q _3589_/A2 _3589_/B1 _6046_/Q _5929_/B2 vssd1 vssd1 vccd1 vccd1 _3429_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__3478__A2 _3477_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5872__B1 _5638_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6148_ _6180_/CLK _6148_/D vssd1 vssd1 vccd1 vccd1 _6148_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6079_ _6079_/CLK _6079_/D vssd1 vssd1 vccd1 vccd1 _6079_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5624__B1 _3025_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4525__A _4540_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5927__A1 _5936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3402__A2 _3500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5075__B _5075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4902__A2 _5561_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4410__D _4410_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5615__A0 _4659_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4969__A2 _5871_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3626__C1 _3145_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5091__A1 _6198_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5379__C1 _5470_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5918__A1 _5870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3780_ _4663_/B _3816_/B _3779_/X vssd1 vssd1 vccd1 vccd1 _3780_/X sky130_fd_sc_hd__o21a_1
XFILLER_9_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_14_clk_A _6233_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5450_ _5599_/B _5450_/B vssd1 vssd1 vccd1 vccd1 _5451_/B sky130_fd_sc_hd__or2_1
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4401_ _4401_/A _4401_/B vssd1 vssd1 vccd1 vccd1 _4402_/B sky130_fd_sc_hd__and2_1
X_5381_ _5442_/A _5380_/Y _5376_/X vssd1 vssd1 vccd1 vccd1 _5381_/X sky130_fd_sc_hd__o21a_1
XANTENNA_clkbuf_leaf_29_clk_A clkbuf_3_5__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4332_ _6110_/Q _4296_/Y _4331_/X _4437_/A1 vssd1 vssd1 vccd1 vccd1 _4332_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_113_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout208 _3054_/Y vssd1 vssd1 vccd1 vccd1 _4022_/C sky130_fd_sc_hd__buf_6
XFILLER_114_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout219 _5742_/A vssd1 vssd1 vccd1 vccd1 _5767_/A sky130_fd_sc_hd__buf_8
XFILLER_87_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4263_ _4362_/A _4309_/B _4342_/B _4334_/A vssd1 vssd1 vccd1 vccd1 _4266_/A sky130_fd_sc_hd__a22oi_4
XFILLER_87_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6002_ _6148_/Q vssd1 vssd1 vccd1 vccd1 _6148_/D sky130_fd_sc_hd__clkbuf_2
X_3214_ _3948_/A _5512_/A vssd1 vssd1 vccd1 vccd1 _5464_/A sky130_fd_sc_hd__nand2_8
XFILLER_101_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4194_ _4214_/A _4173_/B _4178_/B _4176_/X vssd1 vssd1 vccd1 vccd1 _4225_/A sky130_fd_sc_hd__a31o_2
XANTENNA__3233__B _3706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3145_ _3880_/A _5883_/A _3145_/C vssd1 vssd1 vccd1 vccd1 _3867_/A sky130_fd_sc_hd__and3b_4
XANTENNA__4409__A1 _4410_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4409__B2 _4426_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3076_ _5218_/B _5244_/A vssd1 vssd1 vccd1 vccd1 _3076_/X sky130_fd_sc_hd__or2_2
XFILLER_54_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout259_A _3943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3978_ _4643_/A _3978_/B vssd1 vssd1 vccd1 vccd1 _5647_/C sky130_fd_sc_hd__or2_2
XFILLER_50_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5717_ _4202_/A _5649_/X _5716_/X _5799_/A vssd1 vssd1 vccd1 vccd1 _6239_/D sky130_fd_sc_hd__o211a_1
XFILLER_109_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5648_ _5052_/A _5648_/B _5648_/C _5648_/D vssd1 vssd1 vccd1 vccd1 _5649_/C sky130_fd_sc_hd__and4b_1
XFILLER_136_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5579_ _5598_/B _5579_/B vssd1 vssd1 vccd1 vccd1 _5595_/B sky130_fd_sc_hd__nand2_2
XFILLER_104_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3143__B _3881_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3320__B2 _3960_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5073__A1 _5244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4887__A1 _3740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5836__B1 _5638_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5300__A2 _5360_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3053__B _3869_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput8 io_in[7] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__buf_8
XFILLER_37_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5064__A1 _3019_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4950_ _4949_/X _4946_/Y _4944_/X _4948_/X vssd1 vssd1 vccd1 vccd1 _4950_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_64_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3901_ _5767_/A _3901_/B _5743_/C vssd1 vssd1 vccd1 vccd1 _4439_/S sky130_fd_sc_hd__or3_4
XANTENNA__3500__C _3500_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4881_ _4879_/Y _4880_/X _3029_/Y _4806_/S vssd1 vssd1 vccd1 vccd1 _4881_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_32_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3832_ _4202_/A _3832_/A2 _3536_/X _3765_/X _3772_/X vssd1 vssd1 vccd1 vccd1 _3832_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_32_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3763_ _3793_/B _3761_/Y _3762_/Y vssd1 vssd1 vccd1 vccd1 _4069_/A sky130_fd_sc_hd__a21o_2
X_5502_ _3060_/A _4961_/Y _5261_/Y _5513_/B _4644_/B vssd1 vssd1 vccd1 vccd1 _5503_/C
+ sky130_fd_sc_hd__a32o_1
X_3694_ _3942_/D _3693_/X _3705_/A vssd1 vssd1 vccd1 vccd1 _6022_/D sky130_fd_sc_hd__mux2_1
XANTENNA__3228__B _5617_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5433_ _5312_/B _5421_/Y _5417_/X _3122_/A vssd1 vssd1 vccd1 vccd1 _5433_/X sky130_fd_sc_hd__o211a_1
XFILLER_133_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5364_ _5367_/A _5476_/A vssd1 vssd1 vccd1 vccd1 _5364_/Y sky130_fd_sc_hd__nand2_1
XFILLER_126_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4315_ _4315_/A _4315_/B vssd1 vssd1 vccd1 vccd1 _4318_/A sky130_fd_sc_hd__xor2_4
X_5295_ _5296_/A _5296_/B vssd1 vssd1 vccd1 vccd1 _5295_/Y sky130_fd_sc_hd__nand2_4
XFILLER_87_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5162__C _5258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4246_ _6093_/Q _3730_/X _4246_/S vssd1 vssd1 vccd1 vccd1 _6093_/D sky130_fd_sc_hd__mux2_1
XFILLER_113_196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4177_ _4177_/A _4177_/B vssd1 vssd1 vccd1 vccd1 _4178_/B sky130_fd_sc_hd__xnor2_4
XFILLER_110_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3128_ _4633_/B _4974_/A _3135_/S vssd1 vssd1 vccd1 vccd1 _6003_/D sky130_fd_sc_hd__mux2_1
XANTENNA__5055__A1 _5072_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4075__A _4197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3059_ _4646_/A _5227_/A vssd1 vssd1 vccd1 vccd1 _3059_/Y sky130_fd_sc_hd__nor2_8
XFILLER_35_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4803__A _5392_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3138__B _3257_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3154__A _3922_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4097__A2 _4111_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5597__A2 _5250_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5349__A2 _4234_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4021__A2 _3975_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3780__A1 _4663_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5263__B _5263_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4100_ _4083_/Y _4087_/A _4099_/X vssd1 vssd1 vccd1 vccd1 _4123_/A sky130_fd_sc_hd__o21ai_4
XFILLER_69_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5080_ _5080_/A _5080_/B _5878_/A vssd1 vssd1 vccd1 vccd1 _5080_/X sky130_fd_sc_hd__or3b_1
XANTENNA__5285__A1 _5512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4031_ _4027_/X _4030_/X _3984_/X vssd1 vssd1 vccd1 vccd1 _4031_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_111_689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5037__A1 _6196_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5588__A2 _5454_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5982_ _5982_/A _5985_/B _5985_/C vssd1 vssd1 vccd1 vccd1 _5982_/X sky130_fd_sc_hd__or3_1
XFILLER_80_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4933_ _4934_/B _4934_/A vssd1 vssd1 vccd1 vccd1 _4987_/A sky130_fd_sc_hd__nand2b_1
XFILLER_33_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4864_ _5330_/B _4864_/B vssd1 vssd1 vccd1 vccd1 _4864_/Y sky130_fd_sc_hd__nand2_1
XFILLER_60_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3815_ _4772_/B _3740_/X _3749_/X _3814_/X vssd1 vssd1 vccd1 vccd1 _3815_/X sky130_fd_sc_hd__a211o_1
XANTENNA__4342__B _4342_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4795_ _3122_/Y _4793_/Y _4794_/X _4788_/X vssd1 vssd1 vccd1 vccd1 _4795_/X sky130_fd_sc_hd__a31o_1
XANTENNA__4012__A2 _5848_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3746_ _3746_/A vssd1 vssd1 vccd1 vccd1 _3812_/S sky130_fd_sc_hd__inv_2
XANTENNA_fanout124_A _4604_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3677_ _3881_/B _3677_/B vssd1 vssd1 vccd1 vccd1 _3678_/C sky130_fd_sc_hd__nand2b_2
XFILLER_118_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5454__A _5454_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5416_ _5446_/B _5446_/C vssd1 vssd1 vccd1 vccd1 _5416_/X sky130_fd_sc_hd__or2_1
XFILLER_106_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5347_ _5347_/A _5347_/B _5338_/Y vssd1 vssd1 vccd1 vccd1 _5347_/X sky130_fd_sc_hd__or3b_2
XANTENNA__3523__B2 _3312_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5278_ _6174_/Q _4234_/B _4058_/B _6134_/Q vssd1 vssd1 vccd1 vccd1 _5278_/X sky130_fd_sc_hd__o22a_1
XANTENNA__5276__A1 _5227_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4229_ _4229_/A _4229_/B vssd1 vssd1 vccd1 vccd1 _4231_/B sky130_fd_sc_hd__nand2_1
XFILLER_101_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3826__A2 _3777_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5028__A1 _4745_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5028__B2 _4744_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5200__A1 _5218_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3149__A _3948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3246__A_N _3236_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4679__S _5041_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5364__A _5367_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4711__B1 _4701_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5303__S _5360_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5019__B2 _4753_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4778__B1 _4753_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output18_A _6192_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5258__B _5507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4162__B _4162_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3059__A _4646_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3600_ _3595_/Y _3596_/X _3599_/X vssd1 vssd1 vccd1 vccd1 _5721_/B sky130_fd_sc_hd__o21ba_2
XFILLER_128_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4580_ _5239_/B _5238_/C _4580_/C vssd1 vssd1 vccd1 vccd1 _4580_/X sky130_fd_sc_hd__or3_1
X_3531_ _6015_/Q _3231_/Y _3530_/X vssd1 vssd1 vccd1 vccd1 _6015_/D sky130_fd_sc_hd__o21a_1
XFILLER_116_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6250_ _6250_/CLK _6250_/D vssd1 vssd1 vccd1 vccd1 _6250_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3462_ _3926_/C _3462_/B vssd1 vssd1 vccd1 vccd1 _3462_/X sky130_fd_sc_hd__or2_1
X_5201_ _5191_/A _6216_/Q _5199_/X _5200_/X _5071_/A vssd1 vssd1 vccd1 vccd1 _6216_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_131_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6181_ _6214_/CLK _6181_/D vssd1 vssd1 vccd1 vccd1 _6181_/Q sky130_fd_sc_hd__dfxtp_1
X_3393_ _6276_/Q _6112_/Q _3551_/S vssd1 vssd1 vccd1 vccd1 _5341_/B sky130_fd_sc_hd__mux2_4
XFILLER_124_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5132_ _5221_/B _5132_/B vssd1 vssd1 vccd1 vccd1 _5603_/S sky130_fd_sc_hd__or2_4
XFILLER_69_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5063_ _5063_/A _5250_/A _5063_/C vssd1 vssd1 vccd1 vccd1 _5070_/S sky130_fd_sc_hd__and3_2
XFILLER_96_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5213__S _5561_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4014_ _3029_/Y _3986_/B _4008_/Y _4011_/X _4013_/X vssd1 vssd1 vccd1 vccd1 _4014_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_65_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3241__B _3241_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4056__C _5767_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5965_ _4767_/A _5934_/A _4023_/A _5120_/Y vssd1 vssd1 vccd1 vccd1 _5966_/B sky130_fd_sc_hd__o31a_1
XFILLER_40_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5449__A _5599_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4916_ _6192_/Q _6191_/Q _4916_/C vssd1 vssd1 vccd1 vccd1 _4952_/B sky130_fd_sc_hd__and3_1
XANTENNA_fanout241_A _5128_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5896_ _5887_/Y _5895_/X _5888_/Y vssd1 vssd1 vccd1 vccd1 _5896_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout339_A input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4847_ _4847_/A _4847_/B vssd1 vssd1 vccd1 vccd1 _4849_/A sky130_fd_sc_hd__nand2_1
X_4778_ _4705_/A _4777_/Y _4753_/A vssd1 vssd1 vccd1 vccd1 _4778_/X sky130_fd_sc_hd__o21a_1
XFILLER_5_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3729_ _4167_/D _3684_/X _3708_/Y _6233_/Q vssd1 vssd1 vccd1 vccd1 _3729_/X sky130_fd_sc_hd__o22a_1
XFILLER_107_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4528__A _4539_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5123__S _5129_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3432__A _3432_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4247__B _5436_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3680__B1 _4462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3578__S _3658_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5793__S _5798_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5185__B1 _5158_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4160__A1 _4202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3996__B _3996_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3488__S _3709_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5750_ _5305_/A _5763_/B _5742_/Y vssd1 vssd1 vccd1 vccd1 _5750_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__4173__A _4214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4604__C _4604_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4701_ _4972_/A _4694_/X _4700_/X _3740_/A vssd1 vssd1 vccd1 vccd1 _4701_/X sky130_fd_sc_hd__a22o_4
X_5681_ _6302_/Q _4615_/A _5680_/X vssd1 vssd1 vccd1 vccd1 _5681_/X sky130_fd_sc_hd__a21o_1
X_4632_ _5255_/B _4633_/B vssd1 vssd1 vccd1 vccd1 _4678_/A sky130_fd_sc_hd__nand2_2
XANTENNA__5176__B1 _5071_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3726__A1 _3488_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4563_ _4891_/A _4252_/A _4239_/B vssd1 vssd1 vccd1 vccd1 _4563_/X sky130_fd_sc_hd__o21a_1
XANTENNA__3726__B2 _6232_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6302_ _6302_/CLK _6302_/D vssd1 vssd1 vccd1 vccd1 _6302_/Q sky130_fd_sc_hd__dfxtp_2
X_3514_ _3571_/B _3514_/B vssd1 vssd1 vccd1 vccd1 _3935_/C sky130_fd_sc_hd__nor2_4
X_4494_ _5385_/A _4239_/A _4059_/B vssd1 vssd1 vccd1 vccd1 _4494_/X sky130_fd_sc_hd__o21a_1
X_6233_ _6233_/CLK _6233_/D vssd1 vssd1 vccd1 vccd1 _6233_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_104_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3445_ _3398_/A _5707_/B _3498_/S vssd1 vssd1 vccd1 vccd1 _3445_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_116_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6164_ _6279_/CLK _6164_/D vssd1 vssd1 vccd1 vccd1 _6164_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3376_ _3631_/A _3375_/X _3332_/X _3592_/A vssd1 vssd1 vccd1 vccd1 _3376_/X sky130_fd_sc_hd__a211o_1
XFILLER_97_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5115_ _6237_/Q _5158_/A vssd1 vssd1 vccd1 vccd1 _5115_/Y sky130_fd_sc_hd__nand2_1
XFILLER_97_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout191_A _3241_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6095_ _6098_/CLK _6095_/D vssd1 vssd1 vccd1 vccd1 _6095_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3252__A _3960_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5046_ _6196_/Q _5046_/B vssd1 vssd1 vccd1 vccd1 _5046_/X sky130_fd_sc_hd__or2_1
XFILLER_57_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5100__B1 _5097_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4067__B _4294_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4454__A2 _3900_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5651__A1 _5733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4191__A1_N _3842_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3662__B1 _3422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5948_ _5948_/A _5948_/B vssd1 vssd1 vccd1 vccd1 _6295_/D sky130_fd_sc_hd__and2_1
XFILLER_43_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5879_ _4819_/B _5911_/C _3972_/Y _5878_/X vssd1 vssd1 vccd1 vccd1 _5879_/X sky130_fd_sc_hd__o31a_1
XFILLER_138_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3717__A1 _4111_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3717__B2 _5540_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5118__S _5129_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4390__A1 _4426_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3146__B _5065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4142__A1 _4270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3162__A _3575_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4445__A2 _3900_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5945__A2 _5108_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3956__A1 _5090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4440__B _4458_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3056__B _3312_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3230_ _4539_/A _3255_/A _3231_/C vssd1 vssd1 vccd1 vccd1 _3592_/A sky130_fd_sc_hd__and3_4
XFILLER_113_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3161_ _4642_/A _3163_/B vssd1 vssd1 vccd1 vccd1 _5903_/A sky130_fd_sc_hd__or2_2
XFILLER_67_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3092_ _5179_/A _3092_/B _3111_/B vssd1 vssd1 vccd1 vccd1 _5051_/C sky130_fd_sc_hd__or3_4
XFILLER_54_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5094__C1 _5071_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5397__A0 _5385_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5802_ _4136_/A _5817_/A1 _4173_/B _5801_/B _3322_/X vssd1 vssd1 vccd1 vccd1 _5802_/X
+ sky130_fd_sc_hd__a32o_1
X_3994_ _5207_/S _3996_/B vssd1 vssd1 vccd1 vccd1 _5738_/A sky130_fd_sc_hd__nand2_1
X_5733_ _5733_/A _5733_/B vssd1 vssd1 vccd1 vccd1 _5740_/B sky130_fd_sc_hd__nor2_1
XFILLER_30_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5664_ _4096_/A _5649_/X _5663_/X _5956_/A vssd1 vssd1 vccd1 vccd1 _6235_/D sky130_fd_sc_hd__o211a_1
XFILLER_108_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5446__B _5446_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4615_ _4615_/A _4615_/B _5634_/C vssd1 vssd1 vccd1 vccd1 _4615_/Y sky130_fd_sc_hd__nor3_1
X_5595_ _5595_/A _5595_/B vssd1 vssd1 vccd1 vccd1 _5595_/Y sky130_fd_sc_hd__nor2_1
XFILLER_117_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4546_ _5935_/A0 _4564_/A2 _4544_/X _4545_/X vssd1 vssd1 vccd1 vccd1 _6174_/D sky130_fd_sc_hd__a22o_1
XANTENNA__5165__C _5634_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4477_ _5790_/A1 _4476_/X _4477_/S vssd1 vssd1 vccd1 vccd1 _6132_/D sky130_fd_sc_hd__mux2_1
XFILLER_104_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3428_ _6097_/Q _3589_/A2 _5743_/B _6075_/Q _3427_/X vssd1 vssd1 vccd1 vccd1 _3428_/X
+ sky130_fd_sc_hd__o221a_2
X_6216_ _6217_/CLK _6216_/D vssd1 vssd1 vccd1 vccd1 _6216_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__5872__A1 _4577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input9_A rst vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6147_ _6180_/CLK _6147_/D vssd1 vssd1 vccd1 vccd1 _6147_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3359_ _3316_/A _3316_/B _3303_/X _5889_/A vssd1 vssd1 vccd1 vccd1 _3361_/B sky130_fd_sc_hd__o2bb2a_2
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6078_ _6093_/CLK _6078_/D vssd1 vssd1 vccd1 vccd1 _6078_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5624__A1 _5048_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5029_ _5567_/A _5029_/B vssd1 vssd1 vccd1 vccd1 _5040_/A sky130_fd_sc_hd__xor2_4
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5388__B1 _5387_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5927__A2 _5943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3157__A _5883_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5075__C _5075_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5457__A1_N _4644_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5863__A1 _3607_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_635 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5615__A1 _4665_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4716__A _5330_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4823__C1 _4753_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5091__A2 _5870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5379__B1 _4058_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5918__A2 _3883_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5547__A _5547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4400_ _4401_/A _4401_/B vssd1 vssd1 vccd1 vccd1 _4419_/A sky130_fd_sc_hd__nor2_1
X_5380_ _5929_/B2 _5377_/X _5378_/X _5379_/X vssd1 vssd1 vccd1 vccd1 _5380_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_132_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4331_ _4358_/B _4331_/B vssd1 vssd1 vccd1 vccd1 _4331_/X sky130_fd_sc_hd__and2_1
XFILLER_125_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5303__A0 _4707_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4106__A1 _4162_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4262_ _4325_/A _4262_/B vssd1 vssd1 vccd1 vccd1 _4283_/A sky130_fd_sc_hd__nor2_1
Xfanout209 _3053_/X vssd1 vssd1 vccd1 vccd1 _3885_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_113_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6001_ _6147_/Q vssd1 vssd1 vccd1 vccd1 _6147_/D sky130_fd_sc_hd__clkbuf_2
X_3213_ _4638_/A _5570_/A vssd1 vssd1 vccd1 vccd1 _4596_/D sky130_fd_sc_hd__nor2_4
XFILLER_113_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4193_ _4193_/A _4193_/B vssd1 vssd1 vccd1 vccd1 _4231_/A sky130_fd_sc_hd__nor2_1
XFILLER_79_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3233__C _5734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3144_ _3974_/B _3365_/B vssd1 vssd1 vccd1 vccd1 _3960_/B sky130_fd_sc_hd__nand2_8
XFILLER_94_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4409__A2 _4426_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5606__A1 _5227_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3075_ _5218_/B _5244_/A vssd1 vssd1 vccd1 vccd1 _3123_/A sky130_fd_sc_hd__nor2_8
XFILLER_36_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout154_A _3069_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3977_ _5191_/A _4596_/B vssd1 vssd1 vccd1 vccd1 _4577_/D sky130_fd_sc_hd__nand2_1
XANTENNA_fanout321_A _3028_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5716_ _3593_/A _3958_/Y _5705_/X _5715_/X vssd1 vssd1 vccd1 vccd1 _5716_/X sky130_fd_sc_hd__a211o_2
X_5647_ _3127_/A _5647_/B _5647_/C _5647_/D vssd1 vssd1 vccd1 vccd1 _5648_/D sky130_fd_sc_hd__and4b_1
X_5578_ _6232_/Q _5578_/B vssd1 vssd1 vccd1 vccd1 _5579_/B sky130_fd_sc_hd__or2_1
XFILLER_117_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4529_ _4540_/A _6165_/Q vssd1 vssd1 vccd1 vccd1 _6164_/D sky130_fd_sc_hd__or2_1
XFILLER_2_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3705__A _3705_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5192__A _5192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout67_A _5513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5073__A2 _4638_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5367__A _5367_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4702__C _6184_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5533__B1 _5251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5836__A1 _5165_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput9 rst vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__buf_8
XFILLER_76_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5041__S _5041_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5064__A2 _5143_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3900_ _5767_/A _3901_/B _5743_/C vssd1 vssd1 vccd1 vccd1 _3900_/Y sky130_fd_sc_hd__nor3_4
XFILLER_45_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3500__D _3513_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4880_ _4879_/A _4879_/B _4806_/S vssd1 vssd1 vccd1 vccd1 _4880_/X sky130_fd_sc_hd__o21a_1
X_3831_ _3855_/S _3831_/B vssd1 vssd1 vccd1 vccd1 _3831_/Y sky130_fd_sc_hd__nor2_1
XFILLER_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5979__A1_N _4846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5277__A _5436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3762_ _5889_/B _3841_/S vssd1 vssd1 vccd1 vccd1 _3762_/Y sky130_fd_sc_hd__nor2_1
X_5501_ _5540_/C _5501_/B vssd1 vssd1 vccd1 vccd1 _5513_/B sky130_fd_sc_hd__or2_4
XFILLER_9_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3693_ _5333_/A _6022_/Q _3902_/A vssd1 vssd1 vccd1 vccd1 _3693_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5524__B1 _3060_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5432_ _5424_/Y _5431_/X _5936_/A vssd1 vssd1 vccd1 vccd1 _5432_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_105_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5363_ _5498_/A _5359_/X _5362_/X vssd1 vssd1 vccd1 vccd1 _5363_/X sky130_fd_sc_hd__o21a_1
XFILLER_99_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4314_ _4315_/A _4315_/B vssd1 vssd1 vccd1 vccd1 _4347_/B sky130_fd_sc_hd__nor2_1
XANTENNA__3550__A2 _5706_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5294_ _5326_/B _5293_/Y _5291_/Y vssd1 vssd1 vccd1 vccd1 _5294_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5827__A1 _3477_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4245_ _6092_/Q _3727_/X _4246_/S vssd1 vssd1 vccd1 vccd1 _6092_/D sky130_fd_sc_hd__mux2_1
XFILLER_99_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_17 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4176_ _4202_/A _4176_/B _4177_/A vssd1 vssd1 vccd1 vccd1 _4176_/X sky130_fd_sc_hd__and3_1
X_3127_ _3127_/A _4462_/A _3127_/C _3104_/X vssd1 vssd1 vccd1 vccd1 _3135_/S sky130_fd_sc_hd__or4b_4
XFILLER_110_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout271_A _5540_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5055__A2 _5870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3058_ _5218_/B _3058_/B vssd1 vssd1 vccd1 vccd1 _3058_/Y sky130_fd_sc_hd__nand2_2
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4075__B _4173_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4263__B1 _4342_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4803__B _5703_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5212__C1 _3060_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5634__B _5634_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5126__S _5128_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3435__A _3450_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5796__S _5798_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_28_clk_A _6084_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_53_clk _6133_/CLK vssd1 vssd1 vccd1 vccd1 _6179_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4006__B1 _5714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5097__A _5097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4557__A1 _5385_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3532__A2 _5439_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5809__A1 _5835_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4030_ _5934_/A _4029_/X _4028_/X _5883_/A vssd1 vssd1 vccd1 vccd1 _4030_/X sky130_fd_sc_hd__a211o_1
XFILLER_111_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4176__A _4202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5037__A2 _4647_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5981_ _5119_/Y _5985_/C _6301_/Q vssd1 vssd1 vccd1 vccd1 _5981_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__5588__A3 _5072_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4932_ _4828_/B _4926_/A _4924_/X vssd1 vssd1 vccd1 vccd1 _4934_/B sky130_fd_sc_hd__o21ba_1
XFILLER_52_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4796__A1 _5358_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_44_clk clkbuf_3_4__f_clk/X vssd1 vssd1 vccd1 vccd1 _6295_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_45_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4796__B2 _4643_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4863_ _5034_/A _4862_/X _4856_/Y _4852_/X vssd1 vssd1 vccd1 vccd1 _4863_/X sky130_fd_sc_hd__a211o_1
XFILLER_20_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5745__A0 _3943_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4548__A1 _5305_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3814_ _4163_/A _3777_/S _3813_/X _3751_/A vssd1 vssd1 vccd1 vccd1 _3814_/X sky130_fd_sc_hd__o211a_1
X_4794_ _6188_/Q _5041_/S vssd1 vssd1 vccd1 vccd1 _4794_/X sky130_fd_sc_hd__or2_1
XANTENNA__3239__B _3241_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3745_ _5503_/A _3745_/B _3745_/C vssd1 vssd1 vccd1 vccd1 _3746_/A sky130_fd_sc_hd__and3_4
XFILLER_118_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3676_ _3948_/A _5075_/C vssd1 vssd1 vccd1 vccd1 _3678_/B sky130_fd_sc_hd__nand2_2
XFILLER_106_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5454__B _5454_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5415_ _5446_/B _5446_/C vssd1 vssd1 vccd1 vccd1 _5415_/Y sky130_fd_sc_hd__nand2_1
XFILLER_133_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4720__A1 _5051_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5346_ _5507_/A _5227_/B _5354_/B _5345_/X vssd1 vssd1 vccd1 vccd1 _5347_/A sky130_fd_sc_hd__a31o_1
XFILLER_88_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5277_ _5436_/A _6150_/Q _5436_/C vssd1 vssd1 vccd1 vccd1 _5277_/X sky130_fd_sc_hd__and3_1
XFILLER_88_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4228_ _4224_/Y _4225_/X _4185_/B _4185_/Y vssd1 vssd1 vccd1 vccd1 _4229_/B sky130_fd_sc_hd__o211ai_2
XFILLER_68_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4159_ _4233_/A1 _4157_/X _4158_/X vssd1 vssd1 vccd1 vccd1 _6084_/D sky130_fd_sc_hd__a21o_1
XFILLER_46_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5433__C1 _3122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4814__A _6189_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5984__B1 _6302_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_35_clk clkbuf_3_5__f_clk/X vssd1 vssd1 vccd1 vccd1 _6264_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_62_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3149__B _5936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5364__B _5476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3165__A _5840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4711__A1 _5034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4711__B2 _3116_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4475__A0 _3942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5672__C1 _3996_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4778__A1 _4705_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4724__A _5114_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5975__B1 _3960_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_26_clk _6084_/CLK vssd1 vssd1 vccd1 vccd1 _6278_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4443__B _4458_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5727__B1 _3615_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4162__C _4309_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3059__B _5227_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3530_ _3631_/A _3529_/X _3485_/X _3592_/A vssd1 vssd1 vccd1 vccd1 _3530_/X sky130_fd_sc_hd__a211o_1
XFILLER_128_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3461_ _3412_/Y _3414_/B _3926_/B _3926_/A vssd1 vssd1 vccd1 vccd1 _3462_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_115_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3075__A _5218_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5200_ _5218_/B _5050_/C _4596_/D _5052_/B _5097_/A vssd1 vssd1 vccd1 vccd1 _5200_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3505__A2 _3513_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6180_ _6180_/CLK _6180_/D vssd1 vssd1 vccd1 vccd1 _6180_/Q sky130_fd_sc_hd__dfxtp_1
X_3392_ _4697_/A _3636_/A _3211_/Y _3391_/Y vssd1 vssd1 vccd1 vccd1 _3392_/X sky130_fd_sc_hd__a211o_1
XFILLER_97_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5131_ _5131_/A _5131_/B vssd1 vssd1 vccd1 vccd1 _5131_/Y sky130_fd_sc_hd__nand2_1
XFILLER_97_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5290__A _5512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5062_ _5062_/A _5062_/B _5062_/C _5249_/D vssd1 vssd1 vccd1 vccd1 _5063_/C sky130_fd_sc_hd__and4_1
XFILLER_97_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4466__A0 _6221_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_3_6__f_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4013_ _5108_/A _3274_/X _3615_/B _4850_/A _4012_/X vssd1 vssd1 vccd1 vccd1 _4013_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_38_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5964_ _5119_/Y _5970_/A _3766_/A vssd1 vssd1 vccd1 vccd1 _5964_/Y sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_17_clk _6084_/CLK vssd1 vssd1 vccd1 vccd1 _6241_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__5449__B _5450_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4915_ _5731_/S _4910_/Y _4914_/Y _3101_/A vssd1 vssd1 vccd1 vccd1 _4915_/X sky130_fd_sc_hd__o22a_1
XANTENNA__3441__A1 _6015_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5895_ _3571_/A _3937_/D _5893_/X _5894_/X vssd1 vssd1 vccd1 vccd1 _5895_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_33_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4846_ _4846_/A _4846_/B vssd1 vssd1 vccd1 vccd1 _4847_/B sky130_fd_sc_hd__or2_2
XANTENNA_fanout234_A _6290_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4072__C _4072_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4777_ _6188_/Q _4814_/C vssd1 vssd1 vccd1 vccd1 _4777_/Y sky130_fd_sc_hd__xnor2_1
X_3728_ _6032_/Q _3727_/X _3731_/S vssd1 vssd1 vccd1 vccd1 _6032_/D sky130_fd_sc_hd__mux2_1
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3659_ _3313_/Y _3657_/Y _3658_/X _4003_/C _3365_/Y vssd1 vssd1 vccd1 vccd1 _3659_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_134_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5329_ _5329_/A vssd1 vssd1 vccd1 vccd1 _5329_/Y sky130_fd_sc_hd__inv_2
XFILLER_102_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5709__A0 _5409_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5185__A1 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3607__B _3607_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3326__C _5436_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3499__A1 _4163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4160__A2 _4173_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5660__A2 _3388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4173__B _4173_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3423__A1 _3511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4700_ _4697_/A _4699_/Y _4812_/S vssd1 vssd1 vccd1 vccd1 _4700_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4604__D _5928_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5680_ _6298_/Q _5692_/B _3772_/B vssd1 vssd1 vccd1 vccd1 _5680_/X sky130_fd_sc_hd__a21o_1
XFILLER_30_441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4631_ _4626_/Y _4627_/X _4630_/Y vssd1 vssd1 vccd1 vccd1 _4631_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__5176__A1 _5191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4562_ _6180_/Q _4562_/B vssd1 vssd1 vccd1 vccd1 _4562_/X sky130_fd_sc_hd__or2_1
X_6301_ _6301_/CLK _6301_/D vssd1 vssd1 vccd1 vccd1 _6301_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_116_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3513_ _6205_/Q _3513_/B vssd1 vssd1 vccd1 vccd1 _3514_/B sky130_fd_sc_hd__nor2_1
X_4493_ _6138_/Q _4499_/B vssd1 vssd1 vccd1 vccd1 _4493_/X sky130_fd_sc_hd__or2_1
XFILLER_131_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6232_ _6232_/CLK _6232_/D vssd1 vssd1 vccd1 vccd1 _6232_/Q sky130_fd_sc_hd__dfxtp_4
X_3444_ _3444_/A _3444_/B vssd1 vssd1 vccd1 vccd1 _3513_/B sky130_fd_sc_hd__or2_4
Xclkbuf_leaf_6_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _6217_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_69_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6163_ _6279_/CLK _6163_/D vssd1 vssd1 vccd1 vccd1 _6163_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3375_ _3583_/S _5653_/B _3355_/Y vssd1 vssd1 vccd1 vccd1 _3375_/X sky130_fd_sc_hd__a21bo_4
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5532__A2_N _5522_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5114_ _5114_/A _5957_/B vssd1 vssd1 vccd1 vccd1 _5114_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__4439__A0 _3943_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6094_ _6260_/CLK _6094_/D vssd1 vssd1 vccd1 vccd1 _6094_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5100__A1 _6009_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5045_ _5567_/A _4872_/B _5044_/X _4931_/B vssd1 vssd1 vccd1 vccd1 _5045_/X sky130_fd_sc_hd__o22a_1
XANTENNA_fanout184_A _4112_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5947_ _6295_/Q _5946_/X _5947_/S vssd1 vssd1 vccd1 vccd1 _5948_/B sky130_fd_sc_hd__mux2_1
XFILLER_34_780 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5878_ _5878_/A _5951_/B _5878_/C _5878_/D vssd1 vssd1 vccd1 vccd1 _5878_/X sky130_fd_sc_hd__and4_1
XANTENNA__5167__A1 _3112_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4829_ _4925_/A _4829_/B vssd1 vssd1 vccd1 vccd1 _4829_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_138_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3708__A _3732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3717__A2 _5743_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4390__A2 _4389_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3146__C _3960_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5875__C1 _5911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4142__A2 _4111_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4539__A _4539_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4602__B1 _5097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5945__A3 _5934_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3056__C _4022_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3160_ _3880_/A _3163_/B vssd1 vssd1 vccd1 vccd1 _3867_/B sky130_fd_sc_hd__nor2_4
XFILLER_94_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3091_ _6217_/Q _3170_/B vssd1 vssd1 vccd1 vccd1 _3091_/Y sky130_fd_sc_hd__nand2_1
XFILLER_66_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4584__B1_N _6183_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5633__A2 _5065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5801_ _5819_/A _5801_/B vssd1 vssd1 vccd1 vccd1 _5801_/Y sky130_fd_sc_hd__nor2_4
XFILLER_62_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3993_ _3993_/A _3993_/B vssd1 vssd1 vccd1 vccd1 _3999_/C sky130_fd_sc_hd__nand2_1
X_5732_ _5718_/A _5731_/X _5730_/X _5732_/C1 vssd1 vssd1 vccd1 vccd1 _5740_/A sky130_fd_sc_hd__o211a_1
XANTENNA__4912__A _5617_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5663_ _5075_/A _4619_/A _5655_/X _5662_/X vssd1 vssd1 vccd1 vccd1 _5663_/X sky130_fd_sc_hd__a211o_1
XANTENNA__5149__B2 _3958_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4614_ _4614_/A _4614_/B vssd1 vssd1 vccd1 vccd1 _5919_/A sky130_fd_sc_hd__or2_4
XFILLER_129_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5594_ _5588_/X _5591_/X _5593_/X _5581_/X vssd1 vssd1 vccd1 vccd1 _5594_/X sky130_fd_sc_hd__a31o_1
XFILLER_117_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4545_ _4672_/A _4252_/A _4239_/B vssd1 vssd1 vccd1 vccd1 _4545_/X sky130_fd_sc_hd__o21a_1
XANTENNA__5743__A _5767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4476_ _4891_/A _6132_/Q _4476_/S vssd1 vssd1 vccd1 vccd1 _4476_/X sky130_fd_sc_hd__mux2_1
XFILLER_116_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5471__A2_N _5734_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5857__C1 _5867_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6215_ _6217_/CLK _6215_/D vssd1 vssd1 vccd1 vccd1 _6215_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_104_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5321__A1 _5929_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3427_ _6062_/Q _5439_/A2 _3589_/B1 _6090_/Q vssd1 vssd1 vccd1 vccd1 _3427_/X sky130_fd_sc_hd__o22a_1
XANTENNA__3263__A _5800_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5872__A2 _4577_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6146_ _6180_/CLK _6146_/D vssd1 vssd1 vccd1 vccd1 _6146_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3358_ _3358_/A _3358_/B vssd1 vssd1 vccd1 vccd1 _3935_/B sky130_fd_sc_hd__nor2_8
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6077_ _6264_/CLK _6077_/D vssd1 vssd1 vccd1 vccd1 _6077_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3289_ _4136_/A _3210_/B _3210_/C _3288_/X vssd1 vssd1 vccd1 vccd1 _3289_/X sky130_fd_sc_hd__o211a_1
XFILLER_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5028_ _4745_/A _5023_/X _5026_/Y _5036_/B _4744_/B vssd1 vssd1 vccd1 vccd1 _5028_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_57_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4832__B1 _5058_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4094__A _4162_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3399__B1 _3500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4060__A1 _3711_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5129__S _5129_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3157__B _4622_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5653__A _5653_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4269__A _4270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3173__A _3741_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3901__A _5767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5076__B1 _5238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3626__B2 _3312_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4732__A _5114_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4051__A1 _3869_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5547__B _5547_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3348__A _3388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4330_ _4330_/A _4330_/B _4330_/C vssd1 vssd1 vccd1 vccd1 _4331_/B sky130_fd_sc_hd__nand3_1
XFILLER_114_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4106__A2 _4176_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4261_ _4216_/A _4214_/B _4205_/B _4206_/X vssd1 vssd1 vccd1 vccd1 _4262_/B sky130_fd_sc_hd__a211oi_1
XFILLER_113_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3083__A _5075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6000_ _6146_/Q vssd1 vssd1 vccd1 vccd1 _6146_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_113_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3314__B1 _3312_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3212_ _3212_/A _3738_/A vssd1 vssd1 vccd1 vccd1 _3398_/A sky130_fd_sc_hd__or2_4
X_4192_ _4233_/A1 _4190_/Y _4191_/X vssd1 vssd1 vccd1 vccd1 _6085_/D sky130_fd_sc_hd__a21o_1
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3143_ _4003_/B _3881_/A vssd1 vssd1 vccd1 vccd1 _3145_/C sky130_fd_sc_hd__nor2_8
XFILLER_121_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3074_ _3060_/B _5244_/B _5169_/C _3060_/Y _3062_/Y vssd1 vssd1 vccd1 vccd1 _3085_/A
+ sky130_fd_sc_hd__o32a_1
XFILLER_95_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4642__A _4642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout147_A _5605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3976_ _5097_/A _5096_/C vssd1 vssd1 vccd1 vccd1 _3979_/B sky130_fd_sc_hd__nor2_2
X_5715_ _3974_/C _5713_/X _5714_/Y _5728_/A _5706_/Y vssd1 vssd1 vccd1 vccd1 _5715_/X
+ sky130_fd_sc_hd__a311o_1
XANTENNA__5790__A1 _5790_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3258__A _3766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout314_A _5556_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5646_ _4577_/A _5128_/S _4614_/B _3955_/X vssd1 vssd1 vccd1 vccd1 _5648_/C sky130_fd_sc_hd__o31a_1
XANTENNA__3692__S _3705_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5577_ _6232_/Q _5578_/B vssd1 vssd1 vccd1 vccd1 _5598_/B sky130_fd_sc_hd__nand2_4
XFILLER_117_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4528_ _4539_/A _6164_/Q vssd1 vssd1 vccd1 vccd1 _6163_/D sky130_fd_sc_hd__and2_1
XFILLER_2_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4459_ _4891_/A _4438_/S _4439_/S vssd1 vssd1 vccd1 vccd1 _4459_/X sky130_fd_sc_hd__o21a_1
XFILLER_49_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6129_ _6154_/CLK _6129_/D vssd1 vssd1 vccd1 vccd1 _6129_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5073__A3 _4644_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5230__B1 _4644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5367__B _5367_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5781__A1 _5856_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3168__A _4648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_775 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5533__A1 _5595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3615__B _3615_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5836__A2 _3974_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3847__A1 _3987_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_723 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4446__B _4458_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3777__S _3777_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4462__A _4462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3830_ _3841_/S _3828_/Y _3829_/Y vssd1 vssd1 vccd1 vccd1 _3831_/B sky130_fd_sc_hd__a21o_2
XFILLER_20_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5772__A1 _5935_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3761_ _4665_/B _3816_/B _3760_/X vssd1 vssd1 vccd1 vccd1 _3761_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__3078__A _3105_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5500_ _6228_/Q _5500_/B vssd1 vssd1 vccd1 vccd1 _5501_/B sky130_fd_sc_hd__nor2_1
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3692_ _5926_/A0 _3691_/X _3705_/A vssd1 vssd1 vccd1 vccd1 _6021_/D sky130_fd_sc_hd__mux2_1
XFILLER_118_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5431_ _5605_/B _5429_/Y _5452_/B _5425_/Y _3059_/Y vssd1 vssd1 vccd1 vccd1 _5431_/X
+ sky130_fd_sc_hd__o311a_1
XANTENNA__5524__A1 _3121_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3535__B1 _3589_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5362_ _4642_/Y _5358_/Y _5361_/Y _4646_/A _5227_/A vssd1 vssd1 vccd1 vccd1 _5362_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_126_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4313_ _4313_/A _4313_/B vssd1 vssd1 vccd1 vccd1 _4315_/B sky130_fd_sc_hd__or2_4
XFILLER_114_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5293_ _5292_/B _5292_/C _6221_/Q vssd1 vssd1 vccd1 vccd1 _5293_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__5288__B1 _5250_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4244_ _6091_/Q _3724_/X _4246_/S vssd1 vssd1 vccd1 vccd1 _6091_/D sky130_fd_sc_hd__mux2_1
XFILLER_87_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3838__A1 _4214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4175_ _4202_/A _4176_/B vssd1 vssd1 vccd1 vccd1 _4177_/B sky130_fd_sc_hd__nand2_2
XFILLER_67_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3541__A _3541_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3126_ _3126_/A _5647_/B _3126_/C vssd1 vssd1 vccd1 vccd1 _3127_/C sky130_fd_sc_hd__nand3_1
XFILLER_83_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5055__A3 _5075_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3057_ _5218_/B _3058_/B vssd1 vssd1 vccd1 vccd1 _3057_/X sky130_fd_sc_hd__and2_1
XFILLER_24_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4263__A1 _4362_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4263__B2 _4334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5212__B1 _5456_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3959_ _5148_/A _5634_/C _5203_/A _5635_/A vssd1 vssd1 vccd1 vccd1 _5105_/A sky130_fd_sc_hd__a22o_1
XANTENNA__3774__A0 _4657_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4971__C1 _5071_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5515__A1 _3331_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5629_ _5710_/S _3709_/X _5236_/Y _5734_/A _3950_/C vssd1 vssd1 vccd1 vccd1 _5629_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__5515__B2 _5943_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4723__C1 _5866_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4254__A1 _3715_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4006__A1 _3766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5754__A1 _3942_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4557__A2 _4252_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3517__B1 _3312_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4176__B _4176_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3080__B _5227_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5980_ _5985_/C _5979_/X _5978_/X _4576_/A vssd1 vssd1 vccd1 vccd1 _6300_/D sky130_fd_sc_hd__o211a_1
XANTENNA__4245__A1 _3727_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4931_ _5051_/D _4931_/B _4931_/C _4931_/D vssd1 vssd1 vccd1 vccd1 _4931_/X sky130_fd_sc_hd__or4_1
XFILLER_17_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4862_ _4867_/A _4862_/B vssd1 vssd1 vccd1 vccd1 _4862_/X sky130_fd_sc_hd__xor2_2
XFILLER_32_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3813_ _3849_/B _3813_/B vssd1 vssd1 vccd1 vccd1 _3813_/X sky130_fd_sc_hd__or2_1
X_4793_ _4990_/A _4793_/B vssd1 vssd1 vccd1 vccd1 _4793_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__4920__A _5488_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3744_ _5124_/S _3744_/B _3744_/C vssd1 vssd1 vccd1 vccd1 _3777_/S sky130_fd_sc_hd__or3_4
X_3675_ _4638_/A _5403_/A vssd1 vssd1 vccd1 vccd1 _5072_/C sky130_fd_sc_hd__nor2_4
XFILLER_133_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5414_ _5385_/A _5556_/A2 _5413_/X _5556_/C1 vssd1 vssd1 vccd1 vccd1 _6224_/D sky130_fd_sc_hd__o211a_1
XFILLER_133_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5345_ _5653_/A _5342_/X _5343_/Y _5344_/Y _5227_/Y vssd1 vssd1 vccd1 vccd1 _5345_/X
+ sky130_fd_sc_hd__o311a_2
XFILLER_114_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5276_ _5227_/B _5275_/X _5272_/Y _5607_/B1 vssd1 vssd1 vccd1 vccd1 _5276_/X sky130_fd_sc_hd__a211o_1
XFILLER_101_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4227_ _4185_/B _4185_/Y _4224_/Y _4225_/X vssd1 vssd1 vccd1 vccd1 _4229_/A sky130_fd_sc_hd__a211o_1
XFILLER_75_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3271__A _4022_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4158_ _3831_/B _4069_/B _4072_/C _6084_/Q vssd1 vssd1 vccd1 vccd1 _4158_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_110_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3109_ _5096_/C _3114_/B vssd1 vssd1 vccd1 vccd1 _3109_/Y sky130_fd_sc_hd__nor2_1
XFILLER_55_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4089_ _4089_/A _4089_/B vssd1 vssd1 vccd1 vccd1 _4090_/B sky130_fd_sc_hd__or2_1
XFILLER_83_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_664 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5736__A1 _5710_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5736__B2 _3772_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5200__A3 _4596_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4830__A _6189_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3149__C _5712_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4041__S _4044_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3165__B _4462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3142__A_N _3970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3181__A _4638_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5672__B1 _3458_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4724__B _4726_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5727__A1 _3974_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5727__B2 _3958_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4162__D _4342_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3460_ _6203_/Q _3410_/B _3575_/B vssd1 vssd1 vccd1 vccd1 _3460_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3075__B _5244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3391_ _3636_/A _4620_/B vssd1 vssd1 vccd1 vccd1 _3391_/Y sky130_fd_sc_hd__nor2_1
X_5130_ _5191_/A _5647_/C _5986_/B1 vssd1 vssd1 vccd1 vccd1 _6209_/D sky130_fd_sc_hd__a21oi_1
XFILLER_69_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5061_ _4604_/A _4615_/Y _5060_/X _5640_/B vssd1 vssd1 vccd1 vccd1 _5249_/D sky130_fd_sc_hd__o211a_1
XFILLER_38_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4012_ _3032_/Y _5848_/A0 _3513_/B _4767_/A vssd1 vssd1 vccd1 vccd1 _4012_/X sky130_fd_sc_hd__o22a_1
XFILLER_84_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5963_ _5970_/A vssd1 vssd1 vccd1 vccd1 _5963_/Y sky130_fd_sc_hd__inv_2
XFILLER_92_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4914_ _4974_/A _4914_/B vssd1 vssd1 vccd1 vccd1 _4914_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_80_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5894_ _3518_/B _5677_/B _3510_/Y _3526_/B vssd1 vssd1 vccd1 vccd1 _5894_/X sky130_fd_sc_hd__o22a_1
XFILLER_33_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4845_ _4847_/A vssd1 vssd1 vccd1 vccd1 _4845_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4776_ _3101_/A _4770_/X _4775_/X _4946_/A vssd1 vssd1 vccd1 vccd1 _4776_/X sky130_fd_sc_hd__a2bb2o_2
XANTENNA_fanout227_A _6293_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_12_clk_A _6219_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3727_ _6016_/Q _3706_/Y _3726_/X vssd1 vssd1 vccd1 vccd1 _3727_/X sky130_fd_sc_hd__a21o_4
XANTENNA__3266__A _3266_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3658_ _3649_/A _3649_/B _3658_/S vssd1 vssd1 vccd1 vccd1 _3658_/X sky130_fd_sc_hd__mux2_1
XFILLER_106_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3589_ _6100_/Q _3589_/A2 _3589_/B1 _6093_/Q _5470_/S vssd1 vssd1 vccd1 vccd1 _3589_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_27_clk_A _6084_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5328_ _6222_/Q _4755_/X _5561_/S vssd1 vssd1 vccd1 vccd1 _5329_/A sky130_fd_sc_hd__mux2_1
XFILLER_88_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5259_ _5292_/B _5292_/C vssd1 vssd1 vccd1 vccd1 _5259_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__4457__A1 _3942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_870 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5654__A0 _4658_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5406__B1 _4058_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5656__A _5656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5185__A2 _5050_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3176__A _3880_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4448__A1 _3942_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout190 _3241_/Y vssd1 vssd1 vccd1 vccd1 _5742_/B sky130_fd_sc_hd__buf_6
XFILLER_93_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output23_A _6196_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3959__B1 _5203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5566__A _5567_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4630_ _4628_/X _4629_/Y _4972_/A vssd1 vssd1 vccd1 vccd1 _4630_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_30_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4561_ _3942_/A _4564_/A2 _4559_/X _4560_/X vssd1 vssd1 vccd1 vccd1 _6179_/D sky130_fd_sc_hd__a22o_1
XFILLER_128_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6300_ _6302_/CLK _6300_/D vssd1 vssd1 vccd1 vccd1 _6300_/Q sky130_fd_sc_hd__dfxtp_4
X_3512_ _3512_/A _5707_/B vssd1 vssd1 vccd1 vccd1 _3571_/B sky130_fd_sc_hd__nor2_4
X_4492_ _5856_/A _4501_/A2 _4490_/X _4491_/Y vssd1 vssd1 vccd1 vccd1 _6137_/D sky130_fd_sc_hd__a22o_1
X_6231_ _6232_/CLK _6231_/D vssd1 vssd1 vccd1 vccd1 _6231_/Q sky130_fd_sc_hd__dfxtp_1
X_3443_ _3444_/A _3444_/B vssd1 vssd1 vccd1 vccd1 _3443_/Y sky130_fd_sc_hd__nor2_8
XFILLER_131_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6162_ _6279_/CLK _6162_/D vssd1 vssd1 vccd1 vccd1 _6162_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3374_ _3374_/A _3374_/B vssd1 vssd1 vccd1 vccd1 _5653_/B sky130_fd_sc_hd__xnor2_4
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5113_ _5112_/X _6203_/Q _5129_/S vssd1 vssd1 vccd1 vccd1 _6203_/D sky130_fd_sc_hd__mux2_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6093_ _6093_/CLK _6093_/D vssd1 vssd1 vccd1 vccd1 _6093_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5044_ _5051_/D _5035_/Y _5043_/X _4963_/A vssd1 vssd1 vccd1 vccd1 _5044_/X sky130_fd_sc_hd__o22a_1
XFILLER_111_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5100__A2 _3111_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4645__A _5463_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout177_A _3709_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3662__A2 _3145_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5939__A1 _3948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5946_ _3240_/A _4586_/Y _5943_/X _5945_/X _4586_/B vssd1 vssd1 vccd1 vccd1 _5946_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout344_A input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4611__A1 _5712_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5877_ _6298_/Q _3972_/Y _3164_/C vssd1 vssd1 vccd1 vccd1 _5878_/D sky130_fd_sc_hd__a21o_1
XANTENNA__3695__S _3902_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5476__A _5476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4828_ _4860_/A _4828_/B vssd1 vssd1 vccd1 vccd1 _4829_/B sky130_fd_sc_hd__nand2_2
XANTENNA__5167__A2 _3950_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3708__B _3734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4759_ _4759_/A _4759_/B vssd1 vssd1 vccd1 vccd1 _4759_/X sky130_fd_sc_hd__or2_1
XFILLER_107_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5324__C1 _5556_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5875__B1 _5712_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4602__A1 _5075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5563__C1 _5507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_366 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5866__B1 _5866_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4449__B _4458_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5618__B1 _3940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3090_ _3170_/A _5143_/A vssd1 vssd1 vccd1 vccd1 _3090_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__5094__A1 _6198_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5633__A3 _4744_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_692 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5800_ _5800_/A _5818_/B vssd1 vssd1 vccd1 vccd1 _5801_/B sky130_fd_sc_hd__nor2_8
XFILLER_23_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3992_ _3868_/Y _3991_/X _3987_/X _3179_/X vssd1 vssd1 vccd1 vccd1 _3993_/B sky130_fd_sc_hd__o211a_1
XFILLER_16_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5731_ _4883_/B _4877_/B _5731_/S vssd1 vssd1 vccd1 vccd1 _5731_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5296__A _5296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5662_ _3388_/B _5203_/A _5728_/A _5661_/X vssd1 vssd1 vccd1 vccd1 _5662_/X sky130_fd_sc_hd__a211o_1
X_4613_ _4577_/C _3879_/X _5638_/B _5095_/A _3109_/Y vssd1 vssd1 vccd1 vccd1 _4613_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_30_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5593_ _5605_/C _5592_/X _5590_/Y _5227_/A vssd1 vssd1 vccd1 vccd1 _5593_/X sky130_fd_sc_hd__a211o_1
XFILLER_116_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4544_ _6174_/Q _4562_/B vssd1 vssd1 vccd1 vccd1 _4544_/X sky130_fd_sc_hd__or2_1
XANTENNA__5743__B _5743_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4475_ _3942_/A _4474_/X _4475_/S vssd1 vssd1 vccd1 vccd1 _6131_/D sky130_fd_sc_hd__mux2_1
XFILLER_117_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6214_ _6214_/CLK _6214_/D vssd1 vssd1 vccd1 vccd1 _6214_/Q sky130_fd_sc_hd__dfxtp_2
X_3426_ _6013_/Q _3231_/Y _3384_/X _3425_/X vssd1 vssd1 vccd1 vccd1 _6013_/D sky130_fd_sc_hd__o22a_1
XANTENNA__3332__A1 _5109_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3263__B _6067_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6145_ _6180_/CLK _6145_/D vssd1 vssd1 vccd1 vccd1 _6145_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3357_ _6202_/Q _3388_/B vssd1 vssd1 vccd1 vccd1 _3358_/B sky130_fd_sc_hd__nor2_4
XANTENNA_fanout294_A _5960_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6076_ _6259_/CLK _6076_/D vssd1 vssd1 vccd1 vccd1 _6076_/Q sky130_fd_sc_hd__dfxtp_1
X_3288_ _3164_/Y _3287_/A _3276_/X _3560_/S vssd1 vssd1 vccd1 vccd1 _3288_/X sky130_fd_sc_hd__a211o_1
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5027_ _6196_/Q _5027_/B vssd1 vssd1 vccd1 vccd1 _5036_/B sky130_fd_sc_hd__xnor2_1
XFILLER_54_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4094__B _4162_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3399__A1 _3388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5929_ _5928_/B _5927_/X _5928_/Y _5929_/B2 _4638_/A vssd1 vssd1 vccd1 vccd1 _5929_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_70_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5545__C1 _3060_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5934__A _5934_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3157__C _3970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5653__B _5653_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5848__A0 _5848_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4269__B _4426_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_751 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4520__A0 _4891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3173__B _4842_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3901__B _3901_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4823__A1 _3116_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5379__A2 _4234_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4732__B _4734_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3348__B _3986_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5000__A1 _4946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4260_ _4205_/B _4206_/X _4216_/A _4214_/B vssd1 vssd1 vccd1 vccd1 _4325_/A sky130_fd_sc_hd__o211a_2
XFILLER_4_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3211_ _3212_/A _3738_/A vssd1 vssd1 vccd1 vccd1 _3211_/Y sky130_fd_sc_hd__nor2_4
XFILLER_69_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4191_ _3842_/B _4069_/B _4072_/C _6085_/Q vssd1 vssd1 vccd1 vccd1 _4191_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_122_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3142_ _3970_/A _6070_/Q vssd1 vssd1 vccd1 vccd1 _3881_/A sky130_fd_sc_hd__nand2b_4
XFILLER_39_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4621__A_N _3495_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5067__A1 _6197_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4195__A _4270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3073_ _3121_/B _5330_/B vssd1 vssd1 vccd1 vccd1 _5169_/C sky130_fd_sc_hd__nand2_4
XFILLER_82_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_670 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4578__A0 _4622_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4642__B _4646_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3975_ _5976_/A _5870_/A _3975_/C vssd1 vssd1 vccd1 vccd1 _5206_/B sky130_fd_sc_hd__or3_4
XFILLER_51_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3539__A _3567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5714_ _5714_/A _5714_/B vssd1 vssd1 vccd1 vccd1 _5714_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__3258__B _3555_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5645_ _5645_/A _5645_/B vssd1 vssd1 vccd1 vccd1 _5648_/B sky130_fd_sc_hd__nor2_1
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5576_ _5567_/A _5250_/X _5575_/X _5948_/A vssd1 vssd1 vccd1 vccd1 _6231_/D sky130_fd_sc_hd__o211a_1
XANTENNA_fanout307_A _5800_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4527_ _4540_/A _6163_/Q vssd1 vssd1 vccd1 vccd1 _6162_/D sky130_fd_sc_hd__or2_1
XFILLER_116_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4458_ _6124_/Q _4458_/B vssd1 vssd1 vccd1 vccd1 _4458_/X sky130_fd_sc_hd__or2_1
XANTENNA__4502__A0 _5255_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3305__A1 _3575_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3409_ _6203_/Q _3410_/B vssd1 vssd1 vccd1 vccd1 _3465_/A sky130_fd_sc_hd__and2_2
X_4389_ _4426_/A _4389_/B _4389_/C vssd1 vssd1 vccd1 vccd1 _4391_/A sky130_fd_sc_hd__and3_1
XFILLER_86_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6128_ _6177_/CLK _6128_/D vssd1 vssd1 vccd1 vccd1 _6128_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6059_ _6260_/CLK _6059_/D vssd1 vssd1 vccd1 vccd1 _6059_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3449__A _3500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4044__S _4044_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3168__B _4946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3792__A1 _4690_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5518__C1 _5948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_787 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5533__A2 _5522_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3631__B _3631_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4833__A1_N _5385_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4462__B _4462_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4024__A2 _5207_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5277__C _5436_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3760_ _4659_/B _3740_/X _3749_/X _3759_/X vssd1 vssd1 vccd1 vccd1 _3760_/X sky130_fd_sc_hd__a211o_1
XFILLER_9_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3078__B _5239_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3691_ _6221_/Q _6021_/Q _3902_/A vssd1 vssd1 vccd1 vccd1 _3691_/X sky130_fd_sc_hd__mux2_1
X_5430_ _5391_/Y _5393_/X _5427_/Y _5428_/X vssd1 vssd1 vccd1 vccd1 _5452_/B sky130_fd_sc_hd__o211a_1
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5361_ _5361_/A vssd1 vssd1 vccd1 vccd1 _5361_/Y sky130_fd_sc_hd__inv_2
X_4312_ _4426_/A _4311_/B _4311_/C vssd1 vssd1 vccd1 vccd1 _4313_/B sky130_fd_sc_hd__a21oi_1
XFILLER_113_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5292_ _6221_/Q _5292_/B _5292_/C vssd1 vssd1 vccd1 vccd1 _5326_/B sky130_fd_sc_hd__and3_1
XFILLER_114_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5288__A1 _5595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_667 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4243_ _6090_/Q _3721_/X _4246_/S vssd1 vssd1 vccd1 vccd1 _6090_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3838__A2 _3777_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3822__A _5706_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4174_ _4135_/A _4135_/B _4135_/C vssd1 vssd1 vccd1 vccd1 _4177_/A sky130_fd_sc_hd__a21bo_4
XFILLER_67_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3125_ _5075_/C _4643_/A _5498_/A _5239_/A vssd1 vssd1 vccd1 vccd1 _3126_/C sky130_fd_sc_hd__a31o_1
XFILLER_55_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3056_ _5239_/A _3312_/B _4022_/C vssd1 vssd1 vccd1 vccd1 _5638_/A sky130_fd_sc_hd__or3_4
XANTENNA__5460__A1 _5454_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4263__A2 _4309_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout257_A _3943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5212__A1 _4633_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5212__B2 _4974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3958_ _3958_/A _4604_/A vssd1 vssd1 vccd1 vccd1 _3958_/Y sky130_fd_sc_hd__nor2_8
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3889_ _5911_/B _5911_/C _5911_/D _3888_/Y _3864_/X vssd1 vssd1 vccd1 vccd1 _3889_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_109_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5515__A2 _5442_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5628_ _6295_/Q _4615_/A _5627_/X _3772_/B vssd1 vssd1 vccd1 vccd1 _5628_/X sky130_fd_sc_hd__a211o_1
XFILLER_105_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5559_ _5578_/B _5559_/B vssd1 vssd1 vccd1 vccd1 _5572_/B sky130_fd_sc_hd__nor2_2
XANTENNA__5279__B2 _3236_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3732__A _3732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4039__S _4044_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_779 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5739__C1 _5728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4006__A2 _4767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3179__A _6071_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_551 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3642__A _3649_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4930_ _5034_/A _4983_/A _4930_/C vssd1 vssd1 vccd1 vccd1 _4931_/D sky130_fd_sc_hd__and3_1
XFILLER_52_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4787__A1_N _5360_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4861_ _4783_/Y _4860_/Y _4820_/B vssd1 vssd1 vccd1 vccd1 _4862_/B sky130_fd_sc_hd__o21a_2
XFILLER_60_451 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3812_ _3450_/D _3811_/X _3812_/S vssd1 vssd1 vccd1 vccd1 _3813_/B sky130_fd_sc_hd__mux2_1
X_4792_ _4828_/B _4792_/B vssd1 vssd1 vccd1 vccd1 _4793_/B sky130_fd_sc_hd__nand2_1
XFILLER_32_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3756__A1 _5226_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3743_ _5503_/A _3980_/B _3745_/C vssd1 vssd1 vccd1 vccd1 _3849_/B sky130_fd_sc_hd__and3_4
XANTENNA__4920__B _4979_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3674_ _5072_/A _5498_/A _3673_/Y _5238_/A vssd1 vssd1 vccd1 vccd1 _3678_/A sky130_fd_sc_hd__o22a_1
XFILLER_106_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5413_ _5058_/C _5389_/Y _5412_/Y _5251_/Y vssd1 vssd1 vccd1 vccd1 _5413_/X sky130_fd_sc_hd__a211o_1
XFILLER_133_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5344_ _5344_/A _5653_/A vssd1 vssd1 vccd1 vccd1 _5344_/Y sky130_fd_sc_hd__nand2_1
XFILLER_88_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5275_ _5603_/S _5258_/Y _5260_/Y _5274_/Y _5257_/Y vssd1 vssd1 vccd1 vccd1 _5275_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__4648__A _4648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4226_ _4185_/B _4185_/Y _4224_/Y _4225_/X vssd1 vssd1 vccd1 vccd1 _4226_/Y sky130_fd_sc_hd__a211oi_4
XANTENNA__5681__A1 _6302_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3271__B _5622_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4157_ _4157_/A _4157_/B vssd1 vssd1 vccd1 vccd1 _4157_/X sky130_fd_sc_hd__and2_1
XFILLER_96_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3692__A0 _5926_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3108_ _3958_/A _3669_/B vssd1 vssd1 vccd1 vccd1 _3114_/B sky130_fd_sc_hd__nor2_2
X_4088_ _4089_/A _4089_/B vssd1 vssd1 vccd1 vccd1 _4103_/A sky130_fd_sc_hd__nand2_2
XANTENNA__3698__S _3705_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3039_ _4974_/A vssd1 vssd1 vccd1 vccd1 _4943_/A sky130_fd_sc_hd__inv_2
XFILLER_70_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5736__A2 _3280_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4944__B1 _4972_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4830__B _5539_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5418__S _5539_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3181__B _5840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5424__A1 _5072_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5328__S _5561_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3356__B _3388_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5360__A0 _5367_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3390_ _4620_/B vssd1 vssd1 vccd1 vccd1 _3390_/Y sky130_fd_sc_hd__inv_2
XFILLER_130_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5112__A0 _3943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5060_ _5065_/A _5244_/B _5712_/S _3879_/X vssd1 vssd1 vccd1 vccd1 _5060_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4011_ _3033_/Y _3500_/C _3593_/A _5714_/A _4010_/Y vssd1 vssd1 vccd1 vccd1 _4011_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__5663__A1 _5075_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5962_ _5934_/A _3954_/Y _5961_/X vssd1 vssd1 vccd1 vccd1 _5970_/A sky130_fd_sc_hd__a21o_4
X_4913_ _4972_/B _4972_/C vssd1 vssd1 vccd1 vccd1 _4914_/B sky130_fd_sc_hd__nand2_1
X_5893_ _3518_/B _5677_/B _5891_/Y _3460_/X _5892_/X vssd1 vssd1 vccd1 vccd1 _5893_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4931__A _5051_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4844_ _4846_/A _4846_/B vssd1 vssd1 vccd1 vccd1 _4847_/A sky130_fd_sc_hd__nand2_1
XFILLER_32_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3729__A1 _4167_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3729__B2 _6233_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4775_ _5119_/A _4774_/X _4812_/S vssd1 vssd1 vccd1 vccd1 _4775_/X sky130_fd_sc_hd__mux2_1
XFILLER_119_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout122_A _3245_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3726_ _3488_/X _3684_/X _3708_/Y _6232_/Q vssd1 vssd1 vccd1 vccd1 _3726_/X sky130_fd_sc_hd__o22a_1
XANTENNA__3266__B _3266_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3657_ _3923_/B _3657_/B vssd1 vssd1 vccd1 vccd1 _3657_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__5351__B1 _4058_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3588_ _6065_/Q _5439_/A2 _5743_/B _6078_/Q vssd1 vssd1 vccd1 vccd1 _3588_/X sky130_fd_sc_hd__o22a_1
X_5327_ _5327_/A _5385_/C _5327_/C vssd1 vssd1 vccd1 vccd1 _5338_/A sky130_fd_sc_hd__or3_1
XANTENNA__3282__A _5818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5258_ _5258_/A _5507_/A vssd1 vssd1 vccd1 vccd1 _5258_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__4457__A2 _3900_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5654__A1 _4663_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4209_ _4209_/A _4209_/B _4209_/C vssd1 vssd1 vccd1 vccd1 _4210_/C sky130_fd_sc_hd__and3_2
XFILLER_75_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5189_ _5191_/A _5179_/A _5181_/Y _5188_/X _5071_/A vssd1 vssd1 vccd1 vccd1 _6213_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_56_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5002__A _6195_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4917__B1 _6192_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3192__A _5840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4448__A2 _3900_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout180 _4167_/C vssd1 vssd1 vccd1 vccd1 _4389_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_47_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout191 _3241_/Y vssd1 vssd1 vccd1 vccd1 _5743_/B sky130_fd_sc_hd__buf_6
XFILLER_75_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3131__S _3135_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3959__A1 _5148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3959__B2 _5635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4081__B1 _4176_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output16_A _6190_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4908__B1 _4812_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4560_ _4872_/A _4252_/A _4239_/B vssd1 vssd1 vccd1 vccd1 _4560_/X sky130_fd_sc_hd__o21a_1
XFILLER_129_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3511_ _3511_/A _3571_/A vssd1 vssd1 vccd1 vccd1 _3526_/A sky130_fd_sc_hd__nor2_2
X_4491_ _3010_/Y _4499_/B _4501_/A2 vssd1 vssd1 vccd1 vccd1 _4491_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__5582__A _6232_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6230_ _6230_/CLK _6230_/D vssd1 vssd1 vccd1 vccd1 _6230_/Q sky130_fd_sc_hd__dfxtp_2
X_3442_ _5818_/A _3555_/B _3442_/C vssd1 vssd1 vccd1 vccd1 _3444_/B sky130_fd_sc_hd__and3_4
XANTENNA__5884__A1 _3941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6161_ _6263_/CLK _6161_/D vssd1 vssd1 vccd1 vccd1 _6161_/Q sky130_fd_sc_hd__dfxtp_1
X_3373_ _3511_/A _3373_/B vssd1 vssd1 vccd1 vccd1 _3374_/B sky130_fd_sc_hd__or2_4
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5112_ _3943_/A _4697_/A _5124_/S vssd1 vssd1 vccd1 vccd1 _5112_/X sky130_fd_sc_hd__mux2_1
X_6092_ _6260_/CLK _6092_/D vssd1 vssd1 vccd1 vccd1 _6092_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5043_ _5567_/A _5463_/A _5042_/X _4638_/A vssd1 vssd1 vccd1 vccd1 _5043_/X sky130_fd_sc_hd__o22a_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5521__S _5539_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4645__B _4645_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3662__A3 _3986_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5945_ _5264_/A _5108_/B _5934_/B _5944_/X vssd1 vssd1 vccd1 vccd1 _5945_/X sky130_fd_sc_hd__a31o_1
XFILLER_80_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout337_A input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5876_ _5876_/A _5876_/B _5876_/C vssd1 vssd1 vccd1 vccd1 _5878_/C sky130_fd_sc_hd__and3_1
XFILLER_21_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5476__B _5476_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4827_ _5385_/A _4644_/Y _4825_/X _4826_/Y vssd1 vssd1 vccd1 vccd1 _4827_/X sky130_fd_sc_hd__o22a_1
XFILLER_21_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3708__C _4462_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4758_ _6187_/Q _4647_/B _4648_/Y _5344_/A vssd1 vssd1 vccd1 vccd1 _4759_/B sky130_fd_sc_hd__a22o_1
XFILLER_119_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3709_ _6011_/Q _6034_/Q _3709_/S vssd1 vssd1 vccd1 vccd1 _3709_/X sky130_fd_sc_hd__mux2_8
X_4689_ _4707_/B _4690_/B vssd1 vssd1 vccd1 vccd1 _4691_/A sky130_fd_sc_hd__or2_2
XFILLER_107_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5875__A1 _6298_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4836__A _5428_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3740__A _3740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3810__A0 _5119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5012__C1 _5227_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3187__A _5622_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5618__A1 _5622_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5618__B2 _5456_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_11_clk_A _6219_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3991_ _3878_/A _5241_/A _3975_/C _3988_/X _3990_/Y vssd1 vssd1 vccd1 vccd1 _3991_/X
+ sky130_fd_sc_hd__o41a_1
XFILLER_50_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5577__A _6232_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_26_clk_A _6084_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5730_ _5730_/A _5900_/A vssd1 vssd1 vccd1 vccd1 _5730_/X sky130_fd_sc_hd__or2_1
XFILLER_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5296__B _5296_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5661_ input2/X _3179_/X _5659_/X _5660_/X _3974_/C vssd1 vssd1 vccd1 vccd1 _5661_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_31_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3097__A _4946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4612_ _5239_/A _4612_/B _5095_/A vssd1 vssd1 vccd1 vccd1 _4618_/B sky130_fd_sc_hd__nor3_1
XANTENNA__5554__B1 _5058_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5592_ _6008_/Q _5360_/S _5560_/B _6007_/Q vssd1 vssd1 vccd1 vccd1 _5592_/X sky130_fd_sc_hd__a22o_1
XFILLER_129_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4543_ _3943_/C _4564_/A2 _4541_/X _4542_/Y vssd1 vssd1 vccd1 vccd1 _6173_/D sky130_fd_sc_hd__a22o_1
XFILLER_132_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5743__C _5743_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4474_ _5446_/B _6131_/Q _4476_/S vssd1 vssd1 vccd1 vccd1 _4474_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5857__A1 _3443_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6213_ _6214_/CLK _6213_/D vssd1 vssd1 vccd1 vccd1 _6213_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3425_ _3631_/A _3425_/B vssd1 vssd1 vccd1 vccd1 _3425_/X sky130_fd_sc_hd__and2_1
XFILLER_131_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6144_ _6144_/CLK _6144_/D vssd1 vssd1 vccd1 vccd1 _6144_/Q sky130_fd_sc_hd__dfxtp_1
X_3356_ _6202_/Q _3388_/B vssd1 vssd1 vccd1 vccd1 _3358_/A sky130_fd_sc_hd__and2_4
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5609__A1 _5058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6075_ _6260_/CLK _6075_/D vssd1 vssd1 vccd1 vccd1 _6075_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3287_ _3287_/A vssd1 vssd1 vccd1 vccd1 _5626_/B sky130_fd_sc_hd__inv_2
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4817__C1 _5034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout287_A _5768_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5026_ _4999_/B _5537_/A _4947_/Y _3041_/Y vssd1 vssd1 vccd1 vccd1 _5026_/Y sky130_fd_sc_hd__o211ai_2
XFILLER_38_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4094__C _4216_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4045__B1 _5075_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3399__A2 _3388_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5928_ _5928_/A _5928_/B vssd1 vssd1 vccd1 vccd1 _5928_/Y sky130_fd_sc_hd__nor2_2
X_5859_ _5859_/A _5862_/B vssd1 vssd1 vccd1 vccd1 _5859_/Y sky130_fd_sc_hd__nand2_1
XFILLER_21_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5934__B _5934_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3735__A _3736_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5848__A1 _5926_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3323__A2 _3322_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3901__C _5743_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5233__C1 _5470_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4240__S _4246_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3562__A2 _3567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3210_ _3549_/B _3210_/B _3210_/C _3210_/D vssd1 vssd1 vccd1 vccd1 _3218_/B sky130_fd_sc_hd__and4_1
XANTENNA__4511__A1 _3942_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4190_ _4193_/B _4190_/B vssd1 vssd1 vccd1 vccd1 _4190_/Y sky130_fd_sc_hd__nor2_2
XFILLER_79_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3141_ _3970_/A _6070_/Q vssd1 vssd1 vccd1 vccd1 _3365_/B sky130_fd_sc_hd__and2b_4
XFILLER_122_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5067__A2 _4604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3072_ _3072_/A _3111_/B vssd1 vssd1 vccd1 vccd1 _5605_/B sky130_fd_sc_hd__or2_4
XANTENNA__4195__B _4389_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5224__C1 _3060_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4578__A1 _6182_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3974_ _3886_/X _3974_/B _3974_/C vssd1 vssd1 vccd1 vccd1 _3984_/C sky130_fd_sc_hd__and3b_1
X_5713_ _5714_/B _5713_/B vssd1 vssd1 vccd1 vccd1 _5713_/X sky130_fd_sc_hd__or2_1
XANTENNA__3250__A1 _3590_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5644_ _5644_/A _5644_/B _5644_/C vssd1 vssd1 vccd1 vccd1 _5649_/B sky130_fd_sc_hd__and3_1
XFILLER_129_470 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5575_ _4586_/B _5572_/B _5572_/X _5574_/X _5251_/Y vssd1 vssd1 vccd1 vccd1 _5575_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3555__A _5818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4526_ _4539_/A _6162_/Q vssd1 vssd1 vccd1 vccd1 _6161_/D sky130_fd_sc_hd__and2_1
XFILLER_117_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4457_ _3942_/A _3900_/Y _4455_/X _4456_/X vssd1 vssd1 vccd1 vccd1 _6123_/D sky130_fd_sc_hd__a22o_1
XFILLER_116_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3305__A2 _3266_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3408_ _3564_/S _4690_/B _3407_/X vssd1 vssd1 vccd1 vccd1 _3408_/X sky130_fd_sc_hd__o21a_1
XFILLER_131_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4388_ _4388_/A _4426_/C vssd1 vssd1 vccd1 vccd1 _4389_/C sky130_fd_sc_hd__xor2_1
XFILLER_105_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6127_ _6177_/CLK _6127_/D vssd1 vssd1 vccd1 vccd1 _6127_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input7_A io_in[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3339_ _5818_/A _3555_/B _3339_/C vssd1 vssd1 vccd1 vccd1 _3339_/X sky130_fd_sc_hd__and3_1
XFILLER_112_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6058_ _6301_/CLK _6058_/D vssd1 vssd1 vccd1 vccd1 _6058_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5009_ _5015_/A _5009_/B vssd1 vssd1 vccd1 vccd1 _5009_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_45_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4018__B1 _5714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5230__A2 _5464_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3449__B _3458_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4060__S _4066_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3184__B _3736_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3912__B _5742_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4296__A _4296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_56_clk _6133_/CLK vssd1 vssd1 vccd1 vccd1 _6286_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_92_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4462__C _5925_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4024__A3 _3883_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3690_ _5935_/A0 _3689_/X _3705_/A vssd1 vssd1 vccd1 vccd1 _6020_/D sky130_fd_sc_hd__mux2_1
XFILLER_118_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3535__A2 _3589_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5360_ _5367_/A _6007_/Q _5360_/S vssd1 vssd1 vccd1 vccd1 _5361_/A sky130_fd_sc_hd__mux2_1
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4311_ _4426_/A _4311_/B _4311_/C vssd1 vssd1 vccd1 vccd1 _4313_/A sky130_fd_sc_hd__and3_1
XFILLER_114_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5291_ _5507_/A _5327_/A vssd1 vssd1 vccd1 vccd1 _5291_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__5590__A _5605_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4242_ _6089_/Q _3718_/X _4246_/S vssd1 vssd1 vccd1 vccd1 _6089_/D sky130_fd_sc_hd__mux2_1
XFILLER_99_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5693__C1 _3194_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4173_ _4214_/A _4173_/B vssd1 vssd1 vccd1 vccd1 _4178_/A sky130_fd_sc_hd__nand2_2
XFILLER_67_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3124_ _5097_/A _5192_/A vssd1 vssd1 vccd1 vccd1 _3734_/A sky130_fd_sc_hd__or2_4
XFILLER_27_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5445__C1 _5948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3055_ _5075_/A _4003_/C _3885_/A vssd1 vssd1 vccd1 vccd1 _3058_/B sky130_fd_sc_hd__and3_4
XFILLER_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_47_clk _6230_/CLK vssd1 vssd1 vccd1 vccd1 _6254_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_36_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5212__A2 _5330_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3957_ _5104_/A _3960_/C vssd1 vssd1 vccd1 vccd1 _5634_/C sky130_fd_sc_hd__nor2_2
XFILLER_50_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4971__A1 _4625_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3888_ _5241_/A _4608_/C _3887_/X _5138_/A _5943_/B vssd1 vssd1 vccd1 vccd1 _3888_/Y
+ sky130_fd_sc_hd__a2111oi_1
X_5627_ _6292_/Q _5692_/B vssd1 vssd1 vccd1 vccd1 _5627_/X sky130_fd_sc_hd__and2_1
XANTENNA__3285__A _6298_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4723__A1 _4625_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5558_ _6231_/Q _5558_/B vssd1 vssd1 vccd1 vccd1 _5559_/B sky130_fd_sc_hd__nor2_1
XFILLER_3_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4509_ _6152_/Q _4515_/B vssd1 vssd1 vccd1 vccd1 _4509_/X sky130_fd_sc_hd__or2_1
XFILLER_105_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5489_ _5291_/Y _5487_/Y _5488_/X _5607_/B1 vssd1 vssd1 vccd1 vccd1 _5489_/X sky130_fd_sc_hd__a31o_1
XANTENNA__5279__A2 _5767_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3732__B _5936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout65_A _4601_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4844__A _4846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_38_clk clkbuf_3_4__f_clk/X vssd1 vssd1 vccd1 vccd1 _6248_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3179__B _4577_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4962__A1 _5504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_563 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3195__A _3960_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3134__S _3135_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_29_clk clkbuf_3_5__f_clk/X vssd1 vssd1 vccd1 vccd1 _6279_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__4650__B1 _5172_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4860_ _4860_/A _4860_/B vssd1 vssd1 vccd1 vccd1 _4860_/Y sky130_fd_sc_hd__nand2_1
XFILLER_32_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3811_ _3593_/A _3810_/X _3811_/S vssd1 vssd1 vccd1 vccd1 _3811_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4791_ _4791_/A _4791_/B _4791_/C vssd1 vssd1 vccd1 vccd1 _4792_/B sky130_fd_sc_hd__nand3_1
XFILLER_21_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3742_ _3948_/A _5124_/S _5712_/S _3744_/C vssd1 vssd1 vccd1 vccd1 _3811_/S sky130_fd_sc_hd__or4_2
XFILLER_119_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3673_ _5158_/B _4647_/B vssd1 vssd1 vccd1 vccd1 _3673_/Y sky130_fd_sc_hd__nor2_1
X_5412_ _5412_/A _5412_/B vssd1 vssd1 vccd1 vccd1 _5412_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__3508__A2 _3513_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5902__B1 _3883_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5343_ _5295_/Y _5297_/Y _5340_/X _5341_/Y vssd1 vssd1 vccd1 vccd1 _5343_/Y sky130_fd_sc_hd__a211oi_4
XFILLER_99_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4469__A0 _3942_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5274_ _5311_/B vssd1 vssd1 vccd1 vccd1 _5274_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4648__B _5330_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4225_ _4225_/A _4225_/B _4225_/C vssd1 vssd1 vccd1 vccd1 _4225_/X sky130_fd_sc_hd__and3_2
XANTENNA__5130__A1 _5191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5681__A2 _4615_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4156_ _4153_/X _4154_/Y _4123_/Y _4126_/A vssd1 vssd1 vccd1 vccd1 _4157_/B sky130_fd_sc_hd__a211o_1
XFILLER_95_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3107_ _3107_/A _3107_/B vssd1 vssd1 vccd1 vccd1 _4596_/B sky130_fd_sc_hd__or2_4
XFILLER_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4087_ _4087_/A _4087_/B vssd1 vssd1 vccd1 vccd1 _4089_/B sky130_fd_sc_hd__nor2_1
XFILLER_24_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3038_ _6208_/Q vssd1 vssd1 vccd1 vccd1 _3649_/A sky130_fd_sc_hd__inv_2
XFILLER_102_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4989_ _4989_/A _4989_/B vssd1 vssd1 vccd1 vccd1 _4990_/B sky130_fd_sc_hd__xnor2_1
XFILLER_11_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3743__A _5503_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5121__A1 _4767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout340 input4/X vssd1 vssd1 vccd1 vccd1 _5114_/A sky130_fd_sc_hd__buf_6
XANTENNA__3132__A0 _5119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5672__A2 _3388_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4880__B1 _4806_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5424__A2 _5418_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5188__A1 _5075_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4935__A1 _6192_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3129__S _3135_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5112__A1 _4697_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4010_ _5226_/A _4010_/B vssd1 vssd1 vccd1 vccd1 _4010_/Y sky130_fd_sc_hd__nand2_1
XFILLER_84_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3674__A1 _5072_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4871__B1 _4931_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3674__B2 _5238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3426__A1 _6013_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5961_ _5961_/A _5961_/B _5961_/C _5961_/D vssd1 vssd1 vccd1 vccd1 _5961_/X sky130_fd_sc_hd__or4_1
XFILLER_52_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4912_ _5617_/B _4912_/B vssd1 vssd1 vccd1 vccd1 _4972_/C sky130_fd_sc_hd__and2_1
XFILLER_80_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5892_ _3460_/X _5891_/Y _3937_/C vssd1 vssd1 vccd1 vccd1 _5892_/X sky130_fd_sc_hd__o21ba_1
X_4843_ _4842_/B _4841_/X _4842_/Y _4972_/A vssd1 vssd1 vccd1 vccd1 _4843_/X sky130_fd_sc_hd__o211a_1
XFILLER_61_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4931__B _4931_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4774_ _4774_/A _4774_/B vssd1 vssd1 vccd1 vccd1 _4774_/X sky130_fd_sc_hd__xor2_1
X_3725_ _6031_/Q _3724_/X _3731_/S vssd1 vssd1 vccd1 vccd1 _6031_/D sky130_fd_sc_hd__mux2_1
XFILLER_119_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_9_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _6209_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_fanout115_A _3410_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3656_ _3619_/B _3623_/B _3652_/A vssd1 vssd1 vccd1 vccd1 _3657_/B sky130_fd_sc_hd__a21boi_1
XANTENNA__4659__A _5226_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3587_ _6056_/Q _3589_/A2 _3589_/B1 _6049_/Q _3586_/X vssd1 vssd1 vccd1 vccd1 _3587_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__3362__B1 _3621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5326_ _6222_/Q _5326_/B vssd1 vssd1 vccd1 vccd1 _5327_/C sky130_fd_sc_hd__nor2_1
XFILLER_114_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3282__B _3555_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5103__A1 _5870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5257_ _5305_/B _5257_/B vssd1 vssd1 vccd1 vccd1 _5257_/Y sky130_fd_sc_hd__nand2_2
XFILLER_87_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4208_ _4209_/A _4209_/B _4209_/C vssd1 vssd1 vccd1 vccd1 _4210_/B sky130_fd_sc_hd__a21oi_4
XFILLER_87_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5188_ _5075_/A _5187_/X _5186_/Y _3014_/A vssd1 vssd1 vccd1 vccd1 _5188_/X sky130_fd_sc_hd__a211o_1
XFILLER_29_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4139_ _4138_/A _4138_/B _4138_/C vssd1 vssd1 vccd1 vccd1 _4140_/B sky130_fd_sc_hd__a21oi_1
XFILLER_84_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5406__A2 _4234_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3417__A1 _3410_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5002__B _6194_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3457__B _3458_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_527 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4569__A _5928_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5893__A2 _5677_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3192__B _3952_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout170 _3239_/X vssd1 vssd1 vccd1 vccd1 _3901_/B sky130_fd_sc_hd__buf_6
Xfanout181 _3488_/X vssd1 vssd1 vccd1 vccd1 _4167_/C sky130_fd_sc_hd__buf_4
XFILLER_93_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout192 _3241_/Y vssd1 vssd1 vccd1 vccd1 _5924_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_47_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_750 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4081__A1 _4162_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4081__B2 _4096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_4__f_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_3_4__f_clk/X sky130_fd_sc_hd__clkbuf_16
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4243__S _4246_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4908__A1 _5454_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5030__B1 _5029_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5581__A1 _3536_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5581__B2 _4586_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3510_ _3571_/A vssd1 vssd1 vccd1 vccd1 _3510_/Y sky130_fd_sc_hd__inv_2
XFILLER_128_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4490_ _6137_/Q _4490_/B vssd1 vssd1 vccd1 vccd1 _4490_/X sky130_fd_sc_hd__or2_1
XFILLER_7_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3441_ _6269_/Q _6015_/Q _6083_/Q _6038_/Q _4067_/A _3551_/S vssd1 vssd1 vccd1 vccd1
+ _3442_/C sky130_fd_sc_hd__mux4_1
XFILLER_6_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5884__A2 _3937_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6160_ _6263_/CLK _6160_/D vssd1 vssd1 vccd1 vccd1 _6160_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3372_ _3658_/S _3388_/B _3371_/X vssd1 vssd1 vccd1 vccd1 _3373_/B sky130_fd_sc_hd__o21ai_4
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3895__A1 _5934_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5111_ _5110_/X _6202_/Q _5129_/S vssd1 vssd1 vccd1 vccd1 _6202_/D sky130_fd_sc_hd__mux2_1
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6091_ _6248_/CLK _6091_/D vssd1 vssd1 vccd1 vccd1 _6091_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5042_ _5551_/A _4640_/A _5041_/X _5038_/X _5403_/A vssd1 vssd1 vccd1 vccd1 _5042_/X
+ sky130_fd_sc_hd__o32a_1
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3647__A1 _3541_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5944_ _3869_/A _3575_/B _3893_/B _5934_/A _3943_/C vssd1 vssd1 vccd1 vccd1 _5944_/X
+ sky130_fd_sc_hd__o311a_2
XFILLER_34_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5875_ _6298_/Q _5957_/B _5712_/S _5911_/A vssd1 vssd1 vccd1 vccd1 _5876_/C sky130_fd_sc_hd__a211o_1
X_4826_ _5605_/C _5072_/C vssd1 vssd1 vccd1 vccd1 _4826_/Y sky130_fd_sc_hd__nand2_4
XANTENNA_fanout232_A _6290_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3277__B _6298_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4757_ _5543_/S _4743_/X _4646_/Y vssd1 vssd1 vccd1 vccd1 _4759_/A sky130_fd_sc_hd__o21ai_1
X_3708_ _3732_/A _3734_/A _4462_/B vssd1 vssd1 vccd1 vccd1 _3708_/Y sky130_fd_sc_hd__nor3_4
XFILLER_107_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4688_ _4664_/B _4666_/B _4662_/X vssd1 vssd1 vccd1 vccd1 _4692_/A sky130_fd_sc_hd__a21o_1
XANTENNA__5324__A1 _6221_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4389__A _4426_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3639_ _3398_/A _3987_/B _3637_/X _3498_/S vssd1 vssd1 vccd1 vccd1 _3639_/X sky130_fd_sc_hd__o211a_1
XFILLER_134_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3293__A _4010_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5875__A2 _5957_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5309_ _5551_/A _5308_/X _3122_/A vssd1 vssd1 vccd1 vccd1 _5309_/X sky130_fd_sc_hd__o21a_1
X_6289_ _6290_/CLK _6289_/D vssd1 vssd1 vccd1 vccd1 _6289_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5088__B1 _5072_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5712__S _5712_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3638__A1 _6298_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4836__B _4837_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_20 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5948__A _5948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_878 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4063__A1 _3721_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3810__A1 _3495_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4063__S _4066_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5012__B1 _4648_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3187__B _5635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5563__A1 _4644_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5563__B2 _3121_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5866__A2 _5867_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3931__A _5656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5618__A2 _4592_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3629__A1 _3511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3990_ _3942_/A _4608_/C _3989_/Y vssd1 vssd1 vccd1 vccd1 _3990_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_90_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4054__A1 _6070_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4054__B2 _4846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3378__A _5924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5660_ _3867_/B _3388_/A _3410_/B _3867_/A _3996_/B vssd1 vssd1 vccd1 vccd1 _5660_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5003__B1 _6195_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4611_ _5712_/S _3879_/X _5048_/B vssd1 vssd1 vccd1 vccd1 _5083_/A sky130_fd_sc_hd__o21a_1
XFILLER_129_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5591_ _6232_/Q _5454_/A _4638_/Y _5589_/X _3948_/A vssd1 vssd1 vccd1 vccd1 _5591_/X
+ sky130_fd_sc_hd__a32o_1
X_4542_ _5221_/A _4562_/B _4564_/A2 vssd1 vssd1 vccd1 vccd1 _4542_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_129_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4473_ _3942_/B _4472_/X _4475_/S vssd1 vssd1 vccd1 vccd1 _6130_/D sky130_fd_sc_hd__mux2_1
XFILLER_116_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6212_ _6214_/CLK _6212_/D vssd1 vssd1 vccd1 vccd1 _6212_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_131_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3424_ _3408_/X _3937_/C _3583_/S vssd1 vssd1 vccd1 vccd1 _3425_/B sky130_fd_sc_hd__mux2_4
XFILLER_89_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6143_ _6143_/CLK _6143_/D vssd1 vssd1 vccd1 vccd1 _6143_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3355_ _3227_/X _3351_/X _3354_/X vssd1 vssd1 vccd1 vccd1 _3355_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_112_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6074_ _6098_/CLK _6074_/D vssd1 vssd1 vccd1 vccd1 _6074_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3286_ _6298_/Q _3643_/A _3316_/A vssd1 vssd1 vccd1 vccd1 _3287_/A sky130_fd_sc_hd__o21a_2
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5025_ _5025_/A vssd1 vssd1 vccd1 vccd1 _5537_/A sky130_fd_sc_hd__inv_2
XFILLER_100_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout182_A _4112_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4094__D _4214_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4672__A _4672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4045__A1 _5561_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4045__B2 _4596_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5793__A1 _3715_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5927_ _5936_/A _5943_/A _5926_/X _5923_/X vssd1 vssd1 vccd1 vccd1 _5927_/X sky130_fd_sc_hd__o31a_1
X_5858_ _6285_/Q _5854_/A _5857_/Y _5866_/B1 vssd1 vssd1 vccd1 vccd1 _6285_/D sky130_fd_sc_hd__o211a_1
XANTENNA__5545__A1 _5072_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4809_ _4807_/X _4809_/B vssd1 vssd1 vccd1 vccd1 _4811_/A sky130_fd_sc_hd__and2b_1
X_5789_ _5480_/B _5791_/B _5769_/S vssd1 vssd1 vccd1 vccd1 _5789_/X sky130_fd_sc_hd__o21a_1
XFILLER_119_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout95_A _5148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5233__B1 _4058_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5784__A1 _3942_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3198__A _5635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3140_ _4462_/A _3228_/A vssd1 vssd1 vccd1 vccd1 _3212_/A sky130_fd_sc_hd__or2_4
XFILLER_121_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5067__A3 _3996_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3071_ _3072_/A _3111_/B vssd1 vssd1 vccd1 vccd1 _5456_/S sky130_fd_sc_hd__nor2_8
XANTENNA__5472__B1 _5058_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5775__A1 _5926_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3973_ _4577_/A _5158_/A _3950_/C _4580_/C vssd1 vssd1 vccd1 vccd1 _5644_/A sky130_fd_sc_hd__o31a_1
X_5712_ _3615_/B _5711_/X _5712_/S vssd1 vssd1 vccd1 vccd1 _5713_/B sky130_fd_sc_hd__mux2_1
XFILLER_50_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5643_ _3103_/Y _3188_/X _5617_/X _5632_/D _5839_/B vssd1 vssd1 vccd1 vccd1 _5649_/A
+ sky130_fd_sc_hd__o2111a_1
XFILLER_136_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5574_ _3484_/X _5909_/B _5573_/X vssd1 vssd1 vccd1 vccd1 _5574_/X sky130_fd_sc_hd__a21o_1
XFILLER_129_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3555__B _3555_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4525_ _4540_/A _6161_/Q vssd1 vssd1 vccd1 vccd1 _6160_/D sky130_fd_sc_hd__or2_1
XFILLER_116_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4456_ _5446_/B _4438_/S _4439_/S vssd1 vssd1 vccd1 vccd1 _4456_/X sky130_fd_sc_hd__o21a_1
XFILLER_131_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3407_ _3563_/S _4697_/B _3404_/X _3227_/X vssd1 vssd1 vccd1 vccd1 _3407_/X sky130_fd_sc_hd__a211o_1
XFILLER_132_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3305__A3 _3266_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4387_ _4410_/B _4410_/D vssd1 vssd1 vccd1 vccd1 _4426_/C sky130_fd_sc_hd__nand2_2
XFILLER_86_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6126_ _6155_/CLK _6126_/D vssd1 vssd1 vccd1 vccd1 _6126_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3710__B1 _3709_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3338_ _6267_/Q _6013_/Q _6081_/Q _6036_/Q _4067_/A _3713_/S vssd1 vssd1 vccd1 vccd1
+ _3339_/C sky130_fd_sc_hd__mux4_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3290__B _6008_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6057_ _6206_/CLK _6057_/D vssd1 vssd1 vccd1 vccd1 _6057_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_105_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3269_ _3636_/A _4620_/A vssd1 vssd1 vccd1 vccd1 _3269_/Y sky130_fd_sc_hd__nor2_1
X_5008_ _5547_/B _5029_/B _4984_/Y vssd1 vssd1 vccd1 vccd1 _5009_/B sky130_fd_sc_hd__a21oi_1
XTAP_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5498__A _5498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3777__A0 _4096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_10_clk_A _6219_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3145__A_N _3880_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5377__S0 _3241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4577__A _4577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_25_clk_A clkbuf_3_5__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3701__A0 _4891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5757__A1 _5856_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5270__A1_N _4645_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4310_ _4310_/A _4343_/A vssd1 vssd1 vccd1 vccd1 _4311_/C sky130_fd_sc_hd__xor2_1
XFILLER_99_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5290_ _5512_/A _5603_/S vssd1 vssd1 vccd1 vccd1 _5327_/A sky130_fd_sc_hd__nand2_4
XFILLER_113_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4241_ _6088_/Q _3715_/X _4246_/S vssd1 vssd1 vccd1 vccd1 _6088_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4172_ _4210_/A _4171_/C _4171_/A vssd1 vssd1 vccd1 vccd1 _4180_/B sky130_fd_sc_hd__a21o_1
XFILLER_67_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3123_ _3123_/A _5072_/B vssd1 vssd1 vccd1 vccd1 _4640_/A sky130_fd_sc_hd__nor2_8
XFILLER_95_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3054_ _5800_/A _3869_/A vssd1 vssd1 vccd1 vccd1 _3054_/Y sky130_fd_sc_hd__nand2_1
XFILLER_36_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5748__A1 _5935_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3956_ _5090_/A _5909_/A _5637_/B _3954_/Y vssd1 vssd1 vccd1 vccd1 _5874_/A sky130_fd_sc_hd__a22oi_4
XFILLER_32_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4971__A2 _5093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3887_ _5097_/A _5131_/B _3887_/C _3886_/X vssd1 vssd1 vccd1 vccd1 _3887_/X sky130_fd_sc_hd__or4b_1
X_5626_ _5707_/A _5626_/B vssd1 vssd1 vccd1 vccd1 _5626_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_fanout312_A _3029_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3285__B _6292_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4723__A2 _5093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5557_ _5567_/A _5558_/B vssd1 vssd1 vccd1 vccd1 _5578_/B sky130_fd_sc_hd__and2_2
XFILLER_105_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4508_ _5926_/A0 _3912_/Y _4506_/X _4507_/Y vssd1 vssd1 vccd1 vccd1 _6151_/D sky130_fd_sc_hd__a22o_1
XFILLER_2_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5488_ _5488_/A _5504_/C vssd1 vssd1 vccd1 vccd1 _5488_/X sky130_fd_sc_hd__or2_1
XFILLER_132_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4439_ _3943_/C _4438_/X _4439_/S vssd1 vssd1 vccd1 vccd1 _6117_/D sky130_fd_sc_hd__mux2_1
XFILLER_132_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6109_ _6274_/CLK _6109_/D vssd1 vssd1 vccd1 vccd1 _6109_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4844__B _4846_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5739__A1 _3986_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5739__B2 _3180_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5956__A _5956_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4962__A2 _4644_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5372__C1 _5607_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4246__S _4246_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3989__B1 _3205_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4650__A1 _6184_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3453__A2 _3450_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4650__B2 _3030_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3810_ _5119_/A _3495_/B _3810_/S vssd1 vssd1 vccd1 vccd1 _3810_/X sky130_fd_sc_hd__mux2_1
X_4790_ _4791_/A _4791_/C _4791_/B vssd1 vssd1 vccd1 vccd1 _4828_/B sky130_fd_sc_hd__a21o_1
XFILLER_14_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3741_ _5703_/A _3741_/B _4886_/B _3750_/C vssd1 vssd1 vccd1 vccd1 _3751_/A sky130_fd_sc_hd__or4_4
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3672_ _5543_/S _5158_/B vssd1 vssd1 vccd1 vccd1 _3672_/Y sky130_fd_sc_hd__nor2_2
X_5411_ _5403_/X _5404_/X _5410_/X vssd1 vssd1 vccd1 vccd1 _5412_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__4166__B1 _4167_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5902__A1 _4085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5342_ _5340_/X _5341_/Y _5295_/Y _5297_/Y vssd1 vssd1 vccd1 vccd1 _5342_/X sky130_fd_sc_hd__o211a_1
XFILLER_114_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5273_ _5258_/A _5603_/S _5227_/A vssd1 vssd1 vccd1 vccd1 _5311_/B sky130_fd_sc_hd__o21a_2
XFILLER_99_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4224_ _4225_/B _4225_/C _4225_/A vssd1 vssd1 vccd1 vccd1 _4224_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__4010__A _5226_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4155_ _4123_/A _4125_/A _4122_/A _4122_/B _4154_/B vssd1 vssd1 vccd1 vccd1 _4157_/A
+ sky130_fd_sc_hd__a2111o_4
XANTENNA__5418__A0 _4872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4945__A _4945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3106_ _3107_/A _3107_/B vssd1 vssd1 vccd1 vccd1 _5096_/C sky130_fd_sc_hd__nor2_8
XFILLER_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3429__C1 _5929_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4086_ _4136_/A _4311_/B _4085_/C _4085_/D vssd1 vssd1 vccd1 vccd1 _4087_/B sky130_fd_sc_hd__a22oi_1
XANTENNA__5969__A1 _3033_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3037_ _5428_/A vssd1 vssd1 vccd1 vccd1 _4850_/A sky130_fd_sc_hd__clkinv_4
XFILLER_71_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout262_A _4096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4988_ _4988_/A _4988_/B vssd1 vssd1 vccd1 vccd1 _4989_/B sky130_fd_sc_hd__nand2_1
XFILLER_23_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3939_ _5677_/B _5898_/B _3938_/Y _5900_/A vssd1 vssd1 vccd1 vccd1 _3940_/B sky130_fd_sc_hd__a31o_1
XFILLER_137_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5609_ _5058_/A _5598_/Y _5608_/X vssd1 vssd1 vccd1 vccd1 _5611_/A sky130_fd_sc_hd__a21o_1
XFILLER_3_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3743__B _3980_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3380__B2 _3236_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5657__B1 _3772_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout330 _5207_/S vssd1 vssd1 vccd1 vccd1 _5599_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_59_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5121__A2 _5241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout341 input4/X vssd1 vssd1 vccd1 vccd1 _5344_/A sky130_fd_sc_hd__buf_12
XFILLER_59_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_759 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4066__S _4066_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4590__A _4604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4935__A2 _4990_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5593__C1 _5227_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5345__C1 _5227_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4954__A1_N _4705_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5360__S _5360_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3674__A2 _5498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5960_ _3112_/B _3975_/C _5131_/B _5960_/C1 vssd1 vssd1 vccd1 vccd1 _5961_/D sky130_fd_sc_hd__a211o_1
XFILLER_80_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4911_ _4840_/A _4838_/B _4840_/B _4876_/X _4836_/X vssd1 vssd1 vccd1 vccd1 _4972_/B
+ sky130_fd_sc_hd__a311o_4
X_5891_ _5653_/B _5889_/X _5890_/X vssd1 vssd1 vccd1 vccd1 _5891_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_33_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4842_ _4850_/A _4842_/B vssd1 vssd1 vccd1 vccd1 _4842_/Y sky130_fd_sc_hd__nand2_1
XFILLER_60_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4773_ _4698_/A _4725_/X _4728_/X _4727_/B vssd1 vssd1 vccd1 vccd1 _4774_/B sky130_fd_sc_hd__a31oi_4
XFILLER_119_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3724_ _6015_/Q _3706_/Y _3723_/X vssd1 vssd1 vccd1 vccd1 _3724_/X sky130_fd_sc_hd__a21o_4
X_3655_ _3653_/X _3654_/Y _3621_/A vssd1 vssd1 vccd1 vccd1 _3655_/X sky130_fd_sc_hd__a21o_1
XFILLER_106_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3586_ _6264_/Q _5439_/A2 _5743_/B _6033_/Q vssd1 vssd1 vccd1 vccd1 _3586_/X sky130_fd_sc_hd__o22a_1
XANTENNA__5351__A2 _4234_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4659__B _4659_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout108_A _3593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5544__A2_N _5542_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5325_ _5333_/A _5326_/B vssd1 vssd1 vccd1 vccd1 _5385_/C sky130_fd_sc_hd__and2_2
XFILLER_130_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5256_ _5292_/B _5256_/B vssd1 vssd1 vccd1 vccd1 _5257_/B sky130_fd_sc_hd__or2_1
X_4207_ _4207_/A _4207_/B vssd1 vssd1 vccd1 vccd1 _4209_/C sky130_fd_sc_hd__xnor2_4
XFILLER_69_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5187_ _3050_/B _5244_/A _4648_/Y _5072_/B input8/X vssd1 vssd1 vccd1 vccd1 _5187_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__3665__A2 _4877_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4138_ _4138_/A _4138_/B _4138_/C vssd1 vssd1 vccd1 vccd1 _4171_/A sky130_fd_sc_hd__and3_2
XFILLER_28_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4069_ _4069_/A _4069_/B vssd1 vssd1 vccd1 vccd1 _4069_/Y sky130_fd_sc_hd__nor2_1
XFILLER_71_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5575__C1 _5251_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3754__A _6067_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout160 _3049_/Y vssd1 vssd1 vccd1 vccd1 _4646_/A sky130_fd_sc_hd__buf_12
XFILLER_87_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout171 _3180_/Y vssd1 vssd1 vccd1 vccd1 _3974_/C sky130_fd_sc_hd__buf_6
XFILLER_120_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout182 _4112_/D vssd1 vssd1 vccd1 vccd1 _4342_/B sky130_fd_sc_hd__clkbuf_16
XFILLER_75_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout193 _3235_/X vssd1 vssd1 vccd1 vccd1 _3243_/A sky130_fd_sc_hd__buf_6
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3408__A2 _4690_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4081__A2 _4173_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3648__B _3986_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4908__A2 _4883_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5030__A1 _5547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5581__A2 _5909_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5869__A0 _3958_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3440_ _6015_/Q _6038_/Q _3551_/S vssd1 vssd1 vccd1 vccd1 _3440_/X sky130_fd_sc_hd__mux2_2
XFILLER_6_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3371_ _6202_/Q _3575_/B vssd1 vssd1 vccd1 vccd1 _3371_/X sky130_fd_sc_hd__or2_2
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5110_ _5110_/A _5110_/B vssd1 vssd1 vccd1 vccd1 _5110_/X sky130_fd_sc_hd__and2_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6090_ _6093_/CLK _6090_/D vssd1 vssd1 vccd1 vccd1 _6090_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5041_ _6196_/Q _5040_/Y _5041_/S vssd1 vssd1 vccd1 vccd1 _5041_/X sky130_fd_sc_hd__mux2_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_832 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5943_ _5943_/A _5943_/B _5943_/C vssd1 vssd1 vccd1 vccd1 _5943_/X sky130_fd_sc_hd__or3_1
XFILLER_53_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5874_ _5874_/A _5874_/B _5874_/C vssd1 vssd1 vccd1 vccd1 _5951_/B sky130_fd_sc_hd__and3_1
XFILLER_34_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4825_ _6189_/Q _4647_/B _4648_/Y _4819_/B _4824_/Y vssd1 vssd1 vccd1 vccd1 _4825_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_21_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout225_A _5940_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4756_ _6187_/Q _4755_/X _5041_/S vssd1 vssd1 vccd1 vccd1 _4756_/X sky130_fd_sc_hd__mux2_1
XFILLER_119_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3583__A1 _5888_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3707_ _3732_/A _4462_/A vssd1 vssd1 vccd1 vccd1 _4072_/B sky130_fd_sc_hd__or2_4
X_4687_ _6185_/Q _4721_/B _4686_/Y _5047_/C1 vssd1 vssd1 vccd1 vccd1 _6185_/D sky130_fd_sc_hd__o211a_1
XANTENNA__3574__A _3621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3638_ _6298_/Q _3388_/A _3316_/A vssd1 vssd1 vccd1 vccd1 _3987_/B sky130_fd_sc_hd__o21a_2
XANTENNA__5324__A2 _5556_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4389__B _4389_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4532__B1 _4540_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3569_ _3935_/C _3516_/B _3571_/B vssd1 vssd1 vccd1 vccd1 _3570_/B sky130_fd_sc_hd__a21oi_2
XFILLER_1_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5308_ _3060_/Y _5300_/Y _5302_/Y _5307_/X vssd1 vssd1 vccd1 vccd1 _5308_/X sky130_fd_sc_hd__o22a_1
XFILLER_130_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6288_ _6288_/CLK _6288_/D vssd1 vssd1 vccd1 vccd1 _6288_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5088__A1 _6198_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5088__B2 _5403_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5239_ _5239_/A _5239_/B _5403_/A _5239_/D vssd1 vssd1 vccd1 vccd1 _5248_/B sky130_fd_sc_hd__or4_1
XANTENNA__4835__A1 _6189_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3638__A2 _3388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3740__C _4812_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5260__A1 _4642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3749__A _4592_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5012__A1 _6195_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output21_A _6195_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3051__A_N _4622_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5003__A1 _6194_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4610_ _5095_/A _3164_/C _5876_/B vssd1 vssd1 vccd1 vccd1 _5048_/B sky130_fd_sc_hd__o21a_1
X_5590_ _5605_/C _5595_/B vssd1 vssd1 vccd1 vccd1 _5590_/Y sky130_fd_sc_hd__nor2_1
XFILLER_129_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4541_ _6173_/Q _4562_/B vssd1 vssd1 vccd1 vccd1 _4541_/X sky130_fd_sc_hd__or2_1
XFILLER_128_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4472_ _5387_/A _6130_/Q _4476_/S vssd1 vssd1 vccd1 vccd1 _4472_/X sky130_fd_sc_hd__mux2_1
XFILLER_116_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6211_ _6214_/CLK _6211_/D vssd1 vssd1 vccd1 vccd1 _6211_/Q sky130_fd_sc_hd__dfxtp_1
X_3423_ _3511_/A _3412_/Y _3422_/X vssd1 vssd1 vccd1 vccd1 _3937_/C sky130_fd_sc_hd__o21ai_4
XFILLER_131_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6142_ _6180_/CLK _6142_/D vssd1 vssd1 vccd1 vccd1 _6142_/Q sky130_fd_sc_hd__dfxtp_1
X_3354_ _3564_/S _4663_/B _3476_/A vssd1 vssd1 vccd1 vccd1 _3354_/X sky130_fd_sc_hd__o21a_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_391 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6073_ _6248_/CLK _6073_/D vssd1 vssd1 vccd1 vccd1 _6073_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3285_ _6298_/Q _6292_/Q vssd1 vssd1 vccd1 vccd1 _3285_/Y sky130_fd_sc_hd__nand2_2
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4817__A1 _4745_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4817__B2 _4744_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5114__A _5114_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5024_ _6005_/Q _6006_/Q vssd1 vssd1 vccd1 vccd1 _5025_/A sky130_fd_sc_hd__nand2_1
XFILLER_38_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout175_A _3713_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4672__B _5263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4045__A2 _3112_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout342_A input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5926_ _5926_/A0 _5925_/Y _5943_/B vssd1 vssd1 vccd1 vccd1 _5926_/X sky130_fd_sc_hd__mux2_1
XFILLER_53_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5857_ _3443_/Y _5862_/B _5856_/Y _5867_/A1 vssd1 vssd1 vccd1 vccd1 _5857_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_21_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4808_ input6/X _4808_/B vssd1 vssd1 vccd1 vccd1 _4809_/B sky130_fd_sc_hd__or2_1
X_5788_ _6257_/Q _5788_/B vssd1 vssd1 vccd1 vccd1 _5788_/X sky130_fd_sc_hd__or2_1
XFILLER_119_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4739_ _3033_/Y _4806_/S _4737_/Y _4738_/X vssd1 vssd1 vccd1 vccd1 _4739_/X sky130_fd_sc_hd__o22a_1
XFILLER_107_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4505__A0 _5935_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5702__C1 _5956_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout88_A _5570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5481__A1 _5480_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3244__B1 _3589_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3547__A1 _3387_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3942__A _3942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3070_ _3107_/A _3126_/A vssd1 vssd1 vccd1 vccd1 _3070_/X sky130_fd_sc_hd__or2_2
XFILLER_36_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5224__A1 _4643_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3389__A _3500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3972_ _5883_/A _5124_/S vssd1 vssd1 vccd1 vccd1 _3972_/Y sky130_fd_sc_hd__nand2_2
XFILLER_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5711_ _5707_/A _5710_/X _5707_/Y vssd1 vssd1 vccd1 vccd1 _5711_/X sky130_fd_sc_hd__a21o_1
XFILLER_31_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5642_ _5645_/A _5642_/B _5641_/X vssd1 vssd1 vccd1 vccd1 _5728_/A sky130_fd_sc_hd__or3b_4
X_5573_ _5412_/A _5569_/X _5571_/X _5312_/B _5572_/B vssd1 vssd1 vccd1 vccd1 _5573_/X
+ sky130_fd_sc_hd__o32a_1
XANTENNA__5109__A _5109_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4524_ _4539_/A _6160_/Q vssd1 vssd1 vccd1 vccd1 _6159_/D sky130_fd_sc_hd__and2_1
XFILLER_116_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4455_ _6123_/Q _4458_/B vssd1 vssd1 vccd1 vccd1 _4455_/X sky130_fd_sc_hd__or2_1
XFILLER_104_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5543__S _5543_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3406_ _3646_/B _3500_/A _3400_/X _3541_/A _3405_/X vssd1 vssd1 vccd1 vccd1 _4690_/B
+ sky130_fd_sc_hd__o221a_4
X_4386_ _3807_/B _4295_/A _4385_/Y vssd1 vssd1 vccd1 vccd1 _6112_/D sky130_fd_sc_hd__o21ai_1
XFILLER_131_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3710__A1 _5488_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6125_ _6227_/CLK _6125_/D vssd1 vssd1 vccd1 vccd1 _6125_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3710__B2 _5743_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3337_ _6013_/Q _6036_/Q _3551_/S vssd1 vssd1 vccd1 vccd1 _3337_/X sky130_fd_sc_hd__mux2_2
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6056_ _6260_/CLK _6056_/D vssd1 vssd1 vccd1 vccd1 _6056_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_640 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3268_ _3268_/A _3388_/A vssd1 vssd1 vccd1 vccd1 _4620_/A sky130_fd_sc_hd__xnor2_4
X_5007_ _5007_/A vssd1 vssd1 vccd1 vccd1 _5015_/A sky130_fd_sc_hd__clkinv_2
XFILLER_39_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3199_ _5734_/A _5710_/S vssd1 vssd1 vccd1 vccd1 _3324_/A sky130_fd_sc_hd__and2_2
XTAP_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5498__B _5512_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4018__A2 _3029_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3299__A _4010_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5909_ _5909_/A _5909_/B vssd1 vssd1 vccd1 vccd1 _5909_/Y sky130_fd_sc_hd__nor2_1
XFILLER_22_551 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5518__A2 _5251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4858__A _4872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5377__S1 _3241_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3762__A _5889_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4577__B _4643_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_746 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3701__S _3902_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3002__A _3766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3937__A _5889_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4717__B1 _5172_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5914__C1 _5191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3672__A _5543_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4240_ _6087_/Q _3711_/X _4246_/S vssd1 vssd1 vccd1 vccd1 _6087_/D sky130_fd_sc_hd__mux2_1
XFILLER_113_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5142__B1 _5075_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5693__A1 _3732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4171_ _4171_/A _4210_/A _4171_/C vssd1 vssd1 vccd1 vccd1 _4180_/A sky130_fd_sc_hd__nand3_4
XFILLER_67_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3122_ _3122_/A _5498_/A vssd1 vssd1 vccd1 vccd1 _3122_/Y sky130_fd_sc_hd__nand2_2
XFILLER_68_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5445__A1 _4872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5599__A _6233_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3053_ _5800_/A _3869_/A vssd1 vssd1 vccd1 vccd1 _3053_/X sky130_fd_sc_hd__and2_4
XFILLER_48_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4008__A _6066_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3759__A1 _4136_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3955_ _5128_/S _5911_/B _5911_/C _3955_/D vssd1 vssd1 vccd1 vccd1 _3955_/X sky130_fd_sc_hd__or4_1
XFILLER_50_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3886_ _5870_/A _5911_/B _5911_/C _3886_/D vssd1 vssd1 vccd1 vccd1 _3886_/X sky130_fd_sc_hd__or4_2
XANTENNA_fanout138_A _5503_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5625_ _5625_/A _5625_/B _5625_/C vssd1 vssd1 vccd1 vccd1 _5839_/B sky130_fd_sc_hd__or3_2
XANTENNA__5905__C1 _5065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5556_ _5547_/A _5556_/A2 _5554_/Y _5555_/Y _5556_/C1 vssd1 vssd1 vccd1 vccd1 _6230_/D
+ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout305_A _3873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4507_ _5305_/A _4515_/B _3912_/Y vssd1 vssd1 vccd1 vccd1 _4507_/Y sky130_fd_sc_hd__a21oi_1
X_5487_ _6227_/Q _5504_/C vssd1 vssd1 vccd1 vccd1 _5487_/Y sky130_fd_sc_hd__nand2_1
XFILLER_132_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4438_ _5768_/A0 _6117_/Q _4438_/S vssd1 vssd1 vccd1 vccd1 _4438_/X sky130_fd_sc_hd__mux2_1
XFILLER_104_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3695__A0 _5358_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4369_ _4335_/A _4363_/A _4338_/A vssd1 vssd1 vccd1 vccd1 _4370_/B sky130_fd_sc_hd__o21ba_4
XFILLER_86_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6108_ _6144_/CLK _6108_/D vssd1 vssd1 vccd1 vccd1 _6108_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6039_ _6041_/CLK _6039_/D vssd1 vssd1 vccd1 vccd1 _6039_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5302__A _5498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_698 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5739__A2 _3958_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5372__B1 _5359_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3922__A1 _3649_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4588__A _5090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5124__A0 _5859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_775 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3686__A0 _5768_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_47 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4635__C1 _5051_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4650__A2 _5543_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3740_ _3740_/A _3740_/B _4812_/S _3749_/C vssd1 vssd1 vccd1 vccd1 _3740_/X sky130_fd_sc_hd__and4_4
XFILLER_9_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3386__B _3500_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3671_ _4648_/A _5509_/C vssd1 vssd1 vccd1 vccd1 _3671_/Y sky130_fd_sc_hd__nand2_4
X_5410_ _4586_/B _5389_/Y _5409_/X _5909_/B vssd1 vssd1 vccd1 vccd1 _5410_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4166__A1 _4197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4166__B2 _4197_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5902__A2 _5957_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5341_ _5344_/A _5341_/B vssd1 vssd1 vccd1 vccd1 _5341_/Y sky130_fd_sc_hd__nor2_2
X_5272_ _5267_/Y _5271_/X _5512_/A vssd1 vssd1 vccd1 vccd1 _5272_/Y sky130_fd_sc_hd__a21oi_1
X_4223_ _4180_/A _4181_/C _4219_/Y _4220_/X vssd1 vssd1 vccd1 vccd1 _4225_/C sky130_fd_sc_hd__a211o_2
XANTENNA__4010__B _4010_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4154_ _4154_/A _4154_/B vssd1 vssd1 vccd1 vccd1 _4154_/Y sky130_fd_sc_hd__nand2_1
XFILLER_83_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3105_ _3105_/A _5075_/B vssd1 vssd1 vccd1 vccd1 _5095_/A sky130_fd_sc_hd__nor2_8
XFILLER_110_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3429__B1 _3589_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4085_ _4085_/A _4311_/B _4085_/C _4085_/D vssd1 vssd1 vccd1 vccd1 _4087_/A sky130_fd_sc_hd__and4_4
XANTENNA__5969__A2 _5158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3036_ _5392_/A vssd1 vssd1 vccd1 vccd1 _5714_/A sky130_fd_sc_hd__inv_2
XFILLER_83_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4961__A _6004_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout255_A _4301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4987_ _4987_/A _4987_/B vssd1 vssd1 vccd1 vccd1 _4988_/B sky130_fd_sc_hd__or2_1
XFILLER_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5268__S _5561_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_24_clk_A _6233_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3938_ _5888_/B _3938_/B vssd1 vssd1 vccd1 vccd1 _3938_/Y sky130_fd_sc_hd__nor2_1
X_3869_ _3869_/A _3869_/B vssd1 vssd1 vccd1 vccd1 _3893_/C sky130_fd_sc_hd__nand2_2
XFILLER_137_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5608_ _6233_/Q _5599_/B _5108_/B _3122_/A vssd1 vssd1 vccd1 vccd1 _5608_/X sky130_fd_sc_hd__a31o_1
XANTENNA__3904__A1 _3715_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_39_clk_A clkbuf_3_4__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5539_ _5547_/A _5015_/Y _5539_/S vssd1 vssd1 vccd1 vccd1 _5551_/B sky130_fd_sc_hd__mux2_1
XFILLER_117_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5106__A0 _4085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3380__A2 _5743_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5657__A1 _5940_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout320 _5799_/A vssd1 vssd1 vccd1 vccd1 _5956_/A sky130_fd_sc_hd__buf_6
Xfanout331 input8/X vssd1 vssd1 vccd1 vccd1 _5207_/S sky130_fd_sc_hd__buf_6
XANTENNA__5731__S _5731_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout342 input3/X vssd1 vssd1 vccd1 vccd1 _4707_/B sky130_fd_sc_hd__buf_8
XFILLER_87_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5409__A1 _5929_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4590__B _5635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4111__A _4270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3950__A _5131_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5820__A1 _5835_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4910_ _4974_/A _4910_/B vssd1 vssd1 vccd1 vccd1 _4910_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5890_ _3374_/A _5889_/X _3373_/B vssd1 vssd1 vccd1 vccd1 _5890_/X sky130_fd_sc_hd__o21a_1
XFILLER_45_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4841_ _4841_/A _4841_/B vssd1 vssd1 vccd1 vccd1 _4841_/X sky130_fd_sc_hd__xor2_2
XFILLER_61_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4772_ _5119_/A _4772_/B vssd1 vssd1 vccd1 vccd1 _4774_/A sky130_fd_sc_hd__xnor2_2
X_3723_ _4112_/D _5742_/C _3708_/Y _5567_/A vssd1 vssd1 vccd1 vccd1 _3723_/X sky130_fd_sc_hd__o22a_1
X_3654_ _3653_/A _3653_/C _3931_/B vssd1 vssd1 vccd1 vccd1 _3654_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_115_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3585_ _6016_/Q _3231_/Y _3584_/X vssd1 vssd1 vccd1 vccd1 _6016_/D sky130_fd_sc_hd__o21a_1
XANTENNA__3336__S _3551_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3898__B1 _5192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5324_ _6221_/Q _5556_/A2 _5323_/X _5556_/C1 vssd1 vssd1 vccd1 vccd1 _6221_/D sky130_fd_sc_hd__o211a_1
XFILLER_115_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5255_ _5292_/B _5255_/B vssd1 vssd1 vccd1 vccd1 _5305_/B sky130_fd_sc_hd__nand2_2
XFILLER_114_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4206_ _4362_/A _4311_/B _4207_/B vssd1 vssd1 vccd1 vccd1 _4206_/X sky130_fd_sc_hd__and3_1
XFILLER_84_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5186_ _5186_/A _5186_/B vssd1 vssd1 vccd1 vccd1 _5186_/Y sky130_fd_sc_hd__nor2_1
XFILLER_56_502 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4137_ _4137_/A vssd1 vssd1 vccd1 vccd1 _4138_/C sky130_fd_sc_hd__inv_2
X_4068_ _4069_/B vssd1 vssd1 vccd1 vccd1 _4071_/A sky130_fd_sc_hd__inv_2
XFILLER_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3019_ _6197_/Q vssd1 vssd1 vccd1 vccd1 _3019_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3100__A _5238_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3754__B _4294_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5027__A _6196_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout150 _5476_/A vssd1 vssd1 vccd1 vccd1 _5653_/A sky130_fd_sc_hd__buf_6
XFILLER_47_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout161 _3049_/Y vssd1 vssd1 vccd1 vccd1 _3112_/B sky130_fd_sc_hd__buf_4
Xfanout172 _5638_/A vssd1 vssd1 vccd1 vccd1 _5244_/A sky130_fd_sc_hd__buf_6
Xfanout183 _3440_/X vssd1 vssd1 vccd1 vccd1 _4112_/D sky130_fd_sc_hd__buf_8
XFILLER_120_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout194 _3235_/X vssd1 vssd1 vccd1 vccd1 _5439_/A2 sky130_fd_sc_hd__buf_4
XFILLER_47_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_866 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5802__A1 _4136_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5802__B2 _3322_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3010__A _5358_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5030__A2 _5547_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3945__A _5634_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5869__A1 _5119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3344__A2 _3388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3370_ _3960_/B _3358_/A _3369_/X vssd1 vssd1 vccd1 vccd1 _3374_/A sky130_fd_sc_hd__o21a_4
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5040_ _5040_/A _5040_/B vssd1 vssd1 vccd1 vccd1 _5040_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_844 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5942_ _5264_/A _4586_/Y _5921_/X vssd1 vssd1 vccd1 vccd1 _5947_/S sky130_fd_sc_hd__o21a_1
XFILLER_53_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5873_ _4003_/C _4605_/B _5872_/X _3969_/X vssd1 vssd1 vccd1 vccd1 _5874_/C sky130_fd_sc_hd__o211a_1
XFILLER_61_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4824_ _5509_/C _4824_/B vssd1 vssd1 vccd1 vccd1 _4824_/Y sky130_fd_sc_hd__nor2_1
XFILLER_21_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4755_ _4755_/A _4755_/B vssd1 vssd1 vccd1 vccd1 _4755_/X sky130_fd_sc_hd__xor2_4
XFILLER_119_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3706_ _3706_/A _5048_/C vssd1 vssd1 vccd1 vccd1 _3706_/Y sky130_fd_sc_hd__nor2_8
XANTENNA__5309__B1 _3122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout120_A _3274_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4686_ _5046_/B _4686_/B vssd1 vssd1 vccd1 vccd1 _4686_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_fanout218_A _5210_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3637_ _5207_/S _3636_/A _3211_/Y _3636_/Y vssd1 vssd1 vccd1 vccd1 _3637_/X sky130_fd_sc_hd__a211o_1
X_3568_ _3568_/A _3568_/B vssd1 vssd1 vccd1 vccd1 _3935_/D sky130_fd_sc_hd__nor2_4
XFILLER_0_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5307_ _3121_/B _5303_/X _5312_/A _4644_/B _3060_/B vssd1 vssd1 vccd1 vccd1 _5307_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_102_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6287_ _6288_/CLK _6287_/D vssd1 vssd1 vccd1 vccd1 _6287_/Q sky130_fd_sc_hd__dfxtp_1
X_3499_ _3498_/X _4163_/A _3560_/S vssd1 vssd1 vccd1 vccd1 _3499_/X sky130_fd_sc_hd__mux2_1
X_5238_ _5238_/A _5238_/B _5238_/C vssd1 vssd1 vccd1 vccd1 _5239_/D sky130_fd_sc_hd__or3_1
XFILLER_69_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5169_ _3971_/B _5169_/B _5169_/C vssd1 vssd1 vccd1 vccd1 _5169_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_96_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4599__A1 _5734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5310__A _5605_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5548__B1 _5547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5012__A2 _4647_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5456__S _5456_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3765__A _5108_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4596__A _5244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5484__C1 _5227_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3005__A _5924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5539__A0 _5547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3378__C _5436_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3675__A _4638_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4540_ _4540_/A _6157_/Q vssd1 vssd1 vccd1 vccd1 _6172_/D sky130_fd_sc_hd__or2_1
XANTENNA__4762__A1 _6222_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4762__B2 _5239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_10_clk _6219_/CLK vssd1 vssd1 vccd1 vccd1 _6302_/CLK sky130_fd_sc_hd__clkbuf_16
X_4471_ _5856_/A _4470_/X _4475_/S vssd1 vssd1 vccd1 vccd1 _6129_/D sky130_fd_sc_hd__mux2_1
XFILLER_128_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6210_ _6214_/CLK _6210_/D vssd1 vssd1 vccd1 vccd1 _6210_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4514__A1 _5856_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3422_ _3422_/A _3422_/B _3422_/C vssd1 vssd1 vccd1 vccd1 _3422_/X sky130_fd_sc_hd__or3_2
XFILLER_131_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6141_ _6144_/CLK _6141_/D vssd1 vssd1 vccd1 vccd1 _6141_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3353_ _3353_/A _3353_/B vssd1 vssd1 vccd1 vccd1 _4663_/B sky130_fd_sc_hd__xor2_4
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6072_ _6260_/CLK _6072_/D vssd1 vssd1 vccd1 vccd1 _6072_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3284_ _3284_/A _3284_/B vssd1 vssd1 vccd1 vccd1 _3643_/A sky130_fd_sc_hd__or2_4
XFILLER_112_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4817__A2 _4813_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5023_ _6006_/Q _4973_/Y _4974_/X _3041_/Y vssd1 vssd1 vccd1 vccd1 _5023_/X sky130_fd_sc_hd__a31o_1
XANTENNA__5114__B _5957_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5490__A2 _5482_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout168_A _3239_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5925_ _5925_/A _5925_/B vssd1 vssd1 vccd1 vccd1 _5925_/Y sky130_fd_sc_hd__nand2_1
XFILLER_53_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4450__B1 _3900_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5856_ _5856_/A _5862_/B vssd1 vssd1 vccd1 vccd1 _5856_/Y sky130_fd_sc_hd__nand2_1
XFILLER_61_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout335_A input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4807_ input6/X _4808_/B vssd1 vssd1 vccd1 vccd1 _4807_/X sky130_fd_sc_hd__and2_1
X_5787_ _3942_/A _4250_/Y _5785_/X _5786_/X vssd1 vssd1 vccd1 vccd1 _6256_/D sky130_fd_sc_hd__a22o_1
X_4738_ _4691_/A _4735_/Y _4736_/X _4842_/B vssd1 vssd1 vccd1 vccd1 _4738_/X sky130_fd_sc_hd__a31o_1
XFILLER_108_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4669_ _6185_/Q _6184_/Q vssd1 vssd1 vccd1 vccd1 _4669_/X sky130_fd_sc_hd__xor2_1
XFILLER_107_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5305__A _5305_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5769__A0 _3943_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5233__A2 _4234_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3942__B _3942_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5215__A _5255_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3971_ _4577_/A _3971_/B vssd1 vssd1 vccd1 vccd1 _4580_/C sky130_fd_sc_hd__or2_2
XFILLER_90_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5710_ _3488_/X _5709_/X _5710_/S vssd1 vssd1 vccd1 vccd1 _5710_/X sky130_fd_sc_hd__mux2_1
XFILLER_43_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5641_ _5051_/D _3188_/X _5617_/X _5839_/B _5640_/X vssd1 vssd1 vccd1 vccd1 _5641_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_31_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5572_ _5595_/A _5572_/B vssd1 vssd1 vccd1 vccd1 _5572_/X sky130_fd_sc_hd__or2_1
X_4523_ _4540_/A _6159_/Q vssd1 vssd1 vccd1 vccd1 _6158_/D sky130_fd_sc_hd__or2_1
XFILLER_8_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5109__B _5124_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4454_ _3942_/B _3900_/Y _4452_/X _4453_/X vssd1 vssd1 vccd1 vccd1 _6122_/D sky130_fd_sc_hd__a22o_1
XFILLER_104_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3405_ _3611_/A _3405_/B _3405_/C vssd1 vssd1 vccd1 vccd1 _3405_/X sky130_fd_sc_hd__or3_1
XFILLER_131_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4385_ _6112_/Q _4296_/Y _4384_/Y _4437_/A1 vssd1 vssd1 vccd1 vccd1 _4385_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_98_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6124_ _6257_/CLK _6124_/D vssd1 vssd1 vccd1 vccd1 _6124_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3336_ _6275_/Q _6111_/Q _3551_/S vssd1 vssd1 vccd1 vccd1 _5296_/B sky130_fd_sc_hd__mux2_8
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6055_ _6258_/CLK _6055_/D vssd1 vssd1 vccd1 vccd1 _6055_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3267_ _3267_/A _3267_/B vssd1 vssd1 vccd1 vccd1 _3450_/A sky130_fd_sc_hd__nand2_8
XANTENNA_fanout285_A _6220_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5006_ _5547_/A _5029_/B vssd1 vssd1 vccd1 vccd1 _5007_/A sky130_fd_sc_hd__xor2_1
XFILLER_73_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3474__A1 _4726_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3198_ _5635_/A _3951_/C _3883_/A vssd1 vssd1 vccd1 vccd1 _3198_/X sky130_fd_sc_hd__or3_1
XTAP_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5908_ _5908_/A _5908_/B vssd1 vssd1 vccd1 vccd1 _6292_/D sky130_fd_sc_hd__nor2_1
XFILLER_14_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_563 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5839_ _5839_/A _5839_/B _5839_/C _5839_/D vssd1 vssd1 vccd1 vccd1 _5839_/X sky130_fd_sc_hd__and4_4
XFILLER_10_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3529__A2 _3937_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5923__B1 _5503_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4204__A _4334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4858__B _4979_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4577__C _4577_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4593__B _5258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3217__B2 _3706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_872 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3937__B _5653_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4717__B2 _4707_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5914__B1 _5635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5871__C _5871_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3672__B _5158_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4170_ _4169_/A _4169_/B _4169_/C vssd1 vssd1 vccd1 vccd1 _4171_/C sky130_fd_sc_hd__a21o_2
XFILLER_110_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3121_ _5218_/B _3121_/B vssd1 vssd1 vccd1 vccd1 _3121_/X sky130_fd_sc_hd__or2_4
XFILLER_121_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5445__A2 _5251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5599__B _5599_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3052_ _4622_/B _3970_/A vssd1 vssd1 vccd1 vccd1 _3312_/B sky130_fd_sc_hd__nand2b_4
XFILLER_36_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4653__B1 _5069_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3759__A2 _3777_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3954_ _5959_/B _4615_/B vssd1 vssd1 vccd1 vccd1 _3954_/Y sky130_fd_sc_hd__nor2_2
X_3885_ _3885_/A _3975_/C vssd1 vssd1 vccd1 vccd1 _3886_/D sky130_fd_sc_hd__nor2_1
XFILLER_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5624_ _5048_/C _5623_/X _3025_/Y vssd1 vssd1 vccd1 vccd1 _5632_/D sky130_fd_sc_hd__a21o_1
XFILLER_117_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5381__A1 _5442_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5555_ _5494_/A _5542_/X _5556_/A2 vssd1 vssd1 vccd1 vccd1 _5555_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__4959__A _5509_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4506_ _6151_/Q _4515_/B vssd1 vssd1 vccd1 vccd1 _4506_/X sky130_fd_sc_hd__or2_1
X_5486_ _5478_/Y _5485_/X _5551_/A vssd1 vssd1 vccd1 vccd1 _5486_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_132_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4437_ _4437_/A1 _4436_/Y _4434_/X vssd1 vssd1 vccd1 vccd1 _6116_/D sky130_fd_sc_hd__a21o_1
XFILLER_104_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4368_ _4393_/B _4368_/B vssd1 vssd1 vccd1 vccd1 _4370_/A sky130_fd_sc_hd__or2_4
XFILLER_86_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6107_ _6143_/CLK _6107_/D vssd1 vssd1 vccd1 vccd1 _6107_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_input5_A io_in[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_758 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3319_ _3312_/B _3310_/A _3308_/Y _3365_/B _3145_/C vssd1 vssd1 vccd1 vccd1 _3319_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4299_ _4266_/A _4268_/B _4266_/B vssd1 vssd1 vccd1 vccd1 _4320_/A sky130_fd_sc_hd__o21ba_4
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6038_ _6280_/CLK _6038_/D vssd1 vssd1 vccd1 vccd1 _6038_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3447__A1 _4162_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3103__A _4963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4947__A1 _4946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5372__A1 _5464_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5372__B2 _4644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5124__A1 _4819_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3135__A0 _5072_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_787 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3712__S _3731_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_59 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4635__B1 _5050_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4109__A _4163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3013__A _5255_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3948__A _3948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4938__A1 _5543_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5060__B1 _5712_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3670_ _5054_/A _5330_/B vssd1 vssd1 vccd1 vccd1 _4647_/B sky130_fd_sc_hd__nor2_8
XANTENNA__5363__A1 _5498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4166__A2 _4167_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4779__A _5358_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3683__A _5512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5340_ _5344_/A _5341_/B vssd1 vssd1 vccd1 vccd1 _5340_/X sky130_fd_sc_hd__and2_2
XFILLER_126_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5271_ _5072_/B _5284_/B _5270_/X _5507_/A vssd1 vssd1 vccd1 vccd1 _5271_/X sky130_fd_sc_hd__a211o_1
XFILLER_99_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4222_ _4219_/Y _4220_/X _4180_/A _4181_/C vssd1 vssd1 vccd1 vccd1 _4225_/B sky130_fd_sc_hd__o211ai_4
XFILLER_68_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4153_ _4154_/A _4154_/B vssd1 vssd1 vccd1 vccd1 _4153_/X sky130_fd_sc_hd__or2_2
XFILLER_110_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5403__A _5403_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3104_ _5731_/S _4592_/A _4753_/A _4612_/B _5075_/A vssd1 vssd1 vccd1 vccd1 _3104_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_95_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4084_ _4084_/A _4084_/B vssd1 vssd1 vccd1 vccd1 _4085_/D sky130_fd_sc_hd__or2_1
XFILLER_95_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4626__B1 _3030_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3035_ _6205_/Q vssd1 vssd1 vccd1 vccd1 _3512_/A sky130_fd_sc_hd__inv_2
XFILLER_71_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4961__B _5454_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout150_A _5476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4986_ _4984_/Y _4985_/X _4753_/A _5069_/A _4977_/X vssd1 vssd1 vccd1 vccd1 _4986_/X
+ sky130_fd_sc_hd__o2111a_1
XANTENNA_fanout248_A _4362_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3937_ _5889_/B _5653_/B _3937_/C _3937_/D vssd1 vssd1 vccd1 vccd1 _3938_/B sky130_fd_sc_hd__or4_1
XFILLER_137_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3868_ _5712_/S _5707_/A vssd1 vssd1 vccd1 vccd1 _3868_/Y sky130_fd_sc_hd__nand2_2
XFILLER_109_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5607_ _5604_/X _5606_/X _5607_/B1 vssd1 vssd1 vccd1 vccd1 _5607_/X sky130_fd_sc_hd__a21o_1
XANTENNA__4689__A _4707_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3799_ _3033_/Y _3845_/B _3737_/Y _3798_/Y vssd1 vssd1 vccd1 vccd1 _3799_/X sky130_fd_sc_hd__a211o_1
XANTENNA__3593__A _3593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5538_ _5536_/Y _5560_/B _3059_/Y vssd1 vssd1 vccd1 vccd1 _5538_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5106__A1 _5264_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5469_ _6156_/Q _3243_/A _5767_/B _6132_/Q _5468_/X vssd1 vssd1 vccd1 vccd1 _5469_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_87_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5657__A2 _4615_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout310 _6003_/Q vssd1 vssd1 vccd1 vccd1 _4974_/A sky130_fd_sc_hd__buf_6
Xfanout321 _3028_/Y vssd1 vssd1 vccd1 vccd1 _5799_/A sky130_fd_sc_hd__buf_8
Xfanout332 _5029_/B vssd1 vssd1 vccd1 vccd1 _4979_/B sky130_fd_sc_hd__buf_8
XANTENNA__4865__B1 _5172_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout343 input3/X vssd1 vssd1 vccd1 vccd1 _5296_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_87_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout63_A _4642_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_636 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3840__A1 _4837_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5593__A1 _5605_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5345__A1 _5653_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4111__B _4111_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3008__A _5547_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4856__B1 _4753_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3659__B2 _4003_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3950__B _4577_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5281__B1 _3704_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4840_ _4840_/A _4840_/B vssd1 vssd1 vccd1 vccd1 _4841_/B sky130_fd_sc_hd__nand2_1
XFILLER_61_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4771_ _5119_/A _4772_/B vssd1 vssd1 vccd1 vccd1 _4771_/Y sky130_fd_sc_hd__nand2_1
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3722_ _6030_/Q _3721_/X _3731_/S vssd1 vssd1 vccd1 vccd1 _6030_/D sky130_fd_sc_hd__mux2_1
XANTENNA__3595__B1 _3594_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5336__A1 _5072_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3653_ _3653_/A _3931_/B _3653_/C vssd1 vssd1 vccd1 vccd1 _3653_/X sky130_fd_sc_hd__or3_1
XFILLER_9_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3584_ _3631_/A _3583_/X _3537_/X _3592_/A vssd1 vssd1 vccd1 vccd1 _3584_/X sky130_fd_sc_hd__a211o_1
X_5323_ _5412_/A _5312_/A _5315_/X _5322_/X _5251_/Y vssd1 vssd1 vccd1 vccd1 _5323_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_114_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5254_ _5556_/A2 _5252_/X _5253_/Y vssd1 vssd1 vccd1 vccd1 _6219_/D sky130_fd_sc_hd__a21oi_1
XFILLER_69_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4205_ _4205_/A _4205_/B vssd1 vssd1 vccd1 vccd1 _4207_/B sky130_fd_sc_hd__nor2_4
XANTENNA__3860__B _5976_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5185_ input8/X _5050_/B _5158_/B _5147_/C _3958_/A vssd1 vssd1 vccd1 vccd1 _5186_/B
+ sky130_fd_sc_hd__a2111o_1
XFILLER_29_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5133__A _5570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout198_A _3922_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4136_ _4136_/A _4167_/C vssd1 vssd1 vccd1 vccd1 _4137_/A sky130_fd_sc_hd__nand2_1
XFILLER_96_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4972__A _4972_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4067_ _4067_/A _4294_/B vssd1 vssd1 vccd1 vccd1 _4069_/B sky130_fd_sc_hd__or2_4
XANTENNA__5272__B1 _5512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3018_ _6199_/Q vssd1 vssd1 vccd1 vccd1 _3297_/B sky130_fd_sc_hd__clkinv_4
XFILLER_52_720 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5575__A1 _4586_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4969_ _5504_/A _5871_/C _4968_/X _4931_/B vssd1 vssd1 vccd1 vccd1 _4969_/X sky130_fd_sc_hd__o22a_1
XFILLER_51_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3100__B _5169_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3586__B1 _5743_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout140 _3083_/Y vssd1 vssd1 vccd1 vccd1 _5957_/B sky130_fd_sc_hd__buf_6
Xfanout151 _5476_/A vssd1 vssd1 vccd1 vccd1 _5730_/A sky130_fd_sc_hd__clkbuf_4
Xfanout162 _5865_/S vssd1 vssd1 vccd1 vccd1 _5862_/B sky130_fd_sc_hd__clkbuf_16
Xfanout173 _3043_/Y vssd1 vssd1 vccd1 vccd1 _5075_/A sky130_fd_sc_hd__buf_8
Xfanout184 _4112_/C vssd1 vssd1 vccd1 vccd1 _4309_/B sky130_fd_sc_hd__buf_8
Xfanout195 _3236_/B vssd1 vssd1 vccd1 vccd1 _5436_/C sky130_fd_sc_hd__clkbuf_16
XFILLER_86_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5978__A _6300_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_878 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4066__A1 _3730_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5030__A3 _5504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5318__B2 _3236_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5218__A _5255_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3961__A _5158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3501__B1 _3513_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_38_clk_A clkbuf_3_4__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5941_ _5948_/A _5941_/B vssd1 vssd1 vccd1 vccd1 _6294_/D sky130_fd_sc_hd__and2_1
XFILLER_80_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3804__A1 _4726_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5872_ _4577_/A _4577_/C _5638_/B _5206_/B vssd1 vssd1 vccd1 vccd1 _5872_/X sky130_fd_sc_hd__o211a_1
XANTENNA__3201__A _5936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4823_ _3116_/X _4822_/X _4817_/X _4753_/A vssd1 vssd1 vccd1 vccd1 _4823_/X sky130_fd_sc_hd__o211a_1
X_4754_ _4713_/A _4713_/B _4750_/A vssd1 vssd1 vccd1 vccd1 _4755_/B sky130_fd_sc_hd__o21a_2
XANTENNA__4765__C1 _5866_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3705_ _3705_/A _5761_/S vssd1 vssd1 vccd1 vccd1 _3731_/S sky130_fd_sc_hd__nand2_8
XANTENNA__5309__A1 _5551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4685_ _4672_/A _4872_/B _4684_/Y _5069_/A vssd1 vssd1 vccd1 vccd1 _4686_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_135_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3636_ _3636_/A _5733_/B vssd1 vssd1 vccd1 vccd1 _3636_/Y sky130_fd_sc_hd__nor2_1
XFILLER_108_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3567_ _6206_/Q _3567_/B vssd1 vssd1 vccd1 vccd1 _3568_/B sky130_fd_sc_hd__nor2_2
XFILLER_68_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5306_ _5333_/B _5306_/B vssd1 vssd1 vccd1 vccd1 _5312_/A sky130_fd_sc_hd__nor2_2
X_6286_ _6286_/CLK _6286_/D vssd1 vssd1 vccd1 vccd1 _6286_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3498_ _3450_/D _3497_/X _3498_/S vssd1 vssd1 vccd1 vccd1 _3498_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5237_ _5256_/B _3949_/Y _5638_/B _5236_/A _5231_/X vssd1 vssd1 vccd1 vccd1 _5237_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_88_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5493__B1 _5482_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5168_ _3970_/A _5169_/C _4604_/B _5169_/B vssd1 vssd1 vccd1 vccd1 _5168_/X sky130_fd_sc_hd__a31o_1
XFILLER_29_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4119_ _4121_/A _4121_/B vssd1 vssd1 vccd1 vccd1 _4154_/A sky130_fd_sc_hd__nand2_1
XFILLER_17_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5099_ _3297_/B _5097_/X _5098_/Y _5192_/A vssd1 vssd1 vccd1 vccd1 _6199_/D sky130_fd_sc_hd__a211oi_1
XFILLER_16_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4599__A2 _4604_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3111__A _5075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5548__A1 _5540_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3765__B _3765_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4877__A _5454_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5181__C1 _5065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3781__A _5653_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4596__B _4596_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4039__A1 _3715_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5787__A1 _3942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4995__C1 _5058_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3675__B _5403_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4762__A2 _4587_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4470_ _5358_/A _6129_/Q _4476_/S vssd1 vssd1 vccd1 vccd1 _4470_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3421_ _3960_/B _3465_/A vssd1 vssd1 vccd1 vccd1 _3422_/C sky130_fd_sc_hd__nor2_1
XFILLER_98_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6140_ _6180_/CLK _6140_/D vssd1 vssd1 vccd1 vccd1 _6140_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3352_ _4010_/B _3507_/A _3611_/A vssd1 vssd1 vccd1 vccd1 _3353_/B sky130_fd_sc_hd__o21a_2
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6071_ _6209_/CLK _6071_/D vssd1 vssd1 vccd1 vccd1 _6071_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3283_ _3284_/A _3284_/B vssd1 vssd1 vccd1 vccd1 _3649_/B sky130_fd_sc_hd__nor2_8
XFILLER_39_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5022_ _6195_/Q _5046_/B _5021_/Y _5047_/C1 vssd1 vssd1 vccd1 vccd1 _6195_/D sky130_fd_sc_hd__o211a_1
XFILLER_57_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5020__A2_N _4872_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5778__A1 _3942_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4986__C1 _5069_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5924_ _5924_/A _5924_/B vssd1 vssd1 vccd1 vccd1 _5925_/B sky130_fd_sc_hd__nand2_1
XFILLER_41_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4450__A1 _3010_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5855_ _6284_/Q _5854_/A _5854_/Y _5866_/B1 vssd1 vssd1 vccd1 vccd1 _6284_/D sky130_fd_sc_hd__o211a_1
XFILLER_21_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3866__A _4577_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4806_ _5714_/A _4805_/Y _4806_/S vssd1 vssd1 vccd1 vccd1 _4806_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout230_A _5625_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout328_A input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5786_ _5446_/B _5791_/B _5769_/S vssd1 vssd1 vccd1 vccd1 _5786_/X sky130_fd_sc_hd__o21a_1
X_4737_ _4691_/A _4736_/X _4735_/Y vssd1 vssd1 vccd1 vccd1 _4737_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__5950__A1 _5911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5950__B2 _4697_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4668_ _3740_/A _4661_/X _4667_/X _4972_/A vssd1 vssd1 vccd1 vccd1 _4668_/X sky130_fd_sc_hd__a22o_2
XFILLER_119_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3619_ _3619_/A _3619_/B _3619_/C vssd1 vssd1 vccd1 vccd1 _3621_/B sky130_fd_sc_hd__and3_1
XANTENNA__4697__A _4697_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5702__A1 _4163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4599_ _5734_/A _4604_/C _5959_/A vssd1 vssd1 vccd1 vccd1 _5871_/A sky130_fd_sc_hd__a21o_1
XFILLER_116_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3713__A0 _6012_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6269_ _6272_/CLK _6269_/D vssd1 vssd1 vccd1 vccd1 _6269_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5466__B1 _5742_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4977__C1 _5034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3244__A2 _3589_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4441__A1 _5292_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3495__B _3495_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4901__C1 _4638_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3942__C _5856_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5215__B _5218_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3016__A _5258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_363 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4680__A1 _5263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3970_ _3970_/A _4604_/B vssd1 vssd1 vccd1 vccd1 _3971_/B sky130_fd_sc_hd__nand2_4
XFILLER_50_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5640_ _3127_/A _5640_/B _5919_/A _5640_/D vssd1 vssd1 vccd1 vccd1 _5640_/X sky130_fd_sc_hd__and4b_1
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4196__B1 _4167_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5571_ _5551_/A _5561_/X _5570_/X _5403_/A vssd1 vssd1 vccd1 vccd1 _5571_/X sky130_fd_sc_hd__o211a_1
X_4522_ _4539_/A _6158_/Q vssd1 vssd1 vccd1 vccd1 _6157_/D sky130_fd_sc_hd__and2_1
XFILLER_8_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4453_ _5387_/A _4438_/S _4439_/S vssd1 vssd1 vccd1 vccd1 _4453_/X sky130_fd_sc_hd__o21a_1
XFILLER_105_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3625__S _3658_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3404_ _4162_/B _3210_/B _3560_/S _3403_/X _3210_/C vssd1 vssd1 vccd1 vccd1 _3404_/X
+ sky130_fd_sc_hd__o221a_1
X_4384_ _4384_/A _4384_/B vssd1 vssd1 vccd1 vccd1 _4384_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_131_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6123_ _6248_/CLK _6123_/D vssd1 vssd1 vccd1 vccd1 _6123_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3335_ _3986_/A _3335_/B vssd1 vssd1 vccd1 vccd1 _4619_/A sky130_fd_sc_hd__xor2_4
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6054_ _6259_/CLK _6054_/D vssd1 vssd1 vccd1 vccd1 _6054_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3266_ _3266_/A _3266_/B vssd1 vssd1 vccd1 vccd1 _4010_/B sky130_fd_sc_hd__nor2_8
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5005_ _4745_/A _5000_/X _5001_/X _5011_/B _4744_/B vssd1 vssd1 vccd1 vccd1 _5005_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout180_A _4167_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3197_ _3873_/A _3197_/B vssd1 vssd1 vccd1 vccd1 _3883_/A sky130_fd_sc_hd__nand2_4
XFILLER_66_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5620__B1 _3941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5907_ _6292_/Q _5901_/X _4576_/A vssd1 vssd1 vccd1 vccd1 _5908_/B sky130_fd_sc_hd__o21ai_1
XFILLER_50_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5838_ _5838_/A _5838_/B vssd1 vssd1 vccd1 vccd1 _5839_/D sky130_fd_sc_hd__nor2_1
XFILLER_22_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5384__C1 _5556_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5923__A1 _5296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5769_ _3943_/C _5768_/X _5769_/S vssd1 vssd1 vccd1 vccd1 _6250_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4204__B _4301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3934__B1 _5241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5316__A _5436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout93_A _5058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5439__B1 _5743_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4890__A _4891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3217__A2 _3156_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3937__C _3937_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5914__A1 _3105_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5870__C_N _3975_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5678__A0 _4726_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5226__A _5226_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_691 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3120_ _4642_/A _3121_/B vssd1 vssd1 vccd1 vccd1 _5072_/B sky130_fd_sc_hd__nor2_8
XFILLER_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3051_ _4622_/B _3970_/A vssd1 vssd1 vccd1 vccd1 _4003_/C sky130_fd_sc_hd__and2b_4
XFILLER_83_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3953_ _3953_/A _3955_/D vssd1 vssd1 vccd1 vccd1 _5637_/B sky130_fd_sc_hd__nor2_2
XFILLER_16_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3884_ _3112_/B _4023_/A _3879_/X _5911_/C _4604_/B vssd1 vssd1 vccd1 vccd1 _3887_/C
+ sky130_fd_sc_hd__a2111o_1
XFILLER_137_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5623_ _4622_/B _5058_/A _3257_/B _3678_/B vssd1 vssd1 vccd1 vccd1 _5623_/X sky130_fd_sc_hd__a31o_1
X_5554_ _5552_/X _5553_/X _5058_/C vssd1 vssd1 vccd1 vccd1 _5554_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__5381__A2 _5380_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3863__B _5227_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3392__A1 _4697_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4505_ _5935_/A0 _4504_/X _4521_/S vssd1 vssd1 vccd1 vccd1 _6150_/D sky130_fd_sc_hd__mux2_1
X_5485_ _5072_/B _5491_/B _5484_/X vssd1 vssd1 vccd1 vccd1 _5485_/X sky130_fd_sc_hd__a21bo_1
XFILLER_105_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5669__B1 _3772_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4436_ _4429_/A _4429_/B _4435_/Y _4425_/Y _4432_/A vssd1 vssd1 vccd1 vccd1 _4436_/Y
+ sky130_fd_sc_hd__o221ai_4
XFILLER_116_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4341__B1 _4342_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4367_ _4410_/B _4389_/B _4366_/C vssd1 vssd1 vccd1 vccd1 _4368_/B sky130_fd_sc_hd__a21oi_2
XFILLER_98_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6106_ _6143_/CLK _6106_/D vssd1 vssd1 vccd1 vccd1 _6106_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3318_ _3316_/A _3316_/B _3316_/Y _4003_/C _4003_/B vssd1 vssd1 vccd1 vccd1 _3318_/X
+ sky130_fd_sc_hd__o2111a_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4298_ _4069_/A _4295_/A _4297_/Y vssd1 vssd1 vccd1 vccd1 _6109_/D sky130_fd_sc_hd__o21ai_1
XFILLER_100_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3249_ _6050_/Q _3589_/A2 _3589_/B1 _6043_/Q vssd1 vssd1 vccd1 vccd1 _3249_/X sky130_fd_sc_hd__o22a_1
X_6037_ _6278_/CLK _6037_/D vssd1 vssd1 vccd1 vccd1 _6037_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5841__A0 _4010_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3103__B _5128_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5357__C1 _5556_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3383__A1 _4270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3383__B2 _3382_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5046__A _6196_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3135__A1 _5054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4635__A1 _6184_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4635__B2 _4634_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4109__B _4173_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3948__B _5928_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3610__A2 _4846_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3964__A _5911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5363__A2 _5359_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4779__B _5367_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3683__B _5943_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4571__B1 _5203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5270_ _4645_/B _5257_/Y _5269_/X _3121_/B vssd1 vssd1 vccd1 vccd1 _5270_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4221_ _4221_/A _4221_/B _4221_/C vssd1 vssd1 vccd1 vccd1 _4221_/Y sky130_fd_sc_hd__nand3_2
XFILLER_99_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4874__A1 _6190_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4152_ _4152_/A _4152_/B vssd1 vssd1 vccd1 vccd1 _4154_/B sky130_fd_sc_hd__xnor2_2
XFILLER_110_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3103_ _4963_/A _5128_/S vssd1 vssd1 vccd1 vccd1 _3103_/Y sky130_fd_sc_hd__nand2_2
XFILLER_110_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5403__B _5403_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4083_ _4084_/A _4084_/B vssd1 vssd1 vccd1 vccd1 _4083_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__3429__A2 _3589_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4626__A1 _4812_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3034_ _5119_/A vssd1 vssd1 vccd1 vccd1 _4767_/A sky130_fd_sc_hd__inv_6
XFILLER_48_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3858__B _3869_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4985_ _4981_/A _4988_/A _4983_/X _3116_/X vssd1 vssd1 vccd1 vccd1 _4985_/X sky130_fd_sc_hd__a31o_1
XFILLER_23_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4035__A _5767_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3936_ _3311_/Y _3923_/Y _3925_/X _3935_/X _3934_/X vssd1 vssd1 vccd1 vccd1 _3936_/X
+ sky130_fd_sc_hd__o41a_1
XFILLER_32_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5339__C1 _5607_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3867_ _3867_/A _3867_/B vssd1 vssd1 vccd1 vccd1 _3867_/Y sky130_fd_sc_hd__nor2_2
X_5606_ _5227_/B _5598_/Y _5605_/X _5227_/A vssd1 vssd1 vccd1 vccd1 _5606_/X sky130_fd_sc_hd__a211o_1
XANTENNA_fanout310_A _6003_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5892__B1_N _3937_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4689__B _4690_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3798_ _4619_/B _3845_/B vssd1 vssd1 vccd1 vccd1 _3798_/Y sky130_fd_sc_hd__nor2_1
X_5537_ _5537_/A _5537_/B vssd1 vssd1 vccd1 vccd1 _5560_/B sky130_fd_sc_hd__and2_1
XFILLER_105_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5468_ _6180_/Q _4234_/B _4058_/B _6140_/Q vssd1 vssd1 vccd1 vccd1 _5468_/X sky130_fd_sc_hd__o22a_1
XFILLER_105_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4419_ _4419_/A _4419_/B _4419_/C vssd1 vssd1 vccd1 vccd1 _4420_/B sky130_fd_sc_hd__or3_1
Xfanout300 _6069_/Q vssd1 vssd1 vccd1 vccd1 _4003_/B sky130_fd_sc_hd__buf_8
Xfanout311 _5561_/S vssd1 vssd1 vccd1 vccd1 _5539_/S sky130_fd_sc_hd__buf_6
XFILLER_59_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4865__A1 _6190_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5399_ _4645_/B _5389_/Y _5398_/X _5570_/A vssd1 vssd1 vccd1 vccd1 _5399_/X sky130_fd_sc_hd__o211a_1
XFILLER_87_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4865__B2 _5029_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout322 input9/X vssd1 vssd1 vccd1 vccd1 _5192_/A sky130_fd_sc_hd__buf_8
Xfanout333 _4846_/A vssd1 vssd1 vccd1 vccd1 _5029_/B sky130_fd_sc_hd__buf_6
Xfanout344 input3/X vssd1 vssd1 vccd1 vccd1 _4697_/A sky130_fd_sc_hd__buf_8
XFILLER_87_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3114__A _5096_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5042__A1 _5551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5042__B2 _5403_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4002__C1 _3179_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5504__A _5504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4856__A1 _4705_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3950__C _3950_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3024__A _3948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4770_ _4767_/A _4769_/Y _4806_/S vssd1 vssd1 vccd1 vccd1 _4770_/X sky130_fd_sc_hd__mux2_1
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3595__A1 _3387_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3721_ _6014_/Q _3706_/Y _3720_/X vssd1 vssd1 vccd1 vccd1 _3721_/X sky130_fd_sc_hd__a21o_4
XFILLER_119_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3652_ _3652_/A _5898_/A vssd1 vssd1 vccd1 vccd1 _3653_/C sky130_fd_sc_hd__and2_1
X_3583_ _3564_/X _5888_/B _3583_/S vssd1 vssd1 vccd1 vccd1 _3583_/X sky130_fd_sc_hd__mux2_4
XANTENNA__5741__C1 _5956_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5322_ _5943_/C _5312_/A _5321_/X _5442_/A _5595_/A vssd1 vssd1 vccd1 vccd1 _5322_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_114_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5253_ _5256_/B _5556_/A2 _4576_/A vssd1 vssd1 vccd1 vccd1 _5253_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_88_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4204_ _4334_/A _4301_/A _4309_/B _4342_/B vssd1 vssd1 vccd1 vccd1 _4205_/B sky130_fd_sc_hd__and4_2
XFILLER_87_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5184_ _3116_/X _5143_/B _5182_/X _5183_/X vssd1 vssd1 vccd1 vccd1 _5186_/A sky130_fd_sc_hd__o22a_1
XFILLER_96_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4135_ _4135_/A _4135_/B _4135_/C vssd1 vssd1 vccd1 vccd1 _4138_/B sky130_fd_sc_hd__nand3_1
XFILLER_84_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_494 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4066_ _6078_/Q _3730_/X _4066_/S vssd1 vssd1 vccd1 vccd1 _6078_/D sky130_fd_sc_hd__mux2_1
XFILLER_83_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4972__B _4972_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3869__A _3869_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3017_ _6200_/Q vssd1 vssd1 vccd1 vccd1 _3296_/A sky130_fd_sc_hd__inv_2
XFILLER_36_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4968_ _5051_/D _4958_/X _4963_/X _4967_/X vssd1 vssd1 vccd1 vccd1 _4968_/X sky130_fd_sc_hd__o211a_1
X_3919_ _6054_/Q _3724_/X _3921_/S vssd1 vssd1 vccd1 vccd1 _6054_/D sky130_fd_sc_hd__mux2_1
XANTENNA__5980__C1 _4576_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4899_ _4867_/A _4867_/B _4925_/B vssd1 vssd1 vccd1 vccd1 _4900_/B sky130_fd_sc_hd__a21oi_4
XANTENNA_clkbuf_3_2__f_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3338__A1 _6013_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4535__B1 _4540_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3109__A _5096_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout130 _4654_/A vssd1 vssd1 vccd1 vccd1 _4931_/B sky130_fd_sc_hd__buf_6
Xfanout141 _3078_/Y vssd1 vssd1 vccd1 vccd1 _5605_/C sky130_fd_sc_hd__buf_8
Xfanout152 _3070_/X vssd1 vssd1 vccd1 vccd1 _5476_/A sky130_fd_sc_hd__buf_6
XFILLER_59_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout163 _3856_/X vssd1 vssd1 vccd1 vccd1 _5928_/B sky130_fd_sc_hd__buf_8
Xfanout174 _4214_/B vssd1 vssd1 vccd1 vccd1 _4176_/B sky130_fd_sc_hd__buf_4
XFILLER_87_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout185 _3394_/X vssd1 vssd1 vccd1 vccd1 _4112_/C sky130_fd_sc_hd__buf_6
XFILLER_87_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout196 _5617_/B vssd1 vssd1 vccd1 vccd1 _4806_/S sky130_fd_sc_hd__buf_4
XFILLER_86_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5802__A3 _4173_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3577__A1 _3658_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5030__A4 _5488_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_640 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5318__A2 _5767_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5218__B _5218_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5723__C1 _3950_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3019__A _6197_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5888__B _5888_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5254__A1 _5556_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5940_ _5940_/A0 _5939_/X _5940_/S vssd1 vssd1 vccd1 vccd1 _5941_/B sky130_fd_sc_hd__mux2_1
XFILLER_46_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3804__A2 _3740_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5871_ _5871_/A _5919_/A _5871_/C _5871_/D vssd1 vssd1 vccd1 vccd1 _5874_/B sky130_fd_sc_hd__and4_1
XFILLER_34_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3201__B _3706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4822_ _4925_/A _4822_/B vssd1 vssd1 vccd1 vccd1 _4822_/X sky130_fd_sc_hd__xor2_2
XFILLER_33_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4753_ _4753_/A _4753_/B _4753_/C vssd1 vssd1 vccd1 vccd1 _4753_/Y sky130_fd_sc_hd__nand3_1
X_3704_ _5767_/A _3704_/B _5767_/C vssd1 vssd1 vccd1 vccd1 _5761_/S sky130_fd_sc_hd__or3_4
X_4684_ _5051_/D _4677_/X _4683_/X vssd1 vssd1 vccd1 vccd1 _4684_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_107_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3635_ _3986_/B _3635_/B vssd1 vssd1 vccd1 vccd1 _5733_/B sky130_fd_sc_hd__xnor2_4
XFILLER_128_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout106_A _3557_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3566_ _3618_/A vssd1 vssd1 vccd1 vccd1 _3568_/A sky130_fd_sc_hd__inv_2
XFILLER_1_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5305_ _5305_/A _5305_/B vssd1 vssd1 vccd1 vccd1 _5306_/B sky130_fd_sc_hd__and2_1
XFILLER_130_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6285_ _6286_/CLK _6285_/D vssd1 vssd1 vccd1 vccd1 _6285_/Q sky130_fd_sc_hd__dfxtp_1
X_3497_ _3211_/Y _3593_/A _3495_/X _3496_/Y vssd1 vssd1 vccd1 vccd1 _3497_/X sky130_fd_sc_hd__a22o_1
XFILLER_102_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5236_ _5236_/A vssd1 vssd1 vccd1 vccd1 _5236_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5493__A1 _3250_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5493__B2 _5943_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5167_ _3112_/B _3950_/C _5179_/B _5164_/C vssd1 vssd1 vccd1 vccd1 _5169_/B sky130_fd_sc_hd__a211o_1
XANTENNA__5895__A2_N _3937_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4118_ _4099_/A _4099_/B _4094_/X vssd1 vssd1 vccd1 vccd1 _4121_/B sky130_fd_sc_hd__o21bai_1
XFILLER_84_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5098_ _6008_/Q _3111_/X _5097_/X vssd1 vssd1 vccd1 vccd1 _5098_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__5245__A1 _5911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3599__A _3599_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4049_ _3873_/A _4051_/S _5869_/S _4633_/B _4048_/Y vssd1 vssd1 vccd1 vccd1 _6066_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5650__D1 _5728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4877__B _4877_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3731__A1 _3730_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4596__C _5069_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5054__A _5054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5484__A1 _4645_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5484__B2 _4646_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_816 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3247__B1 _5743_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3302__A _3312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5944__C1 _3943_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4133__A _4162_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3972__A _5883_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3420_ _3365_/Y _3926_/A _3419_/Y _3960_/B vssd1 vssd1 vccd1 vccd1 _3422_/B sky130_fd_sc_hd__o211a_1
XANTENNA__3722__A1 _3721_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3351_ _3345_/X _4658_/B _3563_/S vssd1 vssd1 vccd1 vccd1 _3351_/X sky130_fd_sc_hd__mux2_1
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3282_ _5818_/A _3555_/B _3282_/C vssd1 vssd1 vccd1 vccd1 _3284_/B sky130_fd_sc_hd__and3_4
X_6070_ _6290_/CLK _6070_/D vssd1 vssd1 vccd1 vccd1 _6070_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5021_ _5046_/B _5021_/B vssd1 vssd1 vccd1 vccd1 _5021_/Y sky130_fd_sc_hd__nand2_1
XFILLER_100_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4683__C1 _4963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3789__A1 _3986_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4986__B1 _4753_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5923_ _5296_/A _5934_/B _5503_/A vssd1 vssd1 vccd1 vccd1 _5923_/X sky130_fd_sc_hd__a21o_1
XANTENNA__4450__A2 _4458_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_724 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5854_ _5854_/A _5854_/B vssd1 vssd1 vccd1 vccd1 _5854_/Y sky130_fd_sc_hd__nand2_1
XFILLER_22_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3866__B _3964_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4805_ _4805_/A _4805_/B vssd1 vssd1 vccd1 vccd1 _4805_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__4738__B1 _4842_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5785_ _6256_/Q _5788_/B vssd1 vssd1 vccd1 vccd1 _5785_/X sky130_fd_sc_hd__or2_1
XFILLER_119_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4736_ _5296_/A _4690_/B _4664_/B _4666_/B _4662_/X vssd1 vssd1 vccd1 vccd1 _4736_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5950__A2 _3867_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4978__A _5547_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4667_ _5263_/A _4666_/Y _4806_/S vssd1 vssd1 vccd1 vccd1 _4667_/X sky130_fd_sc_hd__mux2_1
X_3618_ _3618_/A _3618_/B vssd1 vssd1 vccd1 vccd1 _3619_/C sky130_fd_sc_hd__nand2_1
XANTENNA__4697__B _4697_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5702__A2 _5649_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4598_ _5148_/A _5096_/C _3118_/Y _5625_/C _4597_/Y vssd1 vssd1 vccd1 vccd1 _5062_/A
+ sky130_fd_sc_hd__o41a_1
XFILLER_122_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3549_ _5392_/A _3549_/B vssd1 vssd1 vccd1 vccd1 _3549_/Y sky130_fd_sc_hd__nor2_1
XFILLER_88_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6268_ _6274_/CLK _6268_/D vssd1 vssd1 vccd1 vccd1 _6268_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5219_ _5219_/A _5292_/C vssd1 vssd1 vccd1 vccd1 _5219_/X sky130_fd_sc_hd__and2_1
XFILLER_88_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6199_ _6302_/CLK _6199_/D vssd1 vssd1 vccd1 vccd1 _6199_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__5602__A _6233_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3122__A _3122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4441__A2 _4438_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_22_clk_A _6233_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5483__S _5543_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5154__B1 _5065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_37_clk_A clkbuf_3_4__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4901__B1 _4640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3942__D _3942_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5457__B2 _4646_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3731__S _3731_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5512__A _5512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5209__A1 _5206_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3032__A _4707_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3967__A _5138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4196__A1 _4197_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5570_ _5570_/A _5572_/B vssd1 vssd1 vccd1 vccd1 _5570_/X sky130_fd_sc_hd__or2_1
XANTENNA__4196__B2 _4197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4521_ _5790_/A1 _4520_/X _4521_/S vssd1 vssd1 vccd1 vccd1 _6156_/D sky130_fd_sc_hd__mux2_1
XANTENNA__5145__B1 _3116_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4452_ _6122_/Q _4458_/B vssd1 vssd1 vccd1 vccd1 _4452_/X sky130_fd_sc_hd__or2_1
XFILLER_104_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3403_ _3498_/S _3392_/X _3398_/X _3225_/X _3986_/A vssd1 vssd1 vccd1 vccd1 _3403_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__5696__B2 _3500_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4383_ _4382_/Y _4382_/A _4383_/S vssd1 vssd1 vccd1 vccd1 _4384_/B sky130_fd_sc_hd__mux2_1
XFILLER_113_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3207__A _5054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6122_ _6250_/CLK _6122_/D vssd1 vssd1 vccd1 vccd1 _6122_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3334_ _3387_/A _3599_/A _4010_/B vssd1 vssd1 vccd1 vccd1 _3335_/B sky130_fd_sc_hd__mux2_4
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6053_ _6264_/CLK _6053_/D vssd1 vssd1 vccd1 vccd1 _6053_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3265_ _5818_/A _5622_/A _3259_/X _3263_/Y vssd1 vssd1 vccd1 vccd1 _3266_/B sky130_fd_sc_hd__a31o_4
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4656__C1 _5071_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5004_ _5027_/B _5004_/B vssd1 vssd1 vccd1 vccd1 _5011_/B sky130_fd_sc_hd__or2_1
XFILLER_85_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3554__S0 _4067_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_559 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3196_ _3941_/A _4003_/B _3312_/B vssd1 vssd1 vccd1 vccd1 _3951_/C sky130_fd_sc_hd__or3_4
XFILLER_26_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout173_A _3043_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5509__A_N _5476_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3877__A _5976_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5906_ _5883_/A _5899_/X _5949_/B _5901_/X _5905_/X vssd1 vssd1 vccd1 vccd1 _5908_/A
+ sky130_fd_sc_hd__o311a_1
XANTENNA_fanout340_A input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5837_ _5158_/A _3971_/B _4572_/C _5836_/X _3109_/Y vssd1 vssd1 vccd1 vccd1 _5839_/C
+ sky130_fd_sc_hd__o2111a_1
XFILLER_14_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5768_ _5768_/A0 _6250_/Q _5791_/B vssd1 vssd1 vccd1 vccd1 _5768_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5923__A2 _5934_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4204__C _4309_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3934__A1 _3940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4719_ _6221_/Q _4645_/Y _4718_/X _5463_/A _4963_/A vssd1 vssd1 vccd1 vccd1 _4719_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_30_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5699_ _4767_/A _5714_/B _4587_/B vssd1 vssd1 vccd1 vccd1 _5699_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_30_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3698__A0 _3942_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4895__C1 _4753_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3117__A _3958_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout86_A _3090_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3551__S _3551_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5332__A _5333_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4890__B _4979_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3217__A3 _5464_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3937__D _3937_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_587 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5914__A2 _5075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5507__A _5507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5678__A1 _4734_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5226__B _5454_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3689__A0 _5292_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3027__A _5054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3050_ _3107_/A _3050_/B vssd1 vssd1 vccd1 vccd1 _3050_/X sky130_fd_sc_hd__or2_2
XFILLER_83_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_476 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3952_ _4587_/B _3952_/B _4604_/C _4614_/B vssd1 vssd1 vccd1 vccd1 _3955_/D sky130_fd_sc_hd__or4bb_1
XFILLER_32_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3883_ _3883_/A _3975_/C vssd1 vssd1 vccd1 vccd1 _3883_/X sky130_fd_sc_hd__or2_4
XFILLER_31_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5622_ _5622_/A _5622_/B vssd1 vssd1 vccd1 vccd1 _5644_/C sky130_fd_sc_hd__nand2_1
XANTENNA__5905__A2 _4010_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3916__A1 _3715_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5553_ _3432_/A _5442_/A _5542_/X _5943_/C _5550_/X vssd1 vssd1 vccd1 vccd1 _5553_/X
+ sky130_fd_sc_hd__o221a_1
X_4504_ _4672_/A _6150_/Q _4520_/S vssd1 vssd1 vccd1 vccd1 _4504_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3863__C _4594_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5484_ _4645_/B _5482_/Y _5483_/X _4646_/A _5227_/A vssd1 vssd1 vccd1 vccd1 _5484_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_117_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5669__A1 _6293_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_478 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4435_ _4410_/B _4410_/D _4428_/B vssd1 vssd1 vccd1 vccd1 _4435_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_99_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4341__A1 _4426_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4341__B2 _4410_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4366_ _4410_/B _4389_/B _4366_/C vssd1 vssd1 vccd1 vccd1 _4393_/B sky130_fd_sc_hd__and3_2
X_6105_ _6143_/CLK _6105_/D vssd1 vssd1 vccd1 vccd1 _6105_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4467__S _4477_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3317_ _4003_/B _4003_/C vssd1 vssd1 vccd1 vccd1 _3621_/A sky130_fd_sc_hd__nand2_4
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4297_ _4437_/A1 _4293_/X _4296_/Y _6109_/Q vssd1 vssd1 vccd1 vccd1 _4297_/Y sky130_fd_sc_hd__a22oi_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6036_ _6278_/CLK _6036_/D vssd1 vssd1 vccd1 vccd1 _6036_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3248_ _6258_/Q _5439_/A2 _5924_/B _6027_/Q vssd1 vssd1 vccd1 vccd1 _3248_/X sky130_fd_sc_hd__o22a_1
XFILLER_132_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5841__A1 _3251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3179_ _6071_/Q _4577_/C vssd1 vssd1 vccd1 vccd1 _3179_/X sky130_fd_sc_hd__or2_4
XTAP_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3400__A _3500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4332__B2 _4437_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5832__A1 _3631_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4635__A2 _4744_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3843__B1 _3590_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5596__B1 _5251_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5348__B1 _5742_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3964__B _3964_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5899__A1 _5900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4141__A _4202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4571__A1 _3974_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4220_ _4221_/A _4221_/B _4221_/C vssd1 vssd1 vccd1 vccd1 _4220_/X sky130_fd_sc_hd__and3_2
XFILLER_96_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4151_ _4152_/A _4152_/B vssd1 vssd1 vccd1 vccd1 _4151_/Y sky130_fd_sc_hd__nand2_2
XFILLER_122_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3102_ _5090_/A _4638_/B vssd1 vssd1 vccd1 vccd1 _3102_/Y sky130_fd_sc_hd__nor2_4
XFILLER_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4082_ _4162_/B _4176_/B vssd1 vssd1 vccd1 vccd1 _4084_/B sky130_fd_sc_hd__nand2_2
XFILLER_83_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5823__A1 _3375_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4626__A2 _4659_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3033_ _5344_/A vssd1 vssd1 vccd1 vccd1 _3033_/Y sky130_fd_sc_hd__inv_8
XFILLER_95_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4984_ _4988_/A _4983_/X _4981_/A vssd1 vssd1 vccd1 vccd1 _4984_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_63_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3935_ _5241_/A _3935_/B _3935_/C _3935_/D vssd1 vssd1 vccd1 vccd1 _3935_/X sky130_fd_sc_hd__or4_1
XANTENNA__4035__B _5925_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout136_A _4638_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3866_ _4577_/C _3964_/B vssd1 vssd1 vccd1 vccd1 _5911_/B sky130_fd_sc_hd__nand2_4
XFILLER_137_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5605_ _6009_/Q _5605_/B _5605_/C vssd1 vssd1 vccd1 vccd1 _5605_/X sky130_fd_sc_hd__and3_1
XANTENNA__4011__B1 _3593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3797_ _6036_/Q _3771_/X _3795_/Y _3796_/X vssd1 vssd1 vccd1 vccd1 _6036_/D sky130_fd_sc_hd__a211o_1
XANTENNA__3366__S _3658_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5147__A _5543_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3593__C _3594_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5536_ _6005_/Q _5537_/B _6006_/Q vssd1 vssd1 vccd1 vccd1 _5536_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_127_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5467_ _6124_/Q _3901_/B _3704_/B _6026_/Q _5466_/X vssd1 vssd1 vccd1 vccd1 _5467_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__3890__A _5138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4418_ _4419_/A _4419_/B _4419_/C vssd1 vssd1 vccd1 vccd1 _4431_/B sky130_fd_sc_hd__o21ai_2
X_5398_ _4819_/B _5509_/C _5360_/S _6008_/Q _4646_/A vssd1 vssd1 vccd1 vccd1 _5398_/X
+ sky130_fd_sc_hd__a221o_1
Xfanout301 _4642_/A vssd1 vssd1 vccd1 vccd1 _5218_/B sky130_fd_sc_hd__buf_6
Xfanout312 _3029_/Y vssd1 vssd1 vccd1 vccd1 _5561_/S sky130_fd_sc_hd__buf_8
XFILLER_99_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout323 input9/X vssd1 vssd1 vccd1 vccd1 _5986_/B1 sky130_fd_sc_hd__buf_2
XFILLER_132_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout334 _4846_/A vssd1 vssd1 vccd1 vccd1 _5428_/A sky130_fd_sc_hd__buf_8
XFILLER_87_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4349_ _4310_/A _4343_/A _4313_/A vssd1 vssd1 vccd1 vccd1 _4350_/B sky130_fd_sc_hd__o21ba_2
Xfanout345 _4657_/A vssd1 vssd1 vccd1 vccd1 _5263_/A sky130_fd_sc_hd__buf_8
XFILLER_98_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5814__A1 _3631_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6019_ _6293_/CLK _6019_/D vssd1 vssd1 vccd1 vccd1 _6019_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout49_A _5766_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5042__A2 _4640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3589__C1 _5470_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_619 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4002__B1 _3987_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5057__A _5136_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4896__A _5509_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3950__D _4586_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5281__A2 _3901_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3678__C _3678_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4136__A _4136_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3040__A _6004_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5019__A1_N _4963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3975__A _5976_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3720_ _4112_/C _5743_/C _3708_/Y _6230_/Q vssd1 vssd1 vccd1 vccd1 _3720_/X sky130_fd_sc_hd__o22a_1
Xclkbuf_leaf_40_clk clkbuf_3_4__f_clk/X vssd1 vssd1 vccd1 vccd1 _6250_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_13_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3651_ _3651_/A _3651_/B vssd1 vssd1 vccd1 vccd1 _3923_/B sky130_fd_sc_hd__nand2_2
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3582_ _3580_/X _3581_/X _3422_/A _3935_/D vssd1 vssd1 vccd1 vccd1 _5888_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_127_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5321_ _5929_/B2 _5319_/X _5320_/X _5318_/X vssd1 vssd1 vccd1 vccd1 _5321_/X sky130_fd_sc_hd__a31o_4
XFILLER_6_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5252_ _5256_/B _5237_/X _5513_/A vssd1 vssd1 vccd1 vccd1 _5252_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4203_ _4334_/A _4309_/B _4342_/B _4162_/A vssd1 vssd1 vccd1 vccd1 _4205_/A sky130_fd_sc_hd__a22oi_4
XFILLER_102_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5183_ _5054_/A _5143_/B _4946_/A vssd1 vssd1 vccd1 vccd1 _5183_/X sky130_fd_sc_hd__o21a_1
XANTENNA__3215__A _3940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4134_ _4135_/B _4135_/C _4135_/A vssd1 vssd1 vccd1 vccd1 _4138_/A sky130_fd_sc_hd__a21o_1
XFILLER_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_451 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4065_ _6077_/Q _3727_/X _4066_/S vssd1 vssd1 vccd1 vccd1 _6077_/D sky130_fd_sc_hd__mux2_1
XFILLER_113_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3869__B _3869_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3016_ _5258_/A vssd1 vssd1 vccd1 vccd1 _5131_/A sky130_fd_sc_hd__inv_2
XFILLER_37_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout253_A _6238_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4967_ _6193_/Q _5561_/S _5239_/A _4966_/X vssd1 vssd1 vccd1 vccd1 _4967_/X sky130_fd_sc_hd__a211o_1
XANTENNA__4232__B1 _4072_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3885__A _3885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3918_ _6053_/Q _3721_/X _3921_/S vssd1 vssd1 vccd1 vccd1 _6053_/D sky130_fd_sc_hd__mux2_1
XANTENNA__3586__A2 _5439_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_31_clk clkbuf_3_5__f_clk/X vssd1 vssd1 vccd1 vccd1 _6170_/CLK sky130_fd_sc_hd__clkbuf_16
X_4898_ _5480_/B _4644_/Y _4896_/Y _4897_/X vssd1 vssd1 vccd1 vccd1 _4898_/X sky130_fd_sc_hd__o22a_1
X_3849_ _3944_/A _3849_/B vssd1 vssd1 vccd1 vccd1 _3849_/Y sky130_fd_sc_hd__nand2_1
XFILLER_138_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5519_ _6005_/Q _5537_/B vssd1 vssd1 vccd1 vccd1 _5519_/Y sky130_fd_sc_hd__nor2_1
XFILLER_106_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5605__A _6009_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5496__C1 _5556_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout120 _3274_/X vssd1 vssd1 vccd1 vccd1 _3388_/B sky130_fd_sc_hd__buf_12
XFILLER_59_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout131 _3093_/Y vssd1 vssd1 vccd1 vccd1 _4744_/B sky130_fd_sc_hd__buf_8
Xfanout142 _3078_/Y vssd1 vssd1 vccd1 vccd1 _5131_/B sky130_fd_sc_hd__buf_4
XFILLER_59_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout153 _3069_/Y vssd1 vssd1 vccd1 vccd1 _5509_/C sky130_fd_sc_hd__buf_12
XFILLER_75_803 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout164 _5349_/B1 vssd1 vssd1 vccd1 vccd1 _4058_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout175 _3713_/X vssd1 vssd1 vccd1 vccd1 _4214_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_47_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout186 _4111_/B vssd1 vssd1 vccd1 vccd1 _4311_/B sky130_fd_sc_hd__buf_6
Xfanout197 _3172_/X vssd1 vssd1 vccd1 vccd1 _5617_/B sky130_fd_sc_hd__buf_4
XFILLER_47_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5340__A _5344_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4471__A0 _5856_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3577__A2 _3567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_22_clk _6233_/CLK vssd1 vssd1 vccd1 vccd1 _6079_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_11_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5723__B1 _5442_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3501__A2 _3500_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3265__A1 _5818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5870_ _5870_/A _5870_/B _3975_/C vssd1 vssd1 vccd1 vccd1 _5871_/D sky130_fd_sc_hd__or3b_1
XFILLER_73_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4821_ _5358_/A _5367_/A _4783_/Y vssd1 vssd1 vccd1 vccd1 _4822_/B sky130_fd_sc_hd__a21o_1
XTAP_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4752_ _4750_/A _4750_/B _4755_/A _4751_/X vssd1 vssd1 vccd1 vccd1 _4753_/C sky130_fd_sc_hd__a31o_1
XFILLER_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4765__A1 _4625_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3703_ _5742_/A _3704_/B _5767_/C vssd1 vssd1 vccd1 vccd1 _5763_/B sky130_fd_sc_hd__nor3_4
X_4683_ _4672_/A _4645_/Y _4682_/X _5463_/A _4963_/A vssd1 vssd1 vccd1 vccd1 _4683_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_119_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4517__A1 _3942_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3634_ _3387_/A _3594_/A _3594_/B _3599_/X vssd1 vssd1 vccd1 vccd1 _3635_/B sky130_fd_sc_hd__a31o_2
XFILLER_134_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5190__A1 _5191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3565_ _6206_/Q _3567_/B vssd1 vssd1 vccd1 vccd1 _3618_/A sky130_fd_sc_hd__nand2_2
XANTENNA__5425__A _5428_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5304_ _5305_/A _5305_/B vssd1 vssd1 vccd1 vccd1 _5333_/B sky130_fd_sc_hd__nor2_1
X_6284_ _6284_/CLK _6284_/D vssd1 vssd1 vccd1 vccd1 _6284_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3496_ _4767_/A _3636_/A _3211_/Y vssd1 vssd1 vccd1 vccd1 _3496_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_130_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5235_ _5232_/X _5233_/X _5234_/X _5929_/B2 vssd1 vssd1 vccd1 vccd1 _5236_/A sky130_fd_sc_hd__a22oi_4
XFILLER_130_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5493__A2 _5442_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5166_ _5164_/Y _5166_/B vssd1 vssd1 vccd1 vccd1 _5166_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_29_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4117_ _4117_/A _4117_/B vssd1 vssd1 vccd1 vccd1 _4121_/A sky130_fd_sc_hd__xnor2_1
XFILLER_29_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5097_ _5097_/A _5097_/B _5095_/X vssd1 vssd1 vccd1 vccd1 _5097_/X sky130_fd_sc_hd__or3b_4
XANTENNA__5245__A2 _5244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4048_ _5733_/A _5096_/C _4051_/S vssd1 vssd1 vccd1 vccd1 _4048_/Y sky130_fd_sc_hd__nor3_1
XFILLER_84_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5999_ _6145_/Q vssd1 vssd1 vccd1 vccd1 _6145_/D sky130_fd_sc_hd__clkbuf_2
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3559__A2 _3443_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4508__A1 _5926_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5181__A1 _5136_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4596__D _4596_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5484__A2 _5482_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3247__A1 _3236_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4444__B1 _3900_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3302__B _3952_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4995__A1 _5547_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5944__B1 _5934_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4133__B _4197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3972__B _5124_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3350_ _3353_/A _3350_/B vssd1 vssd1 vccd1 vccd1 _4658_/B sky130_fd_sc_hd__xnor2_4
XFILLER_98_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3281_ _6272_/Q _6018_/Q _6086_/Q _6041_/Q _4067_/A _3709_/S vssd1 vssd1 vccd1 vccd1
+ _3282_/C sky130_fd_sc_hd__mux4_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5020_ _5547_/A _4872_/B _5019_/X _5069_/A vssd1 vssd1 vccd1 vccd1 _5021_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5922_ _5296_/A _4586_/Y _5921_/X vssd1 vssd1 vccd1 vccd1 _5931_/S sky130_fd_sc_hd__o21a_1
XFILLER_80_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5853_ _5853_/A vssd1 vssd1 vccd1 vccd1 _5854_/B sky130_fd_sc_hd__inv_2
XFILLER_110_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5935__A0 _5935_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4804_ _4840_/A _4804_/B vssd1 vssd1 vccd1 vccd1 _4805_/B sky130_fd_sc_hd__nand2_1
XFILLER_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5784_ _3942_/B _4250_/Y _5782_/X _5783_/X vssd1 vssd1 vccd1 vccd1 _6255_/D sky130_fd_sc_hd__a22o_1
XFILLER_21_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3946__C1 _5124_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4735_ _4735_/A _4735_/B vssd1 vssd1 vccd1 vccd1 _4735_/Y sky130_fd_sc_hd__nor2_1
X_4666_ _4666_/A _4666_/B vssd1 vssd1 vccd1 vccd1 _4666_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_119_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4978__B _4979_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout216_A _3024_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3882__B _3975_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3617_ _3652_/A _3617_/B vssd1 vssd1 vccd1 vccd1 _3923_/A sky130_fd_sc_hd__nand2_2
X_4597_ _5221_/B _4623_/A vssd1 vssd1 vccd1 vccd1 _4597_/Y sky130_fd_sc_hd__nand2_1
X_3548_ _3567_/B _3548_/B vssd1 vssd1 vccd1 vccd1 _5706_/B sky130_fd_sc_hd__xnor2_4
XFILLER_115_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4091__A1_N _3795_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6267_ _6274_/CLK _6267_/D vssd1 vssd1 vccd1 vccd1 _6267_/Q sky130_fd_sc_hd__dfxtp_1
X_3479_ _6014_/Q _3231_/Y _3478_/X vssd1 vssd1 vccd1 vccd1 _6014_/D sky130_fd_sc_hd__o21a_1
XFILLER_131_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5466__A2 _3243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5218_ _5255_/B _5218_/B vssd1 vssd1 vccd1 vccd1 _5292_/C sky130_fd_sc_hd__or2_2
XFILLER_130_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6198_ _6217_/CLK _6198_/D vssd1 vssd1 vccd1 vccd1 _6198_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_56_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5149_ _4589_/Y _5147_/X _5148_/Y _5142_/Y _3958_/A vssd1 vssd1 vccd1 vccd1 _5149_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_56_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3122__B _5498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4977__A1 _4745_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4977__B2 _4744_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4234__A _5436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5926__A0 _5926_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5049__B _5051_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5065__A _5065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4901__A1 _5041_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3468__A1 _3458_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5512__B _5512_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3313__A _3974_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4968__A1 _5051_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3967__B _5943_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5917__B1 _5172_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4144__A _4163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4196__A2 _3280_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4520_ _4891_/A _6156_/Q _4520_/S vssd1 vssd1 vccd1 vccd1 _4520_/X sky130_fd_sc_hd__mux2_1
X_4451_ _5856_/A _3900_/Y _4449_/X _4450_/Y vssd1 vssd1 vccd1 vccd1 _6121_/D sky130_fd_sc_hd__a22o_1
XANTENNA__5145__A1 _5561_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3402_ _3644_/B _3500_/A _3401_/X vssd1 vssd1 vccd1 vccd1 _4697_/B sky130_fd_sc_hd__o21a_4
XANTENNA__5550__D1 _5607_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4382_ _4382_/A _4382_/B vssd1 vssd1 vccd1 vccd1 _4382_/Y sky130_fd_sc_hd__nor2_1
XFILLER_125_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6121_ _6254_/CLK _6121_/D vssd1 vssd1 vccd1 vccd1 _6121_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3333_ _3677_/B _3881_/B vssd1 vssd1 vccd1 vccd1 _3599_/A sky130_fd_sc_hd__nor2_8
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3922__S _3922_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5703__A _5703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6052_ _6259_/CLK _6052_/D vssd1 vssd1 vccd1 vccd1 _6052_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_18 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3264_ _5818_/A _5622_/A _3259_/X _3263_/Y vssd1 vssd1 vccd1 vccd1 _3267_/B sky130_fd_sc_hd__a31oi_4
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5003_ _6194_/Q _5002_/C _6195_/Q vssd1 vssd1 vccd1 vccd1 _5004_/B sky130_fd_sc_hd__a21oi_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3195_ _3960_/C _3893_/B vssd1 vssd1 vccd1 vccd1 _3195_/X sky130_fd_sc_hd__or2_2
XANTENNA__3223__A _3706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout166_A _5349_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5081__B1 _4642_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5905_ _3867_/A _4010_/B _5903_/Y _5904_/Y _5065_/A vssd1 vssd1 vccd1 vccd1 _5905_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_22_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout333_A _4846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5836_ _5165_/B _3974_/C _5638_/B _5638_/C vssd1 vssd1 vccd1 vccd1 _5836_/X sky130_fd_sc_hd__o211a_1
XFILLER_14_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5767_ _5767_/A _5767_/B _5767_/C vssd1 vssd1 vccd1 vccd1 _5791_/B sky130_fd_sc_hd__or3_4
XANTENNA__3893__A _5124_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4204__D _4342_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4718_ _4646_/Y _4716_/Y _4717_/X _4715_/X vssd1 vssd1 vccd1 vccd1 _4718_/X sky130_fd_sc_hd__a31o_1
X_5698_ _5714_/B _5698_/B vssd1 vssd1 vccd1 vccd1 _5698_/X sky130_fd_sc_hd__or2_1
XFILLER_108_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4649_ _5054_/A _5509_/C vssd1 vssd1 vccd1 vccd1 _5172_/B sky130_fd_sc_hd__nand2_8
XFILLER_30_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5316__C _5436_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3117__B _4654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5439__A2 _5439_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout79_A _3115_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5375__A1 _3122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5226__C _5264_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3043__A _3880_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3978__A _4643_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3951_ _4022_/C _5635_/A _3951_/C vssd1 vssd1 vccd1 vccd1 _4615_/B sky130_fd_sc_hd__nor3_4
XFILLER_91_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3882_ _3883_/A _3975_/C vssd1 vssd1 vccd1 vccd1 _4023_/A sky130_fd_sc_hd__nor2_2
X_5621_ _4614_/A _3950_/C _3736_/A vssd1 vssd1 vccd1 vccd1 _5622_/B sky130_fd_sc_hd__o21ai_1
XFILLER_31_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3917__S _3921_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5552_ _5551_/A _5542_/X _5551_/Y _3122_/A vssd1 vssd1 vccd1 vccd1 _5552_/X sky130_fd_sc_hd__a211o_1
XFILLER_129_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4503_ _3943_/C _4502_/X _4521_/S vssd1 vssd1 vccd1 vccd1 _6149_/D sky130_fd_sc_hd__mux2_1
XFILLER_8_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5483_ _4633_/B _6003_/Q _5543_/S vssd1 vssd1 vccd1 vccd1 _5483_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3129__A0 _4657_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5669__A2 _4615_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4434_ _3853_/X _4296_/B _4296_/Y _6116_/Q vssd1 vssd1 vccd1 vccd1 _4434_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5136__C _5136_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4365_ _4363_/A _4388_/A _4364_/X vssd1 vssd1 vccd1 vccd1 _4366_/C sky130_fd_sc_hd__o21a_1
XANTENNA__4341__A2 _4309_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6104_ _6143_/CLK _6104_/D vssd1 vssd1 vccd1 vccd1 _6104_/Q sky130_fd_sc_hd__dfxtp_1
X_3316_ _3316_/A _3316_/B vssd1 vssd1 vccd1 vccd1 _3316_/Y sky130_fd_sc_hd__nand2_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4296_ _4296_/A _4296_/B vssd1 vssd1 vccd1 vccd1 _4296_/Y sky130_fd_sc_hd__nor2_4
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4629__B1 _5226_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6035_ _6265_/CLK _6035_/D vssd1 vssd1 vccd1 vccd1 _6035_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_112_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3247_ _3236_/Y _3238_/X _5743_/B _6072_/Q _3244_/X vssd1 vssd1 vccd1 vccd1 _3247_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout283_A _6222_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_21_clk_A _6084_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3178_ _3970_/A _4577_/C vssd1 vssd1 vccd1 vccd1 _5714_/B sky130_fd_sc_hd__nor2_4
XANTENNA__3852__A1 _4877_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_36_clk_A clkbuf_3_4__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3400__B _3500_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5357__A1 _5333_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5819_ _5819_/A _5819_/B vssd1 vssd1 vccd1 vccd1 _5819_/Y sky130_fd_sc_hd__nor2_8
XANTENNA__3368__B1 _3881_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4868__A0 _6190_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5293__B1 _6221_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3843__A1 _4214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5596__A1 _5595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4141__B _4173_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3980__B _3980_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4150_ _4150_/A _4150_/B vssd1 vssd1 vccd1 vccd1 _4152_/B sky130_fd_sc_hd__xnor2_4
X_3101_ _3101_/A _5096_/B vssd1 vssd1 vccd1 vccd1 _4592_/A sky130_fd_sc_hd__or2_1
XFILLER_96_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4081_ _4162_/B _4173_/B _4176_/B _4096_/A vssd1 vssd1 vccd1 vccd1 _4085_/C sky130_fd_sc_hd__a22o_1
XFILLER_55_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3032_ _4707_/B vssd1 vssd1 vccd1 vccd1 _3032_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_83_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5587__A1 _5512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4983_ _4983_/A _4987_/B vssd1 vssd1 vccd1 vccd1 _4983_/X sky130_fd_sc_hd__or2_2
X_3934_ _3940_/A _3933_/X _5241_/A vssd1 vssd1 vccd1 vccd1 _3934_/X sky130_fd_sc_hd__a21o_1
XANTENNA__5339__A1 _4644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5339__B2 _5464_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3865_ _4604_/B _5928_/B vssd1 vssd1 vccd1 vccd1 _3865_/Y sky130_fd_sc_hd__nor2_1
XFILLER_31_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5428__A _5428_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5604_ _4638_/B _5603_/X _5601_/X _3060_/B vssd1 vssd1 vccd1 vccd1 _5604_/X sky130_fd_sc_hd__a211o_1
XANTENNA__4011__A1 _3033_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3796_ _4270_/A _3832_/A2 _3382_/X _3765_/X _3772_/X vssd1 vssd1 vccd1 vccd1 _3796_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__4011__B2 _5714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout129_A _3111_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5147__B _5158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5535_ _5540_/B _5251_/A _5534_/X _5948_/A vssd1 vssd1 vccd1 vccd1 _6229_/D sky130_fd_sc_hd__o211a_1
XFILLER_118_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3770__B1 _3250_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5466_ _6257_/Q _3243_/A _5742_/B _6249_/Q vssd1 vssd1 vccd1 vccd1 _5466_/X sky130_fd_sc_hd__o22a_1
X_4417_ _4417_/A _4417_/B vssd1 vssd1 vccd1 vccd1 _4419_/C sky130_fd_sc_hd__xnor2_1
XFILLER_105_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5397_ _5385_/A _4829_/Y _5539_/S vssd1 vssd1 vccd1 vccd1 _5397_/X sky130_fd_sc_hd__mux2_1
Xfanout302 _4642_/A vssd1 vssd1 vccd1 vccd1 _3880_/A sky130_fd_sc_hd__buf_8
Xfanout313 _5556_/C1 vssd1 vssd1 vccd1 vccd1 _5866_/B1 sky130_fd_sc_hd__buf_4
Xfanout324 _5932_/A vssd1 vssd1 vccd1 vccd1 _4540_/A sky130_fd_sc_hd__buf_4
X_4348_ _4348_/A _4348_/B vssd1 vssd1 vccd1 vccd1 _4350_/A sky130_fd_sc_hd__nor2_1
XFILLER_86_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout335 input7/X vssd1 vssd1 vccd1 vccd1 _4846_/A sky130_fd_sc_hd__clkbuf_16
Xfanout346 input2/X vssd1 vssd1 vccd1 vccd1 _4657_/A sky130_fd_sc_hd__buf_12
XFILLER_113_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input3_A io_in[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4279_ _4209_/B _4209_/C _4209_/A vssd1 vssd1 vccd1 vccd1 _4281_/B sky130_fd_sc_hd__a21boi_4
XFILLER_87_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6018_ _6041_/CLK _6018_/D vssd1 vssd1 vccd1 vccd1 _6018_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3825__A1 _3513_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3589__B1 _3589_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4002__B2 _5712_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5057__B _5638_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5750__A1 _5305_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5502__A1 _3060_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5502__B2 _4644_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5266__B1 _5653_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_786 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5569__A1 _4638_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4136__B _4167_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4241__A1 _3715_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3975__B _5870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3467__S _3575_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3650_ _3651_/A _3651_/B vssd1 vssd1 vccd1 vccd1 _3931_/B sky130_fd_sc_hd__and2_2
XANTENNA__5741__A1 _4216_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3581_ _3145_/C _3618_/A _3422_/A vssd1 vssd1 vccd1 vccd1 _3581_/X sky130_fd_sc_hd__a21o_1
XFILLER_127_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5320_ _6252_/Q _3243_/A _3239_/X _6119_/Q vssd1 vssd1 vccd1 vccd1 _5320_/X sky130_fd_sc_hd__o22a_1
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5251_ _5251_/A vssd1 vssd1 vccd1 vccd1 _5251_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_114_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4202_ _4202_/A _4311_/B vssd1 vssd1 vccd1 vccd1 _4207_/A sky130_fd_sc_hd__nand2_2
XFILLER_69_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5182_ _5143_/B _5617_/A _5180_/X _5731_/S vssd1 vssd1 vccd1 vccd1 _5182_/X sky130_fd_sc_hd__o211a_1
X_4133_ _4162_/B _4197_/A _4309_/B _4342_/B vssd1 vssd1 vccd1 vccd1 _4135_/C sky130_fd_sc_hd__nand4_2
XFILLER_95_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4064_ _6076_/Q _3724_/X _4066_/S vssd1 vssd1 vccd1 vccd1 _6076_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3015_ _6217_/Q vssd1 vssd1 vccd1 vccd1 _3170_/A sky130_fd_sc_hd__inv_6
XANTENNA__4480__A1 _3943_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3231__A _5799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4046__B _5075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4966_ _4990_/A _4965_/Y _4640_/A _4638_/B vssd1 vssd1 vccd1 vccd1 _4966_/X sky130_fd_sc_hd__a211o_1
XANTENNA__4232__A1 _3853_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3885__B _3975_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3917_ _6052_/Q _3718_/X _3921_/S vssd1 vssd1 vccd1 vccd1 _6052_/D sky130_fd_sc_hd__mux2_1
X_4897_ _6191_/Q _4647_/B _4648_/Y _5072_/A _4826_/Y vssd1 vssd1 vccd1 vccd1 _4897_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_22_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5158__A _5158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3848_ _3594_/B _3746_/A _3847_/X _3849_/B vssd1 vssd1 vccd1 vccd1 _3848_/X sky130_fd_sc_hd__a211o_1
XFILLER_137_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3779_ _3751_/A _3777_/X _3778_/X vssd1 vssd1 vccd1 vccd1 _3779_/X sky130_fd_sc_hd__a21o_1
X_5518_ _6228_/Q _5251_/A _5513_/Y _5517_/X _5948_/A vssd1 vssd1 vccd1 vccd1 _6228_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_3_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5605__B _5605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5449_ _5599_/B _5450_/B vssd1 vssd1 vccd1 vccd1 _5451_/A sky130_fd_sc_hd__nand2_1
Xfanout110 _3443_/Y vssd1 vssd1 vccd1 vccd1 _5707_/B sky130_fd_sc_hd__buf_12
Xfanout121 _3450_/A vssd1 vssd1 vccd1 vccd1 _3388_/A sky130_fd_sc_hd__buf_12
Xfanout132 _3084_/X vssd1 vssd1 vccd1 vccd1 _4643_/A sky130_fd_sc_hd__buf_12
Xfanout143 _5625_/B vssd1 vssd1 vccd1 vccd1 _5227_/B sky130_fd_sc_hd__buf_6
Xfanout154 _3069_/Y vssd1 vssd1 vccd1 vccd1 _5238_/C sky130_fd_sc_hd__clkbuf_4
Xfanout165 _3704_/B vssd1 vssd1 vccd1 vccd1 _3589_/B1 sky130_fd_sc_hd__buf_6
XFILLER_47_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout176 _4216_/B vssd1 vssd1 vccd1 vccd1 _4173_/B sky130_fd_sc_hd__buf_6
XFILLER_19_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout187 _3337_/X vssd1 vssd1 vccd1 vccd1 _4111_/B sky130_fd_sc_hd__buf_6
XFILLER_86_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout198 _3922_/S vssd1 vssd1 vccd1 vccd1 _5635_/A sky130_fd_sc_hd__buf_8
XFILLER_75_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5340__B _5341_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4237__A _5742_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3795__B _3795_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5723__A1 _5710_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5723__B2 _5734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3501__A3 _3458_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3265__A2 _5622_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3986__A _3986_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4820_ _4860_/B _4820_/B vssd1 vssd1 vccd1 vccd1 _4925_/A sky130_fd_sc_hd__nand2_4
XTAP_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4751_ _4782_/A _4791_/A _4782_/B _3116_/X vssd1 vssd1 vccd1 vccd1 _4751_/X sky130_fd_sc_hd__a31o_1
XANTENNA__4765__A2 _5093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5962__A1 _5934_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3702_ _5790_/A1 _3701_/X _3705_/A vssd1 vssd1 vccd1 vccd1 _6026_/D sky130_fd_sc_hd__mux2_1
XFILLER_119_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4682_ _3122_/Y _4679_/X _4681_/X _4646_/Y vssd1 vssd1 vccd1 vccd1 _4682_/X sky130_fd_sc_hd__a22o_1
XFILLER_135_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3633_ _4216_/A _3765_/B _3255_/Y _3592_/A vssd1 vssd1 vccd1 vccd1 _3633_/X sky130_fd_sc_hd__a31o_1
XFILLER_128_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5706__A _5733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3564_ _5703_/B _3563_/X _3564_/S vssd1 vssd1 vccd1 vccd1 _3564_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5425__B _5653_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5303_ _4707_/B _6005_/Q _5360_/S vssd1 vssd1 vccd1 vccd1 _5303_/X sky130_fd_sc_hd__mux2_1
X_6283_ _6284_/CLK _6283_/D vssd1 vssd1 vccd1 vccd1 _6283_/Q sky130_fd_sc_hd__dfxtp_1
X_3495_ _3495_/A _3495_/B vssd1 vssd1 vccd1 vccd1 _3495_/X sky130_fd_sc_hd__or2_1
XANTENNA__3226__A _4946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5234_ _6250_/Q _6117_/Q _6019_/Q _6242_/Q _3241_/A _3241_/B vssd1 vssd1 vccd1 vccd1
+ _5234_/X sky130_fd_sc_hd__mux4_2
XFILLER_115_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4756__S _5041_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5165_ _5635_/A _5165_/B _5634_/B _5634_/D vssd1 vssd1 vccd1 vccd1 _5166_/B sky130_fd_sc_hd__or4_2
XFILLER_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout196_A _5617_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4116_ _4117_/A _4117_/B vssd1 vssd1 vccd1 vccd1 _4150_/A sky130_fd_sc_hd__nand2b_4
XFILLER_111_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5096_ _5148_/A _5096_/B _5096_/C vssd1 vssd1 vccd1 vccd1 _5097_/B sky130_fd_sc_hd__or3_1
XFILLER_84_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5245__A3 _4648_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4047_ _4596_/B _4462_/A vssd1 vssd1 vccd1 vccd1 _5869_/S sky130_fd_sc_hd__nor2_4
XANTENNA__4057__A _5436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4453__A1 _5387_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3256__A2 _3250_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5998_ _6144_/Q vssd1 vssd1 vccd1 vccd1 _6144_/D sky130_fd_sc_hd__clkbuf_2
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5953__A1 _5883_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4949_ _4943_/A _4910_/B _4943_/B vssd1 vssd1 vccd1 vccd1 _4949_/X sky130_fd_sc_hd__o21a_1
XFILLER_137_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5705__A1 _5730_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5469__B1 _5767_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3136__A _4067_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4444__A1 _5305_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4995__A2 _4644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5497__S _5539_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5944__A1 _3869_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4133__C _4309_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3280_ _6018_/Q _6041_/Q _3709_/S vssd1 vssd1 vccd1 vccd1 _3280_/X sky130_fd_sc_hd__mux2_8
XFILLER_97_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4132__B1 _4112_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4683__A1 _4672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5261__A _5263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4683__B2 _5463_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5880__B1 _3883_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4435__A1 _4410_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5921_ _5921_/A _5921_/B _5921_/C vssd1 vssd1 vccd1 vccd1 _5921_/X sky130_fd_sc_hd__and3_4
XFILLER_0_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5852_ _3500_/C _3942_/D _5862_/B vssd1 vssd1 vccd1 vccd1 _5853_/A sky130_fd_sc_hd__mux2_8
XFILLER_62_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4605__A _4605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4803_ _5392_/A _5703_/B vssd1 vssd1 vccd1 vccd1 _4804_/B sky130_fd_sc_hd__nand2_1
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5783_ _5387_/A _5791_/B _5769_/S vssd1 vssd1 vccd1 vccd1 _5783_/X sky130_fd_sc_hd__o21a_1
X_4734_ _5114_/A _4734_/B vssd1 vssd1 vccd1 vccd1 _4735_/B sky130_fd_sc_hd__and2_1
XFILLER_119_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4665_ _5264_/A _4665_/B vssd1 vssd1 vccd1 vccd1 _4666_/B sky130_fd_sc_hd__and2_1
XFILLER_135_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5436__A _5436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5699__B1 _4587_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout111_A _3458_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3616_ _3652_/A _3617_/B vssd1 vssd1 vccd1 vccd1 _3619_/B sky130_fd_sc_hd__and2_1
X_4596_ _5244_/A _4596_/B _5069_/A _4596_/D vssd1 vssd1 vccd1 vccd1 _4623_/A sky130_fd_sc_hd__and4_2
XANTENNA_fanout209_A _3053_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3547_ _3387_/A _3593_/B _3546_/X vssd1 vssd1 vccd1 vccd1 _3548_/B sky130_fd_sc_hd__a21o_2
XFILLER_88_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3478_ _3631_/A _3477_/Y _3433_/X _3592_/A vssd1 vssd1 vccd1 vccd1 _3478_/X sky130_fd_sc_hd__a211o_1
X_6266_ _6272_/CLK _6266_/D vssd1 vssd1 vccd1 vccd1 _6266_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5217_ _5217_/A _5217_/B vssd1 vssd1 vccd1 vccd1 _5217_/Y sky130_fd_sc_hd__nor2_1
XFILLER_131_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3477__A2 _5677_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6197_ _6290_/CLK _6197_/D vssd1 vssd1 vccd1 vccd1 _6197_/Q sky130_fd_sc_hd__dfxtp_2
X_5148_ _5148_/A _5241_/B vssd1 vssd1 vccd1 vccd1 _5148_/Y sky130_fd_sc_hd__nand2_1
XFILLER_111_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5079_ _5079_/A _5079_/B _5919_/A vssd1 vssd1 vccd1 vccd1 _5080_/B sky130_fd_sc_hd__or3b_2
XFILLER_72_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4831__D1 _4644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4234__B _4234_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4250__A _5743_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5154__A2 _5909_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4901__A2 _4900_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3313__B _4003_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_829 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4425__A _4426_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3640__A2 _3594_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5917__A1 _4577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4144__B _4176_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5256__A _5292_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4450_ _3010_/Y _4458_/B _3900_/Y vssd1 vssd1 vccd1 vccd1 _4450_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__5145__A2 _5143_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3401_ _3608_/A _3405_/B _3405_/C _3400_/X _3561_/A vssd1 vssd1 vccd1 vccd1 _3401_/X
+ sky130_fd_sc_hd__o32a_1
X_4381_ _4381_/A vssd1 vssd1 vccd1 vccd1 _4384_/A sky130_fd_sc_hd__inv_2
XFILLER_98_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6120_ _6155_/CLK _6120_/D vssd1 vssd1 vccd1 vccd1 _6120_/Q sky130_fd_sc_hd__dfxtp_1
X_3332_ _5109_/A _3832_/A2 _3251_/B _3331_/Y _3255_/Y vssd1 vssd1 vccd1 vccd1 _3332_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5703__B _5703_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6051_ _6293_/CLK _6051_/D vssd1 vssd1 vccd1 vccd1 _6051_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3263_ _5800_/A _6067_/Q _4136_/A vssd1 vssd1 vccd1 vccd1 _3263_/Y sky130_fd_sc_hd__nor3b_4
XFILLER_113_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4656__A1 _6184_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3504__A _5707_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5002_ _6195_/Q _6194_/Q _5002_/C vssd1 vssd1 vccd1 vccd1 _5027_/B sky130_fd_sc_hd__and3_1
XFILLER_78_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3194_ _3960_/C _3893_/B vssd1 vssd1 vccd1 vccd1 _3194_/Y sky130_fd_sc_hd__nor2_2
XFILLER_93_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4104__A1_N _3807_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5081__A1 _5570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5081__B2 _5244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5904_ _3867_/B _3986_/B _3867_/A vssd1 vssd1 vccd1 vccd1 _5904_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_34_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_5__f_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_3_5__f_clk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_50_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5835_ _5835_/A1 _4436_/Y _5834_/X vssd1 vssd1 vccd1 vccd1 _6280_/D sky130_fd_sc_hd__a21o_1
XFILLER_50_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5384__A2 _5251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout326_A _5041_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5766_ _5767_/A _5767_/B _5766_/C vssd1 vssd1 vccd1 vccd1 _5788_/B sky130_fd_sc_hd__nor3_4
X_4717_ _6186_/Q _3671_/Y _5172_/B _4707_/B vssd1 vssd1 vccd1 vccd1 _4717_/X sky130_fd_sc_hd__o22a_1
X_5697_ _3593_/A _5696_/X _5712_/S vssd1 vssd1 vccd1 vccd1 _5698_/B sky130_fd_sc_hd__mux2_1
XFILLER_107_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4648_ _4648_/A _5330_/B vssd1 vssd1 vccd1 vccd1 _4648_/Y sky130_fd_sc_hd__nor2_8
XFILLER_135_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4579_ _5071_/A _4579_/B vssd1 vssd1 vccd1 vccd1 _6182_/D sky130_fd_sc_hd__and2_1
XANTENNA__4895__A1 _3116_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6249_ _6257_/CLK _6249_/D vssd1 vssd1 vccd1 vccd1 _6249_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5844__A0 _3274_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5051__D _5051_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4032__C1 _5932_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3043__B _5065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3950_ _5131_/B _4577_/C _3950_/C _4586_/B vssd1 vssd1 vccd1 vccd1 _5909_/A sky130_fd_sc_hd__and4_2
XFILLER_16_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3613__A2 _4837_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3881_ _3881_/A _3881_/B _5241_/B vssd1 vssd1 vccd1 vccd1 _4022_/D sky130_fd_sc_hd__or3b_4
XANTENNA__3994__A _5207_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5620_ _5618_/X _5619_/X _3941_/A vssd1 vssd1 vccd1 vccd1 _5644_/B sky130_fd_sc_hd__o21ai_1
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3377__A1 _6012_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5551_ _5551_/A _5551_/B vssd1 vssd1 vccd1 vccd1 _5551_/Y sky130_fd_sc_hd__nor2_1
X_4502_ _5255_/B _6149_/Q _4520_/S vssd1 vssd1 vccd1 vccd1 _4502_/X sky130_fd_sc_hd__mux2_1
X_5482_ _5500_/B _5482_/B vssd1 vssd1 vccd1 vccd1 _5482_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__3129__A1 _6004_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5402__A1_N _5507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4433_ _4437_/A1 _4432_/X _4423_/X vssd1 vssd1 vccd1 vccd1 _6115_/D sky130_fd_sc_hd__a21o_1
XFILLER_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5714__A _5714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4364_ _4334_/A _4426_/B _4410_/D _4362_/A vssd1 vssd1 vccd1 vccd1 _4364_/X sky130_fd_sc_hd__a22o_1
XFILLER_113_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6103_ _6180_/CLK _6103_/D vssd1 vssd1 vccd1 vccd1 _6103_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3315_ _3285_/Y _3316_/B _3314_/Y vssd1 vssd1 vccd1 vccd1 _3315_/Y sky130_fd_sc_hd__a21oi_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4295_ _4295_/A vssd1 vssd1 vccd1 vccd1 _4296_/B sky130_fd_sc_hd__inv_2
XFILLER_58_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4629__A1 _4806_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3234__A _3241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3246_ _3236_/Y _3913_/A vssd1 vssd1 vccd1 vccd1 _5470_/S sky130_fd_sc_hd__nand2b_4
X_6034_ _6278_/CLK _6034_/D vssd1 vssd1 vccd1 vccd1 _6034_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3177_ _3880_/A _3881_/B vssd1 vssd1 vccd1 vccd1 _4577_/C sky130_fd_sc_hd__or2_4
XFILLER_26_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3604__A2 _3593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5818_ _5818_/A _5818_/B vssd1 vssd1 vccd1 vccd1 _5819_/B sky130_fd_sc_hd__nor2_8
XANTENNA__5357__A2 _5556_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3368__A1 _4003_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5749_ _6244_/Q _5763_/B vssd1 vssd1 vccd1 vccd1 _5749_/X sky130_fd_sc_hd__or2_1
XFILLER_108_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5514__C1 _5075_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3144__A _3974_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5293__A1 _5292_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3843__A2 _5943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5045__A1 _5567_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5045__B2 _4931_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5348__A2 _3243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3980__C _5634_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3531__A1 _6015_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3054__A _5800_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3100_ _5238_/B _5169_/C _3116_/B vssd1 vssd1 vccd1 vccd1 _5096_/B sky130_fd_sc_hd__or3b_1
XFILLER_95_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4080_ _4233_/A1 _4078_/Y _4079_/X vssd1 vssd1 vccd1 vccd1 _6080_/D sky130_fd_sc_hd__a21o_1
XFILLER_95_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3031_ _4657_/A vssd1 vssd1 vccd1 vccd1 _5108_/A sky130_fd_sc_hd__inv_4
XFILLER_48_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4982_ _5504_/A _5488_/A _4979_/B vssd1 vssd1 vccd1 vccd1 _4988_/A sky130_fd_sc_hd__o21ai_2
XFILLER_17_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3933_ _3931_/Y _3932_/X _3933_/S vssd1 vssd1 vccd1 vccd1 _3933_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3864_ _3312_/A _5158_/A _4594_/B _3964_/B vssd1 vssd1 vccd1 vccd1 _3864_/X sky130_fd_sc_hd__a31o_1
XANTENNA__5428__B _5428_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5603_ _5598_/Y _5602_/Y _5603_/S vssd1 vssd1 vccd1 vccd1 _5603_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3795_ _3855_/S _3795_/B vssd1 vssd1 vccd1 vccd1 _3795_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__4011__A2 _3500_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3229__A _3555_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5534_ _5595_/A _5531_/Y _5532_/X _5533_/Y vssd1 vssd1 vccd1 vccd1 _5534_/X sky130_fd_sc_hd__a31o_1
XFILLER_11_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3770__A1 _4197_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5465_ _5607_/B1 _5463_/Y _5464_/X _5462_/X vssd1 vssd1 vccd1 vccd1 _5465_/X sky130_fd_sc_hd__a31o_1
XFILLER_127_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4416_ _4417_/A _4417_/B vssd1 vssd1 vccd1 vccd1 _4431_/A sky130_fd_sc_hd__nand2b_1
X_5396_ _5392_/A _5454_/B _5227_/Y _5395_/Y vssd1 vssd1 vccd1 vccd1 _5403_/B sky130_fd_sc_hd__o211a_1
Xfanout303 _6068_/Q vssd1 vssd1 vccd1 vccd1 _4642_/A sky130_fd_sc_hd__buf_12
XANTENNA__3522__A1 _3513_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout314 _5556_/C1 vssd1 vssd1 vccd1 vccd1 _5047_/C1 sky130_fd_sc_hd__clkbuf_4
XFILLER_99_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout325 input9/X vssd1 vssd1 vccd1 vccd1 _5932_/A sky130_fd_sc_hd__buf_6
X_4347_ _4347_/A _4347_/B _4347_/C vssd1 vssd1 vccd1 vccd1 _4348_/B sky130_fd_sc_hd__nor3_1
XFILLER_113_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_526 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout336 _4819_/B vssd1 vssd1 vccd1 vccd1 _5392_/A sky130_fd_sc_hd__buf_6
Xfanout347 _5264_/A vssd1 vssd1 vccd1 vccd1 _5226_/A sky130_fd_sc_hd__buf_6
XFILLER_98_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4278_ _4278_/A _4278_/B vssd1 vssd1 vccd1 vccd1 _4281_/A sky130_fd_sc_hd__xor2_4
XFILLER_100_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6017_ _6258_/CLK _6017_/D vssd1 vssd1 vccd1 vccd1 _6017_/Q sky130_fd_sc_hd__dfxtp_2
X_3229_ _3555_/B _3980_/B _3229_/C vssd1 vssd1 vccd1 vccd1 _3560_/S sky130_fd_sc_hd__and3_4
XFILLER_27_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3381__S0 _3241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4786__B1 _4785_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4523__A _4540_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4002__A2 _3615_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3139__A _3732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3761__A1 _4665_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5354__A _5595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5018__A1 _5547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5018__B2 _4638_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5974__C1 _5956_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3975__C _3975_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_20_clk_A _6084_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5741__A2 _5649_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3580_ _3313_/Y _3570_/X _3574_/X _3579_/Y vssd1 vssd1 vccd1 vccd1 _3580_/X sky130_fd_sc_hd__o211a_1
XFILLER_127_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3245__A_N _3236_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3752__A1 _3156_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5264__A _5264_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5250_ _5250_/A _5250_/B _5250_/C _5250_/D vssd1 vssd1 vccd1 vccd1 _5250_/X sky130_fd_sc_hd__and4_4
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_35_clk_A clkbuf_3_5__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4201_ _4200_/B _4275_/B _4200_/A vssd1 vssd1 vccd1 vccd1 _4209_/B sky130_fd_sc_hd__a21o_2
XFILLER_114_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5181_ _5136_/C _5177_/Y _5180_/X _5065_/A vssd1 vssd1 vccd1 vccd1 _5181_/Y sky130_fd_sc_hd__a211oi_1
XFILLER_69_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4132_ _4162_/B _4112_/C _4112_/D _4197_/A vssd1 vssd1 vccd1 vccd1 _4135_/B sky130_fd_sc_hd__a22o_1
XFILLER_95_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4063_ _6075_/Q _3721_/X _4066_/S vssd1 vssd1 vccd1 vccd1 _6075_/D sky130_fd_sc_hd__mux2_1
XFILLER_83_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4608__A _5976_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3014_ _3014_/A vssd1 vssd1 vccd1 vccd1 _5210_/B sky130_fd_sc_hd__inv_4
XFILLER_36_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4046__C _4462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4965_ _4987_/B _4965_/B vssd1 vssd1 vccd1 vccd1 _4965_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_51_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3658__S _3658_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3916_ _6051_/Q _3715_/X _3921_/S vssd1 vssd1 vccd1 vccd1 _6051_/D sky130_fd_sc_hd__mux2_1
XANTENNA__3440__A0 _6015_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4896_ _5509_/C _4896_/B vssd1 vssd1 vccd1 vccd1 _4896_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_fanout239_A _5128_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5158__B _5158_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5717__C1 _5799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3847_ _3987_/B _3738_/X _3801_/B _3846_/X vssd1 vssd1 vccd1 vccd1 _3847_/X sky130_fd_sc_hd__o211a_1
XANTENNA__5193__B1 _5192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3778_ _4658_/B _3740_/X _3749_/X vssd1 vssd1 vccd1 vccd1 _3778_/X sky130_fd_sc_hd__a21o_1
X_5517_ _5595_/A _5516_/Y _5251_/Y vssd1 vssd1 vccd1 vccd1 _5517_/X sky130_fd_sc_hd__a21o_1
XANTENNA__4940__B1 _5488_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3393__S _3551_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5448_ _5480_/B _5480_/C vssd1 vssd1 vccd1 vccd1 _5464_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__5605__C _5605_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5496__A1 _5488_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout100 _5238_/A vssd1 vssd1 vccd1 vccd1 _3060_/B sky130_fd_sc_hd__clkbuf_8
X_5379_ _6177_/Q _4234_/B _4058_/B _6137_/Q _5470_/S vssd1 vssd1 vccd1 vccd1 _5379_/X
+ sky130_fd_sc_hd__o221a_2
Xfanout111 _3458_/B vssd1 vssd1 vccd1 vccd1 _3450_/D sky130_fd_sc_hd__clkbuf_16
XFILLER_114_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout122 _3245_/X vssd1 vssd1 vccd1 vccd1 _5929_/B2 sky130_fd_sc_hd__buf_12
XFILLER_99_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout133 _3084_/X vssd1 vssd1 vccd1 vccd1 _5128_/S sky130_fd_sc_hd__buf_4
XFILLER_59_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout144 _5075_/C vssd1 vssd1 vccd1 vccd1 _3122_/A sky130_fd_sc_hd__buf_6
XFILLER_101_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout155 _3069_/Y vssd1 vssd1 vccd1 vccd1 _5454_/B sky130_fd_sc_hd__buf_6
Xfanout166 _5349_/B1 vssd1 vssd1 vccd1 vccd1 _3704_/B sky130_fd_sc_hd__buf_6
XFILLER_47_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout177 _3709_/X vssd1 vssd1 vccd1 vccd1 _4216_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_86_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout188 _3280_/X vssd1 vssd1 vccd1 vccd1 _4426_/B sky130_fd_sc_hd__buf_8
XFILLER_47_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout199 _3922_/S vssd1 vssd1 vccd1 vccd1 _3575_/B sky130_fd_sc_hd__buf_8
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5113__S _5129_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3422__A _3422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3141__B _6070_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_787 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5723__A2 _4167_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3498__A0 _3450_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3051__B _3970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5169__A_N _3971_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3986__B _3986_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5259__A _5292_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4750_ _4750_/A _4750_/B vssd1 vssd1 vccd1 vccd1 _4782_/B sky130_fd_sc_hd__nand2_1
XANTENNA__4163__A _4163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3701_ _4891_/A _6026_/Q _3902_/A vssd1 vssd1 vccd1 vccd1 _3701_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3973__A1 _4577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4681_ _4669_/X _4680_/X _5543_/S vssd1 vssd1 vccd1 vccd1 _4681_/X sky130_fd_sc_hd__mux2_1
X_3632_ _6017_/Q _3231_/Y _3592_/X _3631_/X vssd1 vssd1 vccd1 vccd1 _6017_/D sky130_fd_sc_hd__o22a_1
XFILLER_134_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5706__B _5706_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3563_ _3560_/X _4808_/B _3563_/S vssd1 vssd1 vccd1 vccd1 _3563_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5302_ _5498_/A _5302_/B vssd1 vssd1 vccd1 vccd1 _5302_/Y sky130_fd_sc_hd__nor2_1
X_6282_ _6284_/CLK _6282_/D vssd1 vssd1 vccd1 vccd1 _6282_/Q sky130_fd_sc_hd__dfxtp_1
X_3494_ _5707_/B _3494_/B vssd1 vssd1 vccd1 vccd1 _3495_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__5478__A1 _4974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5233_ _6173_/Q _4234_/B _4058_/B _6133_/Q _5470_/S vssd1 vssd1 vccd1 vccd1 _5233_/X
+ sky130_fd_sc_hd__o221a_2
XFILLER_102_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5164_ _5238_/C _5179_/B _5164_/C vssd1 vssd1 vccd1 vccd1 _5164_/Y sky130_fd_sc_hd__nor3_1
XFILLER_96_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4115_ _4115_/A _4115_/B vssd1 vssd1 vccd1 vccd1 _4117_/B sky130_fd_sc_hd__xnor2_4
XFILLER_110_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5095_ _5095_/A _5203_/A _5203_/C vssd1 vssd1 vccd1 vccd1 _5095_/X sky130_fd_sc_hd__or3_1
XFILLER_110_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3242__A _3243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout189_A _5742_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4046_ _4046_/A _5075_/B _4462_/A _4046_/D vssd1 vssd1 vccd1 vccd1 _4051_/S sky130_fd_sc_hd__or4_4
XANTENNA__4057__B _4058_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4453__A2 _4438_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5650__A1 _3388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5938__C1 _4638_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5997_ _6143_/Q vssd1 vssd1 vccd1 vccd1 _6143_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_52_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4948_ _4974_/A _4972_/B _4972_/C _6004_/Q vssd1 vssd1 vccd1 vccd1 _4948_/X sky130_fd_sc_hd__a31o_1
XFILLER_20_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4879_ _4879_/A _4879_/B vssd1 vssd1 vccd1 vccd1 _4879_/Y sky130_fd_sc_hd__nand2_1
XFILLER_137_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5705__A2 _5888_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3716__A1 _3715_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3136__B _3869_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4248__A _5767_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3152__A _3958_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4444__A2 _4458_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5641__A1 _5051_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5929__C1 _4638_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5944__A2 _3575_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4133__D _4342_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5157__B1 _3116_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4132__A1 _4162_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4132__B2 _4197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5261__B _5653_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5880__A1 _3942_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4435__A2 _4410_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3997__A _4697_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5920_ _5242_/A _5244_/X _5920_/C _5920_/D vssd1 vssd1 vccd1 vccd1 _5921_/C sky130_fd_sc_hd__and4bb_1
XFILLER_47_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5851_ _6283_/Q _5854_/A _5850_/Y _5866_/B1 vssd1 vssd1 vccd1 vccd1 _6283_/D sky130_fd_sc_hd__o211a_1
X_4802_ _5392_/A _5703_/B vssd1 vssd1 vccd1 vccd1 _4840_/A sky130_fd_sc_hd__or2_2
XANTENNA__5396__B1 _5227_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5782_ _6255_/Q _5788_/B vssd1 vssd1 vccd1 vccd1 _5782_/X sky130_fd_sc_hd__or2_1
XFILLER_21_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3946__A1 _3649_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4733_ _5344_/A _4734_/B vssd1 vssd1 vccd1 vccd1 _4733_/X sky130_fd_sc_hd__or2_1
XFILLER_119_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4664_ _4662_/X _4664_/B vssd1 vssd1 vccd1 vccd1 _4666_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__5699__A1 _4767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3615_ _6207_/Q _3615_/B vssd1 vssd1 vccd1 vccd1 _3617_/B sky130_fd_sc_hd__or2_1
XFILLER_128_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4595_ _5840_/A _4003_/C _3862_/B _5241_/C vssd1 vssd1 vccd1 vccd1 _5221_/B sky130_fd_sc_hd__a31o_2
XANTENNA__3237__A _5436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3546_ _3599_/A _5707_/B _3599_/B vssd1 vssd1 vccd1 vccd1 _3546_/X sky130_fd_sc_hd__and3_1
XFILLER_135_17 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6265_ _6265_/CLK _6265_/D vssd1 vssd1 vccd1 vccd1 _6265_/Q sky130_fd_sc_hd__dfxtp_1
X_3477_ _3476_/A _5677_/B _3476_/Y vssd1 vssd1 vccd1 vccd1 _3477_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_103_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5216_ _5218_/B _5214_/A _5219_/A _4646_/A vssd1 vssd1 vccd1 vccd1 _5217_/B sky130_fd_sc_hd__o211a_1
XANTENNA__5320__B1 _3239_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6196_ _6196_/CLK _6196_/D vssd1 vssd1 vccd1 vccd1 _6196_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_69_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5147_ _5543_/S _5158_/A _5147_/C _5147_/D vssd1 vssd1 vccd1 vccd1 _5147_/X sky130_fd_sc_hd__or4_1
XFILLER_69_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5078_ _5258_/A _3059_/Y _3062_/Y _5928_/A _4603_/Y vssd1 vssd1 vccd1 vccd1 _5079_/A
+ sky130_fd_sc_hd__a311o_1
XANTENNA__5623__A1 _4622_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4029_ _5128_/A0 _3986_/B _5634_/B vssd1 vssd1 vccd1 vccd1 _4029_/X sky130_fd_sc_hd__mux2_1
XFILLER_72_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4831__C1 _4640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5627__A _6292_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4531__A _5932_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5234__S0 _3241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4250__B _4251_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3147__A _3880_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4706__A _6221_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5301__S _5539_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4425__B _4426_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5378__B1 _5767_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5917__A2 _3950_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4050__A0 _4657_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4889__C1 _5050_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3057__A _5218_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3400_ _3500_/A _3500_/B vssd1 vssd1 vccd1 vccd1 _3400_/X sky130_fd_sc_hd__xor2_2
X_4380_ _4401_/A _4380_/B vssd1 vssd1 vccd1 vccd1 _4381_/A sky130_fd_sc_hd__nand2_1
XFILLER_125_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3331_ _3331_/A vssd1 vssd1 vccd1 vccd1 _3331_/Y sky130_fd_sc_hd__inv_2
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4105__A1 _4437_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6050_ _6259_/CLK _6050_/D vssd1 vssd1 vccd1 vccd1 _6050_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3262_ _3885_/A _5264_/B vssd1 vssd1 vccd1 vccd1 _3267_/A sky130_fd_sc_hd__nand2_4
XFILLER_98_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5001_ _4973_/Y _4974_/X _6006_/Q vssd1 vssd1 vccd1 vccd1 _5001_/X sky130_fd_sc_hd__a21bo_1
XFILLER_112_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3193_ _3312_/A _4594_/A vssd1 vssd1 vccd1 vccd1 _3893_/B sky130_fd_sc_hd__or2_4
XANTENNA__3864__B1 _3964_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5081__A2 _4604_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5903_ _5903_/A _5903_/B _5903_/C vssd1 vssd1 vccd1 vccd1 _5903_/Y sky130_fd_sc_hd__nand3_1
XFILLER_34_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5834_ _3666_/X _5819_/B _5819_/Y _6280_/Q vssd1 vssd1 vccd1 vccd1 _5834_/X sky130_fd_sc_hd__a22o_1
XFILLER_50_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5765_ _5790_/A1 _5742_/Y _5763_/X _5764_/X vssd1 vssd1 vccd1 vccd1 _6249_/D sky130_fd_sc_hd__a22o_1
X_4716_ _5330_/B _4716_/B vssd1 vssd1 vccd1 vccd1 _4716_/Y sky130_fd_sc_hd__nand2_1
X_5696_ _5694_/X _5695_/Y _3867_/B _3500_/C vssd1 vssd1 vccd1 vccd1 _5696_/X sky130_fd_sc_hd__a2bb2o_1
XANTENNA_fanout319_A _5799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4647_ _6184_/Q _4647_/B vssd1 vssd1 vccd1 vccd1 _4647_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5541__B1 _5547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4578_ _4622_/B _6182_/Q _4578_/S vssd1 vssd1 vccd1 vccd1 _4579_/B sky130_fd_sc_hd__mux2_1
XANTENNA__4895__A2 _4894_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3529_ _3476_/A _3937_/D _3528_/X vssd1 vssd1 vccd1 vccd1 _3529_/X sky130_fd_sc_hd__o21a_4
XFILLER_115_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6248_ _6248_/CLK _6248_/D vssd1 vssd1 vccd1 vccd1 _6248_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5844__A1 _5935_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6179_ _6179_/CLK _6179_/D vssd1 vssd1 vccd1 vccd1 _6179_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3855__A0 _3853_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4526__A _4539_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4583__B2 _4654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5532__B1 _5442_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5835__A1 _5835_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3324__B _4614_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_774 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3074__A1 _3060_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4271__B1 _4410_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3880_ _3880_/A _3880_/B vssd1 vssd1 vccd1 vccd1 _5241_/B sky130_fd_sc_hd__and2_4
XANTENNA__3994__B _3996_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3486__S _3709_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5550_ _5310_/Y _5542_/X _5546_/Y _5549_/X _5607_/B1 vssd1 vssd1 vccd1 vccd1 _5550_/X
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__4574__A1 _3958_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4501_ _5790_/A1 _4501_/A2 _4499_/X _4500_/X vssd1 vssd1 vccd1 vccd1 _6140_/D sky130_fd_sc_hd__a22o_1
X_5481_ _5480_/B _5480_/C _6227_/Q vssd1 vssd1 vccd1 vccd1 _5482_/B sky130_fd_sc_hd__a21oi_2
XANTENNA__5523__A0 _4707_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4432_ _4432_/A _4432_/B vssd1 vssd1 vccd1 vccd1 _4432_/X sky130_fd_sc_hd__and2_1
XANTENNA__5714__B _5714_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4363_ _4363_/A _4388_/A vssd1 vssd1 vccd1 vccd1 _4393_/A sky130_fd_sc_hd__nor2_2
XFILLER_98_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6102_ _6143_/CLK _6102_/D vssd1 vssd1 vccd1 vccd1 _6102_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3314_ _3285_/Y _3316_/B _3312_/Y vssd1 vssd1 vccd1 vccd1 _3314_/Y sky130_fd_sc_hd__o21ai_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4294_ _5818_/A _4294_/B vssd1 vssd1 vccd1 vccd1 _4295_/A sky130_fd_sc_hd__or2_4
XFILLER_98_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3234__B _3241_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5826__A1 _5835_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4629__A2 _4665_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6033_ _6263_/CLK _6033_/D vssd1 vssd1 vccd1 vccd1 _6033_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3245_ _3236_/Y _3913_/A vssd1 vssd1 vccd1 vccd1 _3245_/X sky130_fd_sc_hd__and2b_4
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5730__A _5730_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_752 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3176_ _3880_/A _3881_/B vssd1 vssd1 vccd1 vccd1 _4604_/B sky130_fd_sc_hd__nor2_4
XFILLER_67_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout171_A _3180_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5817_ _5817_/A1 _4231_/X _5816_/X vssd1 vssd1 vccd1 vccd1 _6272_/D sky130_fd_sc_hd__a21o_1
XANTENNA__5211__C1 _5956_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5762__A0 _3942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5748_ _5935_/A0 _5742_/Y _5746_/X _5747_/X vssd1 vssd1 vccd1 vccd1 _6243_/D sky130_fd_sc_hd__a22o_1
XFILLER_136_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3409__B _3410_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5679_ _5718_/A _5678_/X _5677_/Y _5732_/C1 vssd1 vssd1 vccd1 vccd1 _5687_/B sky130_fd_sc_hd__o211a_1
XFILLER_135_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_5__f_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3160__A _3880_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5045__A2 _4872_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_52_clk _6133_/CLK vssd1 vssd1 vccd1 vccd1 _6176_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__4005__B1 _4850_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5505__B1 _5504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3335__A _3986_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5808__A1 _3477_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3054__B _3869_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3030_ _4633_/B vssd1 vssd1 vccd1 vccd1 _3030_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_110_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4981_ _4981_/A vssd1 vssd1 vccd1 vccd1 _4989_/A sky130_fd_sc_hd__inv_2
XFILLER_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3932_ _3923_/B _3653_/C _3931_/Y vssd1 vssd1 vccd1 vccd1 _3932_/X sky130_fd_sc_hd__a21bo_1
Xclkbuf_leaf_43_clk clkbuf_3_4__f_clk/X vssd1 vssd1 vccd1 vccd1 _6262_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_32_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3863_ _4046_/A _5227_/B _4594_/B vssd1 vssd1 vccd1 vccd1 _3863_/X sky130_fd_sc_hd__and3_1
XFILLER_32_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_9_clk_A clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5602_ _6233_/Q _5602_/B vssd1 vssd1 vccd1 vccd1 _5602_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__5744__A0 _5768_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3794_ _3793_/B _3792_/Y _3793_/Y vssd1 vssd1 vccd1 vccd1 _3795_/B sky130_fd_sc_hd__a21o_2
XFILLER_118_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5533_ _5595_/A _5522_/Y _5251_/A vssd1 vssd1 vccd1 vccd1 _5533_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__3229__B _3980_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5464_ _5464_/A _5464_/B vssd1 vssd1 vccd1 vccd1 _5464_/X sky130_fd_sc_hd__or2_1
XANTENNA__3770__A2 _5943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4415_ _4424_/C _4415_/B vssd1 vssd1 vccd1 vccd1 _4417_/B sky130_fd_sc_hd__xnor2_2
X_5395_ _5393_/X _5394_/Y _5454_/B vssd1 vssd1 vccd1 vccd1 _5395_/Y sky130_fd_sc_hd__o21ai_1
X_4346_ _4347_/A _4347_/B _4347_/C vssd1 vssd1 vccd1 vccd1 _4348_/A sky130_fd_sc_hd__o21a_1
Xfanout304 _6067_/Q vssd1 vssd1 vccd1 vccd1 _3869_/A sky130_fd_sc_hd__buf_12
Xfanout315 _3028_/Y vssd1 vssd1 vccd1 vccd1 _5556_/C1 sky130_fd_sc_hd__buf_4
XFILLER_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout326 _5041_/S vssd1 vssd1 vccd1 vccd1 _4990_/A sky130_fd_sc_hd__buf_6
XFILLER_98_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout337 input6/X vssd1 vssd1 vccd1 vccd1 _4819_/B sky130_fd_sc_hd__buf_12
Xfanout348 _4633_/B vssd1 vssd1 vccd1 vccd1 _5264_/A sky130_fd_sc_hd__buf_6
XFILLER_59_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4775__S _4812_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4277_ _4277_/A _4277_/B vssd1 vssd1 vccd1 vccd1 _4278_/B sky130_fd_sc_hd__xor2_4
XFILLER_101_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6016_ _6258_/CLK _6016_/D vssd1 vssd1 vccd1 vccd1 _6016_/Q sky130_fd_sc_hd__dfxtp_2
X_3228_ _3228_/A _5617_/A _3750_/B vssd1 vssd1 vccd1 vccd1 _3564_/S sky130_fd_sc_hd__or3_4
XANTENNA__3286__A1 _6298_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4076__A _4136_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3381__S1 _3241_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3159_ _3974_/B _3268_/A vssd1 vssd1 vccd1 vccd1 _3163_/B sky130_fd_sc_hd__nand2_4
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3589__A2 _3589_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4786__A1 _3116_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_34_clk clkbuf_3_5__f_clk/X vssd1 vssd1 vccd1 vccd1 _6093_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_23_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3139__B _3555_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5635__A _5635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3155__A _3869_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4474__A0 _5446_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5018__A2 _5463_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5423__C1 _5507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4714__A _4990_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_25_clk clkbuf_3_5__f_clk/X vssd1 vssd1 vccd1 vccd1 _6258_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_60_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3752__A2 _5464_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5264__B _5264_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4200_ _4200_/A _4200_/B _4275_/B vssd1 vssd1 vccd1 vccd1 _4209_/A sky130_fd_sc_hd__nand3_4
XANTENNA__4701__A1 _4972_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4701__B2 _3740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5180_ _5180_/A _5195_/C vssd1 vssd1 vccd1 vccd1 _5180_/X sky130_fd_sc_hd__or2_1
X_4131_ _4301_/A _4311_/B vssd1 vssd1 vccd1 vccd1 _4135_/A sky130_fd_sc_hd__and2_1
XFILLER_68_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4062_ _6074_/Q _3718_/X _4066_/S vssd1 vssd1 vccd1 vccd1 _6074_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4465__A0 _5935_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4608__B _5241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3013_ _5255_/B vssd1 vssd1 vccd1 vccd1 _5221_/A sky130_fd_sc_hd__clkinv_4
XANTENNA__3512__B _5707_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5414__C1 _5556_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4964_ _4964_/A _4987_/A vssd1 vssd1 vccd1 vccd1 _4965_/B sky130_fd_sc_hd__nand2_1
XFILLER_52_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_16_clk _6233_/CLK vssd1 vssd1 vccd1 vccd1 _6234_/CLK sky130_fd_sc_hd__clkbuf_16
X_3915_ _6050_/Q _3711_/X _3921_/S vssd1 vssd1 vccd1 vccd1 _6050_/D sky130_fd_sc_hd__mux2_1
XFILLER_20_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4895_ _3116_/X _4894_/Y _4889_/X _4753_/A vssd1 vssd1 vccd1 vccd1 _4895_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_32_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5717__B1 _5716_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3991__A2 _5241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3846_ _5207_/S _3845_/B _3737_/Y _3845_/Y vssd1 vssd1 vccd1 vccd1 _3846_/X sky130_fd_sc_hd__a211o_1
XANTENNA_fanout134_A _5108_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3777_ _4096_/A _3776_/X _3777_/S vssd1 vssd1 vccd1 vccd1 _3777_/X sky130_fd_sc_hd__mux2_1
X_5516_ _5607_/B1 _5511_/X _5515_/X vssd1 vssd1 vccd1 vccd1 _5516_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout301_A _4642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4940__B2 _4872_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5447_ _4872_/A _5446_/C _5480_/B vssd1 vssd1 vccd1 vccd1 _5447_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_106_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5496__A2 _5556_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5378_ _6153_/Q _3243_/A _5767_/B _6129_/Q vssd1 vssd1 vccd1 vccd1 _5378_/X sky130_fd_sc_hd__o22a_2
Xfanout101 _3057_/X vssd1 vssd1 vccd1 vccd1 _5238_/A sky130_fd_sc_hd__buf_4
XFILLER_99_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout112 _3500_/C vssd1 vssd1 vccd1 vccd1 _3458_/B sky130_fd_sc_hd__buf_6
Xfanout123 _3245_/X vssd1 vssd1 vccd1 vccd1 _3590_/A1 sky130_fd_sc_hd__buf_4
XFILLER_114_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4329_ _4330_/A _4330_/B _4330_/C vssd1 vssd1 vccd1 vccd1 _4358_/B sky130_fd_sc_hd__a21o_2
Xfanout134 _5108_/B vssd1 vssd1 vccd1 vccd1 _5124_/S sky130_fd_sc_hd__buf_6
XFILLER_99_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout145 _3076_/X vssd1 vssd1 vccd1 vccd1 _5075_/C sky130_fd_sc_hd__buf_8
XFILLER_113_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout156 _3069_/Y vssd1 vssd1 vccd1 vccd1 _5718_/A sky130_fd_sc_hd__clkbuf_4
Xfanout167 _3240_/Y vssd1 vssd1 vccd1 vccd1 _5349_/B1 sky130_fd_sc_hd__buf_4
XFILLER_59_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout178 _4167_/D vssd1 vssd1 vccd1 vccd1 _4410_/D sky130_fd_sc_hd__clkbuf_16
Xfanout189 _5742_/B vssd1 vssd1 vccd1 vccd1 _5767_/B sky130_fd_sc_hd__buf_6
XANTENNA__3259__A1 _6011_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4534__A _4540_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3431__A1 _5470_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5184__A1 _3116_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5365__A _5367_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4447__B1 _3900_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4998__A1 _6194_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output28_A _6182_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5947__A0 _6295_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4163__B _4311_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3700_ _3942_/A _3699_/X _3705_/A vssd1 vssd1 vccd1 vccd1 _6025_/D sky130_fd_sc_hd__mux2_1
X_4680_ _6185_/Q _5263_/A _5054_/A vssd1 vssd1 vccd1 vccd1 _4680_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3973__A2 _5158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3631_ _3631_/A _3631_/B vssd1 vssd1 vccd1 vccd1 _3631_/X sky130_fd_sc_hd__and2_1
X_3562_ _3644_/B _3567_/B _3544_/X _3608_/A _3561_/X vssd1 vssd1 vccd1 vccd1 _4808_/B
+ sky130_fd_sc_hd__o221a_4
XFILLER_115_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3281__S0 _4067_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5301_ _5305_/A _4714_/B _5539_/S vssd1 vssd1 vccd1 vccd1 _5302_/B sky130_fd_sc_hd__mux2_2
XFILLER_6_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6281_ _6284_/CLK _6281_/D vssd1 vssd1 vccd1 vccd1 _6281_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3493_ _3387_/X _3450_/D _3599_/B _3599_/A vssd1 vssd1 vccd1 vccd1 _3494_/B sky130_fd_sc_hd__a22o_2
XFILLER_5_191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5232_ _6149_/Q _3243_/A _5767_/B _6125_/Q vssd1 vssd1 vccd1 vccd1 _5232_/X sky130_fd_sc_hd__o22a_1
XFILLER_103_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_5_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _6193_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_102_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5163_ _5162_/B _6210_/Q _3092_/B vssd1 vssd1 vccd1 vccd1 _5164_/C sky130_fd_sc_hd__a21oi_2
XFILLER_96_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4114_ _4112_/X _4114_/B vssd1 vssd1 vccd1 vccd1 _4115_/B sky130_fd_sc_hd__and2b_2
XANTENNA__4438__A0 _5768_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5094_ _6198_/Q _5085_/Y _5093_/X _5071_/A vssd1 vssd1 vccd1 vccd1 _6198_/D sky130_fd_sc_hd__o211a_1
XFILLER_111_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3242__B _5924_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4045_ _5561_/S _3112_/B _5075_/C _4596_/B vssd1 vssd1 vccd1 vccd1 _4046_/D sky130_fd_sc_hd__a22o_1
XFILLER_49_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4057__C _5742_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_703 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5650__A2 _5203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout251_A _6238_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout349_A input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5996_ _6142_/Q vssd1 vssd1 vccd1 vccd1 _6142_/D sky130_fd_sc_hd__clkbuf_2
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4947_ _4946_/A _4946_/B _4944_/X vssd1 vssd1 vccd1 vccd1 _4947_/Y sky130_fd_sc_hd__a21oi_2
X_4878_ _4876_/X _4912_/B vssd1 vssd1 vccd1 vccd1 _4879_/B sky130_fd_sc_hd__and2b_1
XFILLER_137_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3829_ _5888_/B _3841_/S vssd1 vssd1 vccd1 vccd1 _3829_/Y sky130_fd_sc_hd__nor2_1
XFILLER_119_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5469__A2 _3243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4529__A _4540_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5124__S _5124_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4248__B _4251_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3152__B _5143_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4264__A _4362_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_34_clk_A clkbuf_3_5__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3404__A1 _4162_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5794__S _5798_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_49_clk_A _6230_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4904__A1 _5480_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4904__B2 _4931_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4132__A2 _4112_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3340__B1 _5296_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5880__A2 _5934_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3997__B _5114_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5850_ _5854_/A _5850_/B vssd1 vssd1 vccd1 vccd1 _5850_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4801_ _4769_/A _4769_/B _4766_/X vssd1 vssd1 vccd1 vccd1 _4805_/A sky130_fd_sc_hd__a21oi_1
XTAP_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5396__A1 _5392_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5781_ _5856_/A _4250_/Y _5779_/X _5780_/Y vssd1 vssd1 vccd1 vccd1 _6254_/D sky130_fd_sc_hd__a22o_1
X_4732_ _5114_/A _4734_/B vssd1 vssd1 vccd1 vccd1 _4735_/A sky130_fd_sc_hd__nor2_1
XFILLER_30_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4663_ _5263_/A _4663_/B vssd1 vssd1 vccd1 vccd1 _4664_/B sky130_fd_sc_hd__or2_1
XANTENNA__4621__B _5706_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5699__A2 _5714_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3614_ _6207_/Q _3615_/B vssd1 vssd1 vccd1 vccd1 _3652_/A sky130_fd_sc_hd__nand2_2
XANTENNA__5436__C _5436_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4594_ _4594_/A _4594_/B vssd1 vssd1 vccd1 vccd1 _5241_/C sky130_fd_sc_hd__nor2_1
XFILLER_116_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3237__B _5436_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3545_ _3646_/B _3567_/B _3544_/X _3611_/A _3541_/X vssd1 vssd1 vccd1 vccd1 _5703_/B
+ sky130_fd_sc_hd__o221a_4
XFILLER_115_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5733__A _5733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6264_ _6264_/CLK _6264_/D vssd1 vssd1 vccd1 vccd1 _6264_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3476_ _3476_/A _3476_/B vssd1 vssd1 vccd1 vccd1 _3476_/Y sky130_fd_sc_hd__nand2_1
XFILLER_89_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5215_ _5255_/B _5218_/B vssd1 vssd1 vccd1 vccd1 _5219_/A sky130_fd_sc_hd__nand2_1
XFILLER_103_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6195_ _6288_/CLK _6195_/D vssd1 vssd1 vccd1 vccd1 _6195_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_130_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3253__A _5936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout299_A _6069_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5146_ _5258_/A _5143_/A _5144_/X _5158_/C vssd1 vssd1 vccd1 vccd1 _5147_/D sky130_fd_sc_hd__a211o_1
XFILLER_97_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5077_ _3062_/Y _5077_/B _5077_/C vssd1 vssd1 vccd1 vccd1 _5079_/B sky130_fd_sc_hd__and3b_1
XANTENNA__5623__A2 _5058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4028_ _3940_/A _5900_/A _3934_/X vssd1 vssd1 vccd1 vccd1 _4028_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__3634__A1 _3387_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5979_ _4846_/A _5985_/B _5959_/A _5862_/A vssd1 vssd1 vccd1 vccd1 _5979_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_40_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5234__S1 _3241_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3147__B _3948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4958__S _5050_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5847__C1 _5866_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3163__A _3575_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3625__A1 _3615_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4706__B _4707_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5818__A _5818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4050__A1 _5075_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3057__B _3058_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4868__S _4990_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3330_ _3590_/A1 _3329_/X _3328_/X vssd1 vssd1 vccd1 vccd1 _3331_/A sky130_fd_sc_hd__a21oi_4
XFILLER_98_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3261_ _3885_/A _5264_/B vssd1 vssd1 vccd1 vccd1 _3266_/A sky130_fd_sc_hd__and2_4
XFILLER_124_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3073__A _3121_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5000_ _4946_/A _4946_/B _4999_/Y _4944_/X _6006_/Q vssd1 vssd1 vccd1 vccd1 _5000_/X
+ sky130_fd_sc_hd__a2111o_1
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3192_ _5840_/A _3952_/B vssd1 vssd1 vccd1 vccd1 _4594_/A sky130_fd_sc_hd__nand2_1
XANTENNA__3864__A1 _3312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5066__B1 _3974_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5902_ _4085_/A _5957_/B _3883_/X vssd1 vssd1 vccd1 vccd1 _5903_/C sky130_fd_sc_hd__a21o_1
XFILLER_50_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5833_ _5835_/A1 _4432_/X _5832_/X vssd1 vssd1 vccd1 vccd1 _6279_/D sky130_fd_sc_hd__a21o_1
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5728__A _5728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4632__A _5255_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5764_ _4891_/A _5761_/S _5791_/A vssd1 vssd1 vccd1 vccd1 _5764_/X sky130_fd_sc_hd__o21a_1
XANTENNA__4041__A1 _3721_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4715_ _6186_/Q _5041_/S _3122_/Y _4714_/Y vssd1 vssd1 vccd1 vccd1 _4715_/X sky130_fd_sc_hd__o211a_1
X_5695_ _5710_/S _4112_/D _5707_/A vssd1 vssd1 vccd1 vccd1 _5695_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_135_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4646_ _4646_/A _5403_/A vssd1 vssd1 vccd1 vccd1 _4646_/Y sky130_fd_sc_hd__nor2_4
XANTENNA_fanout214_A _3025_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5541__A1 _5540_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4577_ _4577_/A _4643_/A _4577_/C _4577_/D vssd1 vssd1 vccd1 vccd1 _4578_/S sky130_fd_sc_hd__or4_1
XANTENNA__5463__A _5463_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3552__B1 _5428_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3528_ _3564_/S _3506_/X _3527_/X vssd1 vssd1 vccd1 vccd1 _3528_/X sky130_fd_sc_hd__a21o_1
XFILLER_103_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6247_ _6254_/CLK _6247_/D vssd1 vssd1 vccd1 vccd1 _6247_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3459_ _3518_/A _3459_/B vssd1 vssd1 vccd1 vccd1 _3926_/C sky130_fd_sc_hd__and2_4
XFILLER_130_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6178_ _6284_/CLK _6178_/D vssd1 vssd1 vccd1 vccd1 _6178_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5129_ _5128_/X _6208_/Q _5129_/S vssd1 vssd1 vccd1 vccd1 _6208_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4807__A input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4526__B _6162_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_801 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5638__A _5638_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5780__A1 _3010_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3158__A _3941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5139__A1_N _5360_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5532__B2 _3382_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3543__B1 _3597_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3846__A1 _5207_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_786 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3621__A _3621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4271__A1 _5109_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3074__A2 _5244_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4271__B2 _4270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output10_A _3019_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5771__A1 _5292_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4574__A2 _3112_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4500_ _4891_/A _4239_/A _4059_/B vssd1 vssd1 vccd1 vccd1 _4500_/X sky130_fd_sc_hd__o21a_1
X_5480_ _5488_/A _5480_/B _5480_/C vssd1 vssd1 vccd1 vccd1 _5500_/B sky130_fd_sc_hd__and3_2
XFILLER_117_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4431_ _4431_/A _4431_/B _4431_/C vssd1 vssd1 vccd1 vccd1 _4432_/B sky130_fd_sc_hd__nand3_1
XFILLER_117_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5283__A _5283_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3534__B1 _5924_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4362_ _4362_/A _4426_/B vssd1 vssd1 vccd1 vccd1 _4388_/A sky130_fd_sc_hd__nand2_4
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6101_ _6180_/CLK _6101_/D vssd1 vssd1 vccd1 vccd1 _6101_/Q sky130_fd_sc_hd__dfxtp_1
X_3313_ _3974_/B _4003_/C vssd1 vssd1 vccd1 vccd1 _3313_/Y sky130_fd_sc_hd__nand2_2
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4293_ _4330_/B _4293_/B vssd1 vssd1 vccd1 vccd1 _4293_/X sky130_fd_sc_hd__and2_1
XFILLER_113_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5287__B1 _5058_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6032_ _6258_/CLK _6032_/D vssd1 vssd1 vccd1 vccd1 _6032_/Q sky130_fd_sc_hd__dfxtp_1
X_3244_ _6094_/Q _3589_/A2 _3589_/B1 _6087_/Q vssd1 vssd1 vccd1 vccd1 _3244_/X sky130_fd_sc_hd__o22a_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3837__A1 _3593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5730__B _5900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3175_ _5634_/A _3312_/A vssd1 vssd1 vccd1 vccd1 _3881_/B sky130_fd_sc_hd__nand2_8
XFILLER_82_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout164_A _5349_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4362__A _4362_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout331_A input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5816_ _3666_/X _5801_/B _5801_/Y _6272_/Q vssd1 vssd1 vccd1 vccd1 _5816_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4014__A1 _3029_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5747_ _5292_/B _5761_/S _5791_/A vssd1 vssd1 vccd1 vccd1 _5747_/X sky130_fd_sc_hd__o21a_1
XFILLER_108_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5678_ _4726_/B _4734_/B _5703_/A vssd1 vssd1 vccd1 vccd1 _5678_/X sky130_fd_sc_hd__mux2_1
XFILLER_136_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5514__A1 _5503_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4629_ _4806_/S _4665_/B _5226_/A vssd1 vssd1 vccd1 vccd1 _4629_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_123_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3706__A _3706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3425__B _3425_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5278__B1 _4058_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3828__A1 _5703_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout77_A _3121_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4253__A1 _3711_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5753__A1 _3011_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3952__C_N _4604_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5269__A0 _4657_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4492__A1 _5856_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4980_ _4980_/A _4980_/B vssd1 vssd1 vccd1 vccd1 _4981_/A sky130_fd_sc_hd__nand2_2
XFILLER_63_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3931_ _5656_/A _3931_/B vssd1 vssd1 vccd1 vccd1 _3931_/Y sky130_fd_sc_hd__nand2_1
XFILLER_16_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3862_ _3885_/A _3862_/B vssd1 vssd1 vccd1 vccd1 _4594_/B sky130_fd_sc_hd__or2_4
XFILLER_20_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5601_ _4645_/B _5598_/Y _5600_/X vssd1 vssd1 vccd1 vccd1 _5601_/X sky130_fd_sc_hd__o21a_1
XFILLER_31_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3793_ _3937_/C _3793_/B vssd1 vssd1 vccd1 vccd1 _3793_/Y sky130_fd_sc_hd__nor2_1
X_5532_ _4586_/B _5522_/Y _5442_/A _3382_/X vssd1 vssd1 vccd1 vccd1 _5532_/X sky130_fd_sc_hd__o2bb2a_1
XANTENNA__4910__A _4974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5463_ _5463_/A _5463_/B vssd1 vssd1 vccd1 vccd1 _5463_/Y sky130_fd_sc_hd__nand2_1
XFILLER_117_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4414_ _4424_/A _4424_/B _4394_/A vssd1 vssd1 vccd1 vccd1 _4415_/B sky130_fd_sc_hd__o21ai_2
X_5394_ _5391_/A _5392_/X _5365_/X _5370_/A vssd1 vssd1 vccd1 vccd1 _5394_/Y sky130_fd_sc_hd__a211oi_1
XFILLER_99_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4345_ _4345_/A _4345_/B vssd1 vssd1 vccd1 vccd1 _4347_/C sky130_fd_sc_hd__xor2_1
Xfanout305 _3873_/A vssd1 vssd1 vccd1 vccd1 _5976_/A sky130_fd_sc_hd__clkbuf_8
Xfanout316 _4576_/A vssd1 vssd1 vccd1 vccd1 _5071_/A sky130_fd_sc_hd__buf_6
XFILLER_98_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout327 _5072_/A vssd1 vssd1 vccd1 vccd1 _5041_/S sky130_fd_sc_hd__buf_6
XFILLER_101_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout338 input5/X vssd1 vssd1 vccd1 vccd1 _5367_/A sky130_fd_sc_hd__buf_6
Xfanout349 input1/X vssd1 vssd1 vccd1 vccd1 _4633_/B sky130_fd_sc_hd__clkbuf_16
X_4276_ _4277_/B _4277_/A vssd1 vssd1 vccd1 vccd1 _4276_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_98_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6015_ _6258_/CLK _6015_/D vssd1 vssd1 vccd1 vccd1 _6015_/Q sky130_fd_sc_hd__dfxtp_4
X_3227_ _3227_/A _4592_/B _3749_/B vssd1 vssd1 vccd1 vccd1 _3227_/X sky130_fd_sc_hd__and3_4
XFILLER_101_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4483__A1 _5935_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3261__A _3885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3286__A2 _3643_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5680__B1 _3772_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3158_ _3941_/A _5143_/B vssd1 vssd1 vccd1 vccd1 _3387_/A sky130_fd_sc_hd__nor2_8
XANTENNA__4076__B _4176_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3089_ _3107_/B _5051_/B vssd1 vssd1 vccd1 vccd1 _5143_/A sky130_fd_sc_hd__or2_4
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5432__B1 _5936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4786__A2 _4776_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5127__S _5129_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3155__B _5165_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5370__B _5653_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4267__A _4410_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3171__A _6200_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5797__S _5798_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5974__A1 _5970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3985__B1 _3594_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4130_ _4163_/A _4173_/B _4110_/A _4108_/B vssd1 vssd1 vccd1 vccd1 _4152_/A sky130_fd_sc_hd__a31o_2
XANTENNA__3141__A_N _3970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_75 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4061_ _6073_/Q _3715_/X _4066_/S vssd1 vssd1 vccd1 vccd1 _6073_/D sky130_fd_sc_hd__mux2_1
XFILLER_49_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3081__A _5403_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_829 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3012_ _6221_/Q vssd1 vssd1 vccd1 vccd1 _5305_/A sky130_fd_sc_hd__inv_4
XFILLER_49_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5662__B1 _5728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3291__A_N _6008_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4217__A1 _4216_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4963_ _4963_/A _4963_/B vssd1 vssd1 vccd1 vccd1 _4963_/X sky130_fd_sc_hd__or2_1
XANTENNA__5965__A1 _4767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3914_ _4438_/S _4521_/S vssd1 vssd1 vccd1 vccd1 _3921_/S sky130_fd_sc_hd__nand2_8
X_4894_ _4900_/A _4894_/B vssd1 vssd1 vccd1 vccd1 _4894_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_20_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5717__A1 _4202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3845_ _5733_/B _3845_/B vssd1 vssd1 vccd1 vccd1 _3845_/Y sky130_fd_sc_hd__nor2_1
XFILLER_20_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3991__A3 _3975_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4640__A _4640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3776_ _3450_/A _3775_/X _3812_/S vssd1 vssd1 vccd1 vccd1 _3776_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5515_ _3331_/A _5442_/A _5513_/B _5943_/C _5514_/X vssd1 vssd1 vccd1 vccd1 _5515_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_133_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5446_ _5480_/B _5446_/B _5446_/C vssd1 vssd1 vccd1 vccd1 _5504_/C sky130_fd_sc_hd__and3_2
XFILLER_121_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5377_ _6254_/Q _6121_/Q _6023_/Q _6246_/Q _3241_/A _3241_/B vssd1 vssd1 vccd1 vccd1
+ _5377_/X sky130_fd_sc_hd__mux4_2
XANTENNA__3690__S _3705_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout102 _3965_/Y vssd1 vssd1 vccd1 vccd1 _5442_/A sky130_fd_sc_hd__buf_4
XFILLER_59_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout113 _3397_/X vssd1 vssd1 vccd1 vccd1 _3500_/C sky130_fd_sc_hd__buf_6
XFILLER_99_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout124 _4604_/C vssd1 vssd1 vccd1 vccd1 _5710_/S sky130_fd_sc_hd__buf_4
X_4328_ _4328_/A _4328_/B vssd1 vssd1 vccd1 vccd1 _4330_/C sky130_fd_sc_hd__xor2_1
Xfanout135 _3084_/X vssd1 vssd1 vccd1 vccd1 _5108_/B sky130_fd_sc_hd__buf_6
XFILLER_87_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout146 _3123_/A vssd1 vssd1 vccd1 vccd1 _5403_/A sky130_fd_sc_hd__clkbuf_16
XANTENNA_input1_A io_in[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout157 _3060_/A vssd1 vssd1 vccd1 vccd1 _3121_/B sky130_fd_sc_hd__clkbuf_16
XANTENNA__3703__B _3704_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout168 _3239_/X vssd1 vssd1 vccd1 vccd1 _4234_/B sky130_fd_sc_hd__buf_6
Xfanout179 _3553_/X vssd1 vssd1 vccd1 vccd1 _4167_/D sky130_fd_sc_hd__buf_6
X_4259_ _6100_/Q _3730_/X _4259_/S vssd1 vssd1 vccd1 vccd1 _6100_/D sky130_fd_sc_hd__mux2_1
XFILLER_74_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4456__A1 _5446_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5184__A2 _5143_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5365__B _5367_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3166__A _5840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_8_clk_A clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4447__A1 _3011_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4725__A _5114_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3973__A3 _3950_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3630_ _3476_/A _5898_/B _3613_/Y vssd1 vssd1 vccd1 vccd1 _3631_/B sky130_fd_sc_hd__o21ai_4
X_3561_ _3561_/A _3561_/B vssd1 vssd1 vccd1 vccd1 _3561_/X sky130_fd_sc_hd__or2_1
XANTENNA__3076__A _5218_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3281__S1 _3709_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5300_ _3032_/Y _5360_/S _5299_/Y vssd1 vssd1 vccd1 vccd1 _5300_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6280_ _6280_/CLK _6280_/D vssd1 vssd1 vccd1 vccd1 _6280_/Q sky130_fd_sc_hd__dfxtp_1
X_3492_ _3492_/A _3492_/B vssd1 vssd1 vccd1 vccd1 _3492_/X sky130_fd_sc_hd__or2_2
XFILLER_6_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5231_ _5075_/C _5224_/X _5229_/X _5230_/X vssd1 vssd1 vccd1 vccd1 _5231_/X sky130_fd_sc_hd__a31o_1
XANTENNA__3226__D _4812_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5291__A _5507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5162_ _6212_/Q _5162_/B _5258_/A vssd1 vssd1 vccd1 vccd1 _5179_/B sky130_fd_sc_hd__and3_2
XFILLER_57_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4113_ _4197_/A _4112_/C _4112_/D _4197_/B vssd1 vssd1 vccd1 vccd1 _4114_/B sky130_fd_sc_hd__a22o_1
X_5093_ _5093_/A _5093_/B _5093_/C vssd1 vssd1 vccd1 vccd1 _5093_/X sky130_fd_sc_hd__or3_1
XFILLER_56_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6133__CLK _6133_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4044_ _6065_/Q _3730_/X _4044_/S vssd1 vssd1 vccd1 vccd1 _6065_/D sky130_fd_sc_hd__mux2_1
XFILLER_56_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5399__C1 _5570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5995_ _6141_/Q vssd1 vssd1 vccd1 vccd1 _6141_/D sky130_fd_sc_hd__clkbuf_2
XANTENNA__5938__B2 _5928_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5169__C _5169_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout244_A _5862_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4946_ _4946_/A _4946_/B vssd1 vssd1 vccd1 vccd1 _4946_/Y sky130_fd_sc_hd__nand2_1
XFILLER_138_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4877_ _5454_/A _4877_/B vssd1 vssd1 vccd1 vccd1 _4912_/B sky130_fd_sc_hd__or2_2
XFILLER_137_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3828_ _5703_/B _3816_/B _3827_/X vssd1 vssd1 vccd1 vccd1 _3828_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_137_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5571__C1 _5403_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3759_ _4136_/A _3777_/S _3758_/X _3751_/A vssd1 vssd1 vccd1 vccd1 _3759_/X sky130_fd_sc_hd__o211a_1
XFILLER_118_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5323__C1 _5251_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5429_ _5427_/Y _5428_/X _5391_/Y _5393_/X vssd1 vssd1 vccd1 vccd1 _5429_/Y sky130_fd_sc_hd__a211oi_1
XANTENNA__4677__A1 _3116_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4677__B2 _4744_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5929__A1 _5928_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4264__B _4342_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5929__B2 _5929_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5095__B _5203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4904__A2 _5871_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4668__A1 _3740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5865__A0 _3649_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4668__B2 _4972_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3340__A1 _4162_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3340__B2 _3885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3628__C1 _3422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3997__C _5119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4800_ _4625_/A _5093_/A _4798_/X _4799_/X _5071_/A vssd1 vssd1 vccd1 vccd1 _6188_/D
+ sky130_fd_sc_hd__o311a_1
XTAP_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5780_ _3010_/Y _5788_/B _4250_/Y vssd1 vssd1 vccd1 vccd1 _5780_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__5396__A2 _5454_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4731_ _4729_/Y _4730_/X _5114_/A _4886_/B vssd1 vssd1 vccd1 vccd1 _4731_/X sky130_fd_sc_hd__a2bb2o_1
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3946__A3 _5634_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4662_ _5263_/A _4663_/B vssd1 vssd1 vccd1 vccd1 _4662_/X sky130_fd_sc_hd__and2_1
XFILLER_119_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3613_ _3564_/S _4837_/B _3610_/X _3476_/A vssd1 vssd1 vccd1 vccd1 _3613_/Y sky130_fd_sc_hd__o211ai_4
X_4593_ _5162_/B _5258_/A vssd1 vssd1 vccd1 vccd1 _4593_/Y sky130_fd_sc_hd__xnor2_2
X_3544_ _3607_/A _3544_/B vssd1 vssd1 vccd1 vccd1 _3544_/X sky130_fd_sc_hd__or2_2
XFILLER_127_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6263_ _6263_/CLK _6263_/D vssd1 vssd1 vccd1 vccd1 _6263_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3475_ _4734_/B _3474_/X _3564_/S vssd1 vssd1 vccd1 vccd1 _3476_/B sky130_fd_sc_hd__mux2_1
XFILLER_88_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5214_ _5214_/A vssd1 vssd1 vccd1 vccd1 _5214_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5320__A2 _3243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6194_ _6288_/CLK _6194_/D vssd1 vssd1 vccd1 vccd1 _6194_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__3253__B _3706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5145_ _5561_/S _5143_/B _3116_/X vssd1 vssd1 vccd1 vccd1 _5158_/C sky130_fd_sc_hd__a21oi_1
XFILLER_96_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5608__B1 _3122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5076_ _3072_/A _3084_/B _5238_/A vssd1 vssd1 vccd1 vccd1 _5077_/C sky130_fd_sc_hd__o21a_1
XFILLER_56_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5084__A1 _5090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5623__A3 _3257_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4027_ _4002_/X _4026_/X _3995_/Y vssd1 vssd1 vccd1 vccd1 _4027_/X sky130_fd_sc_hd__a21o_1
XFILLER_65_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4831__A1 _4990_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5978_ _6300_/Q _5978_/B vssd1 vssd1 vccd1 vccd1 _5978_/X sky130_fd_sc_hd__or2_1
XFILLER_12_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4929_ _4934_/A _4929_/B vssd1 vssd1 vccd1 vccd1 _4930_/C sky130_fd_sc_hd__or2_1
XFILLER_60_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4898__A1 _5480_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5924__A _5924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3322__A1 _5889_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5378__A2 _3243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5818__B _5818_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5535__C1 _5948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4889__A1 _4745_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5550__A2 _5542_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3260_ _6273_/Q _6109_/Q _3551_/S vssd1 vssd1 vccd1 vccd1 _5264_/B sky130_fd_sc_hd__mux2_8
XFILLER_112_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3073__B _5330_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3191_ _4622_/B _6071_/Q vssd1 vssd1 vccd1 vccd1 _3952_/B sky130_fd_sc_hd__nor2_8
XANTENNA__3864__A2 _5158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5066__A1 _4604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4813__A1 _4972_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4813__B2 _3740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5901_ _5226_/A _5911_/C _3972_/Y _5878_/X vssd1 vssd1 vccd1 vccd1 _5901_/X sky130_fd_sc_hd__o31a_1
XFILLER_34_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5832_ _3631_/B _5819_/B _5819_/Y _6279_/Q vssd1 vssd1 vccd1 vccd1 _5832_/X sky130_fd_sc_hd__a22o_1
XFILLER_50_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4913__A _4972_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5763_ _6249_/Q _5763_/B vssd1 vssd1 vccd1 vccd1 _5763_/X sky130_fd_sc_hd__or2_1
XANTENNA__4632__B _4633_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4714_ _4990_/A _4714_/B vssd1 vssd1 vccd1 vccd1 _4714_/Y sky130_fd_sc_hd__nand2_1
X_5694_ _3765_/B _5380_/Y _5693_/X _5710_/S vssd1 vssd1 vccd1 vccd1 _5694_/X sky130_fd_sc_hd__o211a_1
XFILLER_108_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4645_ _5463_/A _4645_/B vssd1 vssd1 vccd1 vccd1 _4645_/Y sky130_fd_sc_hd__nand2_1
XFILLER_135_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout207_A _4022_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4576_ _4576_/A _4576_/B vssd1 vssd1 vccd1 vccd1 _6181_/D sky130_fd_sc_hd__and2_1
XANTENNA__5463__B _5463_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3552__A1 _4214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3552__B2 _3053_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3527_ _3227_/X _4767_/B _3583_/S vssd1 vssd1 vccd1 vccd1 _3527_/X sky130_fd_sc_hd__a21o_1
XFILLER_89_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6246_ _6254_/CLK _6246_/D vssd1 vssd1 vccd1 vccd1 _6246_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3458_ _6204_/Q _3458_/B vssd1 vssd1 vccd1 vccd1 _3459_/B sky130_fd_sc_hd__or2_1
XFILLER_130_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_33_clk_A clkbuf_3_5__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6177_ _6177_/CLK _6177_/D vssd1 vssd1 vccd1 vccd1 _6177_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3389_ _3500_/A _3389_/B vssd1 vssd1 vccd1 vccd1 _4620_/B sky130_fd_sc_hd__xnor2_4
XFILLER_97_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5128_ _5128_/A0 _5072_/A _5128_/S vssd1 vssd1 vccd1 vccd1 _5128_/X sky130_fd_sc_hd__mux2_1
XFILLER_111_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4807__B _4808_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5059_ _5838_/A _5059_/B _5059_/C _5919_/A vssd1 vssd1 vccd1 vccd1 _5062_/C sky130_fd_sc_hd__and4b_1
XFILLER_84_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_48_clk_A _6230_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_640 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5638__B _5638_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3791__A1 _4697_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3158__B _5143_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3543__A1 _5707_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3902__A _3902_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4271__A2 _3280_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3074__A3 _5169_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3881__C_N _5241_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4733__A _5344_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4452__B _4458_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4430_ _4431_/A _4431_/B _4431_/C vssd1 vssd1 vccd1 vccd1 _4432_/A sky130_fd_sc_hd__a21o_1
XFILLER_6_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4731__B1 _5114_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4361_ _3795_/B _4295_/A _4360_/Y vssd1 vssd1 vccd1 vccd1 _6111_/D sky130_fd_sc_hd__o21ai_1
XANTENNA__3084__A _5075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6100_ _6260_/CLK _6100_/D vssd1 vssd1 vccd1 vccd1 _6100_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3312_ _3312_/A _3312_/B vssd1 vssd1 vccd1 vccd1 _3312_/Y sky130_fd_sc_hd__nor2_4
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4292_ _4330_/A _4290_/X _4226_/Y _4230_/X vssd1 vssd1 vccd1 vccd1 _4293_/B sky130_fd_sc_hd__a211o_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6031_ _6262_/CLK _6031_/D vssd1 vssd1 vccd1 vccd1 _6031_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3243_ _3243_/A _5924_/B vssd1 vssd1 vccd1 vccd1 _3243_/Y sky130_fd_sc_hd__nand2_1
XFILLER_100_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3174_ _3740_/B _5617_/B vssd1 vssd1 vccd1 vccd1 _3750_/B sky130_fd_sc_hd__nand2_1
XFILLER_39_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4643__A _4643_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout157_A _3060_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5815_ _5817_/A1 _4190_/Y _5814_/X vssd1 vssd1 vccd1 vccd1 _6271_/D sky130_fd_sc_hd__a21o_1
XANTENNA__4362__B _4426_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5211__A1 _5960_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4014__A2 _3986_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5746_ _6243_/Q _5763_/B vssd1 vssd1 vccd1 vccd1 _5746_/X sky130_fd_sc_hd__or2_1
XFILLER_10_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout324_A _5932_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5677_ _5718_/A _5677_/B vssd1 vssd1 vccd1 vccd1 _5677_/Y sky130_fd_sc_hd__nand2_1
XFILLER_136_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3693__S _3902_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4628_ _5226_/A _4806_/S _4665_/B vssd1 vssd1 vccd1 vccd1 _4628_/X sky130_fd_sc_hd__and3_1
XANTENNA__3706__B _5048_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3525__A1 _3960_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4559_ _6179_/Q _4562_/B vssd1 vssd1 vccd1 vccd1 _4559_/X sky130_fd_sc_hd__or2_1
XFILLER_89_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6229_ _6295_/CLK _6229_/D vssd1 vssd1 vccd1 vccd1 _6229_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4818__A _5385_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4029__S _5634_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_73 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5269__A1 _6004_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5441__A1 _5929_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3930_ _3651_/B _3658_/X _3923_/Y _3929_/X vssd1 vssd1 vccd1 vccd1 _3933_/S sky130_fd_sc_hd__o2bb2a_1
XFILLER_32_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3861_ _3859_/Y _3860_/X _3858_/X vssd1 vssd1 vccd1 vccd1 _3862_/B sky130_fd_sc_hd__a21oi_2
XANTENNA__5729__C1 _5956_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3079__A _5258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5600_ _6009_/Q _4646_/A _3121_/X _5599_/X _5169_/C vssd1 vssd1 vccd1 vccd1 _5600_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3792_ _4690_/B _3816_/B _3791_/X vssd1 vssd1 vccd1 vccd1 _3792_/Y sky130_fd_sc_hd__o21ai_1
X_5531_ _5531_/A _5531_/B vssd1 vssd1 vccd1 vccd1 _5531_/Y sky130_fd_sc_hd__nand2_1
XFILLER_118_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5462_ _5312_/B _5464_/B _5461_/X vssd1 vssd1 vccd1 vccd1 _5462_/X sky130_fd_sc_hd__o21a_1
XFILLER_133_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4413_ _4413_/A _4413_/B vssd1 vssd1 vccd1 vccd1 _4424_/C sky130_fd_sc_hd__xnor2_4
X_5393_ _5365_/X _5370_/A _5391_/A _5392_/X vssd1 vssd1 vccd1 vccd1 _5393_/X sky130_fd_sc_hd__o211a_1
XFILLER_126_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4344_ _4343_/A _4371_/A _4341_/X vssd1 vssd1 vccd1 vccd1 _4345_/B sky130_fd_sc_hd__o21ai_2
XFILLER_98_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout306 _6066_/Q vssd1 vssd1 vccd1 vccd1 _3873_/A sky130_fd_sc_hd__buf_4
Xfanout317 _3028_/Y vssd1 vssd1 vccd1 vccd1 _4576_/A sky130_fd_sc_hd__buf_6
Xfanout328 input8/X vssd1 vssd1 vccd1 vccd1 _5072_/A sky130_fd_sc_hd__buf_8
XFILLER_99_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout339 input5/X vssd1 vssd1 vccd1 vccd1 _5119_/A sky130_fd_sc_hd__buf_12
X_4275_ _4275_/A _4275_/B vssd1 vssd1 vccd1 vccd1 _4277_/B sky130_fd_sc_hd__and2_2
XANTENNA__4638__A _4638_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3542__A _5707_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6014_ _6258_/CLK _6014_/D vssd1 vssd1 vccd1 vccd1 _6014_/Q sky130_fd_sc_hd__dfxtp_2
X_3226_ _4946_/A _3227_/A _3740_/B _4812_/S vssd1 vssd1 vccd1 vccd1 _3563_/S sky130_fd_sc_hd__and4_4
XFILLER_39_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5680__A1 _6298_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3261__B _5264_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3691__A0 _6221_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3157_ _5883_/A _4622_/B _3970_/A vssd1 vssd1 vccd1 vccd1 _3268_/A sky130_fd_sc_hd__and3_4
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3088_ _3107_/B _5051_/B vssd1 vssd1 vccd1 vccd1 _3170_/B sky130_fd_sc_hd__nor2_4
XANTENNA__3688__S _3705_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5729_ _4214_/A _5649_/X _5728_/X _5956_/A vssd1 vssd1 vccd1 vccd1 _6240_/D sky130_fd_sc_hd__o211a_1
XFILLER_136_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5932__A _5932_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4267__B _4311_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5671__A1 _3765_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_448 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5423__A1 _4644_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5423__B2 _3121_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5187__B1 _5072_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5111__A0 _5110_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4060_ _6072_/Q _3711_/X _4066_/S vssd1 vssd1 vccd1 vccd1 _6072_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3081__B _5512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5662__A1 _3388_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3011_ _5333_/A vssd1 vssd1 vccd1 vccd1 _3011_/Y sky130_fd_sc_hd__inv_4
XFILLER_36_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4870__C1 _4963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5414__A1 _5385_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4217__A2 _4216_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4962_ _5504_/A _4644_/Y _4959_/Y _4960_/X vssd1 vssd1 vccd1 vccd1 _4963_/B sky130_fd_sc_hd__o22a_1
XFILLER_91_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5965__A2 _5934_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3913_ _3913_/A _5742_/C vssd1 vssd1 vccd1 vccd1 _4521_/S sky130_fd_sc_hd__or2_4
X_4893_ _4867_/A _4862_/B _4925_/B vssd1 vssd1 vccd1 vccd1 _4894_/B sky130_fd_sc_hd__a21o_2
XANTENNA__4921__A _5488_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3844_ _6040_/Q _3771_/X _3842_/Y _3843_/X vssd1 vssd1 vccd1 vccd1 _6040_/D sky130_fd_sc_hd__a211o_1
XANTENNA__5717__A2 _5649_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3728__A1 _3727_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4640__B _4644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3775_ _5848_/A0 _3774_/X _3811_/S vssd1 vssd1 vccd1 vccd1 _3775_/X sky130_fd_sc_hd__mux2_1
X_5514_ _5503_/A _5513_/B _5512_/Y _5075_/C vssd1 vssd1 vccd1 vccd1 _5514_/X sky130_fd_sc_hd__a211o_1
XFILLER_118_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5445_ _4872_/A _5251_/A _5444_/X _5948_/A vssd1 vssd1 vccd1 vccd1 _6225_/D sky130_fd_sc_hd__o211a_1
XFILLER_118_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5350__B1 _5767_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5376_ _5310_/Y _5358_/Y _5375_/X _5595_/A vssd1 vssd1 vccd1 vccd1 _5376_/X sky130_fd_sc_hd__a22o_1
XFILLER_99_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout103 _3965_/Y vssd1 vssd1 vccd1 vccd1 _5638_/B sky130_fd_sc_hd__buf_4
XFILLER_120_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4327_ _4328_/A _4328_/B vssd1 vssd1 vccd1 vccd1 _4358_/A sky130_fd_sc_hd__nand2b_2
Xfanout114 _3801_/A vssd1 vssd1 vccd1 vccd1 _3500_/A sky130_fd_sc_hd__buf_12
Xfanout125 _3198_/X vssd1 vssd1 vccd1 vccd1 _4604_/C sky130_fd_sc_hd__buf_6
Xfanout136 _4638_/B vssd1 vssd1 vccd1 vccd1 _5158_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout147 _5605_/B vssd1 vssd1 vccd1 vccd1 _5360_/S sky130_fd_sc_hd__buf_8
Xfanout158 _3060_/A vssd1 vssd1 vccd1 vccd1 _5870_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_87_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3703__C _5767_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5102__B1 _3741_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout169 _3901_/B vssd1 vssd1 vccd1 vccd1 _3589_/A2 sky130_fd_sc_hd__buf_6
X_4258_ _6099_/Q _3727_/X _4259_/S vssd1 vssd1 vccd1 vccd1 _6099_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4456__A2 _4438_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3209_ _3228_/A _5617_/A _3750_/B vssd1 vssd1 vccd1 vccd1 _3210_/D sky130_fd_sc_hd__or3_1
XFILLER_27_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4189_ _4193_/A _4187_/X _4153_/X _4157_/A vssd1 vssd1 vccd1 vccd1 _4190_/B sky130_fd_sc_hd__o211a_1
XANTENNA__3664__B1 _4883_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3719__A1 _3718_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4042__S _4044_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3166__B _4462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3182__A _3880_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4447__A2 _4458_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3655__B1 _3621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4725__B _4726_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3560_ _3559_/Y _4202_/A _3560_/S vssd1 vssd1 vccd1 vccd1 _3560_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3076__B _5244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3491_ _3492_/A _3492_/B vssd1 vssd1 vccd1 vccd1 _3597_/B sky130_fd_sc_hd__nor2_8
XANTENNA__5572__A _5595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5230_ _5256_/B _5464_/A _4644_/A _5214_/Y _3678_/B vssd1 vssd1 vccd1 vccd1 _5230_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5161_ _5192_/A _5161_/B vssd1 vssd1 vccd1 vccd1 _6211_/D sky130_fd_sc_hd__nor2_1
XFILLER_96_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4112_ _4197_/A _4197_/B _4112_/C _4112_/D vssd1 vssd1 vccd1 vccd1 _4112_/X sky130_fd_sc_hd__and4_1
X_5092_ _4596_/B _5090_/Y _5091_/X _4931_/B vssd1 vssd1 vccd1 vccd1 _5093_/C sky130_fd_sc_hd__a31o_1
XFILLER_111_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4043_ _6064_/Q _3727_/X _4044_/S vssd1 vssd1 vccd1 vccd1 _6064_/D sky130_fd_sc_hd__mux2_1
XFILLER_56_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4916__A _6192_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4843__C1 _4972_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_587 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5994_ _6108_/Q vssd1 vssd1 vccd1 vccd1 _6108_/D sky130_fd_sc_hd__clkbuf_2
X_4945_ _4945_/A _4945_/B _5509_/B vssd1 vssd1 vccd1 vccd1 _4946_/B sky130_fd_sc_hd__or3b_4
XANTENNA__4610__A2 _3164_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4876_ _5454_/A _4877_/B vssd1 vssd1 vccd1 vccd1 _4876_/X sky130_fd_sc_hd__and2_1
XFILLER_20_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout237_A _5911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3827_ _4808_/B _3740_/X _3749_/X _3826_/X vssd1 vssd1 vccd1 vccd1 _3827_/X sky130_fd_sc_hd__a211o_1
XFILLER_119_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3758_ _3287_/A _3746_/A _3757_/X _3849_/B vssd1 vssd1 vccd1 vccd1 _3758_/X sky130_fd_sc_hd__a211o_1
XFILLER_119_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3689_ _5292_/B _6020_/Q _3902_/A vssd1 vssd1 vccd1 vccd1 _3689_/X sky130_fd_sc_hd__mux2_1
XFILLER_106_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5428_ _5428_/A _5428_/B vssd1 vssd1 vccd1 vccd1 _5428_/X sky130_fd_sc_hd__or2_1
XFILLER_121_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4677__A2 _4668_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5359_ _3010_/Y _4793_/B _5539_/S vssd1 vssd1 vccd1 vccd1 _5359_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4826__A _5605_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout52_A _5871_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3177__A _3880_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5392__A _5392_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5865__A1 _3944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3340__A2 _3257_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_532 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4455__B _4458_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3997__D _5392_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4053__A0 _3312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5567__A _5567_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4730_ _4698_/A _4727_/Y _4728_/X _4886_/B vssd1 vssd1 vccd1 vccd1 _4730_/X sky130_fd_sc_hd__a31o_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_75 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4661_ input2/X _4660_/X _4812_/S vssd1 vssd1 vccd1 vccd1 _4661_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3612_ _3646_/B _3594_/B _3606_/Y _3541_/A _3611_/X vssd1 vssd1 vccd1 vccd1 _4837_/B
+ sky130_fd_sc_hd__o221a_4
XANTENNA__5553__B1 _5542_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4592_ _4592_/A _4592_/B vssd1 vssd1 vccd1 vccd1 _5625_/C sky130_fd_sc_hd__or2_1
XFILLER_134_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3543_ _5707_/B _3599_/B _3597_/B vssd1 vssd1 vccd1 vccd1 _3544_/B sky130_fd_sc_hd__a21oi_1
XFILLER_127_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6262_ _6262_/CLK _6262_/D vssd1 vssd1 vccd1 vccd1 _6262_/Q sky130_fd_sc_hd__dfxtp_1
X_3474_ _3447_/X _4726_/B _3563_/S vssd1 vssd1 vccd1 vccd1 _3474_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5213_ _5255_/B _4634_/X _5561_/S vssd1 vssd1 vccd1 vccd1 _5214_/A sky130_fd_sc_hd__mux2_2
X_6193_ _6193_/CLK _6193_/D vssd1 vssd1 vccd1 vccd1 _6193_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_97_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3253__C _4614_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5144_ _5054_/A _4946_/A _5143_/Y vssd1 vssd1 vccd1 vccd1 _5144_/X sky130_fd_sc_hd__a21o_1
XFILLER_29_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5608__A1 _6233_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4646__A _4646_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5075_ _5075_/A _5075_/B _5075_/C vssd1 vssd1 vccd1 vccd1 _5077_/B sky130_fd_sc_hd__and3_1
XFILLER_56_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4026_ _5790_/A1 _5148_/A _3868_/Y _4025_/Y vssd1 vssd1 vccd1 vccd1 _4026_/X sky130_fd_sc_hd__a211o_1
XFILLER_37_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3634__A3 _3594_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3696__S _3705_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5977_ _4850_/A _5959_/A _5985_/C vssd1 vssd1 vccd1 vccd1 _5978_/B sky130_fd_sc_hd__a21oi_1
XFILLER_12_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4595__A1 _5840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4928_ _4934_/A _4929_/B vssd1 vssd1 vccd1 vccd1 _4983_/A sky130_fd_sc_hd__nand2_1
XFILLER_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4859_ _4925_/B _4925_/C vssd1 vssd1 vccd1 vccd1 _4867_/A sky130_fd_sc_hd__nor2_8
XFILLER_21_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_7_clk_A clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_0__f_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _6133_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__4898__A2 _4644_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5924__B _5924_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5387__A _5387_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4889__A2 _4887_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3635__A _3986_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_752 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4510__A1 _3011_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3190_ _3257_/B _3869_/B vssd1 vssd1 vccd1 vccd1 _3960_/C sky130_fd_sc_hd__nand2_4
XFILLER_79_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3864__A3 _4594_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5066__A2 _3971_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5900_ _5900_/A _5900_/B vssd1 vssd1 vccd1 vccd1 _5949_/B sky130_fd_sc_hd__and2_1
XFILLER_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5831_ _3583_/X _5819_/B _5830_/X vssd1 vssd1 vccd1 vccd1 _6278_/D sky130_fd_sc_hd__a21o_1
XFILLER_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5223__C1 _4638_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5762_ _3942_/A _5761_/X _5791_/A vssd1 vssd1 vccd1 vccd1 _6248_/D sky130_fd_sc_hd__mux2_1
XFILLER_50_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4713_ _4713_/A _4713_/B vssd1 vssd1 vccd1 vccd1 _4714_/B sky130_fd_sc_hd__xnor2_2
X_5693_ _3732_/A _5692_/B _5692_/Y _3194_/Y vssd1 vssd1 vccd1 vccd1 _5693_/X sky130_fd_sc_hd__a211o_1
XFILLER_30_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4644_ _4644_/A _4644_/B vssd1 vssd1 vccd1 vccd1 _4644_/Y sky130_fd_sc_hd__nor2_4
XFILLER_135_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4575_ _6181_/Q _4574_/X _4575_/S vssd1 vssd1 vccd1 vccd1 _4576_/B sky130_fd_sc_hd__mux2_1
X_3526_ _3526_/A _3526_/B vssd1 vssd1 vccd1 vccd1 _3937_/D sky130_fd_sc_hd__xnor2_4
XFILLER_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5829__A1 _3529_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6245_ _6254_/CLK _6245_/D vssd1 vssd1 vccd1 vccd1 _6245_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3457_ _6204_/Q _3458_/B vssd1 vssd1 vccd1 vccd1 _3518_/A sky130_fd_sc_hd__nand2_1
XFILLER_103_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4501__A1 _5790_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6176_ _6176_/CLK _6176_/D vssd1 vssd1 vccd1 vccd1 _6176_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3388_ _3388_/A _3388_/B _3500_/A vssd1 vssd1 vccd1 vccd1 _3405_/B sky130_fd_sc_hd__nor3_4
XANTENNA__4685__A1_N _4672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5127_ _5126_/X _6207_/Q _5129_/S vssd1 vssd1 vccd1 vccd1 _6207_/D sky130_fd_sc_hd__mux2_1
XFILLER_112_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_468 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5058_ _5058_/A _5096_/C _5058_/C _5058_/D vssd1 vssd1 vccd1 vccd1 _5059_/C sky130_fd_sc_hd__or4_1
XFILLER_55_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4009_ _5976_/A _4009_/B _4009_/C _4009_/D vssd1 vssd1 vccd1 vccd1 _4009_/X sky130_fd_sc_hd__and4_1
XFILLER_38_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4017__B1 _4767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5517__B1 _5251_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3791__A2 _3740_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4050__S _4596_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4740__B2 _4972_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3174__B _5617_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3190__A _3257_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_55_clk _6133_/CLK vssd1 vssd1 vccd1 vccd1 _6284_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_16_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4733__B _4734_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5205__C1 _5192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5845__A _5845_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5508__B1 _6004_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3365__A _4003_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3534__A2 _5439_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4360_ _6111_/Q _4296_/Y _4359_/Y _4437_/A1 vssd1 vssd1 vccd1 vccd1 _4360_/Y sky130_fd_sc_hd__a22oi_1
XANTENNA__4731__B2 _4886_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3311_ _3316_/B vssd1 vssd1 vccd1 vccd1 _3311_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4291_ _4226_/Y _4230_/X _4330_/A _4290_/X vssd1 vssd1 vccd1 vccd1 _4330_/B sky130_fd_sc_hd__o211ai_4
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6030_ _6263_/CLK _6030_/D vssd1 vssd1 vccd1 vccd1 _6030_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3242_ _3243_/A _5924_/B vssd1 vssd1 vccd1 vccd1 _3242_/X sky130_fd_sc_hd__and2_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3173_ _3741_/B _4842_/B vssd1 vssd1 vccd1 vccd1 _3749_/B sky130_fd_sc_hd__nor2_1
XFILLER_39_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5444__C1 _5251_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4798__A1 _5358_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_46_clk _6230_/CLK vssd1 vssd1 vccd1 vccd1 _6227_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__4798__B2 _4931_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4643__B _4645_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3470__A1 _3312_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5814_ _3631_/B _5801_/B _5801_/Y _6271_/Q vssd1 vssd1 vccd1 vccd1 _5814_/X sky130_fd_sc_hd__a22o_1
XFILLER_62_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5745_ _3943_/C _5744_/X _5791_/A vssd1 vssd1 vccd1 vccd1 _6242_/D sky130_fd_sc_hd__mux2_1
XANTENNA_fanout317_A _3028_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5676_ _4270_/A _5649_/X _5675_/X _5956_/A vssd1 vssd1 vccd1 vccd1 _6236_/D sky130_fd_sc_hd__o211a_1
XFILLER_108_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4627_ _3030_/Y _4812_/S _4659_/B _5703_/A vssd1 vssd1 vccd1 vccd1 _4627_/X sky130_fd_sc_hd__a31o_1
XFILLER_135_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4722__A1 _6221_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4558_ _3942_/B _4564_/A2 _4556_/X _4557_/X vssd1 vssd1 vccd1 vccd1 _6178_/D sky130_fd_sc_hd__a22o_1
XANTENNA__4722__B2 _4931_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3509_ _3512_/A _5707_/B _3922_/S vssd1 vssd1 vccd1 vccd1 _3571_/A sky130_fd_sc_hd__mux2_2
X_4489_ _3942_/D _4501_/A2 _4487_/X _4488_/Y vssd1 vssd1 vccd1 vccd1 _6136_/D sky130_fd_sc_hd__a22o_1
XANTENNA__5278__A2 _4234_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6228_ _6295_/CLK _6228_/D vssd1 vssd1 vccd1 vccd1 _6228_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__3289__A1 _4136_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4818__B _4819_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5683__C1 _3996_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6159_ _6263_/CLK _6159_/D vssd1 vssd1 vccd1 vccd1 _6159_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4789__A1 _3011_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_37_clk clkbuf_3_4__f_clk/X vssd1 vssd1 vccd1 vccd1 _6098_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_122_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4477__A0 _5790_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5674__C1 _5728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_28_clk _6084_/CLK vssd1 vssd1 vccd1 vccd1 _6113_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_64_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3860_ _6057_/Q _5976_/A vssd1 vssd1 vccd1 vccd1 _3860_/X sky130_fd_sc_hd__or2_1
XANTENNA__3079__B _5605_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_32_clk_A clkbuf_3_5__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3791_ _4697_/B _3740_/X _3749_/X _3790_/X vssd1 vssd1 vccd1 vccd1 _3791_/X sky130_fd_sc_hd__a211o_1
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5530_ _5463_/A _5521_/X _5522_/Y _4596_/D _5072_/C vssd1 vssd1 vccd1 vccd1 _5531_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3807__B _3807_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5461_ _5507_/A _5459_/X _5460_/X _5454_/Y _3122_/A vssd1 vssd1 vccd1 vccd1 _5461_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_118_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4412_ _4413_/A _4413_/B vssd1 vssd1 vccd1 vccd1 _4412_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_47_clk_A _6230_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5392_ _5392_/A _5392_/B vssd1 vssd1 vccd1 vccd1 _5392_/X sky130_fd_sc_hd__or2_1
XFILLER_126_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4343_ _4343_/A _4371_/A vssd1 vssd1 vccd1 vccd1 _4375_/A sky130_fd_sc_hd__nor2_1
XFILLER_125_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout307 _5800_/A vssd1 vssd1 vccd1 vccd1 _4067_/A sky130_fd_sc_hd__buf_8
XFILLER_113_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout318 _5799_/A vssd1 vssd1 vccd1 vccd1 _4539_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_99_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4468__A0 _5333_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4274_ _4274_/A _4274_/B vssd1 vssd1 vccd1 vccd1 _4277_/A sky130_fd_sc_hd__xnor2_4
Xfanout329 _5599_/B vssd1 vssd1 vccd1 vccd1 _5454_/A sky130_fd_sc_hd__buf_6
XANTENNA__4638__B _4638_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6013_ _6278_/CLK _6013_/D vssd1 vssd1 vccd1 vccd1 _6013_/Q sky130_fd_sc_hd__dfxtp_2
X_3225_ _3555_/B _3745_/B _3229_/C vssd1 vssd1 vccd1 vccd1 _3225_/X sky130_fd_sc_hd__and3_1
XFILLER_39_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3156_ _5840_/A _4622_/B vssd1 vssd1 vccd1 vccd1 _3156_/Y sky130_fd_sc_hd__nand2_4
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4654__A _4654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_19_clk _6084_/CLK vssd1 vssd1 vccd1 vccd1 _6272_/CLK sky130_fd_sc_hd__clkbuf_16
X_3087_ _6215_/Q _6214_/Q _6216_/Q vssd1 vssd1 vccd1 vccd1 _5051_/B sky130_fd_sc_hd__or3b_4
XANTENNA__5968__B1 _6298_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout267_A _4085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3989_ _4608_/C _3945_/B _3205_/A vssd1 vssd1 vccd1 vccd1 _3989_/Y sky130_fd_sc_hd__a21oi_1
X_5728_ _5728_/A _5728_/B _5728_/C _5728_/D vssd1 vssd1 vccd1 vccd1 _5728_/X sky130_fd_sc_hd__or4_2
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5659_ _5734_/A _5283_/A _5656_/Y _5657_/X _5658_/X vssd1 vssd1 vccd1 vccd1 _5659_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_136_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3733__A _3734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout82_A _3102_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3131__A0 _5344_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5671__A2 _5321_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3434__A1 _3599_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5187__B2 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3643__A _3643_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4458__B _4458_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3010_ _5358_/A vssd1 vssd1 vccd1 vccd1 _3010_/Y sky130_fd_sc_hd__clkinv_4
XANTENNA__5662__A2 _5203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5414__A2 _5556_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4961_ _6004_/Q _5454_/B vssd1 vssd1 vccd1 vccd1 _4961_/Y sky130_fd_sc_hd__nand2_1
XFILLER_45_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3912_ _3913_/A _5742_/C vssd1 vssd1 vccd1 vccd1 _3912_/Y sky130_fd_sc_hd__nor2_4
X_4892_ _4924_/A _4892_/B vssd1 vssd1 vccd1 vccd1 _4900_/A sky130_fd_sc_hd__nor2_8
X_3843_ _4214_/A _5943_/A _3590_/X _3765_/X _3772_/X vssd1 vssd1 vccd1 vccd1 _3843_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__4921__B _4979_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3774_ _4657_/A _4619_/A _3810_/S vssd1 vssd1 vccd1 vccd1 _3774_/X sky130_fd_sc_hd__mux2_1
X_5513_ _5513_/A _5513_/B vssd1 vssd1 vccd1 vccd1 _5513_/Y sky130_fd_sc_hd__nor2_1
XFILLER_118_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5444_ _5058_/C _5421_/Y _5435_/X _5443_/X _5251_/Y vssd1 vssd1 vccd1 vccd1 _5444_/X
+ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_8_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _6290_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_105_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5375_ _3122_/A _5291_/Y _5374_/Y _5373_/X vssd1 vssd1 vccd1 vccd1 _5375_/X sky130_fd_sc_hd__a31o_1
XANTENNA__4649__A _5054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout104 _3949_/Y vssd1 vssd1 vccd1 vccd1 _5943_/C sky130_fd_sc_hd__buf_4
X_4326_ _4326_/A _4326_/B vssd1 vssd1 vccd1 vccd1 _4328_/B sky130_fd_sc_hd__nand2_1
Xfanout115 _3410_/B vssd1 vssd1 vccd1 vccd1 _3801_/A sky130_fd_sc_hd__buf_4
Xfanout126 _5714_/B vssd1 vssd1 vccd1 vccd1 _3996_/B sky130_fd_sc_hd__buf_6
XFILLER_113_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout137 _5957_/B vssd1 vssd1 vccd1 vccd1 _4638_/B sky130_fd_sc_hd__clkbuf_16
Xfanout148 _5456_/S vssd1 vssd1 vccd1 vccd1 _5543_/S sky130_fd_sc_hd__buf_6
XANTENNA__5102__A1 _5957_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4257_ _6098_/Q _3724_/X _4259_/S vssd1 vssd1 vccd1 vccd1 _6098_/D sky130_fd_sc_hd__mux2_1
Xfanout159 _3050_/X vssd1 vssd1 vccd1 vccd1 _3060_/A sky130_fd_sc_hd__buf_6
XFILLER_101_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3208_ _5703_/A _3228_/A _3741_/B _4886_/B vssd1 vssd1 vccd1 vccd1 _3210_/C sky130_fd_sc_hd__or4_4
X_4188_ _4153_/X _4157_/A _4193_/A _4187_/X vssd1 vssd1 vccd1 vccd1 _4193_/B sky130_fd_sc_hd__a211oi_4
XANTENNA__3699__S _3902_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3139_ _3732_/A _3555_/B vssd1 vssd1 vccd1 vccd1 _3228_/A sky130_fd_sc_hd__nand2_1
XFILLER_103_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4613__B1 _5638_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5943__A _5943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3888__D1 _5943_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5629__C1 _3950_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3182__B _3996_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4852__B1 _3116_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3910__B _5766_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4294__A _5818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_728 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4907__A1 _5454_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3357__B _3388_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5853__A _5853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3490_ _5818_/A _3555_/B _3490_/C vssd1 vssd1 vccd1 vccd1 _3492_/B sky130_fd_sc_hd__and3_4
XFILLER_5_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3373__A _3511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5160_ _3014_/A _3105_/A _5156_/X _5159_/X vssd1 vssd1 vccd1 vccd1 _5161_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4111_ _4270_/A _4111_/B vssd1 vssd1 vccd1 vccd1 _4115_/A sky130_fd_sc_hd__nand2_2
X_5091_ _6198_/Q _5870_/A _3672_/Y _5051_/D vssd1 vssd1 vccd1 vccd1 _5091_/X sky130_fd_sc_hd__a31o_1
XFILLER_96_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4042_ _6063_/Q _3724_/X _4044_/S vssd1 vssd1 vccd1 vccd1 _6063_/D sky130_fd_sc_hd__mux2_1
XFILLER_56_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5399__A1 _4645_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5993_ _6107_/Q vssd1 vssd1 vccd1 vccd1 _6107_/D sky130_fd_sc_hd__clkbuf_2
X_4944_ _4943_/A _4943_/B _4914_/B _4972_/A vssd1 vssd1 vccd1 vccd1 _4944_/X sky130_fd_sc_hd__o31a_2
XFILLER_33_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4875_ _4840_/A _4838_/B _4840_/B _4836_/X vssd1 vssd1 vccd1 vccd1 _4879_/A sky130_fd_sc_hd__a31o_1
XANTENNA__3548__A _3567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3826_ _4202_/A _3777_/S _3825_/X _3751_/A vssd1 vssd1 vccd1 vccd1 _3826_/X sky130_fd_sc_hd__o211a_1
XANTENNA_fanout132_A _3084_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3267__B _3267_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5571__A1 _5551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3757_ _3986_/A _3738_/X _3801_/B _3756_/X vssd1 vssd1 vccd1 vccd1 _3757_/X sky130_fd_sc_hd__o211a_1
XFILLER_119_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3582__B1 _3422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3688_ _3943_/C _3686_/X _3705_/A vssd1 vssd1 vccd1 vccd1 _6019_/D sky130_fd_sc_hd__mux2_1
XFILLER_133_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5323__A1 _5412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5427_ _5452_/A vssd1 vssd1 vccd1 vccd1 _5427_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3334__A0 _3387_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5358_ _5358_/A _5387_/C vssd1 vssd1 vccd1 vccd1 _5358_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_59_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4309_ _4410_/B _4309_/B vssd1 vssd1 vccd1 vccd1 _4343_/A sky130_fd_sc_hd__nand2_2
XFILLER_59_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5289_ _5292_/B _5251_/A _5287_/Y _5288_/Y _5948_/A vssd1 vssd1 vccd1 vccd1 _6220_/D
+ sky130_fd_sc_hd__o221a_1
XANTENNA__5087__B1 _4648_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3637__A1 _5207_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout45_A _5556_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4842__A _4850_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4062__A1 _3718_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5392__B _5392_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5314__A1 _4638_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3193__A _3312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3628__A1 _3145_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4825__B1 _4648_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3132__S _3135_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4053__A1 _4819_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3800__A1 _3443_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4660_ _4660_/A _4660_/B vssd1 vssd1 vccd1 vccd1 _4660_/X sky130_fd_sc_hd__xor2_1
XFILLER_9_87 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3611_ _3611_/A _3611_/B vssd1 vssd1 vccd1 vccd1 _3611_/X sky130_fd_sc_hd__or2_1
XANTENNA__5553__A1 _3432_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5553__B2 _5943_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4591_ _5095_/A _5870_/B _4589_/A _5104_/B vssd1 vssd1 vccd1 vccd1 _4618_/A sky130_fd_sc_hd__o22ai_2
XANTENNA__5583__A _6232_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3564__A0 _5703_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3542_ _5707_/B _3599_/B _3597_/B vssd1 vssd1 vccd1 vccd1 _3607_/A sky130_fd_sc_hd__and3_2
XFILLER_116_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6261_ _6263_/CLK _6261_/D vssd1 vssd1 vccd1 vccd1 _6261_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3473_ _3422_/A _3926_/C _3472_/X vssd1 vssd1 vccd1 vccd1 _5677_/B sky130_fd_sc_hd__a21oi_4
XFILLER_115_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5212_ _4633_/B _5330_/B _5456_/S _4974_/A _3060_/A vssd1 vssd1 vccd1 vccd1 _5217_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_103_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6192_ _6288_/CLK _6192_/D vssd1 vssd1 vccd1 vccd1 _6192_/Q sky130_fd_sc_hd__dfxtp_4
X_5143_ _5143_/A _5143_/B vssd1 vssd1 vccd1 vccd1 _5143_/Y sky130_fd_sc_hd__nor2_1
XFILLER_97_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5608__A2 _5599_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5074_ _5074_/A vssd1 vssd1 vccd1 vccd1 _5074_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4646__B _5403_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4025_ _5148_/A _4025_/B vssd1 vssd1 vccd1 vccd1 _4025_/Y sky130_fd_sc_hd__nor2_1
XFILLER_65_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4662__A _5263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4044__A1 _3730_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout347_A _5264_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5976_ _5976_/A _5976_/B _5976_/C _5976_/D vssd1 vssd1 vccd1 vccd1 _5985_/C sky130_fd_sc_hd__or4_4
XFILLER_52_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5792__A1 _3711_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4927_ _4783_/Y _4926_/Y _4924_/X vssd1 vssd1 vccd1 vccd1 _4929_/B sky130_fd_sc_hd__a21o_1
XANTENNA__4595__A2 _4003_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4858_ _4872_/A _4979_/B vssd1 vssd1 vccd1 vccd1 _4925_/C sky130_fd_sc_hd__nor2_4
XFILLER_20_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3809_ _6037_/Q _3771_/X _3807_/Y _3808_/X vssd1 vssd1 vccd1 vccd1 _6037_/D sky130_fd_sc_hd__a211o_1
XANTENNA__5544__B2 _3121_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4789_ _3011_/Y _3033_/Y _4755_/B vssd1 vssd1 vccd1 vccd1 _4791_/C sky130_fd_sc_hd__a21o_1
XFILLER_109_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4837__A _5428_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3741__A _5703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5232__B1 _5767_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5783__A1 _5387_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3188__A _5730_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5535__A1 _5540_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5299__B1 _5653_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4747__A _5333_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_723 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5578__A _6232_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5830_ _5835_/A1 _4420_/X _5819_/Y _6278_/Q vssd1 vssd1 vccd1 vccd1 _5830_/X sky130_fd_sc_hd__a22o_1
XFILLER_61_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4026__A1 _5790_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5761_ _5446_/B _6248_/Q _5761_/S vssd1 vssd1 vccd1 vccd1 _5761_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5774__A1 _5305_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3098__A _5731_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4712_ _4678_/A _4673_/B _4710_/A vssd1 vssd1 vccd1 vccd1 _4713_/B sky130_fd_sc_hd__o21a_1
XFILLER_30_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5692_ _6301_/Q _5692_/B vssd1 vssd1 vccd1 vccd1 _5692_/Y sky130_fd_sc_hd__nor2_1
XFILLER_30_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5526__A1 _3059_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4643_ _4643_/A _4645_/B vssd1 vssd1 vccd1 vccd1 _4643_/Y sky130_fd_sc_hd__nand2_1
XFILLER_116_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4574_ _3958_/A _3112_/B _3114_/B _4046_/A vssd1 vssd1 vccd1 vccd1 _4574_/X sky130_fd_sc_hd__a22o_1
X_3525_ _3960_/B _3571_/B _3524_/X vssd1 vssd1 vccd1 vccd1 _3526_/B sky130_fd_sc_hd__o21ai_4
X_6244_ _6254_/CLK _6244_/D vssd1 vssd1 vccd1 vccd1 _6244_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3456_ _6204_/Q _3458_/B vssd1 vssd1 vccd1 vccd1 _3456_/X sky130_fd_sc_hd__and2_1
XFILLER_103_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6175_ _6284_/CLK _6175_/D vssd1 vssd1 vccd1 vccd1 _6175_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4657__A _4657_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3387_ _3387_/A _3500_/A _3500_/B vssd1 vssd1 vccd1 vccd1 _3387_/X sky130_fd_sc_hd__and3_2
XANTENNA__5252__S _5513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout297_A _6071_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5126_ _5862_/A _4846_/A _5128_/S vssd1 vssd1 vccd1 vccd1 _5126_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5057_ _5136_/C _5638_/A vssd1 vssd1 vccd1 vccd1 _5058_/D sky130_fd_sc_hd__nand2_2
XFILLER_72_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4008_ _6066_/Q _4009_/B vssd1 vssd1 vccd1 vccd1 _4008_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5488__A _5488_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4017__A1 _6302_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4017__B2 _6301_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5765__A1 _5790_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5959_ _5959_/A _5959_/B vssd1 vssd1 vccd1 vccd1 _5976_/C sky130_fd_sc_hd__nor2_1
XFILLER_40_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3776__A0 _3450_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5517__A1 _5595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3736__A _3736_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4567__A _5097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3700__A0 _3942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3190__B _3869_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4256__A1 _3721_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5756__A1 _3010_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3767__B1 _5932_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5508__A1 _6003_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3646__A _3986_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4241__S _4246_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3310_ _3310_/A _5889_/A vssd1 vssd1 vccd1 vccd1 _3316_/B sky130_fd_sc_hd__xor2_4
X_4290_ _4326_/B _4289_/B _4289_/C vssd1 vssd1 vccd1 vccd1 _4290_/X sky130_fd_sc_hd__a21o_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3241_ _3241_/A _3241_/B vssd1 vssd1 vccd1 vccd1 _3241_/Y sky130_fd_sc_hd__nand2_4
XFILLER_98_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4495__A1 _3942_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3172_ _6200_/Q _6199_/Q vssd1 vssd1 vccd1 vccd1 _3172_/X sky130_fd_sc_hd__or2_1
XFILLER_67_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_6_clk_A clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4798__A2 _5871_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5813_ _5817_/A1 _4157_/X _5812_/X vssd1 vssd1 vccd1 vccd1 _6270_/D sky130_fd_sc_hd__a21o_1
XFILLER_34_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5747__A1 _5292_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5744_ _5768_/A0 _6242_/Q _5761_/S vssd1 vssd1 vccd1 vccd1 _5744_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5675_ _5675_/A _5675_/B _5675_/C vssd1 vssd1 vccd1 vccd1 _5675_/X sky130_fd_sc_hd__or3_2
XFILLER_135_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4626_ _4812_/S _4659_/B _3030_/Y vssd1 vssd1 vccd1 vccd1 _4626_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA_fanout212_A _3025_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4557_ _5385_/A _4252_/A _4239_/B vssd1 vssd1 vccd1 vccd1 _4557_/X sky130_fd_sc_hd__o21a_1
XANTENNA__4722__A2 _4872_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3508_ _3646_/B _3513_/B _3504_/Y _3611_/A _3507_/Y vssd1 vssd1 vccd1 vccd1 _4767_/B
+ sky130_fd_sc_hd__o221a_4
X_4488_ _3011_/Y _4499_/B _4501_/A2 vssd1 vssd1 vccd1 vccd1 _4488_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_103_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6227_ _6227_/CLK _6227_/D vssd1 vssd1 vccd1 vccd1 _6227_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__4387__A _4410_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3439_ _4163_/A _3257_/B _5367_/B _3885_/A vssd1 vssd1 vccd1 vccd1 _3444_/A sky130_fd_sc_hd__a22o_4
XANTENNA__4486__A1 _5926_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5683__B1 _3513_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6158_ _6263_/CLK _6158_/D vssd1 vssd1 vccd1 vccd1 _6158_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5109_ _5109_/A _5124_/S vssd1 vssd1 vccd1 vccd1 _5110_/B sky130_fd_sc_hd__or2_1
X_6089_ _6098_/CLK _6089_/D vssd1 vssd1 vccd1 vccd1 _6089_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5710__S _5710_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4789__A2 _3033_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5011__A _5509_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4850__A _4850_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4061__S _4066_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3185__B _3736_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5910__A1 _4826_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5910__B2 _5551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput30 _6283_/Q vssd1 vssd1 vccd1 vccd1 io_out[2] sky130_fd_sc_hd__buf_4
XANTENNA__3913__B _5742_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5674__B1 _5203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5977__A1 _4850_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4744__B _4744_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_578 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5729__A1 _4214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5856__A _5856_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3790_ _4162_/B _3777_/S _3789_/X _3751_/A vssd1 vssd1 vccd1 vccd1 _3790_/X sky130_fd_sc_hd__o211a_1
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5460_ _5454_/B _5453_/Y _5227_/Y vssd1 vssd1 vccd1 vccd1 _5460_/X sky130_fd_sc_hd__a21bo_1
XFILLER_8_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3095__B _4705_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4411_ _4411_/A _4411_/B vssd1 vssd1 vccd1 vccd1 _4413_/B sky130_fd_sc_hd__nor2_4
XANTENNA__5362__C1 _5227_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5901__A1 _5226_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5391_ _5391_/A vssd1 vssd1 vccd1 vccd1 _5391_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4342_ _4426_/A _4342_/B vssd1 vssd1 vccd1 vccd1 _4371_/A sky130_fd_sc_hd__nand2_4
XFILLER_125_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout308 _6066_/Q vssd1 vssd1 vccd1 vccd1 _5800_/A sky130_fd_sc_hd__buf_6
Xfanout319 _5799_/A vssd1 vssd1 vccd1 vccd1 _5948_/A sky130_fd_sc_hd__buf_4
XFILLER_59_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4273_ _4301_/A _4389_/B vssd1 vssd1 vccd1 vccd1 _4274_/B sky130_fd_sc_hd__nand2_2
XFILLER_101_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5665__A0 _4697_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6012_ _6041_/CLK _6012_/D vssd1 vssd1 vccd1 vccd1 _6012_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_98_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3224_ _5124_/S _3706_/A vssd1 vssd1 vccd1 vccd1 _3229_/C sky130_fd_sc_hd__nor2_1
XANTENNA__3542__C _3597_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
.ends

